

module kernel0_fsm
(
  ap_clk,
  ap_rst_n,
  ap_start,
  ap_ready,
  ap_done,
  ap_idle,
  A,
  B,
  C,
  A_IO_L2_in_0__ap_start,
  A_IO_L2_in_0__ap_ready,
  A_IO_L2_in_0__ap_done,
  A_IO_L2_in_0__ap_idle,
  A_IO_L2_in_1__ap_start,
  A_IO_L2_in_1__ap_ready,
  A_IO_L2_in_1__ap_done,
  A_IO_L2_in_1__ap_idle,
  A_IO_L2_in_2__ap_start,
  A_IO_L2_in_2__ap_ready,
  A_IO_L2_in_2__ap_done,
  A_IO_L2_in_2__ap_idle,
  A_IO_L2_in_3__ap_start,
  A_IO_L2_in_3__ap_ready,
  A_IO_L2_in_3__ap_done,
  A_IO_L2_in_3__ap_idle,
  A_IO_L2_in_4__ap_start,
  A_IO_L2_in_4__ap_ready,
  A_IO_L2_in_4__ap_done,
  A_IO_L2_in_4__ap_idle,
  A_IO_L2_in_5__ap_start,
  A_IO_L2_in_5__ap_ready,
  A_IO_L2_in_5__ap_done,
  A_IO_L2_in_5__ap_idle,
  A_IO_L2_in_6__ap_start,
  A_IO_L2_in_6__ap_ready,
  A_IO_L2_in_6__ap_done,
  A_IO_L2_in_6__ap_idle,
  A_IO_L2_in_7__ap_start,
  A_IO_L2_in_7__ap_ready,
  A_IO_L2_in_7__ap_done,
  A_IO_L2_in_7__ap_idle,
  A_IO_L2_in_8__ap_start,
  A_IO_L2_in_8__ap_ready,
  A_IO_L2_in_8__ap_done,
  A_IO_L2_in_8__ap_idle,
  A_IO_L2_in_9__ap_start,
  A_IO_L2_in_9__ap_ready,
  A_IO_L2_in_9__ap_done,
  A_IO_L2_in_9__ap_idle,
  A_IO_L2_in_10__ap_start,
  A_IO_L2_in_10__ap_ready,
  A_IO_L2_in_10__ap_done,
  A_IO_L2_in_10__ap_idle,
  A_IO_L2_in_11__ap_start,
  A_IO_L2_in_11__ap_ready,
  A_IO_L2_in_11__ap_done,
  A_IO_L2_in_11__ap_idle,
  A_IO_L2_in_12__ap_start,
  A_IO_L2_in_12__ap_ready,
  A_IO_L2_in_12__ap_done,
  A_IO_L2_in_12__ap_idle,
  A_IO_L2_in_13__ap_start,
  A_IO_L2_in_13__ap_ready,
  A_IO_L2_in_13__ap_done,
  A_IO_L2_in_13__ap_idle,
  A_IO_L2_in_14__ap_start,
  A_IO_L2_in_14__ap_ready,
  A_IO_L2_in_14__ap_done,
  A_IO_L2_in_14__ap_idle,
  A_IO_L2_in_15__ap_start,
  A_IO_L2_in_15__ap_ready,
  A_IO_L2_in_15__ap_done,
  A_IO_L2_in_15__ap_idle,
  A_IO_L2_in_16__ap_start,
  A_IO_L2_in_16__ap_ready,
  A_IO_L2_in_16__ap_done,
  A_IO_L2_in_16__ap_idle,
  A_IO_L2_in_boundary_0__ap_start,
  A_IO_L2_in_boundary_0__ap_ready,
  A_IO_L2_in_boundary_0__ap_done,
  A_IO_L2_in_boundary_0__ap_idle,
  A_IO_L3_in_0__ap_start,
  A_IO_L3_in_0__ap_ready,
  A_IO_L3_in_0__ap_done,
  A_IO_L3_in_0__ap_idle,
  A_IO_L3_in_serialize_0___A__q0,
  A_IO_L3_in_serialize_0__ap_start,
  A_IO_L3_in_serialize_0__ap_ready,
  A_IO_L3_in_serialize_0__ap_done,
  A_IO_L3_in_serialize_0__ap_idle,
  A_PE_dummy_in_0__ap_start,
  A_PE_dummy_in_0__ap_ready,
  A_PE_dummy_in_0__ap_done,
  A_PE_dummy_in_0__ap_idle,
  A_PE_dummy_in_1__ap_start,
  A_PE_dummy_in_1__ap_ready,
  A_PE_dummy_in_1__ap_done,
  A_PE_dummy_in_1__ap_idle,
  A_PE_dummy_in_2__ap_start,
  A_PE_dummy_in_2__ap_ready,
  A_PE_dummy_in_2__ap_done,
  A_PE_dummy_in_2__ap_idle,
  A_PE_dummy_in_3__ap_start,
  A_PE_dummy_in_3__ap_ready,
  A_PE_dummy_in_3__ap_done,
  A_PE_dummy_in_3__ap_idle,
  A_PE_dummy_in_4__ap_start,
  A_PE_dummy_in_4__ap_ready,
  A_PE_dummy_in_4__ap_done,
  A_PE_dummy_in_4__ap_idle,
  A_PE_dummy_in_5__ap_start,
  A_PE_dummy_in_5__ap_ready,
  A_PE_dummy_in_5__ap_done,
  A_PE_dummy_in_5__ap_idle,
  A_PE_dummy_in_6__ap_start,
  A_PE_dummy_in_6__ap_ready,
  A_PE_dummy_in_6__ap_done,
  A_PE_dummy_in_6__ap_idle,
  A_PE_dummy_in_7__ap_start,
  A_PE_dummy_in_7__ap_ready,
  A_PE_dummy_in_7__ap_done,
  A_PE_dummy_in_7__ap_idle,
  A_PE_dummy_in_8__ap_start,
  A_PE_dummy_in_8__ap_ready,
  A_PE_dummy_in_8__ap_done,
  A_PE_dummy_in_8__ap_idle,
  A_PE_dummy_in_9__ap_start,
  A_PE_dummy_in_9__ap_ready,
  A_PE_dummy_in_9__ap_done,
  A_PE_dummy_in_9__ap_idle,
  A_PE_dummy_in_10__ap_start,
  A_PE_dummy_in_10__ap_ready,
  A_PE_dummy_in_10__ap_done,
  A_PE_dummy_in_10__ap_idle,
  A_PE_dummy_in_11__ap_start,
  A_PE_dummy_in_11__ap_ready,
  A_PE_dummy_in_11__ap_done,
  A_PE_dummy_in_11__ap_idle,
  A_PE_dummy_in_12__ap_start,
  A_PE_dummy_in_12__ap_ready,
  A_PE_dummy_in_12__ap_done,
  A_PE_dummy_in_12__ap_idle,
  A_PE_dummy_in_13__ap_start,
  A_PE_dummy_in_13__ap_ready,
  A_PE_dummy_in_13__ap_done,
  A_PE_dummy_in_13__ap_idle,
  A_PE_dummy_in_14__ap_start,
  A_PE_dummy_in_14__ap_ready,
  A_PE_dummy_in_14__ap_done,
  A_PE_dummy_in_14__ap_idle,
  A_PE_dummy_in_15__ap_start,
  A_PE_dummy_in_15__ap_ready,
  A_PE_dummy_in_15__ap_done,
  A_PE_dummy_in_15__ap_idle,
  A_PE_dummy_in_16__ap_start,
  A_PE_dummy_in_16__ap_ready,
  A_PE_dummy_in_16__ap_done,
  A_PE_dummy_in_16__ap_idle,
  A_PE_dummy_in_17__ap_start,
  A_PE_dummy_in_17__ap_ready,
  A_PE_dummy_in_17__ap_done,
  A_PE_dummy_in_17__ap_idle,
  B_IO_L2_in_0__ap_start,
  B_IO_L2_in_0__ap_ready,
  B_IO_L2_in_0__ap_done,
  B_IO_L2_in_0__ap_idle,
  B_IO_L2_in_1__ap_start,
  B_IO_L2_in_1__ap_ready,
  B_IO_L2_in_1__ap_done,
  B_IO_L2_in_1__ap_idle,
  B_IO_L2_in_2__ap_start,
  B_IO_L2_in_2__ap_ready,
  B_IO_L2_in_2__ap_done,
  B_IO_L2_in_2__ap_idle,
  B_IO_L2_in_3__ap_start,
  B_IO_L2_in_3__ap_ready,
  B_IO_L2_in_3__ap_done,
  B_IO_L2_in_3__ap_idle,
  B_IO_L2_in_4__ap_start,
  B_IO_L2_in_4__ap_ready,
  B_IO_L2_in_4__ap_done,
  B_IO_L2_in_4__ap_idle,
  B_IO_L2_in_5__ap_start,
  B_IO_L2_in_5__ap_ready,
  B_IO_L2_in_5__ap_done,
  B_IO_L2_in_5__ap_idle,
  B_IO_L2_in_6__ap_start,
  B_IO_L2_in_6__ap_ready,
  B_IO_L2_in_6__ap_done,
  B_IO_L2_in_6__ap_idle,
  B_IO_L2_in_7__ap_start,
  B_IO_L2_in_7__ap_ready,
  B_IO_L2_in_7__ap_done,
  B_IO_L2_in_7__ap_idle,
  B_IO_L2_in_8__ap_start,
  B_IO_L2_in_8__ap_ready,
  B_IO_L2_in_8__ap_done,
  B_IO_L2_in_8__ap_idle,
  B_IO_L2_in_9__ap_start,
  B_IO_L2_in_9__ap_ready,
  B_IO_L2_in_9__ap_done,
  B_IO_L2_in_9__ap_idle,
  B_IO_L2_in_10__ap_start,
  B_IO_L2_in_10__ap_ready,
  B_IO_L2_in_10__ap_done,
  B_IO_L2_in_10__ap_idle,
  B_IO_L2_in_11__ap_start,
  B_IO_L2_in_11__ap_ready,
  B_IO_L2_in_11__ap_done,
  B_IO_L2_in_11__ap_idle,
  B_IO_L2_in_12__ap_start,
  B_IO_L2_in_12__ap_ready,
  B_IO_L2_in_12__ap_done,
  B_IO_L2_in_12__ap_idle,
  B_IO_L2_in_13__ap_start,
  B_IO_L2_in_13__ap_ready,
  B_IO_L2_in_13__ap_done,
  B_IO_L2_in_13__ap_idle,
  B_IO_L2_in_14__ap_start,
  B_IO_L2_in_14__ap_ready,
  B_IO_L2_in_14__ap_done,
  B_IO_L2_in_14__ap_idle,
  B_IO_L2_in_15__ap_start,
  B_IO_L2_in_15__ap_ready,
  B_IO_L2_in_15__ap_done,
  B_IO_L2_in_15__ap_idle,
  B_IO_L2_in_boundary_0__ap_start,
  B_IO_L2_in_boundary_0__ap_ready,
  B_IO_L2_in_boundary_0__ap_done,
  B_IO_L2_in_boundary_0__ap_idle,
  B_IO_L3_in_0__ap_start,
  B_IO_L3_in_0__ap_ready,
  B_IO_L3_in_0__ap_done,
  B_IO_L3_in_0__ap_idle,
  B_IO_L3_in_serialize_0___B__q0,
  B_IO_L3_in_serialize_0__ap_start,
  B_IO_L3_in_serialize_0__ap_ready,
  B_IO_L3_in_serialize_0__ap_done,
  B_IO_L3_in_serialize_0__ap_idle,
  B_PE_dummy_in_0__ap_start,
  B_PE_dummy_in_0__ap_ready,
  B_PE_dummy_in_0__ap_done,
  B_PE_dummy_in_0__ap_idle,
  B_PE_dummy_in_1__ap_start,
  B_PE_dummy_in_1__ap_ready,
  B_PE_dummy_in_1__ap_done,
  B_PE_dummy_in_1__ap_idle,
  B_PE_dummy_in_2__ap_start,
  B_PE_dummy_in_2__ap_ready,
  B_PE_dummy_in_2__ap_done,
  B_PE_dummy_in_2__ap_idle,
  B_PE_dummy_in_3__ap_start,
  B_PE_dummy_in_3__ap_ready,
  B_PE_dummy_in_3__ap_done,
  B_PE_dummy_in_3__ap_idle,
  B_PE_dummy_in_4__ap_start,
  B_PE_dummy_in_4__ap_ready,
  B_PE_dummy_in_4__ap_done,
  B_PE_dummy_in_4__ap_idle,
  B_PE_dummy_in_5__ap_start,
  B_PE_dummy_in_5__ap_ready,
  B_PE_dummy_in_5__ap_done,
  B_PE_dummy_in_5__ap_idle,
  B_PE_dummy_in_6__ap_start,
  B_PE_dummy_in_6__ap_ready,
  B_PE_dummy_in_6__ap_done,
  B_PE_dummy_in_6__ap_idle,
  B_PE_dummy_in_7__ap_start,
  B_PE_dummy_in_7__ap_ready,
  B_PE_dummy_in_7__ap_done,
  B_PE_dummy_in_7__ap_idle,
  B_PE_dummy_in_8__ap_start,
  B_PE_dummy_in_8__ap_ready,
  B_PE_dummy_in_8__ap_done,
  B_PE_dummy_in_8__ap_idle,
  B_PE_dummy_in_9__ap_start,
  B_PE_dummy_in_9__ap_ready,
  B_PE_dummy_in_9__ap_done,
  B_PE_dummy_in_9__ap_idle,
  B_PE_dummy_in_10__ap_start,
  B_PE_dummy_in_10__ap_ready,
  B_PE_dummy_in_10__ap_done,
  B_PE_dummy_in_10__ap_idle,
  B_PE_dummy_in_11__ap_start,
  B_PE_dummy_in_11__ap_ready,
  B_PE_dummy_in_11__ap_done,
  B_PE_dummy_in_11__ap_idle,
  B_PE_dummy_in_12__ap_start,
  B_PE_dummy_in_12__ap_ready,
  B_PE_dummy_in_12__ap_done,
  B_PE_dummy_in_12__ap_idle,
  B_PE_dummy_in_13__ap_start,
  B_PE_dummy_in_13__ap_ready,
  B_PE_dummy_in_13__ap_done,
  B_PE_dummy_in_13__ap_idle,
  B_PE_dummy_in_14__ap_start,
  B_PE_dummy_in_14__ap_ready,
  B_PE_dummy_in_14__ap_done,
  B_PE_dummy_in_14__ap_idle,
  B_PE_dummy_in_15__ap_start,
  B_PE_dummy_in_15__ap_ready,
  B_PE_dummy_in_15__ap_done,
  B_PE_dummy_in_15__ap_idle,
  B_PE_dummy_in_16__ap_start,
  B_PE_dummy_in_16__ap_ready,
  B_PE_dummy_in_16__ap_done,
  B_PE_dummy_in_16__ap_idle,
  C_drain_IO_L1_out_boundary_wrapper_0__ap_start,
  C_drain_IO_L1_out_boundary_wrapper_0__ap_ready,
  C_drain_IO_L1_out_boundary_wrapper_0__ap_done,
  C_drain_IO_L1_out_boundary_wrapper_0__ap_idle,
  C_drain_IO_L1_out_boundary_wrapper_1__ap_start,
  C_drain_IO_L1_out_boundary_wrapper_1__ap_ready,
  C_drain_IO_L1_out_boundary_wrapper_1__ap_done,
  C_drain_IO_L1_out_boundary_wrapper_1__ap_idle,
  C_drain_IO_L1_out_boundary_wrapper_2__ap_start,
  C_drain_IO_L1_out_boundary_wrapper_2__ap_ready,
  C_drain_IO_L1_out_boundary_wrapper_2__ap_done,
  C_drain_IO_L1_out_boundary_wrapper_2__ap_idle,
  C_drain_IO_L1_out_boundary_wrapper_3__ap_start,
  C_drain_IO_L1_out_boundary_wrapper_3__ap_ready,
  C_drain_IO_L1_out_boundary_wrapper_3__ap_done,
  C_drain_IO_L1_out_boundary_wrapper_3__ap_idle,
  C_drain_IO_L1_out_boundary_wrapper_4__ap_start,
  C_drain_IO_L1_out_boundary_wrapper_4__ap_ready,
  C_drain_IO_L1_out_boundary_wrapper_4__ap_done,
  C_drain_IO_L1_out_boundary_wrapper_4__ap_idle,
  C_drain_IO_L1_out_boundary_wrapper_5__ap_start,
  C_drain_IO_L1_out_boundary_wrapper_5__ap_ready,
  C_drain_IO_L1_out_boundary_wrapper_5__ap_done,
  C_drain_IO_L1_out_boundary_wrapper_5__ap_idle,
  C_drain_IO_L1_out_boundary_wrapper_6__ap_start,
  C_drain_IO_L1_out_boundary_wrapper_6__ap_ready,
  C_drain_IO_L1_out_boundary_wrapper_6__ap_done,
  C_drain_IO_L1_out_boundary_wrapper_6__ap_idle,
  C_drain_IO_L1_out_boundary_wrapper_7__ap_start,
  C_drain_IO_L1_out_boundary_wrapper_7__ap_ready,
  C_drain_IO_L1_out_boundary_wrapper_7__ap_done,
  C_drain_IO_L1_out_boundary_wrapper_7__ap_idle,
  C_drain_IO_L1_out_boundary_wrapper_8__ap_start,
  C_drain_IO_L1_out_boundary_wrapper_8__ap_ready,
  C_drain_IO_L1_out_boundary_wrapper_8__ap_done,
  C_drain_IO_L1_out_boundary_wrapper_8__ap_idle,
  C_drain_IO_L1_out_boundary_wrapper_9__ap_start,
  C_drain_IO_L1_out_boundary_wrapper_9__ap_ready,
  C_drain_IO_L1_out_boundary_wrapper_9__ap_done,
  C_drain_IO_L1_out_boundary_wrapper_9__ap_idle,
  C_drain_IO_L1_out_boundary_wrapper_10__ap_start,
  C_drain_IO_L1_out_boundary_wrapper_10__ap_ready,
  C_drain_IO_L1_out_boundary_wrapper_10__ap_done,
  C_drain_IO_L1_out_boundary_wrapper_10__ap_idle,
  C_drain_IO_L1_out_boundary_wrapper_11__ap_start,
  C_drain_IO_L1_out_boundary_wrapper_11__ap_ready,
  C_drain_IO_L1_out_boundary_wrapper_11__ap_done,
  C_drain_IO_L1_out_boundary_wrapper_11__ap_idle,
  C_drain_IO_L1_out_boundary_wrapper_12__ap_start,
  C_drain_IO_L1_out_boundary_wrapper_12__ap_ready,
  C_drain_IO_L1_out_boundary_wrapper_12__ap_done,
  C_drain_IO_L1_out_boundary_wrapper_12__ap_idle,
  C_drain_IO_L1_out_boundary_wrapper_13__ap_start,
  C_drain_IO_L1_out_boundary_wrapper_13__ap_ready,
  C_drain_IO_L1_out_boundary_wrapper_13__ap_done,
  C_drain_IO_L1_out_boundary_wrapper_13__ap_idle,
  C_drain_IO_L1_out_boundary_wrapper_14__ap_start,
  C_drain_IO_L1_out_boundary_wrapper_14__ap_ready,
  C_drain_IO_L1_out_boundary_wrapper_14__ap_done,
  C_drain_IO_L1_out_boundary_wrapper_14__ap_idle,
  C_drain_IO_L1_out_boundary_wrapper_15__ap_start,
  C_drain_IO_L1_out_boundary_wrapper_15__ap_ready,
  C_drain_IO_L1_out_boundary_wrapper_15__ap_done,
  C_drain_IO_L1_out_boundary_wrapper_15__ap_idle,
  C_drain_IO_L1_out_boundary_wrapper_16__ap_start,
  C_drain_IO_L1_out_boundary_wrapper_16__ap_ready,
  C_drain_IO_L1_out_boundary_wrapper_16__ap_done,
  C_drain_IO_L1_out_boundary_wrapper_16__ap_idle,
  C_drain_IO_L1_out_wrapper_0__ap_start,
  C_drain_IO_L1_out_wrapper_0__ap_ready,
  C_drain_IO_L1_out_wrapper_0__ap_done,
  C_drain_IO_L1_out_wrapper_0__ap_idle,
  C_drain_IO_L1_out_wrapper_1__ap_start,
  C_drain_IO_L1_out_wrapper_1__ap_ready,
  C_drain_IO_L1_out_wrapper_1__ap_done,
  C_drain_IO_L1_out_wrapper_1__ap_idle,
  C_drain_IO_L1_out_wrapper_2__ap_start,
  C_drain_IO_L1_out_wrapper_2__ap_ready,
  C_drain_IO_L1_out_wrapper_2__ap_done,
  C_drain_IO_L1_out_wrapper_2__ap_idle,
  C_drain_IO_L1_out_wrapper_3__ap_start,
  C_drain_IO_L1_out_wrapper_3__ap_ready,
  C_drain_IO_L1_out_wrapper_3__ap_done,
  C_drain_IO_L1_out_wrapper_3__ap_idle,
  C_drain_IO_L1_out_wrapper_4__ap_start,
  C_drain_IO_L1_out_wrapper_4__ap_ready,
  C_drain_IO_L1_out_wrapper_4__ap_done,
  C_drain_IO_L1_out_wrapper_4__ap_idle,
  C_drain_IO_L1_out_wrapper_5__ap_start,
  C_drain_IO_L1_out_wrapper_5__ap_ready,
  C_drain_IO_L1_out_wrapper_5__ap_done,
  C_drain_IO_L1_out_wrapper_5__ap_idle,
  C_drain_IO_L1_out_wrapper_6__ap_start,
  C_drain_IO_L1_out_wrapper_6__ap_ready,
  C_drain_IO_L1_out_wrapper_6__ap_done,
  C_drain_IO_L1_out_wrapper_6__ap_idle,
  C_drain_IO_L1_out_wrapper_7__ap_start,
  C_drain_IO_L1_out_wrapper_7__ap_ready,
  C_drain_IO_L1_out_wrapper_7__ap_done,
  C_drain_IO_L1_out_wrapper_7__ap_idle,
  C_drain_IO_L1_out_wrapper_8__ap_start,
  C_drain_IO_L1_out_wrapper_8__ap_ready,
  C_drain_IO_L1_out_wrapper_8__ap_done,
  C_drain_IO_L1_out_wrapper_8__ap_idle,
  C_drain_IO_L1_out_wrapper_9__ap_start,
  C_drain_IO_L1_out_wrapper_9__ap_ready,
  C_drain_IO_L1_out_wrapper_9__ap_done,
  C_drain_IO_L1_out_wrapper_9__ap_idle,
  C_drain_IO_L1_out_wrapper_10__ap_start,
  C_drain_IO_L1_out_wrapper_10__ap_ready,
  C_drain_IO_L1_out_wrapper_10__ap_done,
  C_drain_IO_L1_out_wrapper_10__ap_idle,
  C_drain_IO_L1_out_wrapper_11__ap_start,
  C_drain_IO_L1_out_wrapper_11__ap_ready,
  C_drain_IO_L1_out_wrapper_11__ap_done,
  C_drain_IO_L1_out_wrapper_11__ap_idle,
  C_drain_IO_L1_out_wrapper_12__ap_start,
  C_drain_IO_L1_out_wrapper_12__ap_ready,
  C_drain_IO_L1_out_wrapper_12__ap_done,
  C_drain_IO_L1_out_wrapper_12__ap_idle,
  C_drain_IO_L1_out_wrapper_13__ap_start,
  C_drain_IO_L1_out_wrapper_13__ap_ready,
  C_drain_IO_L1_out_wrapper_13__ap_done,
  C_drain_IO_L1_out_wrapper_13__ap_idle,
  C_drain_IO_L1_out_wrapper_14__ap_start,
  C_drain_IO_L1_out_wrapper_14__ap_ready,
  C_drain_IO_L1_out_wrapper_14__ap_done,
  C_drain_IO_L1_out_wrapper_14__ap_idle,
  C_drain_IO_L1_out_wrapper_15__ap_start,
  C_drain_IO_L1_out_wrapper_15__ap_ready,
  C_drain_IO_L1_out_wrapper_15__ap_done,
  C_drain_IO_L1_out_wrapper_15__ap_idle,
  C_drain_IO_L1_out_wrapper_16__ap_start,
  C_drain_IO_L1_out_wrapper_16__ap_ready,
  C_drain_IO_L1_out_wrapper_16__ap_done,
  C_drain_IO_L1_out_wrapper_16__ap_idle,
  C_drain_IO_L1_out_wrapper_17__ap_start,
  C_drain_IO_L1_out_wrapper_17__ap_ready,
  C_drain_IO_L1_out_wrapper_17__ap_done,
  C_drain_IO_L1_out_wrapper_17__ap_idle,
  C_drain_IO_L1_out_wrapper_18__ap_start,
  C_drain_IO_L1_out_wrapper_18__ap_ready,
  C_drain_IO_L1_out_wrapper_18__ap_done,
  C_drain_IO_L1_out_wrapper_18__ap_idle,
  C_drain_IO_L1_out_wrapper_19__ap_start,
  C_drain_IO_L1_out_wrapper_19__ap_ready,
  C_drain_IO_L1_out_wrapper_19__ap_done,
  C_drain_IO_L1_out_wrapper_19__ap_idle,
  C_drain_IO_L1_out_wrapper_20__ap_start,
  C_drain_IO_L1_out_wrapper_20__ap_ready,
  C_drain_IO_L1_out_wrapper_20__ap_done,
  C_drain_IO_L1_out_wrapper_20__ap_idle,
  C_drain_IO_L1_out_wrapper_21__ap_start,
  C_drain_IO_L1_out_wrapper_21__ap_ready,
  C_drain_IO_L1_out_wrapper_21__ap_done,
  C_drain_IO_L1_out_wrapper_21__ap_idle,
  C_drain_IO_L1_out_wrapper_22__ap_start,
  C_drain_IO_L1_out_wrapper_22__ap_ready,
  C_drain_IO_L1_out_wrapper_22__ap_done,
  C_drain_IO_L1_out_wrapper_22__ap_idle,
  C_drain_IO_L1_out_wrapper_23__ap_start,
  C_drain_IO_L1_out_wrapper_23__ap_ready,
  C_drain_IO_L1_out_wrapper_23__ap_done,
  C_drain_IO_L1_out_wrapper_23__ap_idle,
  C_drain_IO_L1_out_wrapper_24__ap_start,
  C_drain_IO_L1_out_wrapper_24__ap_ready,
  C_drain_IO_L1_out_wrapper_24__ap_done,
  C_drain_IO_L1_out_wrapper_24__ap_idle,
  C_drain_IO_L1_out_wrapper_25__ap_start,
  C_drain_IO_L1_out_wrapper_25__ap_ready,
  C_drain_IO_L1_out_wrapper_25__ap_done,
  C_drain_IO_L1_out_wrapper_25__ap_idle,
  C_drain_IO_L1_out_wrapper_26__ap_start,
  C_drain_IO_L1_out_wrapper_26__ap_ready,
  C_drain_IO_L1_out_wrapper_26__ap_done,
  C_drain_IO_L1_out_wrapper_26__ap_idle,
  C_drain_IO_L1_out_wrapper_27__ap_start,
  C_drain_IO_L1_out_wrapper_27__ap_ready,
  C_drain_IO_L1_out_wrapper_27__ap_done,
  C_drain_IO_L1_out_wrapper_27__ap_idle,
  C_drain_IO_L1_out_wrapper_28__ap_start,
  C_drain_IO_L1_out_wrapper_28__ap_ready,
  C_drain_IO_L1_out_wrapper_28__ap_done,
  C_drain_IO_L1_out_wrapper_28__ap_idle,
  C_drain_IO_L1_out_wrapper_29__ap_start,
  C_drain_IO_L1_out_wrapper_29__ap_ready,
  C_drain_IO_L1_out_wrapper_29__ap_done,
  C_drain_IO_L1_out_wrapper_29__ap_idle,
  C_drain_IO_L1_out_wrapper_30__ap_start,
  C_drain_IO_L1_out_wrapper_30__ap_ready,
  C_drain_IO_L1_out_wrapper_30__ap_done,
  C_drain_IO_L1_out_wrapper_30__ap_idle,
  C_drain_IO_L1_out_wrapper_31__ap_start,
  C_drain_IO_L1_out_wrapper_31__ap_ready,
  C_drain_IO_L1_out_wrapper_31__ap_done,
  C_drain_IO_L1_out_wrapper_31__ap_idle,
  C_drain_IO_L1_out_wrapper_32__ap_start,
  C_drain_IO_L1_out_wrapper_32__ap_ready,
  C_drain_IO_L1_out_wrapper_32__ap_done,
  C_drain_IO_L1_out_wrapper_32__ap_idle,
  C_drain_IO_L1_out_wrapper_33__ap_start,
  C_drain_IO_L1_out_wrapper_33__ap_ready,
  C_drain_IO_L1_out_wrapper_33__ap_done,
  C_drain_IO_L1_out_wrapper_33__ap_idle,
  C_drain_IO_L1_out_wrapper_34__ap_start,
  C_drain_IO_L1_out_wrapper_34__ap_ready,
  C_drain_IO_L1_out_wrapper_34__ap_done,
  C_drain_IO_L1_out_wrapper_34__ap_idle,
  C_drain_IO_L1_out_wrapper_35__ap_start,
  C_drain_IO_L1_out_wrapper_35__ap_ready,
  C_drain_IO_L1_out_wrapper_35__ap_done,
  C_drain_IO_L1_out_wrapper_35__ap_idle,
  C_drain_IO_L1_out_wrapper_36__ap_start,
  C_drain_IO_L1_out_wrapper_36__ap_ready,
  C_drain_IO_L1_out_wrapper_36__ap_done,
  C_drain_IO_L1_out_wrapper_36__ap_idle,
  C_drain_IO_L1_out_wrapper_37__ap_start,
  C_drain_IO_L1_out_wrapper_37__ap_ready,
  C_drain_IO_L1_out_wrapper_37__ap_done,
  C_drain_IO_L1_out_wrapper_37__ap_idle,
  C_drain_IO_L1_out_wrapper_38__ap_start,
  C_drain_IO_L1_out_wrapper_38__ap_ready,
  C_drain_IO_L1_out_wrapper_38__ap_done,
  C_drain_IO_L1_out_wrapper_38__ap_idle,
  C_drain_IO_L1_out_wrapper_39__ap_start,
  C_drain_IO_L1_out_wrapper_39__ap_ready,
  C_drain_IO_L1_out_wrapper_39__ap_done,
  C_drain_IO_L1_out_wrapper_39__ap_idle,
  C_drain_IO_L1_out_wrapper_40__ap_start,
  C_drain_IO_L1_out_wrapper_40__ap_ready,
  C_drain_IO_L1_out_wrapper_40__ap_done,
  C_drain_IO_L1_out_wrapper_40__ap_idle,
  C_drain_IO_L1_out_wrapper_41__ap_start,
  C_drain_IO_L1_out_wrapper_41__ap_ready,
  C_drain_IO_L1_out_wrapper_41__ap_done,
  C_drain_IO_L1_out_wrapper_41__ap_idle,
  C_drain_IO_L1_out_wrapper_42__ap_start,
  C_drain_IO_L1_out_wrapper_42__ap_ready,
  C_drain_IO_L1_out_wrapper_42__ap_done,
  C_drain_IO_L1_out_wrapper_42__ap_idle,
  C_drain_IO_L1_out_wrapper_43__ap_start,
  C_drain_IO_L1_out_wrapper_43__ap_ready,
  C_drain_IO_L1_out_wrapper_43__ap_done,
  C_drain_IO_L1_out_wrapper_43__ap_idle,
  C_drain_IO_L1_out_wrapper_44__ap_start,
  C_drain_IO_L1_out_wrapper_44__ap_ready,
  C_drain_IO_L1_out_wrapper_44__ap_done,
  C_drain_IO_L1_out_wrapper_44__ap_idle,
  C_drain_IO_L1_out_wrapper_45__ap_start,
  C_drain_IO_L1_out_wrapper_45__ap_ready,
  C_drain_IO_L1_out_wrapper_45__ap_done,
  C_drain_IO_L1_out_wrapper_45__ap_idle,
  C_drain_IO_L1_out_wrapper_46__ap_start,
  C_drain_IO_L1_out_wrapper_46__ap_ready,
  C_drain_IO_L1_out_wrapper_46__ap_done,
  C_drain_IO_L1_out_wrapper_46__ap_idle,
  C_drain_IO_L1_out_wrapper_47__ap_start,
  C_drain_IO_L1_out_wrapper_47__ap_ready,
  C_drain_IO_L1_out_wrapper_47__ap_done,
  C_drain_IO_L1_out_wrapper_47__ap_idle,
  C_drain_IO_L1_out_wrapper_48__ap_start,
  C_drain_IO_L1_out_wrapper_48__ap_ready,
  C_drain_IO_L1_out_wrapper_48__ap_done,
  C_drain_IO_L1_out_wrapper_48__ap_idle,
  C_drain_IO_L1_out_wrapper_49__ap_start,
  C_drain_IO_L1_out_wrapper_49__ap_ready,
  C_drain_IO_L1_out_wrapper_49__ap_done,
  C_drain_IO_L1_out_wrapper_49__ap_idle,
  C_drain_IO_L1_out_wrapper_50__ap_start,
  C_drain_IO_L1_out_wrapper_50__ap_ready,
  C_drain_IO_L1_out_wrapper_50__ap_done,
  C_drain_IO_L1_out_wrapper_50__ap_idle,
  C_drain_IO_L1_out_wrapper_51__ap_start,
  C_drain_IO_L1_out_wrapper_51__ap_ready,
  C_drain_IO_L1_out_wrapper_51__ap_done,
  C_drain_IO_L1_out_wrapper_51__ap_idle,
  C_drain_IO_L1_out_wrapper_52__ap_start,
  C_drain_IO_L1_out_wrapper_52__ap_ready,
  C_drain_IO_L1_out_wrapper_52__ap_done,
  C_drain_IO_L1_out_wrapper_52__ap_idle,
  C_drain_IO_L1_out_wrapper_53__ap_start,
  C_drain_IO_L1_out_wrapper_53__ap_ready,
  C_drain_IO_L1_out_wrapper_53__ap_done,
  C_drain_IO_L1_out_wrapper_53__ap_idle,
  C_drain_IO_L1_out_wrapper_54__ap_start,
  C_drain_IO_L1_out_wrapper_54__ap_ready,
  C_drain_IO_L1_out_wrapper_54__ap_done,
  C_drain_IO_L1_out_wrapper_54__ap_idle,
  C_drain_IO_L1_out_wrapper_55__ap_start,
  C_drain_IO_L1_out_wrapper_55__ap_ready,
  C_drain_IO_L1_out_wrapper_55__ap_done,
  C_drain_IO_L1_out_wrapper_55__ap_idle,
  C_drain_IO_L1_out_wrapper_56__ap_start,
  C_drain_IO_L1_out_wrapper_56__ap_ready,
  C_drain_IO_L1_out_wrapper_56__ap_done,
  C_drain_IO_L1_out_wrapper_56__ap_idle,
  C_drain_IO_L1_out_wrapper_57__ap_start,
  C_drain_IO_L1_out_wrapper_57__ap_ready,
  C_drain_IO_L1_out_wrapper_57__ap_done,
  C_drain_IO_L1_out_wrapper_57__ap_idle,
  C_drain_IO_L1_out_wrapper_58__ap_start,
  C_drain_IO_L1_out_wrapper_58__ap_ready,
  C_drain_IO_L1_out_wrapper_58__ap_done,
  C_drain_IO_L1_out_wrapper_58__ap_idle,
  C_drain_IO_L1_out_wrapper_59__ap_start,
  C_drain_IO_L1_out_wrapper_59__ap_ready,
  C_drain_IO_L1_out_wrapper_59__ap_done,
  C_drain_IO_L1_out_wrapper_59__ap_idle,
  C_drain_IO_L1_out_wrapper_60__ap_start,
  C_drain_IO_L1_out_wrapper_60__ap_ready,
  C_drain_IO_L1_out_wrapper_60__ap_done,
  C_drain_IO_L1_out_wrapper_60__ap_idle,
  C_drain_IO_L1_out_wrapper_61__ap_start,
  C_drain_IO_L1_out_wrapper_61__ap_ready,
  C_drain_IO_L1_out_wrapper_61__ap_done,
  C_drain_IO_L1_out_wrapper_61__ap_idle,
  C_drain_IO_L1_out_wrapper_62__ap_start,
  C_drain_IO_L1_out_wrapper_62__ap_ready,
  C_drain_IO_L1_out_wrapper_62__ap_done,
  C_drain_IO_L1_out_wrapper_62__ap_idle,
  C_drain_IO_L1_out_wrapper_63__ap_start,
  C_drain_IO_L1_out_wrapper_63__ap_ready,
  C_drain_IO_L1_out_wrapper_63__ap_done,
  C_drain_IO_L1_out_wrapper_63__ap_idle,
  C_drain_IO_L1_out_wrapper_64__ap_start,
  C_drain_IO_L1_out_wrapper_64__ap_ready,
  C_drain_IO_L1_out_wrapper_64__ap_done,
  C_drain_IO_L1_out_wrapper_64__ap_idle,
  C_drain_IO_L1_out_wrapper_65__ap_start,
  C_drain_IO_L1_out_wrapper_65__ap_ready,
  C_drain_IO_L1_out_wrapper_65__ap_done,
  C_drain_IO_L1_out_wrapper_65__ap_idle,
  C_drain_IO_L1_out_wrapper_66__ap_start,
  C_drain_IO_L1_out_wrapper_66__ap_ready,
  C_drain_IO_L1_out_wrapper_66__ap_done,
  C_drain_IO_L1_out_wrapper_66__ap_idle,
  C_drain_IO_L1_out_wrapper_67__ap_start,
  C_drain_IO_L1_out_wrapper_67__ap_ready,
  C_drain_IO_L1_out_wrapper_67__ap_done,
  C_drain_IO_L1_out_wrapper_67__ap_idle,
  C_drain_IO_L1_out_wrapper_68__ap_start,
  C_drain_IO_L1_out_wrapper_68__ap_ready,
  C_drain_IO_L1_out_wrapper_68__ap_done,
  C_drain_IO_L1_out_wrapper_68__ap_idle,
  C_drain_IO_L1_out_wrapper_69__ap_start,
  C_drain_IO_L1_out_wrapper_69__ap_ready,
  C_drain_IO_L1_out_wrapper_69__ap_done,
  C_drain_IO_L1_out_wrapper_69__ap_idle,
  C_drain_IO_L1_out_wrapper_70__ap_start,
  C_drain_IO_L1_out_wrapper_70__ap_ready,
  C_drain_IO_L1_out_wrapper_70__ap_done,
  C_drain_IO_L1_out_wrapper_70__ap_idle,
  C_drain_IO_L1_out_wrapper_71__ap_start,
  C_drain_IO_L1_out_wrapper_71__ap_ready,
  C_drain_IO_L1_out_wrapper_71__ap_done,
  C_drain_IO_L1_out_wrapper_71__ap_idle,
  C_drain_IO_L1_out_wrapper_72__ap_start,
  C_drain_IO_L1_out_wrapper_72__ap_ready,
  C_drain_IO_L1_out_wrapper_72__ap_done,
  C_drain_IO_L1_out_wrapper_72__ap_idle,
  C_drain_IO_L1_out_wrapper_73__ap_start,
  C_drain_IO_L1_out_wrapper_73__ap_ready,
  C_drain_IO_L1_out_wrapper_73__ap_done,
  C_drain_IO_L1_out_wrapper_73__ap_idle,
  C_drain_IO_L1_out_wrapper_74__ap_start,
  C_drain_IO_L1_out_wrapper_74__ap_ready,
  C_drain_IO_L1_out_wrapper_74__ap_done,
  C_drain_IO_L1_out_wrapper_74__ap_idle,
  C_drain_IO_L1_out_wrapper_75__ap_start,
  C_drain_IO_L1_out_wrapper_75__ap_ready,
  C_drain_IO_L1_out_wrapper_75__ap_done,
  C_drain_IO_L1_out_wrapper_75__ap_idle,
  C_drain_IO_L1_out_wrapper_76__ap_start,
  C_drain_IO_L1_out_wrapper_76__ap_ready,
  C_drain_IO_L1_out_wrapper_76__ap_done,
  C_drain_IO_L1_out_wrapper_76__ap_idle,
  C_drain_IO_L1_out_wrapper_77__ap_start,
  C_drain_IO_L1_out_wrapper_77__ap_ready,
  C_drain_IO_L1_out_wrapper_77__ap_done,
  C_drain_IO_L1_out_wrapper_77__ap_idle,
  C_drain_IO_L1_out_wrapper_78__ap_start,
  C_drain_IO_L1_out_wrapper_78__ap_ready,
  C_drain_IO_L1_out_wrapper_78__ap_done,
  C_drain_IO_L1_out_wrapper_78__ap_idle,
  C_drain_IO_L1_out_wrapper_79__ap_start,
  C_drain_IO_L1_out_wrapper_79__ap_ready,
  C_drain_IO_L1_out_wrapper_79__ap_done,
  C_drain_IO_L1_out_wrapper_79__ap_idle,
  C_drain_IO_L1_out_wrapper_80__ap_start,
  C_drain_IO_L1_out_wrapper_80__ap_ready,
  C_drain_IO_L1_out_wrapper_80__ap_done,
  C_drain_IO_L1_out_wrapper_80__ap_idle,
  C_drain_IO_L1_out_wrapper_81__ap_start,
  C_drain_IO_L1_out_wrapper_81__ap_ready,
  C_drain_IO_L1_out_wrapper_81__ap_done,
  C_drain_IO_L1_out_wrapper_81__ap_idle,
  C_drain_IO_L1_out_wrapper_82__ap_start,
  C_drain_IO_L1_out_wrapper_82__ap_ready,
  C_drain_IO_L1_out_wrapper_82__ap_done,
  C_drain_IO_L1_out_wrapper_82__ap_idle,
  C_drain_IO_L1_out_wrapper_83__ap_start,
  C_drain_IO_L1_out_wrapper_83__ap_ready,
  C_drain_IO_L1_out_wrapper_83__ap_done,
  C_drain_IO_L1_out_wrapper_83__ap_idle,
  C_drain_IO_L1_out_wrapper_84__ap_start,
  C_drain_IO_L1_out_wrapper_84__ap_ready,
  C_drain_IO_L1_out_wrapper_84__ap_done,
  C_drain_IO_L1_out_wrapper_84__ap_idle,
  C_drain_IO_L1_out_wrapper_85__ap_start,
  C_drain_IO_L1_out_wrapper_85__ap_ready,
  C_drain_IO_L1_out_wrapper_85__ap_done,
  C_drain_IO_L1_out_wrapper_85__ap_idle,
  C_drain_IO_L1_out_wrapper_86__ap_start,
  C_drain_IO_L1_out_wrapper_86__ap_ready,
  C_drain_IO_L1_out_wrapper_86__ap_done,
  C_drain_IO_L1_out_wrapper_86__ap_idle,
  C_drain_IO_L1_out_wrapper_87__ap_start,
  C_drain_IO_L1_out_wrapper_87__ap_ready,
  C_drain_IO_L1_out_wrapper_87__ap_done,
  C_drain_IO_L1_out_wrapper_87__ap_idle,
  C_drain_IO_L1_out_wrapper_88__ap_start,
  C_drain_IO_L1_out_wrapper_88__ap_ready,
  C_drain_IO_L1_out_wrapper_88__ap_done,
  C_drain_IO_L1_out_wrapper_88__ap_idle,
  C_drain_IO_L1_out_wrapper_89__ap_start,
  C_drain_IO_L1_out_wrapper_89__ap_ready,
  C_drain_IO_L1_out_wrapper_89__ap_done,
  C_drain_IO_L1_out_wrapper_89__ap_idle,
  C_drain_IO_L1_out_wrapper_90__ap_start,
  C_drain_IO_L1_out_wrapper_90__ap_ready,
  C_drain_IO_L1_out_wrapper_90__ap_done,
  C_drain_IO_L1_out_wrapper_90__ap_idle,
  C_drain_IO_L1_out_wrapper_91__ap_start,
  C_drain_IO_L1_out_wrapper_91__ap_ready,
  C_drain_IO_L1_out_wrapper_91__ap_done,
  C_drain_IO_L1_out_wrapper_91__ap_idle,
  C_drain_IO_L1_out_wrapper_92__ap_start,
  C_drain_IO_L1_out_wrapper_92__ap_ready,
  C_drain_IO_L1_out_wrapper_92__ap_done,
  C_drain_IO_L1_out_wrapper_92__ap_idle,
  C_drain_IO_L1_out_wrapper_93__ap_start,
  C_drain_IO_L1_out_wrapper_93__ap_ready,
  C_drain_IO_L1_out_wrapper_93__ap_done,
  C_drain_IO_L1_out_wrapper_93__ap_idle,
  C_drain_IO_L1_out_wrapper_94__ap_start,
  C_drain_IO_L1_out_wrapper_94__ap_ready,
  C_drain_IO_L1_out_wrapper_94__ap_done,
  C_drain_IO_L1_out_wrapper_94__ap_idle,
  C_drain_IO_L1_out_wrapper_95__ap_start,
  C_drain_IO_L1_out_wrapper_95__ap_ready,
  C_drain_IO_L1_out_wrapper_95__ap_done,
  C_drain_IO_L1_out_wrapper_95__ap_idle,
  C_drain_IO_L1_out_wrapper_96__ap_start,
  C_drain_IO_L1_out_wrapper_96__ap_ready,
  C_drain_IO_L1_out_wrapper_96__ap_done,
  C_drain_IO_L1_out_wrapper_96__ap_idle,
  C_drain_IO_L1_out_wrapper_97__ap_start,
  C_drain_IO_L1_out_wrapper_97__ap_ready,
  C_drain_IO_L1_out_wrapper_97__ap_done,
  C_drain_IO_L1_out_wrapper_97__ap_idle,
  C_drain_IO_L1_out_wrapper_98__ap_start,
  C_drain_IO_L1_out_wrapper_98__ap_ready,
  C_drain_IO_L1_out_wrapper_98__ap_done,
  C_drain_IO_L1_out_wrapper_98__ap_idle,
  C_drain_IO_L1_out_wrapper_99__ap_start,
  C_drain_IO_L1_out_wrapper_99__ap_ready,
  C_drain_IO_L1_out_wrapper_99__ap_done,
  C_drain_IO_L1_out_wrapper_99__ap_idle,
  C_drain_IO_L1_out_wrapper_100__ap_start,
  C_drain_IO_L1_out_wrapper_100__ap_ready,
  C_drain_IO_L1_out_wrapper_100__ap_done,
  C_drain_IO_L1_out_wrapper_100__ap_idle,
  C_drain_IO_L1_out_wrapper_101__ap_start,
  C_drain_IO_L1_out_wrapper_101__ap_ready,
  C_drain_IO_L1_out_wrapper_101__ap_done,
  C_drain_IO_L1_out_wrapper_101__ap_idle,
  C_drain_IO_L1_out_wrapper_102__ap_start,
  C_drain_IO_L1_out_wrapper_102__ap_ready,
  C_drain_IO_L1_out_wrapper_102__ap_done,
  C_drain_IO_L1_out_wrapper_102__ap_idle,
  C_drain_IO_L1_out_wrapper_103__ap_start,
  C_drain_IO_L1_out_wrapper_103__ap_ready,
  C_drain_IO_L1_out_wrapper_103__ap_done,
  C_drain_IO_L1_out_wrapper_103__ap_idle,
  C_drain_IO_L1_out_wrapper_104__ap_start,
  C_drain_IO_L1_out_wrapper_104__ap_ready,
  C_drain_IO_L1_out_wrapper_104__ap_done,
  C_drain_IO_L1_out_wrapper_104__ap_idle,
  C_drain_IO_L1_out_wrapper_105__ap_start,
  C_drain_IO_L1_out_wrapper_105__ap_ready,
  C_drain_IO_L1_out_wrapper_105__ap_done,
  C_drain_IO_L1_out_wrapper_105__ap_idle,
  C_drain_IO_L1_out_wrapper_106__ap_start,
  C_drain_IO_L1_out_wrapper_106__ap_ready,
  C_drain_IO_L1_out_wrapper_106__ap_done,
  C_drain_IO_L1_out_wrapper_106__ap_idle,
  C_drain_IO_L1_out_wrapper_107__ap_start,
  C_drain_IO_L1_out_wrapper_107__ap_ready,
  C_drain_IO_L1_out_wrapper_107__ap_done,
  C_drain_IO_L1_out_wrapper_107__ap_idle,
  C_drain_IO_L1_out_wrapper_108__ap_start,
  C_drain_IO_L1_out_wrapper_108__ap_ready,
  C_drain_IO_L1_out_wrapper_108__ap_done,
  C_drain_IO_L1_out_wrapper_108__ap_idle,
  C_drain_IO_L1_out_wrapper_109__ap_start,
  C_drain_IO_L1_out_wrapper_109__ap_ready,
  C_drain_IO_L1_out_wrapper_109__ap_done,
  C_drain_IO_L1_out_wrapper_109__ap_idle,
  C_drain_IO_L1_out_wrapper_110__ap_start,
  C_drain_IO_L1_out_wrapper_110__ap_ready,
  C_drain_IO_L1_out_wrapper_110__ap_done,
  C_drain_IO_L1_out_wrapper_110__ap_idle,
  C_drain_IO_L1_out_wrapper_111__ap_start,
  C_drain_IO_L1_out_wrapper_111__ap_ready,
  C_drain_IO_L1_out_wrapper_111__ap_done,
  C_drain_IO_L1_out_wrapper_111__ap_idle,
  C_drain_IO_L1_out_wrapper_112__ap_start,
  C_drain_IO_L1_out_wrapper_112__ap_ready,
  C_drain_IO_L1_out_wrapper_112__ap_done,
  C_drain_IO_L1_out_wrapper_112__ap_idle,
  C_drain_IO_L1_out_wrapper_113__ap_start,
  C_drain_IO_L1_out_wrapper_113__ap_ready,
  C_drain_IO_L1_out_wrapper_113__ap_done,
  C_drain_IO_L1_out_wrapper_113__ap_idle,
  C_drain_IO_L1_out_wrapper_114__ap_start,
  C_drain_IO_L1_out_wrapper_114__ap_ready,
  C_drain_IO_L1_out_wrapper_114__ap_done,
  C_drain_IO_L1_out_wrapper_114__ap_idle,
  C_drain_IO_L1_out_wrapper_115__ap_start,
  C_drain_IO_L1_out_wrapper_115__ap_ready,
  C_drain_IO_L1_out_wrapper_115__ap_done,
  C_drain_IO_L1_out_wrapper_115__ap_idle,
  C_drain_IO_L1_out_wrapper_116__ap_start,
  C_drain_IO_L1_out_wrapper_116__ap_ready,
  C_drain_IO_L1_out_wrapper_116__ap_done,
  C_drain_IO_L1_out_wrapper_116__ap_idle,
  C_drain_IO_L1_out_wrapper_117__ap_start,
  C_drain_IO_L1_out_wrapper_117__ap_ready,
  C_drain_IO_L1_out_wrapper_117__ap_done,
  C_drain_IO_L1_out_wrapper_117__ap_idle,
  C_drain_IO_L1_out_wrapper_118__ap_start,
  C_drain_IO_L1_out_wrapper_118__ap_ready,
  C_drain_IO_L1_out_wrapper_118__ap_done,
  C_drain_IO_L1_out_wrapper_118__ap_idle,
  C_drain_IO_L1_out_wrapper_119__ap_start,
  C_drain_IO_L1_out_wrapper_119__ap_ready,
  C_drain_IO_L1_out_wrapper_119__ap_done,
  C_drain_IO_L1_out_wrapper_119__ap_idle,
  C_drain_IO_L1_out_wrapper_120__ap_start,
  C_drain_IO_L1_out_wrapper_120__ap_ready,
  C_drain_IO_L1_out_wrapper_120__ap_done,
  C_drain_IO_L1_out_wrapper_120__ap_idle,
  C_drain_IO_L1_out_wrapper_121__ap_start,
  C_drain_IO_L1_out_wrapper_121__ap_ready,
  C_drain_IO_L1_out_wrapper_121__ap_done,
  C_drain_IO_L1_out_wrapper_121__ap_idle,
  C_drain_IO_L1_out_wrapper_122__ap_start,
  C_drain_IO_L1_out_wrapper_122__ap_ready,
  C_drain_IO_L1_out_wrapper_122__ap_done,
  C_drain_IO_L1_out_wrapper_122__ap_idle,
  C_drain_IO_L1_out_wrapper_123__ap_start,
  C_drain_IO_L1_out_wrapper_123__ap_ready,
  C_drain_IO_L1_out_wrapper_123__ap_done,
  C_drain_IO_L1_out_wrapper_123__ap_idle,
  C_drain_IO_L1_out_wrapper_124__ap_start,
  C_drain_IO_L1_out_wrapper_124__ap_ready,
  C_drain_IO_L1_out_wrapper_124__ap_done,
  C_drain_IO_L1_out_wrapper_124__ap_idle,
  C_drain_IO_L1_out_wrapper_125__ap_start,
  C_drain_IO_L1_out_wrapper_125__ap_ready,
  C_drain_IO_L1_out_wrapper_125__ap_done,
  C_drain_IO_L1_out_wrapper_125__ap_idle,
  C_drain_IO_L1_out_wrapper_126__ap_start,
  C_drain_IO_L1_out_wrapper_126__ap_ready,
  C_drain_IO_L1_out_wrapper_126__ap_done,
  C_drain_IO_L1_out_wrapper_126__ap_idle,
  C_drain_IO_L1_out_wrapper_127__ap_start,
  C_drain_IO_L1_out_wrapper_127__ap_ready,
  C_drain_IO_L1_out_wrapper_127__ap_done,
  C_drain_IO_L1_out_wrapper_127__ap_idle,
  C_drain_IO_L1_out_wrapper_128__ap_start,
  C_drain_IO_L1_out_wrapper_128__ap_ready,
  C_drain_IO_L1_out_wrapper_128__ap_done,
  C_drain_IO_L1_out_wrapper_128__ap_idle,
  C_drain_IO_L1_out_wrapper_129__ap_start,
  C_drain_IO_L1_out_wrapper_129__ap_ready,
  C_drain_IO_L1_out_wrapper_129__ap_done,
  C_drain_IO_L1_out_wrapper_129__ap_idle,
  C_drain_IO_L1_out_wrapper_130__ap_start,
  C_drain_IO_L1_out_wrapper_130__ap_ready,
  C_drain_IO_L1_out_wrapper_130__ap_done,
  C_drain_IO_L1_out_wrapper_130__ap_idle,
  C_drain_IO_L1_out_wrapper_131__ap_start,
  C_drain_IO_L1_out_wrapper_131__ap_ready,
  C_drain_IO_L1_out_wrapper_131__ap_done,
  C_drain_IO_L1_out_wrapper_131__ap_idle,
  C_drain_IO_L1_out_wrapper_132__ap_start,
  C_drain_IO_L1_out_wrapper_132__ap_ready,
  C_drain_IO_L1_out_wrapper_132__ap_done,
  C_drain_IO_L1_out_wrapper_132__ap_idle,
  C_drain_IO_L1_out_wrapper_133__ap_start,
  C_drain_IO_L1_out_wrapper_133__ap_ready,
  C_drain_IO_L1_out_wrapper_133__ap_done,
  C_drain_IO_L1_out_wrapper_133__ap_idle,
  C_drain_IO_L1_out_wrapper_134__ap_start,
  C_drain_IO_L1_out_wrapper_134__ap_ready,
  C_drain_IO_L1_out_wrapper_134__ap_done,
  C_drain_IO_L1_out_wrapper_134__ap_idle,
  C_drain_IO_L1_out_wrapper_135__ap_start,
  C_drain_IO_L1_out_wrapper_135__ap_ready,
  C_drain_IO_L1_out_wrapper_135__ap_done,
  C_drain_IO_L1_out_wrapper_135__ap_idle,
  C_drain_IO_L1_out_wrapper_136__ap_start,
  C_drain_IO_L1_out_wrapper_136__ap_ready,
  C_drain_IO_L1_out_wrapper_136__ap_done,
  C_drain_IO_L1_out_wrapper_136__ap_idle,
  C_drain_IO_L1_out_wrapper_137__ap_start,
  C_drain_IO_L1_out_wrapper_137__ap_ready,
  C_drain_IO_L1_out_wrapper_137__ap_done,
  C_drain_IO_L1_out_wrapper_137__ap_idle,
  C_drain_IO_L1_out_wrapper_138__ap_start,
  C_drain_IO_L1_out_wrapper_138__ap_ready,
  C_drain_IO_L1_out_wrapper_138__ap_done,
  C_drain_IO_L1_out_wrapper_138__ap_idle,
  C_drain_IO_L1_out_wrapper_139__ap_start,
  C_drain_IO_L1_out_wrapper_139__ap_ready,
  C_drain_IO_L1_out_wrapper_139__ap_done,
  C_drain_IO_L1_out_wrapper_139__ap_idle,
  C_drain_IO_L1_out_wrapper_140__ap_start,
  C_drain_IO_L1_out_wrapper_140__ap_ready,
  C_drain_IO_L1_out_wrapper_140__ap_done,
  C_drain_IO_L1_out_wrapper_140__ap_idle,
  C_drain_IO_L1_out_wrapper_141__ap_start,
  C_drain_IO_L1_out_wrapper_141__ap_ready,
  C_drain_IO_L1_out_wrapper_141__ap_done,
  C_drain_IO_L1_out_wrapper_141__ap_idle,
  C_drain_IO_L1_out_wrapper_142__ap_start,
  C_drain_IO_L1_out_wrapper_142__ap_ready,
  C_drain_IO_L1_out_wrapper_142__ap_done,
  C_drain_IO_L1_out_wrapper_142__ap_idle,
  C_drain_IO_L1_out_wrapper_143__ap_start,
  C_drain_IO_L1_out_wrapper_143__ap_ready,
  C_drain_IO_L1_out_wrapper_143__ap_done,
  C_drain_IO_L1_out_wrapper_143__ap_idle,
  C_drain_IO_L1_out_wrapper_144__ap_start,
  C_drain_IO_L1_out_wrapper_144__ap_ready,
  C_drain_IO_L1_out_wrapper_144__ap_done,
  C_drain_IO_L1_out_wrapper_144__ap_idle,
  C_drain_IO_L1_out_wrapper_145__ap_start,
  C_drain_IO_L1_out_wrapper_145__ap_ready,
  C_drain_IO_L1_out_wrapper_145__ap_done,
  C_drain_IO_L1_out_wrapper_145__ap_idle,
  C_drain_IO_L1_out_wrapper_146__ap_start,
  C_drain_IO_L1_out_wrapper_146__ap_ready,
  C_drain_IO_L1_out_wrapper_146__ap_done,
  C_drain_IO_L1_out_wrapper_146__ap_idle,
  C_drain_IO_L1_out_wrapper_147__ap_start,
  C_drain_IO_L1_out_wrapper_147__ap_ready,
  C_drain_IO_L1_out_wrapper_147__ap_done,
  C_drain_IO_L1_out_wrapper_147__ap_idle,
  C_drain_IO_L1_out_wrapper_148__ap_start,
  C_drain_IO_L1_out_wrapper_148__ap_ready,
  C_drain_IO_L1_out_wrapper_148__ap_done,
  C_drain_IO_L1_out_wrapper_148__ap_idle,
  C_drain_IO_L1_out_wrapper_149__ap_start,
  C_drain_IO_L1_out_wrapper_149__ap_ready,
  C_drain_IO_L1_out_wrapper_149__ap_done,
  C_drain_IO_L1_out_wrapper_149__ap_idle,
  C_drain_IO_L1_out_wrapper_150__ap_start,
  C_drain_IO_L1_out_wrapper_150__ap_ready,
  C_drain_IO_L1_out_wrapper_150__ap_done,
  C_drain_IO_L1_out_wrapper_150__ap_idle,
  C_drain_IO_L1_out_wrapper_151__ap_start,
  C_drain_IO_L1_out_wrapper_151__ap_ready,
  C_drain_IO_L1_out_wrapper_151__ap_done,
  C_drain_IO_L1_out_wrapper_151__ap_idle,
  C_drain_IO_L1_out_wrapper_152__ap_start,
  C_drain_IO_L1_out_wrapper_152__ap_ready,
  C_drain_IO_L1_out_wrapper_152__ap_done,
  C_drain_IO_L1_out_wrapper_152__ap_idle,
  C_drain_IO_L1_out_wrapper_153__ap_start,
  C_drain_IO_L1_out_wrapper_153__ap_ready,
  C_drain_IO_L1_out_wrapper_153__ap_done,
  C_drain_IO_L1_out_wrapper_153__ap_idle,
  C_drain_IO_L1_out_wrapper_154__ap_start,
  C_drain_IO_L1_out_wrapper_154__ap_ready,
  C_drain_IO_L1_out_wrapper_154__ap_done,
  C_drain_IO_L1_out_wrapper_154__ap_idle,
  C_drain_IO_L1_out_wrapper_155__ap_start,
  C_drain_IO_L1_out_wrapper_155__ap_ready,
  C_drain_IO_L1_out_wrapper_155__ap_done,
  C_drain_IO_L1_out_wrapper_155__ap_idle,
  C_drain_IO_L1_out_wrapper_156__ap_start,
  C_drain_IO_L1_out_wrapper_156__ap_ready,
  C_drain_IO_L1_out_wrapper_156__ap_done,
  C_drain_IO_L1_out_wrapper_156__ap_idle,
  C_drain_IO_L1_out_wrapper_157__ap_start,
  C_drain_IO_L1_out_wrapper_157__ap_ready,
  C_drain_IO_L1_out_wrapper_157__ap_done,
  C_drain_IO_L1_out_wrapper_157__ap_idle,
  C_drain_IO_L1_out_wrapper_158__ap_start,
  C_drain_IO_L1_out_wrapper_158__ap_ready,
  C_drain_IO_L1_out_wrapper_158__ap_done,
  C_drain_IO_L1_out_wrapper_158__ap_idle,
  C_drain_IO_L1_out_wrapper_159__ap_start,
  C_drain_IO_L1_out_wrapper_159__ap_ready,
  C_drain_IO_L1_out_wrapper_159__ap_done,
  C_drain_IO_L1_out_wrapper_159__ap_idle,
  C_drain_IO_L1_out_wrapper_160__ap_start,
  C_drain_IO_L1_out_wrapper_160__ap_ready,
  C_drain_IO_L1_out_wrapper_160__ap_done,
  C_drain_IO_L1_out_wrapper_160__ap_idle,
  C_drain_IO_L1_out_wrapper_161__ap_start,
  C_drain_IO_L1_out_wrapper_161__ap_ready,
  C_drain_IO_L1_out_wrapper_161__ap_done,
  C_drain_IO_L1_out_wrapper_161__ap_idle,
  C_drain_IO_L1_out_wrapper_162__ap_start,
  C_drain_IO_L1_out_wrapper_162__ap_ready,
  C_drain_IO_L1_out_wrapper_162__ap_done,
  C_drain_IO_L1_out_wrapper_162__ap_idle,
  C_drain_IO_L1_out_wrapper_163__ap_start,
  C_drain_IO_L1_out_wrapper_163__ap_ready,
  C_drain_IO_L1_out_wrapper_163__ap_done,
  C_drain_IO_L1_out_wrapper_163__ap_idle,
  C_drain_IO_L1_out_wrapper_164__ap_start,
  C_drain_IO_L1_out_wrapper_164__ap_ready,
  C_drain_IO_L1_out_wrapper_164__ap_done,
  C_drain_IO_L1_out_wrapper_164__ap_idle,
  C_drain_IO_L1_out_wrapper_165__ap_start,
  C_drain_IO_L1_out_wrapper_165__ap_ready,
  C_drain_IO_L1_out_wrapper_165__ap_done,
  C_drain_IO_L1_out_wrapper_165__ap_idle,
  C_drain_IO_L1_out_wrapper_166__ap_start,
  C_drain_IO_L1_out_wrapper_166__ap_ready,
  C_drain_IO_L1_out_wrapper_166__ap_done,
  C_drain_IO_L1_out_wrapper_166__ap_idle,
  C_drain_IO_L1_out_wrapper_167__ap_start,
  C_drain_IO_L1_out_wrapper_167__ap_ready,
  C_drain_IO_L1_out_wrapper_167__ap_done,
  C_drain_IO_L1_out_wrapper_167__ap_idle,
  C_drain_IO_L1_out_wrapper_168__ap_start,
  C_drain_IO_L1_out_wrapper_168__ap_ready,
  C_drain_IO_L1_out_wrapper_168__ap_done,
  C_drain_IO_L1_out_wrapper_168__ap_idle,
  C_drain_IO_L1_out_wrapper_169__ap_start,
  C_drain_IO_L1_out_wrapper_169__ap_ready,
  C_drain_IO_L1_out_wrapper_169__ap_done,
  C_drain_IO_L1_out_wrapper_169__ap_idle,
  C_drain_IO_L1_out_wrapper_170__ap_start,
  C_drain_IO_L1_out_wrapper_170__ap_ready,
  C_drain_IO_L1_out_wrapper_170__ap_done,
  C_drain_IO_L1_out_wrapper_170__ap_idle,
  C_drain_IO_L1_out_wrapper_171__ap_start,
  C_drain_IO_L1_out_wrapper_171__ap_ready,
  C_drain_IO_L1_out_wrapper_171__ap_done,
  C_drain_IO_L1_out_wrapper_171__ap_idle,
  C_drain_IO_L1_out_wrapper_172__ap_start,
  C_drain_IO_L1_out_wrapper_172__ap_ready,
  C_drain_IO_L1_out_wrapper_172__ap_done,
  C_drain_IO_L1_out_wrapper_172__ap_idle,
  C_drain_IO_L1_out_wrapper_173__ap_start,
  C_drain_IO_L1_out_wrapper_173__ap_ready,
  C_drain_IO_L1_out_wrapper_173__ap_done,
  C_drain_IO_L1_out_wrapper_173__ap_idle,
  C_drain_IO_L1_out_wrapper_174__ap_start,
  C_drain_IO_L1_out_wrapper_174__ap_ready,
  C_drain_IO_L1_out_wrapper_174__ap_done,
  C_drain_IO_L1_out_wrapper_174__ap_idle,
  C_drain_IO_L1_out_wrapper_175__ap_start,
  C_drain_IO_L1_out_wrapper_175__ap_ready,
  C_drain_IO_L1_out_wrapper_175__ap_done,
  C_drain_IO_L1_out_wrapper_175__ap_idle,
  C_drain_IO_L1_out_wrapper_176__ap_start,
  C_drain_IO_L1_out_wrapper_176__ap_ready,
  C_drain_IO_L1_out_wrapper_176__ap_done,
  C_drain_IO_L1_out_wrapper_176__ap_idle,
  C_drain_IO_L1_out_wrapper_177__ap_start,
  C_drain_IO_L1_out_wrapper_177__ap_ready,
  C_drain_IO_L1_out_wrapper_177__ap_done,
  C_drain_IO_L1_out_wrapper_177__ap_idle,
  C_drain_IO_L1_out_wrapper_178__ap_start,
  C_drain_IO_L1_out_wrapper_178__ap_ready,
  C_drain_IO_L1_out_wrapper_178__ap_done,
  C_drain_IO_L1_out_wrapper_178__ap_idle,
  C_drain_IO_L1_out_wrapper_179__ap_start,
  C_drain_IO_L1_out_wrapper_179__ap_ready,
  C_drain_IO_L1_out_wrapper_179__ap_done,
  C_drain_IO_L1_out_wrapper_179__ap_idle,
  C_drain_IO_L1_out_wrapper_180__ap_start,
  C_drain_IO_L1_out_wrapper_180__ap_ready,
  C_drain_IO_L1_out_wrapper_180__ap_done,
  C_drain_IO_L1_out_wrapper_180__ap_idle,
  C_drain_IO_L1_out_wrapper_181__ap_start,
  C_drain_IO_L1_out_wrapper_181__ap_ready,
  C_drain_IO_L1_out_wrapper_181__ap_done,
  C_drain_IO_L1_out_wrapper_181__ap_idle,
  C_drain_IO_L1_out_wrapper_182__ap_start,
  C_drain_IO_L1_out_wrapper_182__ap_ready,
  C_drain_IO_L1_out_wrapper_182__ap_done,
  C_drain_IO_L1_out_wrapper_182__ap_idle,
  C_drain_IO_L1_out_wrapper_183__ap_start,
  C_drain_IO_L1_out_wrapper_183__ap_ready,
  C_drain_IO_L1_out_wrapper_183__ap_done,
  C_drain_IO_L1_out_wrapper_183__ap_idle,
  C_drain_IO_L1_out_wrapper_184__ap_start,
  C_drain_IO_L1_out_wrapper_184__ap_ready,
  C_drain_IO_L1_out_wrapper_184__ap_done,
  C_drain_IO_L1_out_wrapper_184__ap_idle,
  C_drain_IO_L1_out_wrapper_185__ap_start,
  C_drain_IO_L1_out_wrapper_185__ap_ready,
  C_drain_IO_L1_out_wrapper_185__ap_done,
  C_drain_IO_L1_out_wrapper_185__ap_idle,
  C_drain_IO_L1_out_wrapper_186__ap_start,
  C_drain_IO_L1_out_wrapper_186__ap_ready,
  C_drain_IO_L1_out_wrapper_186__ap_done,
  C_drain_IO_L1_out_wrapper_186__ap_idle,
  C_drain_IO_L1_out_wrapper_187__ap_start,
  C_drain_IO_L1_out_wrapper_187__ap_ready,
  C_drain_IO_L1_out_wrapper_187__ap_done,
  C_drain_IO_L1_out_wrapper_187__ap_idle,
  C_drain_IO_L1_out_wrapper_188__ap_start,
  C_drain_IO_L1_out_wrapper_188__ap_ready,
  C_drain_IO_L1_out_wrapper_188__ap_done,
  C_drain_IO_L1_out_wrapper_188__ap_idle,
  C_drain_IO_L1_out_wrapper_189__ap_start,
  C_drain_IO_L1_out_wrapper_189__ap_ready,
  C_drain_IO_L1_out_wrapper_189__ap_done,
  C_drain_IO_L1_out_wrapper_189__ap_idle,
  C_drain_IO_L1_out_wrapper_190__ap_start,
  C_drain_IO_L1_out_wrapper_190__ap_ready,
  C_drain_IO_L1_out_wrapper_190__ap_done,
  C_drain_IO_L1_out_wrapper_190__ap_idle,
  C_drain_IO_L1_out_wrapper_191__ap_start,
  C_drain_IO_L1_out_wrapper_191__ap_ready,
  C_drain_IO_L1_out_wrapper_191__ap_done,
  C_drain_IO_L1_out_wrapper_191__ap_idle,
  C_drain_IO_L1_out_wrapper_192__ap_start,
  C_drain_IO_L1_out_wrapper_192__ap_ready,
  C_drain_IO_L1_out_wrapper_192__ap_done,
  C_drain_IO_L1_out_wrapper_192__ap_idle,
  C_drain_IO_L1_out_wrapper_193__ap_start,
  C_drain_IO_L1_out_wrapper_193__ap_ready,
  C_drain_IO_L1_out_wrapper_193__ap_done,
  C_drain_IO_L1_out_wrapper_193__ap_idle,
  C_drain_IO_L1_out_wrapper_194__ap_start,
  C_drain_IO_L1_out_wrapper_194__ap_ready,
  C_drain_IO_L1_out_wrapper_194__ap_done,
  C_drain_IO_L1_out_wrapper_194__ap_idle,
  C_drain_IO_L1_out_wrapper_195__ap_start,
  C_drain_IO_L1_out_wrapper_195__ap_ready,
  C_drain_IO_L1_out_wrapper_195__ap_done,
  C_drain_IO_L1_out_wrapper_195__ap_idle,
  C_drain_IO_L1_out_wrapper_196__ap_start,
  C_drain_IO_L1_out_wrapper_196__ap_ready,
  C_drain_IO_L1_out_wrapper_196__ap_done,
  C_drain_IO_L1_out_wrapper_196__ap_idle,
  C_drain_IO_L1_out_wrapper_197__ap_start,
  C_drain_IO_L1_out_wrapper_197__ap_ready,
  C_drain_IO_L1_out_wrapper_197__ap_done,
  C_drain_IO_L1_out_wrapper_197__ap_idle,
  C_drain_IO_L1_out_wrapper_198__ap_start,
  C_drain_IO_L1_out_wrapper_198__ap_ready,
  C_drain_IO_L1_out_wrapper_198__ap_done,
  C_drain_IO_L1_out_wrapper_198__ap_idle,
  C_drain_IO_L1_out_wrapper_199__ap_start,
  C_drain_IO_L1_out_wrapper_199__ap_ready,
  C_drain_IO_L1_out_wrapper_199__ap_done,
  C_drain_IO_L1_out_wrapper_199__ap_idle,
  C_drain_IO_L1_out_wrapper_200__ap_start,
  C_drain_IO_L1_out_wrapper_200__ap_ready,
  C_drain_IO_L1_out_wrapper_200__ap_done,
  C_drain_IO_L1_out_wrapper_200__ap_idle,
  C_drain_IO_L1_out_wrapper_201__ap_start,
  C_drain_IO_L1_out_wrapper_201__ap_ready,
  C_drain_IO_L1_out_wrapper_201__ap_done,
  C_drain_IO_L1_out_wrapper_201__ap_idle,
  C_drain_IO_L1_out_wrapper_202__ap_start,
  C_drain_IO_L1_out_wrapper_202__ap_ready,
  C_drain_IO_L1_out_wrapper_202__ap_done,
  C_drain_IO_L1_out_wrapper_202__ap_idle,
  C_drain_IO_L1_out_wrapper_203__ap_start,
  C_drain_IO_L1_out_wrapper_203__ap_ready,
  C_drain_IO_L1_out_wrapper_203__ap_done,
  C_drain_IO_L1_out_wrapper_203__ap_idle,
  C_drain_IO_L1_out_wrapper_204__ap_start,
  C_drain_IO_L1_out_wrapper_204__ap_ready,
  C_drain_IO_L1_out_wrapper_204__ap_done,
  C_drain_IO_L1_out_wrapper_204__ap_idle,
  C_drain_IO_L1_out_wrapper_205__ap_start,
  C_drain_IO_L1_out_wrapper_205__ap_ready,
  C_drain_IO_L1_out_wrapper_205__ap_done,
  C_drain_IO_L1_out_wrapper_205__ap_idle,
  C_drain_IO_L1_out_wrapper_206__ap_start,
  C_drain_IO_L1_out_wrapper_206__ap_ready,
  C_drain_IO_L1_out_wrapper_206__ap_done,
  C_drain_IO_L1_out_wrapper_206__ap_idle,
  C_drain_IO_L1_out_wrapper_207__ap_start,
  C_drain_IO_L1_out_wrapper_207__ap_ready,
  C_drain_IO_L1_out_wrapper_207__ap_done,
  C_drain_IO_L1_out_wrapper_207__ap_idle,
  C_drain_IO_L1_out_wrapper_208__ap_start,
  C_drain_IO_L1_out_wrapper_208__ap_ready,
  C_drain_IO_L1_out_wrapper_208__ap_done,
  C_drain_IO_L1_out_wrapper_208__ap_idle,
  C_drain_IO_L1_out_wrapper_209__ap_start,
  C_drain_IO_L1_out_wrapper_209__ap_ready,
  C_drain_IO_L1_out_wrapper_209__ap_done,
  C_drain_IO_L1_out_wrapper_209__ap_idle,
  C_drain_IO_L1_out_wrapper_210__ap_start,
  C_drain_IO_L1_out_wrapper_210__ap_ready,
  C_drain_IO_L1_out_wrapper_210__ap_done,
  C_drain_IO_L1_out_wrapper_210__ap_idle,
  C_drain_IO_L1_out_wrapper_211__ap_start,
  C_drain_IO_L1_out_wrapper_211__ap_ready,
  C_drain_IO_L1_out_wrapper_211__ap_done,
  C_drain_IO_L1_out_wrapper_211__ap_idle,
  C_drain_IO_L1_out_wrapper_212__ap_start,
  C_drain_IO_L1_out_wrapper_212__ap_ready,
  C_drain_IO_L1_out_wrapper_212__ap_done,
  C_drain_IO_L1_out_wrapper_212__ap_idle,
  C_drain_IO_L1_out_wrapper_213__ap_start,
  C_drain_IO_L1_out_wrapper_213__ap_ready,
  C_drain_IO_L1_out_wrapper_213__ap_done,
  C_drain_IO_L1_out_wrapper_213__ap_idle,
  C_drain_IO_L1_out_wrapper_214__ap_start,
  C_drain_IO_L1_out_wrapper_214__ap_ready,
  C_drain_IO_L1_out_wrapper_214__ap_done,
  C_drain_IO_L1_out_wrapper_214__ap_idle,
  C_drain_IO_L1_out_wrapper_215__ap_start,
  C_drain_IO_L1_out_wrapper_215__ap_ready,
  C_drain_IO_L1_out_wrapper_215__ap_done,
  C_drain_IO_L1_out_wrapper_215__ap_idle,
  C_drain_IO_L1_out_wrapper_216__ap_start,
  C_drain_IO_L1_out_wrapper_216__ap_ready,
  C_drain_IO_L1_out_wrapper_216__ap_done,
  C_drain_IO_L1_out_wrapper_216__ap_idle,
  C_drain_IO_L1_out_wrapper_217__ap_start,
  C_drain_IO_L1_out_wrapper_217__ap_ready,
  C_drain_IO_L1_out_wrapper_217__ap_done,
  C_drain_IO_L1_out_wrapper_217__ap_idle,
  C_drain_IO_L1_out_wrapper_218__ap_start,
  C_drain_IO_L1_out_wrapper_218__ap_ready,
  C_drain_IO_L1_out_wrapper_218__ap_done,
  C_drain_IO_L1_out_wrapper_218__ap_idle,
  C_drain_IO_L1_out_wrapper_219__ap_start,
  C_drain_IO_L1_out_wrapper_219__ap_ready,
  C_drain_IO_L1_out_wrapper_219__ap_done,
  C_drain_IO_L1_out_wrapper_219__ap_idle,
  C_drain_IO_L1_out_wrapper_220__ap_start,
  C_drain_IO_L1_out_wrapper_220__ap_ready,
  C_drain_IO_L1_out_wrapper_220__ap_done,
  C_drain_IO_L1_out_wrapper_220__ap_idle,
  C_drain_IO_L1_out_wrapper_221__ap_start,
  C_drain_IO_L1_out_wrapper_221__ap_ready,
  C_drain_IO_L1_out_wrapper_221__ap_done,
  C_drain_IO_L1_out_wrapper_221__ap_idle,
  C_drain_IO_L1_out_wrapper_222__ap_start,
  C_drain_IO_L1_out_wrapper_222__ap_ready,
  C_drain_IO_L1_out_wrapper_222__ap_done,
  C_drain_IO_L1_out_wrapper_222__ap_idle,
  C_drain_IO_L1_out_wrapper_223__ap_start,
  C_drain_IO_L1_out_wrapper_223__ap_ready,
  C_drain_IO_L1_out_wrapper_223__ap_done,
  C_drain_IO_L1_out_wrapper_223__ap_idle,
  C_drain_IO_L1_out_wrapper_224__ap_start,
  C_drain_IO_L1_out_wrapper_224__ap_ready,
  C_drain_IO_L1_out_wrapper_224__ap_done,
  C_drain_IO_L1_out_wrapper_224__ap_idle,
  C_drain_IO_L1_out_wrapper_225__ap_start,
  C_drain_IO_L1_out_wrapper_225__ap_ready,
  C_drain_IO_L1_out_wrapper_225__ap_done,
  C_drain_IO_L1_out_wrapper_225__ap_idle,
  C_drain_IO_L1_out_wrapper_226__ap_start,
  C_drain_IO_L1_out_wrapper_226__ap_ready,
  C_drain_IO_L1_out_wrapper_226__ap_done,
  C_drain_IO_L1_out_wrapper_226__ap_idle,
  C_drain_IO_L1_out_wrapper_227__ap_start,
  C_drain_IO_L1_out_wrapper_227__ap_ready,
  C_drain_IO_L1_out_wrapper_227__ap_done,
  C_drain_IO_L1_out_wrapper_227__ap_idle,
  C_drain_IO_L1_out_wrapper_228__ap_start,
  C_drain_IO_L1_out_wrapper_228__ap_ready,
  C_drain_IO_L1_out_wrapper_228__ap_done,
  C_drain_IO_L1_out_wrapper_228__ap_idle,
  C_drain_IO_L1_out_wrapper_229__ap_start,
  C_drain_IO_L1_out_wrapper_229__ap_ready,
  C_drain_IO_L1_out_wrapper_229__ap_done,
  C_drain_IO_L1_out_wrapper_229__ap_idle,
  C_drain_IO_L1_out_wrapper_230__ap_start,
  C_drain_IO_L1_out_wrapper_230__ap_ready,
  C_drain_IO_L1_out_wrapper_230__ap_done,
  C_drain_IO_L1_out_wrapper_230__ap_idle,
  C_drain_IO_L1_out_wrapper_231__ap_start,
  C_drain_IO_L1_out_wrapper_231__ap_ready,
  C_drain_IO_L1_out_wrapper_231__ap_done,
  C_drain_IO_L1_out_wrapper_231__ap_idle,
  C_drain_IO_L1_out_wrapper_232__ap_start,
  C_drain_IO_L1_out_wrapper_232__ap_ready,
  C_drain_IO_L1_out_wrapper_232__ap_done,
  C_drain_IO_L1_out_wrapper_232__ap_idle,
  C_drain_IO_L1_out_wrapper_233__ap_start,
  C_drain_IO_L1_out_wrapper_233__ap_ready,
  C_drain_IO_L1_out_wrapper_233__ap_done,
  C_drain_IO_L1_out_wrapper_233__ap_idle,
  C_drain_IO_L1_out_wrapper_234__ap_start,
  C_drain_IO_L1_out_wrapper_234__ap_ready,
  C_drain_IO_L1_out_wrapper_234__ap_done,
  C_drain_IO_L1_out_wrapper_234__ap_idle,
  C_drain_IO_L1_out_wrapper_235__ap_start,
  C_drain_IO_L1_out_wrapper_235__ap_ready,
  C_drain_IO_L1_out_wrapper_235__ap_done,
  C_drain_IO_L1_out_wrapper_235__ap_idle,
  C_drain_IO_L1_out_wrapper_236__ap_start,
  C_drain_IO_L1_out_wrapper_236__ap_ready,
  C_drain_IO_L1_out_wrapper_236__ap_done,
  C_drain_IO_L1_out_wrapper_236__ap_idle,
  C_drain_IO_L1_out_wrapper_237__ap_start,
  C_drain_IO_L1_out_wrapper_237__ap_ready,
  C_drain_IO_L1_out_wrapper_237__ap_done,
  C_drain_IO_L1_out_wrapper_237__ap_idle,
  C_drain_IO_L1_out_wrapper_238__ap_start,
  C_drain_IO_L1_out_wrapper_238__ap_ready,
  C_drain_IO_L1_out_wrapper_238__ap_done,
  C_drain_IO_L1_out_wrapper_238__ap_idle,
  C_drain_IO_L1_out_wrapper_239__ap_start,
  C_drain_IO_L1_out_wrapper_239__ap_ready,
  C_drain_IO_L1_out_wrapper_239__ap_done,
  C_drain_IO_L1_out_wrapper_239__ap_idle,
  C_drain_IO_L1_out_wrapper_240__ap_start,
  C_drain_IO_L1_out_wrapper_240__ap_ready,
  C_drain_IO_L1_out_wrapper_240__ap_done,
  C_drain_IO_L1_out_wrapper_240__ap_idle,
  C_drain_IO_L1_out_wrapper_241__ap_start,
  C_drain_IO_L1_out_wrapper_241__ap_ready,
  C_drain_IO_L1_out_wrapper_241__ap_done,
  C_drain_IO_L1_out_wrapper_241__ap_idle,
  C_drain_IO_L1_out_wrapper_242__ap_start,
  C_drain_IO_L1_out_wrapper_242__ap_ready,
  C_drain_IO_L1_out_wrapper_242__ap_done,
  C_drain_IO_L1_out_wrapper_242__ap_idle,
  C_drain_IO_L1_out_wrapper_243__ap_start,
  C_drain_IO_L1_out_wrapper_243__ap_ready,
  C_drain_IO_L1_out_wrapper_243__ap_done,
  C_drain_IO_L1_out_wrapper_243__ap_idle,
  C_drain_IO_L1_out_wrapper_244__ap_start,
  C_drain_IO_L1_out_wrapper_244__ap_ready,
  C_drain_IO_L1_out_wrapper_244__ap_done,
  C_drain_IO_L1_out_wrapper_244__ap_idle,
  C_drain_IO_L1_out_wrapper_245__ap_start,
  C_drain_IO_L1_out_wrapper_245__ap_ready,
  C_drain_IO_L1_out_wrapper_245__ap_done,
  C_drain_IO_L1_out_wrapper_245__ap_idle,
  C_drain_IO_L1_out_wrapper_246__ap_start,
  C_drain_IO_L1_out_wrapper_246__ap_ready,
  C_drain_IO_L1_out_wrapper_246__ap_done,
  C_drain_IO_L1_out_wrapper_246__ap_idle,
  C_drain_IO_L1_out_wrapper_247__ap_start,
  C_drain_IO_L1_out_wrapper_247__ap_ready,
  C_drain_IO_L1_out_wrapper_247__ap_done,
  C_drain_IO_L1_out_wrapper_247__ap_idle,
  C_drain_IO_L1_out_wrapper_248__ap_start,
  C_drain_IO_L1_out_wrapper_248__ap_ready,
  C_drain_IO_L1_out_wrapper_248__ap_done,
  C_drain_IO_L1_out_wrapper_248__ap_idle,
  C_drain_IO_L1_out_wrapper_249__ap_start,
  C_drain_IO_L1_out_wrapper_249__ap_ready,
  C_drain_IO_L1_out_wrapper_249__ap_done,
  C_drain_IO_L1_out_wrapper_249__ap_idle,
  C_drain_IO_L1_out_wrapper_250__ap_start,
  C_drain_IO_L1_out_wrapper_250__ap_ready,
  C_drain_IO_L1_out_wrapper_250__ap_done,
  C_drain_IO_L1_out_wrapper_250__ap_idle,
  C_drain_IO_L1_out_wrapper_251__ap_start,
  C_drain_IO_L1_out_wrapper_251__ap_ready,
  C_drain_IO_L1_out_wrapper_251__ap_done,
  C_drain_IO_L1_out_wrapper_251__ap_idle,
  C_drain_IO_L1_out_wrapper_252__ap_start,
  C_drain_IO_L1_out_wrapper_252__ap_ready,
  C_drain_IO_L1_out_wrapper_252__ap_done,
  C_drain_IO_L1_out_wrapper_252__ap_idle,
  C_drain_IO_L1_out_wrapper_253__ap_start,
  C_drain_IO_L1_out_wrapper_253__ap_ready,
  C_drain_IO_L1_out_wrapper_253__ap_done,
  C_drain_IO_L1_out_wrapper_253__ap_idle,
  C_drain_IO_L1_out_wrapper_254__ap_start,
  C_drain_IO_L1_out_wrapper_254__ap_ready,
  C_drain_IO_L1_out_wrapper_254__ap_done,
  C_drain_IO_L1_out_wrapper_254__ap_idle,
  C_drain_IO_L1_out_wrapper_255__ap_start,
  C_drain_IO_L1_out_wrapper_255__ap_ready,
  C_drain_IO_L1_out_wrapper_255__ap_done,
  C_drain_IO_L1_out_wrapper_255__ap_idle,
  C_drain_IO_L1_out_wrapper_256__ap_start,
  C_drain_IO_L1_out_wrapper_256__ap_ready,
  C_drain_IO_L1_out_wrapper_256__ap_done,
  C_drain_IO_L1_out_wrapper_256__ap_idle,
  C_drain_IO_L1_out_wrapper_257__ap_start,
  C_drain_IO_L1_out_wrapper_257__ap_ready,
  C_drain_IO_L1_out_wrapper_257__ap_done,
  C_drain_IO_L1_out_wrapper_257__ap_idle,
  C_drain_IO_L1_out_wrapper_258__ap_start,
  C_drain_IO_L1_out_wrapper_258__ap_ready,
  C_drain_IO_L1_out_wrapper_258__ap_done,
  C_drain_IO_L1_out_wrapper_258__ap_idle,
  C_drain_IO_L1_out_wrapper_259__ap_start,
  C_drain_IO_L1_out_wrapper_259__ap_ready,
  C_drain_IO_L1_out_wrapper_259__ap_done,
  C_drain_IO_L1_out_wrapper_259__ap_idle,
  C_drain_IO_L1_out_wrapper_260__ap_start,
  C_drain_IO_L1_out_wrapper_260__ap_ready,
  C_drain_IO_L1_out_wrapper_260__ap_done,
  C_drain_IO_L1_out_wrapper_260__ap_idle,
  C_drain_IO_L1_out_wrapper_261__ap_start,
  C_drain_IO_L1_out_wrapper_261__ap_ready,
  C_drain_IO_L1_out_wrapper_261__ap_done,
  C_drain_IO_L1_out_wrapper_261__ap_idle,
  C_drain_IO_L1_out_wrapper_262__ap_start,
  C_drain_IO_L1_out_wrapper_262__ap_ready,
  C_drain_IO_L1_out_wrapper_262__ap_done,
  C_drain_IO_L1_out_wrapper_262__ap_idle,
  C_drain_IO_L1_out_wrapper_263__ap_start,
  C_drain_IO_L1_out_wrapper_263__ap_ready,
  C_drain_IO_L1_out_wrapper_263__ap_done,
  C_drain_IO_L1_out_wrapper_263__ap_idle,
  C_drain_IO_L1_out_wrapper_264__ap_start,
  C_drain_IO_L1_out_wrapper_264__ap_ready,
  C_drain_IO_L1_out_wrapper_264__ap_done,
  C_drain_IO_L1_out_wrapper_264__ap_idle,
  C_drain_IO_L1_out_wrapper_265__ap_start,
  C_drain_IO_L1_out_wrapper_265__ap_ready,
  C_drain_IO_L1_out_wrapper_265__ap_done,
  C_drain_IO_L1_out_wrapper_265__ap_idle,
  C_drain_IO_L1_out_wrapper_266__ap_start,
  C_drain_IO_L1_out_wrapper_266__ap_ready,
  C_drain_IO_L1_out_wrapper_266__ap_done,
  C_drain_IO_L1_out_wrapper_266__ap_idle,
  C_drain_IO_L1_out_wrapper_267__ap_start,
  C_drain_IO_L1_out_wrapper_267__ap_ready,
  C_drain_IO_L1_out_wrapper_267__ap_done,
  C_drain_IO_L1_out_wrapper_267__ap_idle,
  C_drain_IO_L1_out_wrapper_268__ap_start,
  C_drain_IO_L1_out_wrapper_268__ap_ready,
  C_drain_IO_L1_out_wrapper_268__ap_done,
  C_drain_IO_L1_out_wrapper_268__ap_idle,
  C_drain_IO_L1_out_wrapper_269__ap_start,
  C_drain_IO_L1_out_wrapper_269__ap_ready,
  C_drain_IO_L1_out_wrapper_269__ap_done,
  C_drain_IO_L1_out_wrapper_269__ap_idle,
  C_drain_IO_L1_out_wrapper_270__ap_start,
  C_drain_IO_L1_out_wrapper_270__ap_ready,
  C_drain_IO_L1_out_wrapper_270__ap_done,
  C_drain_IO_L1_out_wrapper_270__ap_idle,
  C_drain_IO_L1_out_wrapper_271__ap_start,
  C_drain_IO_L1_out_wrapper_271__ap_ready,
  C_drain_IO_L1_out_wrapper_271__ap_done,
  C_drain_IO_L1_out_wrapper_271__ap_idle,
  C_drain_IO_L1_out_wrapper_272__ap_start,
  C_drain_IO_L1_out_wrapper_272__ap_ready,
  C_drain_IO_L1_out_wrapper_272__ap_done,
  C_drain_IO_L1_out_wrapper_272__ap_idle,
  C_drain_IO_L1_out_wrapper_273__ap_start,
  C_drain_IO_L1_out_wrapper_273__ap_ready,
  C_drain_IO_L1_out_wrapper_273__ap_done,
  C_drain_IO_L1_out_wrapper_273__ap_idle,
  C_drain_IO_L1_out_wrapper_274__ap_start,
  C_drain_IO_L1_out_wrapper_274__ap_ready,
  C_drain_IO_L1_out_wrapper_274__ap_done,
  C_drain_IO_L1_out_wrapper_274__ap_idle,
  C_drain_IO_L1_out_wrapper_275__ap_start,
  C_drain_IO_L1_out_wrapper_275__ap_ready,
  C_drain_IO_L1_out_wrapper_275__ap_done,
  C_drain_IO_L1_out_wrapper_275__ap_idle,
  C_drain_IO_L1_out_wrapper_276__ap_start,
  C_drain_IO_L1_out_wrapper_276__ap_ready,
  C_drain_IO_L1_out_wrapper_276__ap_done,
  C_drain_IO_L1_out_wrapper_276__ap_idle,
  C_drain_IO_L1_out_wrapper_277__ap_start,
  C_drain_IO_L1_out_wrapper_277__ap_ready,
  C_drain_IO_L1_out_wrapper_277__ap_done,
  C_drain_IO_L1_out_wrapper_277__ap_idle,
  C_drain_IO_L1_out_wrapper_278__ap_start,
  C_drain_IO_L1_out_wrapper_278__ap_ready,
  C_drain_IO_L1_out_wrapper_278__ap_done,
  C_drain_IO_L1_out_wrapper_278__ap_idle,
  C_drain_IO_L1_out_wrapper_279__ap_start,
  C_drain_IO_L1_out_wrapper_279__ap_ready,
  C_drain_IO_L1_out_wrapper_279__ap_done,
  C_drain_IO_L1_out_wrapper_279__ap_idle,
  C_drain_IO_L1_out_wrapper_280__ap_start,
  C_drain_IO_L1_out_wrapper_280__ap_ready,
  C_drain_IO_L1_out_wrapper_280__ap_done,
  C_drain_IO_L1_out_wrapper_280__ap_idle,
  C_drain_IO_L1_out_wrapper_281__ap_start,
  C_drain_IO_L1_out_wrapper_281__ap_ready,
  C_drain_IO_L1_out_wrapper_281__ap_done,
  C_drain_IO_L1_out_wrapper_281__ap_idle,
  C_drain_IO_L1_out_wrapper_282__ap_start,
  C_drain_IO_L1_out_wrapper_282__ap_ready,
  C_drain_IO_L1_out_wrapper_282__ap_done,
  C_drain_IO_L1_out_wrapper_282__ap_idle,
  C_drain_IO_L1_out_wrapper_283__ap_start,
  C_drain_IO_L1_out_wrapper_283__ap_ready,
  C_drain_IO_L1_out_wrapper_283__ap_done,
  C_drain_IO_L1_out_wrapper_283__ap_idle,
  C_drain_IO_L1_out_wrapper_284__ap_start,
  C_drain_IO_L1_out_wrapper_284__ap_ready,
  C_drain_IO_L1_out_wrapper_284__ap_done,
  C_drain_IO_L1_out_wrapper_284__ap_idle,
  C_drain_IO_L1_out_wrapper_285__ap_start,
  C_drain_IO_L1_out_wrapper_285__ap_ready,
  C_drain_IO_L1_out_wrapper_285__ap_done,
  C_drain_IO_L1_out_wrapper_285__ap_idle,
  C_drain_IO_L1_out_wrapper_286__ap_start,
  C_drain_IO_L1_out_wrapper_286__ap_ready,
  C_drain_IO_L1_out_wrapper_286__ap_done,
  C_drain_IO_L1_out_wrapper_286__ap_idle,
  C_drain_IO_L1_out_wrapper_287__ap_start,
  C_drain_IO_L1_out_wrapper_287__ap_ready,
  C_drain_IO_L1_out_wrapper_287__ap_done,
  C_drain_IO_L1_out_wrapper_287__ap_idle,
  C_drain_IO_L1_out_wrapper_288__ap_start,
  C_drain_IO_L1_out_wrapper_288__ap_ready,
  C_drain_IO_L1_out_wrapper_288__ap_done,
  C_drain_IO_L1_out_wrapper_288__ap_idle,
  C_drain_IO_L2_out_0__ap_start,
  C_drain_IO_L2_out_0__ap_ready,
  C_drain_IO_L2_out_0__ap_done,
  C_drain_IO_L2_out_0__ap_idle,
  C_drain_IO_L2_out_1__ap_start,
  C_drain_IO_L2_out_1__ap_ready,
  C_drain_IO_L2_out_1__ap_done,
  C_drain_IO_L2_out_1__ap_idle,
  C_drain_IO_L2_out_2__ap_start,
  C_drain_IO_L2_out_2__ap_ready,
  C_drain_IO_L2_out_2__ap_done,
  C_drain_IO_L2_out_2__ap_idle,
  C_drain_IO_L2_out_3__ap_start,
  C_drain_IO_L2_out_3__ap_ready,
  C_drain_IO_L2_out_3__ap_done,
  C_drain_IO_L2_out_3__ap_idle,
  C_drain_IO_L2_out_4__ap_start,
  C_drain_IO_L2_out_4__ap_ready,
  C_drain_IO_L2_out_4__ap_done,
  C_drain_IO_L2_out_4__ap_idle,
  C_drain_IO_L2_out_5__ap_start,
  C_drain_IO_L2_out_5__ap_ready,
  C_drain_IO_L2_out_5__ap_done,
  C_drain_IO_L2_out_5__ap_idle,
  C_drain_IO_L2_out_6__ap_start,
  C_drain_IO_L2_out_6__ap_ready,
  C_drain_IO_L2_out_6__ap_done,
  C_drain_IO_L2_out_6__ap_idle,
  C_drain_IO_L2_out_7__ap_start,
  C_drain_IO_L2_out_7__ap_ready,
  C_drain_IO_L2_out_7__ap_done,
  C_drain_IO_L2_out_7__ap_idle,
  C_drain_IO_L2_out_8__ap_start,
  C_drain_IO_L2_out_8__ap_ready,
  C_drain_IO_L2_out_8__ap_done,
  C_drain_IO_L2_out_8__ap_idle,
  C_drain_IO_L2_out_9__ap_start,
  C_drain_IO_L2_out_9__ap_ready,
  C_drain_IO_L2_out_9__ap_done,
  C_drain_IO_L2_out_9__ap_idle,
  C_drain_IO_L2_out_10__ap_start,
  C_drain_IO_L2_out_10__ap_ready,
  C_drain_IO_L2_out_10__ap_done,
  C_drain_IO_L2_out_10__ap_idle,
  C_drain_IO_L2_out_11__ap_start,
  C_drain_IO_L2_out_11__ap_ready,
  C_drain_IO_L2_out_11__ap_done,
  C_drain_IO_L2_out_11__ap_idle,
  C_drain_IO_L2_out_12__ap_start,
  C_drain_IO_L2_out_12__ap_ready,
  C_drain_IO_L2_out_12__ap_done,
  C_drain_IO_L2_out_12__ap_idle,
  C_drain_IO_L2_out_13__ap_start,
  C_drain_IO_L2_out_13__ap_ready,
  C_drain_IO_L2_out_13__ap_done,
  C_drain_IO_L2_out_13__ap_idle,
  C_drain_IO_L2_out_14__ap_start,
  C_drain_IO_L2_out_14__ap_ready,
  C_drain_IO_L2_out_14__ap_done,
  C_drain_IO_L2_out_14__ap_idle,
  C_drain_IO_L2_out_15__ap_start,
  C_drain_IO_L2_out_15__ap_ready,
  C_drain_IO_L2_out_15__ap_done,
  C_drain_IO_L2_out_15__ap_idle,
  C_drain_IO_L2_out_boundary_0__ap_start,
  C_drain_IO_L2_out_boundary_0__ap_ready,
  C_drain_IO_L2_out_boundary_0__ap_done,
  C_drain_IO_L2_out_boundary_0__ap_idle,
  C_drain_IO_L3_out_0__ap_start,
  C_drain_IO_L3_out_0__ap_ready,
  C_drain_IO_L3_out_0__ap_done,
  C_drain_IO_L3_out_0__ap_idle,
  C_drain_IO_L3_out_serialize_0___C__q0,
  C_drain_IO_L3_out_serialize_0__ap_start,
  C_drain_IO_L3_out_serialize_0__ap_ready,
  C_drain_IO_L3_out_serialize_0__ap_done,
  C_drain_IO_L3_out_serialize_0__ap_idle,
  PE_wrapper_0__ap_start,
  PE_wrapper_0__ap_ready,
  PE_wrapper_0__ap_done,
  PE_wrapper_0__ap_idle,
  PE_wrapper_1__ap_start,
  PE_wrapper_1__ap_ready,
  PE_wrapper_1__ap_done,
  PE_wrapper_1__ap_idle,
  PE_wrapper_2__ap_start,
  PE_wrapper_2__ap_ready,
  PE_wrapper_2__ap_done,
  PE_wrapper_2__ap_idle,
  PE_wrapper_3__ap_start,
  PE_wrapper_3__ap_ready,
  PE_wrapper_3__ap_done,
  PE_wrapper_3__ap_idle,
  PE_wrapper_4__ap_start,
  PE_wrapper_4__ap_ready,
  PE_wrapper_4__ap_done,
  PE_wrapper_4__ap_idle,
  PE_wrapper_5__ap_start,
  PE_wrapper_5__ap_ready,
  PE_wrapper_5__ap_done,
  PE_wrapper_5__ap_idle,
  PE_wrapper_6__ap_start,
  PE_wrapper_6__ap_ready,
  PE_wrapper_6__ap_done,
  PE_wrapper_6__ap_idle,
  PE_wrapper_7__ap_start,
  PE_wrapper_7__ap_ready,
  PE_wrapper_7__ap_done,
  PE_wrapper_7__ap_idle,
  PE_wrapper_8__ap_start,
  PE_wrapper_8__ap_ready,
  PE_wrapper_8__ap_done,
  PE_wrapper_8__ap_idle,
  PE_wrapper_9__ap_start,
  PE_wrapper_9__ap_ready,
  PE_wrapper_9__ap_done,
  PE_wrapper_9__ap_idle,
  PE_wrapper_10__ap_start,
  PE_wrapper_10__ap_ready,
  PE_wrapper_10__ap_done,
  PE_wrapper_10__ap_idle,
  PE_wrapper_11__ap_start,
  PE_wrapper_11__ap_ready,
  PE_wrapper_11__ap_done,
  PE_wrapper_11__ap_idle,
  PE_wrapper_12__ap_start,
  PE_wrapper_12__ap_ready,
  PE_wrapper_12__ap_done,
  PE_wrapper_12__ap_idle,
  PE_wrapper_13__ap_start,
  PE_wrapper_13__ap_ready,
  PE_wrapper_13__ap_done,
  PE_wrapper_13__ap_idle,
  PE_wrapper_14__ap_start,
  PE_wrapper_14__ap_ready,
  PE_wrapper_14__ap_done,
  PE_wrapper_14__ap_idle,
  PE_wrapper_15__ap_start,
  PE_wrapper_15__ap_ready,
  PE_wrapper_15__ap_done,
  PE_wrapper_15__ap_idle,
  PE_wrapper_16__ap_start,
  PE_wrapper_16__ap_ready,
  PE_wrapper_16__ap_done,
  PE_wrapper_16__ap_idle,
  PE_wrapper_17__ap_start,
  PE_wrapper_17__ap_ready,
  PE_wrapper_17__ap_done,
  PE_wrapper_17__ap_idle,
  PE_wrapper_18__ap_start,
  PE_wrapper_18__ap_ready,
  PE_wrapper_18__ap_done,
  PE_wrapper_18__ap_idle,
  PE_wrapper_19__ap_start,
  PE_wrapper_19__ap_ready,
  PE_wrapper_19__ap_done,
  PE_wrapper_19__ap_idle,
  PE_wrapper_20__ap_start,
  PE_wrapper_20__ap_ready,
  PE_wrapper_20__ap_done,
  PE_wrapper_20__ap_idle,
  PE_wrapper_21__ap_start,
  PE_wrapper_21__ap_ready,
  PE_wrapper_21__ap_done,
  PE_wrapper_21__ap_idle,
  PE_wrapper_22__ap_start,
  PE_wrapper_22__ap_ready,
  PE_wrapper_22__ap_done,
  PE_wrapper_22__ap_idle,
  PE_wrapper_23__ap_start,
  PE_wrapper_23__ap_ready,
  PE_wrapper_23__ap_done,
  PE_wrapper_23__ap_idle,
  PE_wrapper_24__ap_start,
  PE_wrapper_24__ap_ready,
  PE_wrapper_24__ap_done,
  PE_wrapper_24__ap_idle,
  PE_wrapper_25__ap_start,
  PE_wrapper_25__ap_ready,
  PE_wrapper_25__ap_done,
  PE_wrapper_25__ap_idle,
  PE_wrapper_26__ap_start,
  PE_wrapper_26__ap_ready,
  PE_wrapper_26__ap_done,
  PE_wrapper_26__ap_idle,
  PE_wrapper_27__ap_start,
  PE_wrapper_27__ap_ready,
  PE_wrapper_27__ap_done,
  PE_wrapper_27__ap_idle,
  PE_wrapper_28__ap_start,
  PE_wrapper_28__ap_ready,
  PE_wrapper_28__ap_done,
  PE_wrapper_28__ap_idle,
  PE_wrapper_29__ap_start,
  PE_wrapper_29__ap_ready,
  PE_wrapper_29__ap_done,
  PE_wrapper_29__ap_idle,
  PE_wrapper_30__ap_start,
  PE_wrapper_30__ap_ready,
  PE_wrapper_30__ap_done,
  PE_wrapper_30__ap_idle,
  PE_wrapper_31__ap_start,
  PE_wrapper_31__ap_ready,
  PE_wrapper_31__ap_done,
  PE_wrapper_31__ap_idle,
  PE_wrapper_32__ap_start,
  PE_wrapper_32__ap_ready,
  PE_wrapper_32__ap_done,
  PE_wrapper_32__ap_idle,
  PE_wrapper_33__ap_start,
  PE_wrapper_33__ap_ready,
  PE_wrapper_33__ap_done,
  PE_wrapper_33__ap_idle,
  PE_wrapper_34__ap_start,
  PE_wrapper_34__ap_ready,
  PE_wrapper_34__ap_done,
  PE_wrapper_34__ap_idle,
  PE_wrapper_35__ap_start,
  PE_wrapper_35__ap_ready,
  PE_wrapper_35__ap_done,
  PE_wrapper_35__ap_idle,
  PE_wrapper_36__ap_start,
  PE_wrapper_36__ap_ready,
  PE_wrapper_36__ap_done,
  PE_wrapper_36__ap_idle,
  PE_wrapper_37__ap_start,
  PE_wrapper_37__ap_ready,
  PE_wrapper_37__ap_done,
  PE_wrapper_37__ap_idle,
  PE_wrapper_38__ap_start,
  PE_wrapper_38__ap_ready,
  PE_wrapper_38__ap_done,
  PE_wrapper_38__ap_idle,
  PE_wrapper_39__ap_start,
  PE_wrapper_39__ap_ready,
  PE_wrapper_39__ap_done,
  PE_wrapper_39__ap_idle,
  PE_wrapper_40__ap_start,
  PE_wrapper_40__ap_ready,
  PE_wrapper_40__ap_done,
  PE_wrapper_40__ap_idle,
  PE_wrapper_41__ap_start,
  PE_wrapper_41__ap_ready,
  PE_wrapper_41__ap_done,
  PE_wrapper_41__ap_idle,
  PE_wrapper_42__ap_start,
  PE_wrapper_42__ap_ready,
  PE_wrapper_42__ap_done,
  PE_wrapper_42__ap_idle,
  PE_wrapper_43__ap_start,
  PE_wrapper_43__ap_ready,
  PE_wrapper_43__ap_done,
  PE_wrapper_43__ap_idle,
  PE_wrapper_44__ap_start,
  PE_wrapper_44__ap_ready,
  PE_wrapper_44__ap_done,
  PE_wrapper_44__ap_idle,
  PE_wrapper_45__ap_start,
  PE_wrapper_45__ap_ready,
  PE_wrapper_45__ap_done,
  PE_wrapper_45__ap_idle,
  PE_wrapper_46__ap_start,
  PE_wrapper_46__ap_ready,
  PE_wrapper_46__ap_done,
  PE_wrapper_46__ap_idle,
  PE_wrapper_47__ap_start,
  PE_wrapper_47__ap_ready,
  PE_wrapper_47__ap_done,
  PE_wrapper_47__ap_idle,
  PE_wrapper_48__ap_start,
  PE_wrapper_48__ap_ready,
  PE_wrapper_48__ap_done,
  PE_wrapper_48__ap_idle,
  PE_wrapper_49__ap_start,
  PE_wrapper_49__ap_ready,
  PE_wrapper_49__ap_done,
  PE_wrapper_49__ap_idle,
  PE_wrapper_50__ap_start,
  PE_wrapper_50__ap_ready,
  PE_wrapper_50__ap_done,
  PE_wrapper_50__ap_idle,
  PE_wrapper_51__ap_start,
  PE_wrapper_51__ap_ready,
  PE_wrapper_51__ap_done,
  PE_wrapper_51__ap_idle,
  PE_wrapper_52__ap_start,
  PE_wrapper_52__ap_ready,
  PE_wrapper_52__ap_done,
  PE_wrapper_52__ap_idle,
  PE_wrapper_53__ap_start,
  PE_wrapper_53__ap_ready,
  PE_wrapper_53__ap_done,
  PE_wrapper_53__ap_idle,
  PE_wrapper_54__ap_start,
  PE_wrapper_54__ap_ready,
  PE_wrapper_54__ap_done,
  PE_wrapper_54__ap_idle,
  PE_wrapper_55__ap_start,
  PE_wrapper_55__ap_ready,
  PE_wrapper_55__ap_done,
  PE_wrapper_55__ap_idle,
  PE_wrapper_56__ap_start,
  PE_wrapper_56__ap_ready,
  PE_wrapper_56__ap_done,
  PE_wrapper_56__ap_idle,
  PE_wrapper_57__ap_start,
  PE_wrapper_57__ap_ready,
  PE_wrapper_57__ap_done,
  PE_wrapper_57__ap_idle,
  PE_wrapper_58__ap_start,
  PE_wrapper_58__ap_ready,
  PE_wrapper_58__ap_done,
  PE_wrapper_58__ap_idle,
  PE_wrapper_59__ap_start,
  PE_wrapper_59__ap_ready,
  PE_wrapper_59__ap_done,
  PE_wrapper_59__ap_idle,
  PE_wrapper_60__ap_start,
  PE_wrapper_60__ap_ready,
  PE_wrapper_60__ap_done,
  PE_wrapper_60__ap_idle,
  PE_wrapper_61__ap_start,
  PE_wrapper_61__ap_ready,
  PE_wrapper_61__ap_done,
  PE_wrapper_61__ap_idle,
  PE_wrapper_62__ap_start,
  PE_wrapper_62__ap_ready,
  PE_wrapper_62__ap_done,
  PE_wrapper_62__ap_idle,
  PE_wrapper_63__ap_start,
  PE_wrapper_63__ap_ready,
  PE_wrapper_63__ap_done,
  PE_wrapper_63__ap_idle,
  PE_wrapper_64__ap_start,
  PE_wrapper_64__ap_ready,
  PE_wrapper_64__ap_done,
  PE_wrapper_64__ap_idle,
  PE_wrapper_65__ap_start,
  PE_wrapper_65__ap_ready,
  PE_wrapper_65__ap_done,
  PE_wrapper_65__ap_idle,
  PE_wrapper_66__ap_start,
  PE_wrapper_66__ap_ready,
  PE_wrapper_66__ap_done,
  PE_wrapper_66__ap_idle,
  PE_wrapper_67__ap_start,
  PE_wrapper_67__ap_ready,
  PE_wrapper_67__ap_done,
  PE_wrapper_67__ap_idle,
  PE_wrapper_68__ap_start,
  PE_wrapper_68__ap_ready,
  PE_wrapper_68__ap_done,
  PE_wrapper_68__ap_idle,
  PE_wrapper_69__ap_start,
  PE_wrapper_69__ap_ready,
  PE_wrapper_69__ap_done,
  PE_wrapper_69__ap_idle,
  PE_wrapper_70__ap_start,
  PE_wrapper_70__ap_ready,
  PE_wrapper_70__ap_done,
  PE_wrapper_70__ap_idle,
  PE_wrapper_71__ap_start,
  PE_wrapper_71__ap_ready,
  PE_wrapper_71__ap_done,
  PE_wrapper_71__ap_idle,
  PE_wrapper_72__ap_start,
  PE_wrapper_72__ap_ready,
  PE_wrapper_72__ap_done,
  PE_wrapper_72__ap_idle,
  PE_wrapper_73__ap_start,
  PE_wrapper_73__ap_ready,
  PE_wrapper_73__ap_done,
  PE_wrapper_73__ap_idle,
  PE_wrapper_74__ap_start,
  PE_wrapper_74__ap_ready,
  PE_wrapper_74__ap_done,
  PE_wrapper_74__ap_idle,
  PE_wrapper_75__ap_start,
  PE_wrapper_75__ap_ready,
  PE_wrapper_75__ap_done,
  PE_wrapper_75__ap_idle,
  PE_wrapper_76__ap_start,
  PE_wrapper_76__ap_ready,
  PE_wrapper_76__ap_done,
  PE_wrapper_76__ap_idle,
  PE_wrapper_77__ap_start,
  PE_wrapper_77__ap_ready,
  PE_wrapper_77__ap_done,
  PE_wrapper_77__ap_idle,
  PE_wrapper_78__ap_start,
  PE_wrapper_78__ap_ready,
  PE_wrapper_78__ap_done,
  PE_wrapper_78__ap_idle,
  PE_wrapper_79__ap_start,
  PE_wrapper_79__ap_ready,
  PE_wrapper_79__ap_done,
  PE_wrapper_79__ap_idle,
  PE_wrapper_80__ap_start,
  PE_wrapper_80__ap_ready,
  PE_wrapper_80__ap_done,
  PE_wrapper_80__ap_idle,
  PE_wrapper_81__ap_start,
  PE_wrapper_81__ap_ready,
  PE_wrapper_81__ap_done,
  PE_wrapper_81__ap_idle,
  PE_wrapper_82__ap_start,
  PE_wrapper_82__ap_ready,
  PE_wrapper_82__ap_done,
  PE_wrapper_82__ap_idle,
  PE_wrapper_83__ap_start,
  PE_wrapper_83__ap_ready,
  PE_wrapper_83__ap_done,
  PE_wrapper_83__ap_idle,
  PE_wrapper_84__ap_start,
  PE_wrapper_84__ap_ready,
  PE_wrapper_84__ap_done,
  PE_wrapper_84__ap_idle,
  PE_wrapper_85__ap_start,
  PE_wrapper_85__ap_ready,
  PE_wrapper_85__ap_done,
  PE_wrapper_85__ap_idle,
  PE_wrapper_86__ap_start,
  PE_wrapper_86__ap_ready,
  PE_wrapper_86__ap_done,
  PE_wrapper_86__ap_idle,
  PE_wrapper_87__ap_start,
  PE_wrapper_87__ap_ready,
  PE_wrapper_87__ap_done,
  PE_wrapper_87__ap_idle,
  PE_wrapper_88__ap_start,
  PE_wrapper_88__ap_ready,
  PE_wrapper_88__ap_done,
  PE_wrapper_88__ap_idle,
  PE_wrapper_89__ap_start,
  PE_wrapper_89__ap_ready,
  PE_wrapper_89__ap_done,
  PE_wrapper_89__ap_idle,
  PE_wrapper_90__ap_start,
  PE_wrapper_90__ap_ready,
  PE_wrapper_90__ap_done,
  PE_wrapper_90__ap_idle,
  PE_wrapper_91__ap_start,
  PE_wrapper_91__ap_ready,
  PE_wrapper_91__ap_done,
  PE_wrapper_91__ap_idle,
  PE_wrapper_92__ap_start,
  PE_wrapper_92__ap_ready,
  PE_wrapper_92__ap_done,
  PE_wrapper_92__ap_idle,
  PE_wrapper_93__ap_start,
  PE_wrapper_93__ap_ready,
  PE_wrapper_93__ap_done,
  PE_wrapper_93__ap_idle,
  PE_wrapper_94__ap_start,
  PE_wrapper_94__ap_ready,
  PE_wrapper_94__ap_done,
  PE_wrapper_94__ap_idle,
  PE_wrapper_95__ap_start,
  PE_wrapper_95__ap_ready,
  PE_wrapper_95__ap_done,
  PE_wrapper_95__ap_idle,
  PE_wrapper_96__ap_start,
  PE_wrapper_96__ap_ready,
  PE_wrapper_96__ap_done,
  PE_wrapper_96__ap_idle,
  PE_wrapper_97__ap_start,
  PE_wrapper_97__ap_ready,
  PE_wrapper_97__ap_done,
  PE_wrapper_97__ap_idle,
  PE_wrapper_98__ap_start,
  PE_wrapper_98__ap_ready,
  PE_wrapper_98__ap_done,
  PE_wrapper_98__ap_idle,
  PE_wrapper_99__ap_start,
  PE_wrapper_99__ap_ready,
  PE_wrapper_99__ap_done,
  PE_wrapper_99__ap_idle,
  PE_wrapper_100__ap_start,
  PE_wrapper_100__ap_ready,
  PE_wrapper_100__ap_done,
  PE_wrapper_100__ap_idle,
  PE_wrapper_101__ap_start,
  PE_wrapper_101__ap_ready,
  PE_wrapper_101__ap_done,
  PE_wrapper_101__ap_idle,
  PE_wrapper_102__ap_start,
  PE_wrapper_102__ap_ready,
  PE_wrapper_102__ap_done,
  PE_wrapper_102__ap_idle,
  PE_wrapper_103__ap_start,
  PE_wrapper_103__ap_ready,
  PE_wrapper_103__ap_done,
  PE_wrapper_103__ap_idle,
  PE_wrapper_104__ap_start,
  PE_wrapper_104__ap_ready,
  PE_wrapper_104__ap_done,
  PE_wrapper_104__ap_idle,
  PE_wrapper_105__ap_start,
  PE_wrapper_105__ap_ready,
  PE_wrapper_105__ap_done,
  PE_wrapper_105__ap_idle,
  PE_wrapper_106__ap_start,
  PE_wrapper_106__ap_ready,
  PE_wrapper_106__ap_done,
  PE_wrapper_106__ap_idle,
  PE_wrapper_107__ap_start,
  PE_wrapper_107__ap_ready,
  PE_wrapper_107__ap_done,
  PE_wrapper_107__ap_idle,
  PE_wrapper_108__ap_start,
  PE_wrapper_108__ap_ready,
  PE_wrapper_108__ap_done,
  PE_wrapper_108__ap_idle,
  PE_wrapper_109__ap_start,
  PE_wrapper_109__ap_ready,
  PE_wrapper_109__ap_done,
  PE_wrapper_109__ap_idle,
  PE_wrapper_110__ap_start,
  PE_wrapper_110__ap_ready,
  PE_wrapper_110__ap_done,
  PE_wrapper_110__ap_idle,
  PE_wrapper_111__ap_start,
  PE_wrapper_111__ap_ready,
  PE_wrapper_111__ap_done,
  PE_wrapper_111__ap_idle,
  PE_wrapper_112__ap_start,
  PE_wrapper_112__ap_ready,
  PE_wrapper_112__ap_done,
  PE_wrapper_112__ap_idle,
  PE_wrapper_113__ap_start,
  PE_wrapper_113__ap_ready,
  PE_wrapper_113__ap_done,
  PE_wrapper_113__ap_idle,
  PE_wrapper_114__ap_start,
  PE_wrapper_114__ap_ready,
  PE_wrapper_114__ap_done,
  PE_wrapper_114__ap_idle,
  PE_wrapper_115__ap_start,
  PE_wrapper_115__ap_ready,
  PE_wrapper_115__ap_done,
  PE_wrapper_115__ap_idle,
  PE_wrapper_116__ap_start,
  PE_wrapper_116__ap_ready,
  PE_wrapper_116__ap_done,
  PE_wrapper_116__ap_idle,
  PE_wrapper_117__ap_start,
  PE_wrapper_117__ap_ready,
  PE_wrapper_117__ap_done,
  PE_wrapper_117__ap_idle,
  PE_wrapper_118__ap_start,
  PE_wrapper_118__ap_ready,
  PE_wrapper_118__ap_done,
  PE_wrapper_118__ap_idle,
  PE_wrapper_119__ap_start,
  PE_wrapper_119__ap_ready,
  PE_wrapper_119__ap_done,
  PE_wrapper_119__ap_idle,
  PE_wrapper_120__ap_start,
  PE_wrapper_120__ap_ready,
  PE_wrapper_120__ap_done,
  PE_wrapper_120__ap_idle,
  PE_wrapper_121__ap_start,
  PE_wrapper_121__ap_ready,
  PE_wrapper_121__ap_done,
  PE_wrapper_121__ap_idle,
  PE_wrapper_122__ap_start,
  PE_wrapper_122__ap_ready,
  PE_wrapper_122__ap_done,
  PE_wrapper_122__ap_idle,
  PE_wrapper_123__ap_start,
  PE_wrapper_123__ap_ready,
  PE_wrapper_123__ap_done,
  PE_wrapper_123__ap_idle,
  PE_wrapper_124__ap_start,
  PE_wrapper_124__ap_ready,
  PE_wrapper_124__ap_done,
  PE_wrapper_124__ap_idle,
  PE_wrapper_125__ap_start,
  PE_wrapper_125__ap_ready,
  PE_wrapper_125__ap_done,
  PE_wrapper_125__ap_idle,
  PE_wrapper_126__ap_start,
  PE_wrapper_126__ap_ready,
  PE_wrapper_126__ap_done,
  PE_wrapper_126__ap_idle,
  PE_wrapper_127__ap_start,
  PE_wrapper_127__ap_ready,
  PE_wrapper_127__ap_done,
  PE_wrapper_127__ap_idle,
  PE_wrapper_128__ap_start,
  PE_wrapper_128__ap_ready,
  PE_wrapper_128__ap_done,
  PE_wrapper_128__ap_idle,
  PE_wrapper_129__ap_start,
  PE_wrapper_129__ap_ready,
  PE_wrapper_129__ap_done,
  PE_wrapper_129__ap_idle,
  PE_wrapper_130__ap_start,
  PE_wrapper_130__ap_ready,
  PE_wrapper_130__ap_done,
  PE_wrapper_130__ap_idle,
  PE_wrapper_131__ap_start,
  PE_wrapper_131__ap_ready,
  PE_wrapper_131__ap_done,
  PE_wrapper_131__ap_idle,
  PE_wrapper_132__ap_start,
  PE_wrapper_132__ap_ready,
  PE_wrapper_132__ap_done,
  PE_wrapper_132__ap_idle,
  PE_wrapper_133__ap_start,
  PE_wrapper_133__ap_ready,
  PE_wrapper_133__ap_done,
  PE_wrapper_133__ap_idle,
  PE_wrapper_134__ap_start,
  PE_wrapper_134__ap_ready,
  PE_wrapper_134__ap_done,
  PE_wrapper_134__ap_idle,
  PE_wrapper_135__ap_start,
  PE_wrapper_135__ap_ready,
  PE_wrapper_135__ap_done,
  PE_wrapper_135__ap_idle,
  PE_wrapper_136__ap_start,
  PE_wrapper_136__ap_ready,
  PE_wrapper_136__ap_done,
  PE_wrapper_136__ap_idle,
  PE_wrapper_137__ap_start,
  PE_wrapper_137__ap_ready,
  PE_wrapper_137__ap_done,
  PE_wrapper_137__ap_idle,
  PE_wrapper_138__ap_start,
  PE_wrapper_138__ap_ready,
  PE_wrapper_138__ap_done,
  PE_wrapper_138__ap_idle,
  PE_wrapper_139__ap_start,
  PE_wrapper_139__ap_ready,
  PE_wrapper_139__ap_done,
  PE_wrapper_139__ap_idle,
  PE_wrapper_140__ap_start,
  PE_wrapper_140__ap_ready,
  PE_wrapper_140__ap_done,
  PE_wrapper_140__ap_idle,
  PE_wrapper_141__ap_start,
  PE_wrapper_141__ap_ready,
  PE_wrapper_141__ap_done,
  PE_wrapper_141__ap_idle,
  PE_wrapper_142__ap_start,
  PE_wrapper_142__ap_ready,
  PE_wrapper_142__ap_done,
  PE_wrapper_142__ap_idle,
  PE_wrapper_143__ap_start,
  PE_wrapper_143__ap_ready,
  PE_wrapper_143__ap_done,
  PE_wrapper_143__ap_idle,
  PE_wrapper_144__ap_start,
  PE_wrapper_144__ap_ready,
  PE_wrapper_144__ap_done,
  PE_wrapper_144__ap_idle,
  PE_wrapper_145__ap_start,
  PE_wrapper_145__ap_ready,
  PE_wrapper_145__ap_done,
  PE_wrapper_145__ap_idle,
  PE_wrapper_146__ap_start,
  PE_wrapper_146__ap_ready,
  PE_wrapper_146__ap_done,
  PE_wrapper_146__ap_idle,
  PE_wrapper_147__ap_start,
  PE_wrapper_147__ap_ready,
  PE_wrapper_147__ap_done,
  PE_wrapper_147__ap_idle,
  PE_wrapper_148__ap_start,
  PE_wrapper_148__ap_ready,
  PE_wrapper_148__ap_done,
  PE_wrapper_148__ap_idle,
  PE_wrapper_149__ap_start,
  PE_wrapper_149__ap_ready,
  PE_wrapper_149__ap_done,
  PE_wrapper_149__ap_idle,
  PE_wrapper_150__ap_start,
  PE_wrapper_150__ap_ready,
  PE_wrapper_150__ap_done,
  PE_wrapper_150__ap_idle,
  PE_wrapper_151__ap_start,
  PE_wrapper_151__ap_ready,
  PE_wrapper_151__ap_done,
  PE_wrapper_151__ap_idle,
  PE_wrapper_152__ap_start,
  PE_wrapper_152__ap_ready,
  PE_wrapper_152__ap_done,
  PE_wrapper_152__ap_idle,
  PE_wrapper_153__ap_start,
  PE_wrapper_153__ap_ready,
  PE_wrapper_153__ap_done,
  PE_wrapper_153__ap_idle,
  PE_wrapper_154__ap_start,
  PE_wrapper_154__ap_ready,
  PE_wrapper_154__ap_done,
  PE_wrapper_154__ap_idle,
  PE_wrapper_155__ap_start,
  PE_wrapper_155__ap_ready,
  PE_wrapper_155__ap_done,
  PE_wrapper_155__ap_idle,
  PE_wrapper_156__ap_start,
  PE_wrapper_156__ap_ready,
  PE_wrapper_156__ap_done,
  PE_wrapper_156__ap_idle,
  PE_wrapper_157__ap_start,
  PE_wrapper_157__ap_ready,
  PE_wrapper_157__ap_done,
  PE_wrapper_157__ap_idle,
  PE_wrapper_158__ap_start,
  PE_wrapper_158__ap_ready,
  PE_wrapper_158__ap_done,
  PE_wrapper_158__ap_idle,
  PE_wrapper_159__ap_start,
  PE_wrapper_159__ap_ready,
  PE_wrapper_159__ap_done,
  PE_wrapper_159__ap_idle,
  PE_wrapper_160__ap_start,
  PE_wrapper_160__ap_ready,
  PE_wrapper_160__ap_done,
  PE_wrapper_160__ap_idle,
  PE_wrapper_161__ap_start,
  PE_wrapper_161__ap_ready,
  PE_wrapper_161__ap_done,
  PE_wrapper_161__ap_idle,
  PE_wrapper_162__ap_start,
  PE_wrapper_162__ap_ready,
  PE_wrapper_162__ap_done,
  PE_wrapper_162__ap_idle,
  PE_wrapper_163__ap_start,
  PE_wrapper_163__ap_ready,
  PE_wrapper_163__ap_done,
  PE_wrapper_163__ap_idle,
  PE_wrapper_164__ap_start,
  PE_wrapper_164__ap_ready,
  PE_wrapper_164__ap_done,
  PE_wrapper_164__ap_idle,
  PE_wrapper_165__ap_start,
  PE_wrapper_165__ap_ready,
  PE_wrapper_165__ap_done,
  PE_wrapper_165__ap_idle,
  PE_wrapper_166__ap_start,
  PE_wrapper_166__ap_ready,
  PE_wrapper_166__ap_done,
  PE_wrapper_166__ap_idle,
  PE_wrapper_167__ap_start,
  PE_wrapper_167__ap_ready,
  PE_wrapper_167__ap_done,
  PE_wrapper_167__ap_idle,
  PE_wrapper_168__ap_start,
  PE_wrapper_168__ap_ready,
  PE_wrapper_168__ap_done,
  PE_wrapper_168__ap_idle,
  PE_wrapper_169__ap_start,
  PE_wrapper_169__ap_ready,
  PE_wrapper_169__ap_done,
  PE_wrapper_169__ap_idle,
  PE_wrapper_170__ap_start,
  PE_wrapper_170__ap_ready,
  PE_wrapper_170__ap_done,
  PE_wrapper_170__ap_idle,
  PE_wrapper_171__ap_start,
  PE_wrapper_171__ap_ready,
  PE_wrapper_171__ap_done,
  PE_wrapper_171__ap_idle,
  PE_wrapper_172__ap_start,
  PE_wrapper_172__ap_ready,
  PE_wrapper_172__ap_done,
  PE_wrapper_172__ap_idle,
  PE_wrapper_173__ap_start,
  PE_wrapper_173__ap_ready,
  PE_wrapper_173__ap_done,
  PE_wrapper_173__ap_idle,
  PE_wrapper_174__ap_start,
  PE_wrapper_174__ap_ready,
  PE_wrapper_174__ap_done,
  PE_wrapper_174__ap_idle,
  PE_wrapper_175__ap_start,
  PE_wrapper_175__ap_ready,
  PE_wrapper_175__ap_done,
  PE_wrapper_175__ap_idle,
  PE_wrapper_176__ap_start,
  PE_wrapper_176__ap_ready,
  PE_wrapper_176__ap_done,
  PE_wrapper_176__ap_idle,
  PE_wrapper_177__ap_start,
  PE_wrapper_177__ap_ready,
  PE_wrapper_177__ap_done,
  PE_wrapper_177__ap_idle,
  PE_wrapper_178__ap_start,
  PE_wrapper_178__ap_ready,
  PE_wrapper_178__ap_done,
  PE_wrapper_178__ap_idle,
  PE_wrapper_179__ap_start,
  PE_wrapper_179__ap_ready,
  PE_wrapper_179__ap_done,
  PE_wrapper_179__ap_idle,
  PE_wrapper_180__ap_start,
  PE_wrapper_180__ap_ready,
  PE_wrapper_180__ap_done,
  PE_wrapper_180__ap_idle,
  PE_wrapper_181__ap_start,
  PE_wrapper_181__ap_ready,
  PE_wrapper_181__ap_done,
  PE_wrapper_181__ap_idle,
  PE_wrapper_182__ap_start,
  PE_wrapper_182__ap_ready,
  PE_wrapper_182__ap_done,
  PE_wrapper_182__ap_idle,
  PE_wrapper_183__ap_start,
  PE_wrapper_183__ap_ready,
  PE_wrapper_183__ap_done,
  PE_wrapper_183__ap_idle,
  PE_wrapper_184__ap_start,
  PE_wrapper_184__ap_ready,
  PE_wrapper_184__ap_done,
  PE_wrapper_184__ap_idle,
  PE_wrapper_185__ap_start,
  PE_wrapper_185__ap_ready,
  PE_wrapper_185__ap_done,
  PE_wrapper_185__ap_idle,
  PE_wrapper_186__ap_start,
  PE_wrapper_186__ap_ready,
  PE_wrapper_186__ap_done,
  PE_wrapper_186__ap_idle,
  PE_wrapper_187__ap_start,
  PE_wrapper_187__ap_ready,
  PE_wrapper_187__ap_done,
  PE_wrapper_187__ap_idle,
  PE_wrapper_188__ap_start,
  PE_wrapper_188__ap_ready,
  PE_wrapper_188__ap_done,
  PE_wrapper_188__ap_idle,
  PE_wrapper_189__ap_start,
  PE_wrapper_189__ap_ready,
  PE_wrapper_189__ap_done,
  PE_wrapper_189__ap_idle,
  PE_wrapper_190__ap_start,
  PE_wrapper_190__ap_ready,
  PE_wrapper_190__ap_done,
  PE_wrapper_190__ap_idle,
  PE_wrapper_191__ap_start,
  PE_wrapper_191__ap_ready,
  PE_wrapper_191__ap_done,
  PE_wrapper_191__ap_idle,
  PE_wrapper_192__ap_start,
  PE_wrapper_192__ap_ready,
  PE_wrapper_192__ap_done,
  PE_wrapper_192__ap_idle,
  PE_wrapper_193__ap_start,
  PE_wrapper_193__ap_ready,
  PE_wrapper_193__ap_done,
  PE_wrapper_193__ap_idle,
  PE_wrapper_194__ap_start,
  PE_wrapper_194__ap_ready,
  PE_wrapper_194__ap_done,
  PE_wrapper_194__ap_idle,
  PE_wrapper_195__ap_start,
  PE_wrapper_195__ap_ready,
  PE_wrapper_195__ap_done,
  PE_wrapper_195__ap_idle,
  PE_wrapper_196__ap_start,
  PE_wrapper_196__ap_ready,
  PE_wrapper_196__ap_done,
  PE_wrapper_196__ap_idle,
  PE_wrapper_197__ap_start,
  PE_wrapper_197__ap_ready,
  PE_wrapper_197__ap_done,
  PE_wrapper_197__ap_idle,
  PE_wrapper_198__ap_start,
  PE_wrapper_198__ap_ready,
  PE_wrapper_198__ap_done,
  PE_wrapper_198__ap_idle,
  PE_wrapper_199__ap_start,
  PE_wrapper_199__ap_ready,
  PE_wrapper_199__ap_done,
  PE_wrapper_199__ap_idle,
  PE_wrapper_200__ap_start,
  PE_wrapper_200__ap_ready,
  PE_wrapper_200__ap_done,
  PE_wrapper_200__ap_idle,
  PE_wrapper_201__ap_start,
  PE_wrapper_201__ap_ready,
  PE_wrapper_201__ap_done,
  PE_wrapper_201__ap_idle,
  PE_wrapper_202__ap_start,
  PE_wrapper_202__ap_ready,
  PE_wrapper_202__ap_done,
  PE_wrapper_202__ap_idle,
  PE_wrapper_203__ap_start,
  PE_wrapper_203__ap_ready,
  PE_wrapper_203__ap_done,
  PE_wrapper_203__ap_idle,
  PE_wrapper_204__ap_start,
  PE_wrapper_204__ap_ready,
  PE_wrapper_204__ap_done,
  PE_wrapper_204__ap_idle,
  PE_wrapper_205__ap_start,
  PE_wrapper_205__ap_ready,
  PE_wrapper_205__ap_done,
  PE_wrapper_205__ap_idle,
  PE_wrapper_206__ap_start,
  PE_wrapper_206__ap_ready,
  PE_wrapper_206__ap_done,
  PE_wrapper_206__ap_idle,
  PE_wrapper_207__ap_start,
  PE_wrapper_207__ap_ready,
  PE_wrapper_207__ap_done,
  PE_wrapper_207__ap_idle,
  PE_wrapper_208__ap_start,
  PE_wrapper_208__ap_ready,
  PE_wrapper_208__ap_done,
  PE_wrapper_208__ap_idle,
  PE_wrapper_209__ap_start,
  PE_wrapper_209__ap_ready,
  PE_wrapper_209__ap_done,
  PE_wrapper_209__ap_idle,
  PE_wrapper_210__ap_start,
  PE_wrapper_210__ap_ready,
  PE_wrapper_210__ap_done,
  PE_wrapper_210__ap_idle,
  PE_wrapper_211__ap_start,
  PE_wrapper_211__ap_ready,
  PE_wrapper_211__ap_done,
  PE_wrapper_211__ap_idle,
  PE_wrapper_212__ap_start,
  PE_wrapper_212__ap_ready,
  PE_wrapper_212__ap_done,
  PE_wrapper_212__ap_idle,
  PE_wrapper_213__ap_start,
  PE_wrapper_213__ap_ready,
  PE_wrapper_213__ap_done,
  PE_wrapper_213__ap_idle,
  PE_wrapper_214__ap_start,
  PE_wrapper_214__ap_ready,
  PE_wrapper_214__ap_done,
  PE_wrapper_214__ap_idle,
  PE_wrapper_215__ap_start,
  PE_wrapper_215__ap_ready,
  PE_wrapper_215__ap_done,
  PE_wrapper_215__ap_idle,
  PE_wrapper_216__ap_start,
  PE_wrapper_216__ap_ready,
  PE_wrapper_216__ap_done,
  PE_wrapper_216__ap_idle,
  PE_wrapper_217__ap_start,
  PE_wrapper_217__ap_ready,
  PE_wrapper_217__ap_done,
  PE_wrapper_217__ap_idle,
  PE_wrapper_218__ap_start,
  PE_wrapper_218__ap_ready,
  PE_wrapper_218__ap_done,
  PE_wrapper_218__ap_idle,
  PE_wrapper_219__ap_start,
  PE_wrapper_219__ap_ready,
  PE_wrapper_219__ap_done,
  PE_wrapper_219__ap_idle,
  PE_wrapper_220__ap_start,
  PE_wrapper_220__ap_ready,
  PE_wrapper_220__ap_done,
  PE_wrapper_220__ap_idle,
  PE_wrapper_221__ap_start,
  PE_wrapper_221__ap_ready,
  PE_wrapper_221__ap_done,
  PE_wrapper_221__ap_idle,
  PE_wrapper_222__ap_start,
  PE_wrapper_222__ap_ready,
  PE_wrapper_222__ap_done,
  PE_wrapper_222__ap_idle,
  PE_wrapper_223__ap_start,
  PE_wrapper_223__ap_ready,
  PE_wrapper_223__ap_done,
  PE_wrapper_223__ap_idle,
  PE_wrapper_224__ap_start,
  PE_wrapper_224__ap_ready,
  PE_wrapper_224__ap_done,
  PE_wrapper_224__ap_idle,
  PE_wrapper_225__ap_start,
  PE_wrapper_225__ap_ready,
  PE_wrapper_225__ap_done,
  PE_wrapper_225__ap_idle,
  PE_wrapper_226__ap_start,
  PE_wrapper_226__ap_ready,
  PE_wrapper_226__ap_done,
  PE_wrapper_226__ap_idle,
  PE_wrapper_227__ap_start,
  PE_wrapper_227__ap_ready,
  PE_wrapper_227__ap_done,
  PE_wrapper_227__ap_idle,
  PE_wrapper_228__ap_start,
  PE_wrapper_228__ap_ready,
  PE_wrapper_228__ap_done,
  PE_wrapper_228__ap_idle,
  PE_wrapper_229__ap_start,
  PE_wrapper_229__ap_ready,
  PE_wrapper_229__ap_done,
  PE_wrapper_229__ap_idle,
  PE_wrapper_230__ap_start,
  PE_wrapper_230__ap_ready,
  PE_wrapper_230__ap_done,
  PE_wrapper_230__ap_idle,
  PE_wrapper_231__ap_start,
  PE_wrapper_231__ap_ready,
  PE_wrapper_231__ap_done,
  PE_wrapper_231__ap_idle,
  PE_wrapper_232__ap_start,
  PE_wrapper_232__ap_ready,
  PE_wrapper_232__ap_done,
  PE_wrapper_232__ap_idle,
  PE_wrapper_233__ap_start,
  PE_wrapper_233__ap_ready,
  PE_wrapper_233__ap_done,
  PE_wrapper_233__ap_idle,
  PE_wrapper_234__ap_start,
  PE_wrapper_234__ap_ready,
  PE_wrapper_234__ap_done,
  PE_wrapper_234__ap_idle,
  PE_wrapper_235__ap_start,
  PE_wrapper_235__ap_ready,
  PE_wrapper_235__ap_done,
  PE_wrapper_235__ap_idle,
  PE_wrapper_236__ap_start,
  PE_wrapper_236__ap_ready,
  PE_wrapper_236__ap_done,
  PE_wrapper_236__ap_idle,
  PE_wrapper_237__ap_start,
  PE_wrapper_237__ap_ready,
  PE_wrapper_237__ap_done,
  PE_wrapper_237__ap_idle,
  PE_wrapper_238__ap_start,
  PE_wrapper_238__ap_ready,
  PE_wrapper_238__ap_done,
  PE_wrapper_238__ap_idle,
  PE_wrapper_239__ap_start,
  PE_wrapper_239__ap_ready,
  PE_wrapper_239__ap_done,
  PE_wrapper_239__ap_idle,
  PE_wrapper_240__ap_start,
  PE_wrapper_240__ap_ready,
  PE_wrapper_240__ap_done,
  PE_wrapper_240__ap_idle,
  PE_wrapper_241__ap_start,
  PE_wrapper_241__ap_ready,
  PE_wrapper_241__ap_done,
  PE_wrapper_241__ap_idle,
  PE_wrapper_242__ap_start,
  PE_wrapper_242__ap_ready,
  PE_wrapper_242__ap_done,
  PE_wrapper_242__ap_idle,
  PE_wrapper_243__ap_start,
  PE_wrapper_243__ap_ready,
  PE_wrapper_243__ap_done,
  PE_wrapper_243__ap_idle,
  PE_wrapper_244__ap_start,
  PE_wrapper_244__ap_ready,
  PE_wrapper_244__ap_done,
  PE_wrapper_244__ap_idle,
  PE_wrapper_245__ap_start,
  PE_wrapper_245__ap_ready,
  PE_wrapper_245__ap_done,
  PE_wrapper_245__ap_idle,
  PE_wrapper_246__ap_start,
  PE_wrapper_246__ap_ready,
  PE_wrapper_246__ap_done,
  PE_wrapper_246__ap_idle,
  PE_wrapper_247__ap_start,
  PE_wrapper_247__ap_ready,
  PE_wrapper_247__ap_done,
  PE_wrapper_247__ap_idle,
  PE_wrapper_248__ap_start,
  PE_wrapper_248__ap_ready,
  PE_wrapper_248__ap_done,
  PE_wrapper_248__ap_idle,
  PE_wrapper_249__ap_start,
  PE_wrapper_249__ap_ready,
  PE_wrapper_249__ap_done,
  PE_wrapper_249__ap_idle,
  PE_wrapper_250__ap_start,
  PE_wrapper_250__ap_ready,
  PE_wrapper_250__ap_done,
  PE_wrapper_250__ap_idle,
  PE_wrapper_251__ap_start,
  PE_wrapper_251__ap_ready,
  PE_wrapper_251__ap_done,
  PE_wrapper_251__ap_idle,
  PE_wrapper_252__ap_start,
  PE_wrapper_252__ap_ready,
  PE_wrapper_252__ap_done,
  PE_wrapper_252__ap_idle,
  PE_wrapper_253__ap_start,
  PE_wrapper_253__ap_ready,
  PE_wrapper_253__ap_done,
  PE_wrapper_253__ap_idle,
  PE_wrapper_254__ap_start,
  PE_wrapper_254__ap_ready,
  PE_wrapper_254__ap_done,
  PE_wrapper_254__ap_idle,
  PE_wrapper_255__ap_start,
  PE_wrapper_255__ap_ready,
  PE_wrapper_255__ap_done,
  PE_wrapper_255__ap_idle,
  PE_wrapper_256__ap_start,
  PE_wrapper_256__ap_ready,
  PE_wrapper_256__ap_done,
  PE_wrapper_256__ap_idle,
  PE_wrapper_257__ap_start,
  PE_wrapper_257__ap_ready,
  PE_wrapper_257__ap_done,
  PE_wrapper_257__ap_idle,
  PE_wrapper_258__ap_start,
  PE_wrapper_258__ap_ready,
  PE_wrapper_258__ap_done,
  PE_wrapper_258__ap_idle,
  PE_wrapper_259__ap_start,
  PE_wrapper_259__ap_ready,
  PE_wrapper_259__ap_done,
  PE_wrapper_259__ap_idle,
  PE_wrapper_260__ap_start,
  PE_wrapper_260__ap_ready,
  PE_wrapper_260__ap_done,
  PE_wrapper_260__ap_idle,
  PE_wrapper_261__ap_start,
  PE_wrapper_261__ap_ready,
  PE_wrapper_261__ap_done,
  PE_wrapper_261__ap_idle,
  PE_wrapper_262__ap_start,
  PE_wrapper_262__ap_ready,
  PE_wrapper_262__ap_done,
  PE_wrapper_262__ap_idle,
  PE_wrapper_263__ap_start,
  PE_wrapper_263__ap_ready,
  PE_wrapper_263__ap_done,
  PE_wrapper_263__ap_idle,
  PE_wrapper_264__ap_start,
  PE_wrapper_264__ap_ready,
  PE_wrapper_264__ap_done,
  PE_wrapper_264__ap_idle,
  PE_wrapper_265__ap_start,
  PE_wrapper_265__ap_ready,
  PE_wrapper_265__ap_done,
  PE_wrapper_265__ap_idle,
  PE_wrapper_266__ap_start,
  PE_wrapper_266__ap_ready,
  PE_wrapper_266__ap_done,
  PE_wrapper_266__ap_idle,
  PE_wrapper_267__ap_start,
  PE_wrapper_267__ap_ready,
  PE_wrapper_267__ap_done,
  PE_wrapper_267__ap_idle,
  PE_wrapper_268__ap_start,
  PE_wrapper_268__ap_ready,
  PE_wrapper_268__ap_done,
  PE_wrapper_268__ap_idle,
  PE_wrapper_269__ap_start,
  PE_wrapper_269__ap_ready,
  PE_wrapper_269__ap_done,
  PE_wrapper_269__ap_idle,
  PE_wrapper_270__ap_start,
  PE_wrapper_270__ap_ready,
  PE_wrapper_270__ap_done,
  PE_wrapper_270__ap_idle,
  PE_wrapper_271__ap_start,
  PE_wrapper_271__ap_ready,
  PE_wrapper_271__ap_done,
  PE_wrapper_271__ap_idle,
  PE_wrapper_272__ap_start,
  PE_wrapper_272__ap_ready,
  PE_wrapper_272__ap_done,
  PE_wrapper_272__ap_idle,
  PE_wrapper_273__ap_start,
  PE_wrapper_273__ap_ready,
  PE_wrapper_273__ap_done,
  PE_wrapper_273__ap_idle,
  PE_wrapper_274__ap_start,
  PE_wrapper_274__ap_ready,
  PE_wrapper_274__ap_done,
  PE_wrapper_274__ap_idle,
  PE_wrapper_275__ap_start,
  PE_wrapper_275__ap_ready,
  PE_wrapper_275__ap_done,
  PE_wrapper_275__ap_idle,
  PE_wrapper_276__ap_start,
  PE_wrapper_276__ap_ready,
  PE_wrapper_276__ap_done,
  PE_wrapper_276__ap_idle,
  PE_wrapper_277__ap_start,
  PE_wrapper_277__ap_ready,
  PE_wrapper_277__ap_done,
  PE_wrapper_277__ap_idle,
  PE_wrapper_278__ap_start,
  PE_wrapper_278__ap_ready,
  PE_wrapper_278__ap_done,
  PE_wrapper_278__ap_idle,
  PE_wrapper_279__ap_start,
  PE_wrapper_279__ap_ready,
  PE_wrapper_279__ap_done,
  PE_wrapper_279__ap_idle,
  PE_wrapper_280__ap_start,
  PE_wrapper_280__ap_ready,
  PE_wrapper_280__ap_done,
  PE_wrapper_280__ap_idle,
  PE_wrapper_281__ap_start,
  PE_wrapper_281__ap_ready,
  PE_wrapper_281__ap_done,
  PE_wrapper_281__ap_idle,
  PE_wrapper_282__ap_start,
  PE_wrapper_282__ap_ready,
  PE_wrapper_282__ap_done,
  PE_wrapper_282__ap_idle,
  PE_wrapper_283__ap_start,
  PE_wrapper_283__ap_ready,
  PE_wrapper_283__ap_done,
  PE_wrapper_283__ap_idle,
  PE_wrapper_284__ap_start,
  PE_wrapper_284__ap_ready,
  PE_wrapper_284__ap_done,
  PE_wrapper_284__ap_idle,
  PE_wrapper_285__ap_start,
  PE_wrapper_285__ap_ready,
  PE_wrapper_285__ap_done,
  PE_wrapper_285__ap_idle,
  PE_wrapper_286__ap_start,
  PE_wrapper_286__ap_ready,
  PE_wrapper_286__ap_done,
  PE_wrapper_286__ap_idle,
  PE_wrapper_287__ap_start,
  PE_wrapper_287__ap_ready,
  PE_wrapper_287__ap_done,
  PE_wrapper_287__ap_idle,
  PE_wrapper_288__ap_start,
  PE_wrapper_288__ap_ready,
  PE_wrapper_288__ap_done,
  PE_wrapper_288__ap_idle,
  PE_wrapper_289__ap_start,
  PE_wrapper_289__ap_ready,
  PE_wrapper_289__ap_done,
  PE_wrapper_289__ap_idle,
  PE_wrapper_290__ap_start,
  PE_wrapper_290__ap_ready,
  PE_wrapper_290__ap_done,
  PE_wrapper_290__ap_idle,
  PE_wrapper_291__ap_start,
  PE_wrapper_291__ap_ready,
  PE_wrapper_291__ap_done,
  PE_wrapper_291__ap_idle,
  PE_wrapper_292__ap_start,
  PE_wrapper_292__ap_ready,
  PE_wrapper_292__ap_done,
  PE_wrapper_292__ap_idle,
  PE_wrapper_293__ap_start,
  PE_wrapper_293__ap_ready,
  PE_wrapper_293__ap_done,
  PE_wrapper_293__ap_idle,
  PE_wrapper_294__ap_start,
  PE_wrapper_294__ap_ready,
  PE_wrapper_294__ap_done,
  PE_wrapper_294__ap_idle,
  PE_wrapper_295__ap_start,
  PE_wrapper_295__ap_ready,
  PE_wrapper_295__ap_done,
  PE_wrapper_295__ap_idle,
  PE_wrapper_296__ap_start,
  PE_wrapper_296__ap_ready,
  PE_wrapper_296__ap_done,
  PE_wrapper_296__ap_idle,
  PE_wrapper_297__ap_start,
  PE_wrapper_297__ap_ready,
  PE_wrapper_297__ap_done,
  PE_wrapper_297__ap_idle,
  PE_wrapper_298__ap_start,
  PE_wrapper_298__ap_ready,
  PE_wrapper_298__ap_done,
  PE_wrapper_298__ap_idle,
  PE_wrapper_299__ap_start,
  PE_wrapper_299__ap_ready,
  PE_wrapper_299__ap_done,
  PE_wrapper_299__ap_idle,
  PE_wrapper_300__ap_start,
  PE_wrapper_300__ap_ready,
  PE_wrapper_300__ap_done,
  PE_wrapper_300__ap_idle,
  PE_wrapper_301__ap_start,
  PE_wrapper_301__ap_ready,
  PE_wrapper_301__ap_done,
  PE_wrapper_301__ap_idle,
  PE_wrapper_302__ap_start,
  PE_wrapper_302__ap_ready,
  PE_wrapper_302__ap_done,
  PE_wrapper_302__ap_idle,
  PE_wrapper_303__ap_start,
  PE_wrapper_303__ap_ready,
  PE_wrapper_303__ap_done,
  PE_wrapper_303__ap_idle,
  PE_wrapper_304__ap_start,
  PE_wrapper_304__ap_ready,
  PE_wrapper_304__ap_done,
  PE_wrapper_304__ap_idle,
  PE_wrapper_305__ap_start,
  PE_wrapper_305__ap_ready,
  PE_wrapper_305__ap_done,
  PE_wrapper_305__ap_idle
);

  // pragma RS clk port=ap_clk
  // pragma RS rst port=ap_rst_n active=low
  // pragma RS ap-ctrl ap_start=ap_start ap_done=ap_done ap_idle=ap_idle ap_ready=ap_ready scalar=(A|B|C)
  // pragma RS ap-ctrl ap_start=A_IO_L2_in_0__ap_start ap_done=A_IO_L2_in_0__ap_done ap_idle=A_IO_L2_in_0__ap_idle ap_ready=A_IO_L2_in_0__ap_ready
  // pragma RS ap-ctrl ap_start=A_IO_L2_in_1__ap_start ap_done=A_IO_L2_in_1__ap_done ap_idle=A_IO_L2_in_1__ap_idle ap_ready=A_IO_L2_in_1__ap_ready
  // pragma RS ap-ctrl ap_start=A_IO_L2_in_2__ap_start ap_done=A_IO_L2_in_2__ap_done ap_idle=A_IO_L2_in_2__ap_idle ap_ready=A_IO_L2_in_2__ap_ready
  // pragma RS ap-ctrl ap_start=A_IO_L2_in_3__ap_start ap_done=A_IO_L2_in_3__ap_done ap_idle=A_IO_L2_in_3__ap_idle ap_ready=A_IO_L2_in_3__ap_ready
  // pragma RS ap-ctrl ap_start=A_IO_L2_in_4__ap_start ap_done=A_IO_L2_in_4__ap_done ap_idle=A_IO_L2_in_4__ap_idle ap_ready=A_IO_L2_in_4__ap_ready
  // pragma RS ap-ctrl ap_start=A_IO_L2_in_5__ap_start ap_done=A_IO_L2_in_5__ap_done ap_idle=A_IO_L2_in_5__ap_idle ap_ready=A_IO_L2_in_5__ap_ready
  // pragma RS ap-ctrl ap_start=A_IO_L2_in_6__ap_start ap_done=A_IO_L2_in_6__ap_done ap_idle=A_IO_L2_in_6__ap_idle ap_ready=A_IO_L2_in_6__ap_ready
  // pragma RS ap-ctrl ap_start=A_IO_L2_in_7__ap_start ap_done=A_IO_L2_in_7__ap_done ap_idle=A_IO_L2_in_7__ap_idle ap_ready=A_IO_L2_in_7__ap_ready
  // pragma RS ap-ctrl ap_start=A_IO_L2_in_8__ap_start ap_done=A_IO_L2_in_8__ap_done ap_idle=A_IO_L2_in_8__ap_idle ap_ready=A_IO_L2_in_8__ap_ready
  // pragma RS ap-ctrl ap_start=A_IO_L2_in_9__ap_start ap_done=A_IO_L2_in_9__ap_done ap_idle=A_IO_L2_in_9__ap_idle ap_ready=A_IO_L2_in_9__ap_ready
  // pragma RS ap-ctrl ap_start=A_IO_L2_in_10__ap_start ap_done=A_IO_L2_in_10__ap_done ap_idle=A_IO_L2_in_10__ap_idle ap_ready=A_IO_L2_in_10__ap_ready
  // pragma RS ap-ctrl ap_start=A_IO_L2_in_11__ap_start ap_done=A_IO_L2_in_11__ap_done ap_idle=A_IO_L2_in_11__ap_idle ap_ready=A_IO_L2_in_11__ap_ready
  // pragma RS ap-ctrl ap_start=A_IO_L2_in_12__ap_start ap_done=A_IO_L2_in_12__ap_done ap_idle=A_IO_L2_in_12__ap_idle ap_ready=A_IO_L2_in_12__ap_ready
  // pragma RS ap-ctrl ap_start=A_IO_L2_in_13__ap_start ap_done=A_IO_L2_in_13__ap_done ap_idle=A_IO_L2_in_13__ap_idle ap_ready=A_IO_L2_in_13__ap_ready
  // pragma RS ap-ctrl ap_start=A_IO_L2_in_14__ap_start ap_done=A_IO_L2_in_14__ap_done ap_idle=A_IO_L2_in_14__ap_idle ap_ready=A_IO_L2_in_14__ap_ready
  // pragma RS ap-ctrl ap_start=A_IO_L2_in_15__ap_start ap_done=A_IO_L2_in_15__ap_done ap_idle=A_IO_L2_in_15__ap_idle ap_ready=A_IO_L2_in_15__ap_ready
  // pragma RS ap-ctrl ap_start=A_IO_L2_in_16__ap_start ap_done=A_IO_L2_in_16__ap_done ap_idle=A_IO_L2_in_16__ap_idle ap_ready=A_IO_L2_in_16__ap_ready
  // pragma RS ap-ctrl ap_start=A_IO_L2_in_boundary_0__ap_start ap_done=A_IO_L2_in_boundary_0__ap_done ap_idle=A_IO_L2_in_boundary_0__ap_idle ap_ready=A_IO_L2_in_boundary_0__ap_ready
  // pragma RS ap-ctrl ap_start=A_IO_L3_in_0__ap_start ap_done=A_IO_L3_in_0__ap_done ap_idle=A_IO_L3_in_0__ap_idle ap_ready=A_IO_L3_in_0__ap_ready
  // pragma RS ap-ctrl ap_start=A_IO_L3_in_serialize_0__ap_start ap_done=A_IO_L3_in_serialize_0__ap_done ap_idle=A_IO_L3_in_serialize_0__ap_idle ap_ready=A_IO_L3_in_serialize_0__ap_ready scalar=A_IO_L3_in_serialize_0___.*
  // pragma RS ap-ctrl ap_start=A_PE_dummy_in_0__ap_start ap_done=A_PE_dummy_in_0__ap_done ap_idle=A_PE_dummy_in_0__ap_idle ap_ready=A_PE_dummy_in_0__ap_ready
  // pragma RS ap-ctrl ap_start=A_PE_dummy_in_1__ap_start ap_done=A_PE_dummy_in_1__ap_done ap_idle=A_PE_dummy_in_1__ap_idle ap_ready=A_PE_dummy_in_1__ap_ready
  // pragma RS ap-ctrl ap_start=A_PE_dummy_in_2__ap_start ap_done=A_PE_dummy_in_2__ap_done ap_idle=A_PE_dummy_in_2__ap_idle ap_ready=A_PE_dummy_in_2__ap_ready
  // pragma RS ap-ctrl ap_start=A_PE_dummy_in_3__ap_start ap_done=A_PE_dummy_in_3__ap_done ap_idle=A_PE_dummy_in_3__ap_idle ap_ready=A_PE_dummy_in_3__ap_ready
  // pragma RS ap-ctrl ap_start=A_PE_dummy_in_4__ap_start ap_done=A_PE_dummy_in_4__ap_done ap_idle=A_PE_dummy_in_4__ap_idle ap_ready=A_PE_dummy_in_4__ap_ready
  // pragma RS ap-ctrl ap_start=A_PE_dummy_in_5__ap_start ap_done=A_PE_dummy_in_5__ap_done ap_idle=A_PE_dummy_in_5__ap_idle ap_ready=A_PE_dummy_in_5__ap_ready
  // pragma RS ap-ctrl ap_start=A_PE_dummy_in_6__ap_start ap_done=A_PE_dummy_in_6__ap_done ap_idle=A_PE_dummy_in_6__ap_idle ap_ready=A_PE_dummy_in_6__ap_ready
  // pragma RS ap-ctrl ap_start=A_PE_dummy_in_7__ap_start ap_done=A_PE_dummy_in_7__ap_done ap_idle=A_PE_dummy_in_7__ap_idle ap_ready=A_PE_dummy_in_7__ap_ready
  // pragma RS ap-ctrl ap_start=A_PE_dummy_in_8__ap_start ap_done=A_PE_dummy_in_8__ap_done ap_idle=A_PE_dummy_in_8__ap_idle ap_ready=A_PE_dummy_in_8__ap_ready
  // pragma RS ap-ctrl ap_start=A_PE_dummy_in_9__ap_start ap_done=A_PE_dummy_in_9__ap_done ap_idle=A_PE_dummy_in_9__ap_idle ap_ready=A_PE_dummy_in_9__ap_ready
  // pragma RS ap-ctrl ap_start=A_PE_dummy_in_10__ap_start ap_done=A_PE_dummy_in_10__ap_done ap_idle=A_PE_dummy_in_10__ap_idle ap_ready=A_PE_dummy_in_10__ap_ready
  // pragma RS ap-ctrl ap_start=A_PE_dummy_in_11__ap_start ap_done=A_PE_dummy_in_11__ap_done ap_idle=A_PE_dummy_in_11__ap_idle ap_ready=A_PE_dummy_in_11__ap_ready
  // pragma RS ap-ctrl ap_start=A_PE_dummy_in_12__ap_start ap_done=A_PE_dummy_in_12__ap_done ap_idle=A_PE_dummy_in_12__ap_idle ap_ready=A_PE_dummy_in_12__ap_ready
  // pragma RS ap-ctrl ap_start=A_PE_dummy_in_13__ap_start ap_done=A_PE_dummy_in_13__ap_done ap_idle=A_PE_dummy_in_13__ap_idle ap_ready=A_PE_dummy_in_13__ap_ready
  // pragma RS ap-ctrl ap_start=A_PE_dummy_in_14__ap_start ap_done=A_PE_dummy_in_14__ap_done ap_idle=A_PE_dummy_in_14__ap_idle ap_ready=A_PE_dummy_in_14__ap_ready
  // pragma RS ap-ctrl ap_start=A_PE_dummy_in_15__ap_start ap_done=A_PE_dummy_in_15__ap_done ap_idle=A_PE_dummy_in_15__ap_idle ap_ready=A_PE_dummy_in_15__ap_ready
  // pragma RS ap-ctrl ap_start=A_PE_dummy_in_16__ap_start ap_done=A_PE_dummy_in_16__ap_done ap_idle=A_PE_dummy_in_16__ap_idle ap_ready=A_PE_dummy_in_16__ap_ready
  // pragma RS ap-ctrl ap_start=A_PE_dummy_in_17__ap_start ap_done=A_PE_dummy_in_17__ap_done ap_idle=A_PE_dummy_in_17__ap_idle ap_ready=A_PE_dummy_in_17__ap_ready
  // pragma RS ap-ctrl ap_start=B_IO_L2_in_0__ap_start ap_done=B_IO_L2_in_0__ap_done ap_idle=B_IO_L2_in_0__ap_idle ap_ready=B_IO_L2_in_0__ap_ready
  // pragma RS ap-ctrl ap_start=B_IO_L2_in_1__ap_start ap_done=B_IO_L2_in_1__ap_done ap_idle=B_IO_L2_in_1__ap_idle ap_ready=B_IO_L2_in_1__ap_ready
  // pragma RS ap-ctrl ap_start=B_IO_L2_in_2__ap_start ap_done=B_IO_L2_in_2__ap_done ap_idle=B_IO_L2_in_2__ap_idle ap_ready=B_IO_L2_in_2__ap_ready
  // pragma RS ap-ctrl ap_start=B_IO_L2_in_3__ap_start ap_done=B_IO_L2_in_3__ap_done ap_idle=B_IO_L2_in_3__ap_idle ap_ready=B_IO_L2_in_3__ap_ready
  // pragma RS ap-ctrl ap_start=B_IO_L2_in_4__ap_start ap_done=B_IO_L2_in_4__ap_done ap_idle=B_IO_L2_in_4__ap_idle ap_ready=B_IO_L2_in_4__ap_ready
  // pragma RS ap-ctrl ap_start=B_IO_L2_in_5__ap_start ap_done=B_IO_L2_in_5__ap_done ap_idle=B_IO_L2_in_5__ap_idle ap_ready=B_IO_L2_in_5__ap_ready
  // pragma RS ap-ctrl ap_start=B_IO_L2_in_6__ap_start ap_done=B_IO_L2_in_6__ap_done ap_idle=B_IO_L2_in_6__ap_idle ap_ready=B_IO_L2_in_6__ap_ready
  // pragma RS ap-ctrl ap_start=B_IO_L2_in_7__ap_start ap_done=B_IO_L2_in_7__ap_done ap_idle=B_IO_L2_in_7__ap_idle ap_ready=B_IO_L2_in_7__ap_ready
  // pragma RS ap-ctrl ap_start=B_IO_L2_in_8__ap_start ap_done=B_IO_L2_in_8__ap_done ap_idle=B_IO_L2_in_8__ap_idle ap_ready=B_IO_L2_in_8__ap_ready
  // pragma RS ap-ctrl ap_start=B_IO_L2_in_9__ap_start ap_done=B_IO_L2_in_9__ap_done ap_idle=B_IO_L2_in_9__ap_idle ap_ready=B_IO_L2_in_9__ap_ready
  // pragma RS ap-ctrl ap_start=B_IO_L2_in_10__ap_start ap_done=B_IO_L2_in_10__ap_done ap_idle=B_IO_L2_in_10__ap_idle ap_ready=B_IO_L2_in_10__ap_ready
  // pragma RS ap-ctrl ap_start=B_IO_L2_in_11__ap_start ap_done=B_IO_L2_in_11__ap_done ap_idle=B_IO_L2_in_11__ap_idle ap_ready=B_IO_L2_in_11__ap_ready
  // pragma RS ap-ctrl ap_start=B_IO_L2_in_12__ap_start ap_done=B_IO_L2_in_12__ap_done ap_idle=B_IO_L2_in_12__ap_idle ap_ready=B_IO_L2_in_12__ap_ready
  // pragma RS ap-ctrl ap_start=B_IO_L2_in_13__ap_start ap_done=B_IO_L2_in_13__ap_done ap_idle=B_IO_L2_in_13__ap_idle ap_ready=B_IO_L2_in_13__ap_ready
  // pragma RS ap-ctrl ap_start=B_IO_L2_in_14__ap_start ap_done=B_IO_L2_in_14__ap_done ap_idle=B_IO_L2_in_14__ap_idle ap_ready=B_IO_L2_in_14__ap_ready
  // pragma RS ap-ctrl ap_start=B_IO_L2_in_15__ap_start ap_done=B_IO_L2_in_15__ap_done ap_idle=B_IO_L2_in_15__ap_idle ap_ready=B_IO_L2_in_15__ap_ready
  // pragma RS ap-ctrl ap_start=B_IO_L2_in_boundary_0__ap_start ap_done=B_IO_L2_in_boundary_0__ap_done ap_idle=B_IO_L2_in_boundary_0__ap_idle ap_ready=B_IO_L2_in_boundary_0__ap_ready
  // pragma RS ap-ctrl ap_start=B_IO_L3_in_0__ap_start ap_done=B_IO_L3_in_0__ap_done ap_idle=B_IO_L3_in_0__ap_idle ap_ready=B_IO_L3_in_0__ap_ready
  // pragma RS ap-ctrl ap_start=B_IO_L3_in_serialize_0__ap_start ap_done=B_IO_L3_in_serialize_0__ap_done ap_idle=B_IO_L3_in_serialize_0__ap_idle ap_ready=B_IO_L3_in_serialize_0__ap_ready scalar=B_IO_L3_in_serialize_0___.*
  // pragma RS ap-ctrl ap_start=B_PE_dummy_in_0__ap_start ap_done=B_PE_dummy_in_0__ap_done ap_idle=B_PE_dummy_in_0__ap_idle ap_ready=B_PE_dummy_in_0__ap_ready
  // pragma RS ap-ctrl ap_start=B_PE_dummy_in_1__ap_start ap_done=B_PE_dummy_in_1__ap_done ap_idle=B_PE_dummy_in_1__ap_idle ap_ready=B_PE_dummy_in_1__ap_ready
  // pragma RS ap-ctrl ap_start=B_PE_dummy_in_2__ap_start ap_done=B_PE_dummy_in_2__ap_done ap_idle=B_PE_dummy_in_2__ap_idle ap_ready=B_PE_dummy_in_2__ap_ready
  // pragma RS ap-ctrl ap_start=B_PE_dummy_in_3__ap_start ap_done=B_PE_dummy_in_3__ap_done ap_idle=B_PE_dummy_in_3__ap_idle ap_ready=B_PE_dummy_in_3__ap_ready
  // pragma RS ap-ctrl ap_start=B_PE_dummy_in_4__ap_start ap_done=B_PE_dummy_in_4__ap_done ap_idle=B_PE_dummy_in_4__ap_idle ap_ready=B_PE_dummy_in_4__ap_ready
  // pragma RS ap-ctrl ap_start=B_PE_dummy_in_5__ap_start ap_done=B_PE_dummy_in_5__ap_done ap_idle=B_PE_dummy_in_5__ap_idle ap_ready=B_PE_dummy_in_5__ap_ready
  // pragma RS ap-ctrl ap_start=B_PE_dummy_in_6__ap_start ap_done=B_PE_dummy_in_6__ap_done ap_idle=B_PE_dummy_in_6__ap_idle ap_ready=B_PE_dummy_in_6__ap_ready
  // pragma RS ap-ctrl ap_start=B_PE_dummy_in_7__ap_start ap_done=B_PE_dummy_in_7__ap_done ap_idle=B_PE_dummy_in_7__ap_idle ap_ready=B_PE_dummy_in_7__ap_ready
  // pragma RS ap-ctrl ap_start=B_PE_dummy_in_8__ap_start ap_done=B_PE_dummy_in_8__ap_done ap_idle=B_PE_dummy_in_8__ap_idle ap_ready=B_PE_dummy_in_8__ap_ready
  // pragma RS ap-ctrl ap_start=B_PE_dummy_in_9__ap_start ap_done=B_PE_dummy_in_9__ap_done ap_idle=B_PE_dummy_in_9__ap_idle ap_ready=B_PE_dummy_in_9__ap_ready
  // pragma RS ap-ctrl ap_start=B_PE_dummy_in_10__ap_start ap_done=B_PE_dummy_in_10__ap_done ap_idle=B_PE_dummy_in_10__ap_idle ap_ready=B_PE_dummy_in_10__ap_ready
  // pragma RS ap-ctrl ap_start=B_PE_dummy_in_11__ap_start ap_done=B_PE_dummy_in_11__ap_done ap_idle=B_PE_dummy_in_11__ap_idle ap_ready=B_PE_dummy_in_11__ap_ready
  // pragma RS ap-ctrl ap_start=B_PE_dummy_in_12__ap_start ap_done=B_PE_dummy_in_12__ap_done ap_idle=B_PE_dummy_in_12__ap_idle ap_ready=B_PE_dummy_in_12__ap_ready
  // pragma RS ap-ctrl ap_start=B_PE_dummy_in_13__ap_start ap_done=B_PE_dummy_in_13__ap_done ap_idle=B_PE_dummy_in_13__ap_idle ap_ready=B_PE_dummy_in_13__ap_ready
  // pragma RS ap-ctrl ap_start=B_PE_dummy_in_14__ap_start ap_done=B_PE_dummy_in_14__ap_done ap_idle=B_PE_dummy_in_14__ap_idle ap_ready=B_PE_dummy_in_14__ap_ready
  // pragma RS ap-ctrl ap_start=B_PE_dummy_in_15__ap_start ap_done=B_PE_dummy_in_15__ap_done ap_idle=B_PE_dummy_in_15__ap_idle ap_ready=B_PE_dummy_in_15__ap_ready
  // pragma RS ap-ctrl ap_start=B_PE_dummy_in_16__ap_start ap_done=B_PE_dummy_in_16__ap_done ap_idle=B_PE_dummy_in_16__ap_idle ap_ready=B_PE_dummy_in_16__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_boundary_wrapper_0__ap_start ap_done=C_drain_IO_L1_out_boundary_wrapper_0__ap_done ap_idle=C_drain_IO_L1_out_boundary_wrapper_0__ap_idle ap_ready=C_drain_IO_L1_out_boundary_wrapper_0__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_boundary_wrapper_1__ap_start ap_done=C_drain_IO_L1_out_boundary_wrapper_1__ap_done ap_idle=C_drain_IO_L1_out_boundary_wrapper_1__ap_idle ap_ready=C_drain_IO_L1_out_boundary_wrapper_1__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_boundary_wrapper_2__ap_start ap_done=C_drain_IO_L1_out_boundary_wrapper_2__ap_done ap_idle=C_drain_IO_L1_out_boundary_wrapper_2__ap_idle ap_ready=C_drain_IO_L1_out_boundary_wrapper_2__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_boundary_wrapper_3__ap_start ap_done=C_drain_IO_L1_out_boundary_wrapper_3__ap_done ap_idle=C_drain_IO_L1_out_boundary_wrapper_3__ap_idle ap_ready=C_drain_IO_L1_out_boundary_wrapper_3__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_boundary_wrapper_4__ap_start ap_done=C_drain_IO_L1_out_boundary_wrapper_4__ap_done ap_idle=C_drain_IO_L1_out_boundary_wrapper_4__ap_idle ap_ready=C_drain_IO_L1_out_boundary_wrapper_4__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_boundary_wrapper_5__ap_start ap_done=C_drain_IO_L1_out_boundary_wrapper_5__ap_done ap_idle=C_drain_IO_L1_out_boundary_wrapper_5__ap_idle ap_ready=C_drain_IO_L1_out_boundary_wrapper_5__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_boundary_wrapper_6__ap_start ap_done=C_drain_IO_L1_out_boundary_wrapper_6__ap_done ap_idle=C_drain_IO_L1_out_boundary_wrapper_6__ap_idle ap_ready=C_drain_IO_L1_out_boundary_wrapper_6__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_boundary_wrapper_7__ap_start ap_done=C_drain_IO_L1_out_boundary_wrapper_7__ap_done ap_idle=C_drain_IO_L1_out_boundary_wrapper_7__ap_idle ap_ready=C_drain_IO_L1_out_boundary_wrapper_7__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_boundary_wrapper_8__ap_start ap_done=C_drain_IO_L1_out_boundary_wrapper_8__ap_done ap_idle=C_drain_IO_L1_out_boundary_wrapper_8__ap_idle ap_ready=C_drain_IO_L1_out_boundary_wrapper_8__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_boundary_wrapper_9__ap_start ap_done=C_drain_IO_L1_out_boundary_wrapper_9__ap_done ap_idle=C_drain_IO_L1_out_boundary_wrapper_9__ap_idle ap_ready=C_drain_IO_L1_out_boundary_wrapper_9__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_boundary_wrapper_10__ap_start ap_done=C_drain_IO_L1_out_boundary_wrapper_10__ap_done ap_idle=C_drain_IO_L1_out_boundary_wrapper_10__ap_idle ap_ready=C_drain_IO_L1_out_boundary_wrapper_10__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_boundary_wrapper_11__ap_start ap_done=C_drain_IO_L1_out_boundary_wrapper_11__ap_done ap_idle=C_drain_IO_L1_out_boundary_wrapper_11__ap_idle ap_ready=C_drain_IO_L1_out_boundary_wrapper_11__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_boundary_wrapper_12__ap_start ap_done=C_drain_IO_L1_out_boundary_wrapper_12__ap_done ap_idle=C_drain_IO_L1_out_boundary_wrapper_12__ap_idle ap_ready=C_drain_IO_L1_out_boundary_wrapper_12__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_boundary_wrapper_13__ap_start ap_done=C_drain_IO_L1_out_boundary_wrapper_13__ap_done ap_idle=C_drain_IO_L1_out_boundary_wrapper_13__ap_idle ap_ready=C_drain_IO_L1_out_boundary_wrapper_13__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_boundary_wrapper_14__ap_start ap_done=C_drain_IO_L1_out_boundary_wrapper_14__ap_done ap_idle=C_drain_IO_L1_out_boundary_wrapper_14__ap_idle ap_ready=C_drain_IO_L1_out_boundary_wrapper_14__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_boundary_wrapper_15__ap_start ap_done=C_drain_IO_L1_out_boundary_wrapper_15__ap_done ap_idle=C_drain_IO_L1_out_boundary_wrapper_15__ap_idle ap_ready=C_drain_IO_L1_out_boundary_wrapper_15__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_boundary_wrapper_16__ap_start ap_done=C_drain_IO_L1_out_boundary_wrapper_16__ap_done ap_idle=C_drain_IO_L1_out_boundary_wrapper_16__ap_idle ap_ready=C_drain_IO_L1_out_boundary_wrapper_16__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_0__ap_start ap_done=C_drain_IO_L1_out_wrapper_0__ap_done ap_idle=C_drain_IO_L1_out_wrapper_0__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_0__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_1__ap_start ap_done=C_drain_IO_L1_out_wrapper_1__ap_done ap_idle=C_drain_IO_L1_out_wrapper_1__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_1__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_2__ap_start ap_done=C_drain_IO_L1_out_wrapper_2__ap_done ap_idle=C_drain_IO_L1_out_wrapper_2__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_2__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_3__ap_start ap_done=C_drain_IO_L1_out_wrapper_3__ap_done ap_idle=C_drain_IO_L1_out_wrapper_3__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_3__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_4__ap_start ap_done=C_drain_IO_L1_out_wrapper_4__ap_done ap_idle=C_drain_IO_L1_out_wrapper_4__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_4__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_5__ap_start ap_done=C_drain_IO_L1_out_wrapper_5__ap_done ap_idle=C_drain_IO_L1_out_wrapper_5__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_5__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_6__ap_start ap_done=C_drain_IO_L1_out_wrapper_6__ap_done ap_idle=C_drain_IO_L1_out_wrapper_6__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_6__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_7__ap_start ap_done=C_drain_IO_L1_out_wrapper_7__ap_done ap_idle=C_drain_IO_L1_out_wrapper_7__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_7__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_8__ap_start ap_done=C_drain_IO_L1_out_wrapper_8__ap_done ap_idle=C_drain_IO_L1_out_wrapper_8__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_8__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_9__ap_start ap_done=C_drain_IO_L1_out_wrapper_9__ap_done ap_idle=C_drain_IO_L1_out_wrapper_9__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_9__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_10__ap_start ap_done=C_drain_IO_L1_out_wrapper_10__ap_done ap_idle=C_drain_IO_L1_out_wrapper_10__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_10__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_11__ap_start ap_done=C_drain_IO_L1_out_wrapper_11__ap_done ap_idle=C_drain_IO_L1_out_wrapper_11__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_11__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_12__ap_start ap_done=C_drain_IO_L1_out_wrapper_12__ap_done ap_idle=C_drain_IO_L1_out_wrapper_12__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_12__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_13__ap_start ap_done=C_drain_IO_L1_out_wrapper_13__ap_done ap_idle=C_drain_IO_L1_out_wrapper_13__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_13__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_14__ap_start ap_done=C_drain_IO_L1_out_wrapper_14__ap_done ap_idle=C_drain_IO_L1_out_wrapper_14__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_14__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_15__ap_start ap_done=C_drain_IO_L1_out_wrapper_15__ap_done ap_idle=C_drain_IO_L1_out_wrapper_15__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_15__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_16__ap_start ap_done=C_drain_IO_L1_out_wrapper_16__ap_done ap_idle=C_drain_IO_L1_out_wrapper_16__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_16__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_17__ap_start ap_done=C_drain_IO_L1_out_wrapper_17__ap_done ap_idle=C_drain_IO_L1_out_wrapper_17__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_17__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_18__ap_start ap_done=C_drain_IO_L1_out_wrapper_18__ap_done ap_idle=C_drain_IO_L1_out_wrapper_18__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_18__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_19__ap_start ap_done=C_drain_IO_L1_out_wrapper_19__ap_done ap_idle=C_drain_IO_L1_out_wrapper_19__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_19__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_20__ap_start ap_done=C_drain_IO_L1_out_wrapper_20__ap_done ap_idle=C_drain_IO_L1_out_wrapper_20__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_20__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_21__ap_start ap_done=C_drain_IO_L1_out_wrapper_21__ap_done ap_idle=C_drain_IO_L1_out_wrapper_21__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_21__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_22__ap_start ap_done=C_drain_IO_L1_out_wrapper_22__ap_done ap_idle=C_drain_IO_L1_out_wrapper_22__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_22__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_23__ap_start ap_done=C_drain_IO_L1_out_wrapper_23__ap_done ap_idle=C_drain_IO_L1_out_wrapper_23__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_23__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_24__ap_start ap_done=C_drain_IO_L1_out_wrapper_24__ap_done ap_idle=C_drain_IO_L1_out_wrapper_24__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_24__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_25__ap_start ap_done=C_drain_IO_L1_out_wrapper_25__ap_done ap_idle=C_drain_IO_L1_out_wrapper_25__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_25__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_26__ap_start ap_done=C_drain_IO_L1_out_wrapper_26__ap_done ap_idle=C_drain_IO_L1_out_wrapper_26__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_26__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_27__ap_start ap_done=C_drain_IO_L1_out_wrapper_27__ap_done ap_idle=C_drain_IO_L1_out_wrapper_27__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_27__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_28__ap_start ap_done=C_drain_IO_L1_out_wrapper_28__ap_done ap_idle=C_drain_IO_L1_out_wrapper_28__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_28__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_29__ap_start ap_done=C_drain_IO_L1_out_wrapper_29__ap_done ap_idle=C_drain_IO_L1_out_wrapper_29__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_29__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_30__ap_start ap_done=C_drain_IO_L1_out_wrapper_30__ap_done ap_idle=C_drain_IO_L1_out_wrapper_30__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_30__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_31__ap_start ap_done=C_drain_IO_L1_out_wrapper_31__ap_done ap_idle=C_drain_IO_L1_out_wrapper_31__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_31__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_32__ap_start ap_done=C_drain_IO_L1_out_wrapper_32__ap_done ap_idle=C_drain_IO_L1_out_wrapper_32__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_32__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_33__ap_start ap_done=C_drain_IO_L1_out_wrapper_33__ap_done ap_idle=C_drain_IO_L1_out_wrapper_33__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_33__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_34__ap_start ap_done=C_drain_IO_L1_out_wrapper_34__ap_done ap_idle=C_drain_IO_L1_out_wrapper_34__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_34__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_35__ap_start ap_done=C_drain_IO_L1_out_wrapper_35__ap_done ap_idle=C_drain_IO_L1_out_wrapper_35__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_35__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_36__ap_start ap_done=C_drain_IO_L1_out_wrapper_36__ap_done ap_idle=C_drain_IO_L1_out_wrapper_36__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_36__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_37__ap_start ap_done=C_drain_IO_L1_out_wrapper_37__ap_done ap_idle=C_drain_IO_L1_out_wrapper_37__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_37__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_38__ap_start ap_done=C_drain_IO_L1_out_wrapper_38__ap_done ap_idle=C_drain_IO_L1_out_wrapper_38__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_38__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_39__ap_start ap_done=C_drain_IO_L1_out_wrapper_39__ap_done ap_idle=C_drain_IO_L1_out_wrapper_39__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_39__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_40__ap_start ap_done=C_drain_IO_L1_out_wrapper_40__ap_done ap_idle=C_drain_IO_L1_out_wrapper_40__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_40__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_41__ap_start ap_done=C_drain_IO_L1_out_wrapper_41__ap_done ap_idle=C_drain_IO_L1_out_wrapper_41__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_41__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_42__ap_start ap_done=C_drain_IO_L1_out_wrapper_42__ap_done ap_idle=C_drain_IO_L1_out_wrapper_42__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_42__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_43__ap_start ap_done=C_drain_IO_L1_out_wrapper_43__ap_done ap_idle=C_drain_IO_L1_out_wrapper_43__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_43__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_44__ap_start ap_done=C_drain_IO_L1_out_wrapper_44__ap_done ap_idle=C_drain_IO_L1_out_wrapper_44__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_44__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_45__ap_start ap_done=C_drain_IO_L1_out_wrapper_45__ap_done ap_idle=C_drain_IO_L1_out_wrapper_45__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_45__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_46__ap_start ap_done=C_drain_IO_L1_out_wrapper_46__ap_done ap_idle=C_drain_IO_L1_out_wrapper_46__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_46__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_47__ap_start ap_done=C_drain_IO_L1_out_wrapper_47__ap_done ap_idle=C_drain_IO_L1_out_wrapper_47__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_47__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_48__ap_start ap_done=C_drain_IO_L1_out_wrapper_48__ap_done ap_idle=C_drain_IO_L1_out_wrapper_48__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_48__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_49__ap_start ap_done=C_drain_IO_L1_out_wrapper_49__ap_done ap_idle=C_drain_IO_L1_out_wrapper_49__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_49__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_50__ap_start ap_done=C_drain_IO_L1_out_wrapper_50__ap_done ap_idle=C_drain_IO_L1_out_wrapper_50__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_50__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_51__ap_start ap_done=C_drain_IO_L1_out_wrapper_51__ap_done ap_idle=C_drain_IO_L1_out_wrapper_51__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_51__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_52__ap_start ap_done=C_drain_IO_L1_out_wrapper_52__ap_done ap_idle=C_drain_IO_L1_out_wrapper_52__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_52__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_53__ap_start ap_done=C_drain_IO_L1_out_wrapper_53__ap_done ap_idle=C_drain_IO_L1_out_wrapper_53__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_53__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_54__ap_start ap_done=C_drain_IO_L1_out_wrapper_54__ap_done ap_idle=C_drain_IO_L1_out_wrapper_54__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_54__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_55__ap_start ap_done=C_drain_IO_L1_out_wrapper_55__ap_done ap_idle=C_drain_IO_L1_out_wrapper_55__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_55__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_56__ap_start ap_done=C_drain_IO_L1_out_wrapper_56__ap_done ap_idle=C_drain_IO_L1_out_wrapper_56__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_56__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_57__ap_start ap_done=C_drain_IO_L1_out_wrapper_57__ap_done ap_idle=C_drain_IO_L1_out_wrapper_57__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_57__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_58__ap_start ap_done=C_drain_IO_L1_out_wrapper_58__ap_done ap_idle=C_drain_IO_L1_out_wrapper_58__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_58__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_59__ap_start ap_done=C_drain_IO_L1_out_wrapper_59__ap_done ap_idle=C_drain_IO_L1_out_wrapper_59__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_59__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_60__ap_start ap_done=C_drain_IO_L1_out_wrapper_60__ap_done ap_idle=C_drain_IO_L1_out_wrapper_60__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_60__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_61__ap_start ap_done=C_drain_IO_L1_out_wrapper_61__ap_done ap_idle=C_drain_IO_L1_out_wrapper_61__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_61__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_62__ap_start ap_done=C_drain_IO_L1_out_wrapper_62__ap_done ap_idle=C_drain_IO_L1_out_wrapper_62__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_62__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_63__ap_start ap_done=C_drain_IO_L1_out_wrapper_63__ap_done ap_idle=C_drain_IO_L1_out_wrapper_63__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_63__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_64__ap_start ap_done=C_drain_IO_L1_out_wrapper_64__ap_done ap_idle=C_drain_IO_L1_out_wrapper_64__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_64__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_65__ap_start ap_done=C_drain_IO_L1_out_wrapper_65__ap_done ap_idle=C_drain_IO_L1_out_wrapper_65__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_65__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_66__ap_start ap_done=C_drain_IO_L1_out_wrapper_66__ap_done ap_idle=C_drain_IO_L1_out_wrapper_66__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_66__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_67__ap_start ap_done=C_drain_IO_L1_out_wrapper_67__ap_done ap_idle=C_drain_IO_L1_out_wrapper_67__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_67__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_68__ap_start ap_done=C_drain_IO_L1_out_wrapper_68__ap_done ap_idle=C_drain_IO_L1_out_wrapper_68__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_68__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_69__ap_start ap_done=C_drain_IO_L1_out_wrapper_69__ap_done ap_idle=C_drain_IO_L1_out_wrapper_69__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_69__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_70__ap_start ap_done=C_drain_IO_L1_out_wrapper_70__ap_done ap_idle=C_drain_IO_L1_out_wrapper_70__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_70__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_71__ap_start ap_done=C_drain_IO_L1_out_wrapper_71__ap_done ap_idle=C_drain_IO_L1_out_wrapper_71__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_71__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_72__ap_start ap_done=C_drain_IO_L1_out_wrapper_72__ap_done ap_idle=C_drain_IO_L1_out_wrapper_72__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_72__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_73__ap_start ap_done=C_drain_IO_L1_out_wrapper_73__ap_done ap_idle=C_drain_IO_L1_out_wrapper_73__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_73__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_74__ap_start ap_done=C_drain_IO_L1_out_wrapper_74__ap_done ap_idle=C_drain_IO_L1_out_wrapper_74__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_74__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_75__ap_start ap_done=C_drain_IO_L1_out_wrapper_75__ap_done ap_idle=C_drain_IO_L1_out_wrapper_75__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_75__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_76__ap_start ap_done=C_drain_IO_L1_out_wrapper_76__ap_done ap_idle=C_drain_IO_L1_out_wrapper_76__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_76__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_77__ap_start ap_done=C_drain_IO_L1_out_wrapper_77__ap_done ap_idle=C_drain_IO_L1_out_wrapper_77__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_77__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_78__ap_start ap_done=C_drain_IO_L1_out_wrapper_78__ap_done ap_idle=C_drain_IO_L1_out_wrapper_78__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_78__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_79__ap_start ap_done=C_drain_IO_L1_out_wrapper_79__ap_done ap_idle=C_drain_IO_L1_out_wrapper_79__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_79__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_80__ap_start ap_done=C_drain_IO_L1_out_wrapper_80__ap_done ap_idle=C_drain_IO_L1_out_wrapper_80__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_80__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_81__ap_start ap_done=C_drain_IO_L1_out_wrapper_81__ap_done ap_idle=C_drain_IO_L1_out_wrapper_81__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_81__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_82__ap_start ap_done=C_drain_IO_L1_out_wrapper_82__ap_done ap_idle=C_drain_IO_L1_out_wrapper_82__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_82__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_83__ap_start ap_done=C_drain_IO_L1_out_wrapper_83__ap_done ap_idle=C_drain_IO_L1_out_wrapper_83__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_83__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_84__ap_start ap_done=C_drain_IO_L1_out_wrapper_84__ap_done ap_idle=C_drain_IO_L1_out_wrapper_84__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_84__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_85__ap_start ap_done=C_drain_IO_L1_out_wrapper_85__ap_done ap_idle=C_drain_IO_L1_out_wrapper_85__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_85__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_86__ap_start ap_done=C_drain_IO_L1_out_wrapper_86__ap_done ap_idle=C_drain_IO_L1_out_wrapper_86__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_86__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_87__ap_start ap_done=C_drain_IO_L1_out_wrapper_87__ap_done ap_idle=C_drain_IO_L1_out_wrapper_87__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_87__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_88__ap_start ap_done=C_drain_IO_L1_out_wrapper_88__ap_done ap_idle=C_drain_IO_L1_out_wrapper_88__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_88__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_89__ap_start ap_done=C_drain_IO_L1_out_wrapper_89__ap_done ap_idle=C_drain_IO_L1_out_wrapper_89__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_89__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_90__ap_start ap_done=C_drain_IO_L1_out_wrapper_90__ap_done ap_idle=C_drain_IO_L1_out_wrapper_90__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_90__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_91__ap_start ap_done=C_drain_IO_L1_out_wrapper_91__ap_done ap_idle=C_drain_IO_L1_out_wrapper_91__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_91__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_92__ap_start ap_done=C_drain_IO_L1_out_wrapper_92__ap_done ap_idle=C_drain_IO_L1_out_wrapper_92__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_92__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_93__ap_start ap_done=C_drain_IO_L1_out_wrapper_93__ap_done ap_idle=C_drain_IO_L1_out_wrapper_93__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_93__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_94__ap_start ap_done=C_drain_IO_L1_out_wrapper_94__ap_done ap_idle=C_drain_IO_L1_out_wrapper_94__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_94__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_95__ap_start ap_done=C_drain_IO_L1_out_wrapper_95__ap_done ap_idle=C_drain_IO_L1_out_wrapper_95__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_95__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_96__ap_start ap_done=C_drain_IO_L1_out_wrapper_96__ap_done ap_idle=C_drain_IO_L1_out_wrapper_96__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_96__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_97__ap_start ap_done=C_drain_IO_L1_out_wrapper_97__ap_done ap_idle=C_drain_IO_L1_out_wrapper_97__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_97__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_98__ap_start ap_done=C_drain_IO_L1_out_wrapper_98__ap_done ap_idle=C_drain_IO_L1_out_wrapper_98__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_98__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_99__ap_start ap_done=C_drain_IO_L1_out_wrapper_99__ap_done ap_idle=C_drain_IO_L1_out_wrapper_99__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_99__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_100__ap_start ap_done=C_drain_IO_L1_out_wrapper_100__ap_done ap_idle=C_drain_IO_L1_out_wrapper_100__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_100__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_101__ap_start ap_done=C_drain_IO_L1_out_wrapper_101__ap_done ap_idle=C_drain_IO_L1_out_wrapper_101__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_101__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_102__ap_start ap_done=C_drain_IO_L1_out_wrapper_102__ap_done ap_idle=C_drain_IO_L1_out_wrapper_102__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_102__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_103__ap_start ap_done=C_drain_IO_L1_out_wrapper_103__ap_done ap_idle=C_drain_IO_L1_out_wrapper_103__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_103__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_104__ap_start ap_done=C_drain_IO_L1_out_wrapper_104__ap_done ap_idle=C_drain_IO_L1_out_wrapper_104__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_104__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_105__ap_start ap_done=C_drain_IO_L1_out_wrapper_105__ap_done ap_idle=C_drain_IO_L1_out_wrapper_105__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_105__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_106__ap_start ap_done=C_drain_IO_L1_out_wrapper_106__ap_done ap_idle=C_drain_IO_L1_out_wrapper_106__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_106__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_107__ap_start ap_done=C_drain_IO_L1_out_wrapper_107__ap_done ap_idle=C_drain_IO_L1_out_wrapper_107__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_107__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_108__ap_start ap_done=C_drain_IO_L1_out_wrapper_108__ap_done ap_idle=C_drain_IO_L1_out_wrapper_108__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_108__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_109__ap_start ap_done=C_drain_IO_L1_out_wrapper_109__ap_done ap_idle=C_drain_IO_L1_out_wrapper_109__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_109__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_110__ap_start ap_done=C_drain_IO_L1_out_wrapper_110__ap_done ap_idle=C_drain_IO_L1_out_wrapper_110__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_110__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_111__ap_start ap_done=C_drain_IO_L1_out_wrapper_111__ap_done ap_idle=C_drain_IO_L1_out_wrapper_111__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_111__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_112__ap_start ap_done=C_drain_IO_L1_out_wrapper_112__ap_done ap_idle=C_drain_IO_L1_out_wrapper_112__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_112__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_113__ap_start ap_done=C_drain_IO_L1_out_wrapper_113__ap_done ap_idle=C_drain_IO_L1_out_wrapper_113__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_113__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_114__ap_start ap_done=C_drain_IO_L1_out_wrapper_114__ap_done ap_idle=C_drain_IO_L1_out_wrapper_114__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_114__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_115__ap_start ap_done=C_drain_IO_L1_out_wrapper_115__ap_done ap_idle=C_drain_IO_L1_out_wrapper_115__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_115__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_116__ap_start ap_done=C_drain_IO_L1_out_wrapper_116__ap_done ap_idle=C_drain_IO_L1_out_wrapper_116__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_116__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_117__ap_start ap_done=C_drain_IO_L1_out_wrapper_117__ap_done ap_idle=C_drain_IO_L1_out_wrapper_117__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_117__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_118__ap_start ap_done=C_drain_IO_L1_out_wrapper_118__ap_done ap_idle=C_drain_IO_L1_out_wrapper_118__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_118__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_119__ap_start ap_done=C_drain_IO_L1_out_wrapper_119__ap_done ap_idle=C_drain_IO_L1_out_wrapper_119__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_119__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_120__ap_start ap_done=C_drain_IO_L1_out_wrapper_120__ap_done ap_idle=C_drain_IO_L1_out_wrapper_120__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_120__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_121__ap_start ap_done=C_drain_IO_L1_out_wrapper_121__ap_done ap_idle=C_drain_IO_L1_out_wrapper_121__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_121__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_122__ap_start ap_done=C_drain_IO_L1_out_wrapper_122__ap_done ap_idle=C_drain_IO_L1_out_wrapper_122__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_122__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_123__ap_start ap_done=C_drain_IO_L1_out_wrapper_123__ap_done ap_idle=C_drain_IO_L1_out_wrapper_123__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_123__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_124__ap_start ap_done=C_drain_IO_L1_out_wrapper_124__ap_done ap_idle=C_drain_IO_L1_out_wrapper_124__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_124__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_125__ap_start ap_done=C_drain_IO_L1_out_wrapper_125__ap_done ap_idle=C_drain_IO_L1_out_wrapper_125__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_125__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_126__ap_start ap_done=C_drain_IO_L1_out_wrapper_126__ap_done ap_idle=C_drain_IO_L1_out_wrapper_126__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_126__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_127__ap_start ap_done=C_drain_IO_L1_out_wrapper_127__ap_done ap_idle=C_drain_IO_L1_out_wrapper_127__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_127__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_128__ap_start ap_done=C_drain_IO_L1_out_wrapper_128__ap_done ap_idle=C_drain_IO_L1_out_wrapper_128__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_128__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_129__ap_start ap_done=C_drain_IO_L1_out_wrapper_129__ap_done ap_idle=C_drain_IO_L1_out_wrapper_129__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_129__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_130__ap_start ap_done=C_drain_IO_L1_out_wrapper_130__ap_done ap_idle=C_drain_IO_L1_out_wrapper_130__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_130__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_131__ap_start ap_done=C_drain_IO_L1_out_wrapper_131__ap_done ap_idle=C_drain_IO_L1_out_wrapper_131__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_131__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_132__ap_start ap_done=C_drain_IO_L1_out_wrapper_132__ap_done ap_idle=C_drain_IO_L1_out_wrapper_132__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_132__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_133__ap_start ap_done=C_drain_IO_L1_out_wrapper_133__ap_done ap_idle=C_drain_IO_L1_out_wrapper_133__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_133__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_134__ap_start ap_done=C_drain_IO_L1_out_wrapper_134__ap_done ap_idle=C_drain_IO_L1_out_wrapper_134__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_134__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_135__ap_start ap_done=C_drain_IO_L1_out_wrapper_135__ap_done ap_idle=C_drain_IO_L1_out_wrapper_135__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_135__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_136__ap_start ap_done=C_drain_IO_L1_out_wrapper_136__ap_done ap_idle=C_drain_IO_L1_out_wrapper_136__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_136__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_137__ap_start ap_done=C_drain_IO_L1_out_wrapper_137__ap_done ap_idle=C_drain_IO_L1_out_wrapper_137__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_137__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_138__ap_start ap_done=C_drain_IO_L1_out_wrapper_138__ap_done ap_idle=C_drain_IO_L1_out_wrapper_138__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_138__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_139__ap_start ap_done=C_drain_IO_L1_out_wrapper_139__ap_done ap_idle=C_drain_IO_L1_out_wrapper_139__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_139__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_140__ap_start ap_done=C_drain_IO_L1_out_wrapper_140__ap_done ap_idle=C_drain_IO_L1_out_wrapper_140__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_140__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_141__ap_start ap_done=C_drain_IO_L1_out_wrapper_141__ap_done ap_idle=C_drain_IO_L1_out_wrapper_141__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_141__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_142__ap_start ap_done=C_drain_IO_L1_out_wrapper_142__ap_done ap_idle=C_drain_IO_L1_out_wrapper_142__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_142__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_143__ap_start ap_done=C_drain_IO_L1_out_wrapper_143__ap_done ap_idle=C_drain_IO_L1_out_wrapper_143__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_143__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_144__ap_start ap_done=C_drain_IO_L1_out_wrapper_144__ap_done ap_idle=C_drain_IO_L1_out_wrapper_144__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_144__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_145__ap_start ap_done=C_drain_IO_L1_out_wrapper_145__ap_done ap_idle=C_drain_IO_L1_out_wrapper_145__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_145__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_146__ap_start ap_done=C_drain_IO_L1_out_wrapper_146__ap_done ap_idle=C_drain_IO_L1_out_wrapper_146__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_146__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_147__ap_start ap_done=C_drain_IO_L1_out_wrapper_147__ap_done ap_idle=C_drain_IO_L1_out_wrapper_147__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_147__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_148__ap_start ap_done=C_drain_IO_L1_out_wrapper_148__ap_done ap_idle=C_drain_IO_L1_out_wrapper_148__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_148__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_149__ap_start ap_done=C_drain_IO_L1_out_wrapper_149__ap_done ap_idle=C_drain_IO_L1_out_wrapper_149__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_149__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_150__ap_start ap_done=C_drain_IO_L1_out_wrapper_150__ap_done ap_idle=C_drain_IO_L1_out_wrapper_150__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_150__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_151__ap_start ap_done=C_drain_IO_L1_out_wrapper_151__ap_done ap_idle=C_drain_IO_L1_out_wrapper_151__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_151__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_152__ap_start ap_done=C_drain_IO_L1_out_wrapper_152__ap_done ap_idle=C_drain_IO_L1_out_wrapper_152__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_152__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_153__ap_start ap_done=C_drain_IO_L1_out_wrapper_153__ap_done ap_idle=C_drain_IO_L1_out_wrapper_153__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_153__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_154__ap_start ap_done=C_drain_IO_L1_out_wrapper_154__ap_done ap_idle=C_drain_IO_L1_out_wrapper_154__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_154__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_155__ap_start ap_done=C_drain_IO_L1_out_wrapper_155__ap_done ap_idle=C_drain_IO_L1_out_wrapper_155__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_155__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_156__ap_start ap_done=C_drain_IO_L1_out_wrapper_156__ap_done ap_idle=C_drain_IO_L1_out_wrapper_156__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_156__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_157__ap_start ap_done=C_drain_IO_L1_out_wrapper_157__ap_done ap_idle=C_drain_IO_L1_out_wrapper_157__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_157__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_158__ap_start ap_done=C_drain_IO_L1_out_wrapper_158__ap_done ap_idle=C_drain_IO_L1_out_wrapper_158__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_158__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_159__ap_start ap_done=C_drain_IO_L1_out_wrapper_159__ap_done ap_idle=C_drain_IO_L1_out_wrapper_159__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_159__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_160__ap_start ap_done=C_drain_IO_L1_out_wrapper_160__ap_done ap_idle=C_drain_IO_L1_out_wrapper_160__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_160__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_161__ap_start ap_done=C_drain_IO_L1_out_wrapper_161__ap_done ap_idle=C_drain_IO_L1_out_wrapper_161__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_161__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_162__ap_start ap_done=C_drain_IO_L1_out_wrapper_162__ap_done ap_idle=C_drain_IO_L1_out_wrapper_162__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_162__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_163__ap_start ap_done=C_drain_IO_L1_out_wrapper_163__ap_done ap_idle=C_drain_IO_L1_out_wrapper_163__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_163__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_164__ap_start ap_done=C_drain_IO_L1_out_wrapper_164__ap_done ap_idle=C_drain_IO_L1_out_wrapper_164__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_164__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_165__ap_start ap_done=C_drain_IO_L1_out_wrapper_165__ap_done ap_idle=C_drain_IO_L1_out_wrapper_165__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_165__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_166__ap_start ap_done=C_drain_IO_L1_out_wrapper_166__ap_done ap_idle=C_drain_IO_L1_out_wrapper_166__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_166__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_167__ap_start ap_done=C_drain_IO_L1_out_wrapper_167__ap_done ap_idle=C_drain_IO_L1_out_wrapper_167__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_167__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_168__ap_start ap_done=C_drain_IO_L1_out_wrapper_168__ap_done ap_idle=C_drain_IO_L1_out_wrapper_168__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_168__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_169__ap_start ap_done=C_drain_IO_L1_out_wrapper_169__ap_done ap_idle=C_drain_IO_L1_out_wrapper_169__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_169__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_170__ap_start ap_done=C_drain_IO_L1_out_wrapper_170__ap_done ap_idle=C_drain_IO_L1_out_wrapper_170__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_170__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_171__ap_start ap_done=C_drain_IO_L1_out_wrapper_171__ap_done ap_idle=C_drain_IO_L1_out_wrapper_171__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_171__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_172__ap_start ap_done=C_drain_IO_L1_out_wrapper_172__ap_done ap_idle=C_drain_IO_L1_out_wrapper_172__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_172__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_173__ap_start ap_done=C_drain_IO_L1_out_wrapper_173__ap_done ap_idle=C_drain_IO_L1_out_wrapper_173__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_173__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_174__ap_start ap_done=C_drain_IO_L1_out_wrapper_174__ap_done ap_idle=C_drain_IO_L1_out_wrapper_174__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_174__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_175__ap_start ap_done=C_drain_IO_L1_out_wrapper_175__ap_done ap_idle=C_drain_IO_L1_out_wrapper_175__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_175__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_176__ap_start ap_done=C_drain_IO_L1_out_wrapper_176__ap_done ap_idle=C_drain_IO_L1_out_wrapper_176__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_176__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_177__ap_start ap_done=C_drain_IO_L1_out_wrapper_177__ap_done ap_idle=C_drain_IO_L1_out_wrapper_177__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_177__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_178__ap_start ap_done=C_drain_IO_L1_out_wrapper_178__ap_done ap_idle=C_drain_IO_L1_out_wrapper_178__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_178__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_179__ap_start ap_done=C_drain_IO_L1_out_wrapper_179__ap_done ap_idle=C_drain_IO_L1_out_wrapper_179__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_179__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_180__ap_start ap_done=C_drain_IO_L1_out_wrapper_180__ap_done ap_idle=C_drain_IO_L1_out_wrapper_180__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_180__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_181__ap_start ap_done=C_drain_IO_L1_out_wrapper_181__ap_done ap_idle=C_drain_IO_L1_out_wrapper_181__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_181__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_182__ap_start ap_done=C_drain_IO_L1_out_wrapper_182__ap_done ap_idle=C_drain_IO_L1_out_wrapper_182__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_182__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_183__ap_start ap_done=C_drain_IO_L1_out_wrapper_183__ap_done ap_idle=C_drain_IO_L1_out_wrapper_183__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_183__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_184__ap_start ap_done=C_drain_IO_L1_out_wrapper_184__ap_done ap_idle=C_drain_IO_L1_out_wrapper_184__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_184__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_185__ap_start ap_done=C_drain_IO_L1_out_wrapper_185__ap_done ap_idle=C_drain_IO_L1_out_wrapper_185__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_185__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_186__ap_start ap_done=C_drain_IO_L1_out_wrapper_186__ap_done ap_idle=C_drain_IO_L1_out_wrapper_186__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_186__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_187__ap_start ap_done=C_drain_IO_L1_out_wrapper_187__ap_done ap_idle=C_drain_IO_L1_out_wrapper_187__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_187__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_188__ap_start ap_done=C_drain_IO_L1_out_wrapper_188__ap_done ap_idle=C_drain_IO_L1_out_wrapper_188__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_188__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_189__ap_start ap_done=C_drain_IO_L1_out_wrapper_189__ap_done ap_idle=C_drain_IO_L1_out_wrapper_189__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_189__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_190__ap_start ap_done=C_drain_IO_L1_out_wrapper_190__ap_done ap_idle=C_drain_IO_L1_out_wrapper_190__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_190__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_191__ap_start ap_done=C_drain_IO_L1_out_wrapper_191__ap_done ap_idle=C_drain_IO_L1_out_wrapper_191__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_191__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_192__ap_start ap_done=C_drain_IO_L1_out_wrapper_192__ap_done ap_idle=C_drain_IO_L1_out_wrapper_192__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_192__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_193__ap_start ap_done=C_drain_IO_L1_out_wrapper_193__ap_done ap_idle=C_drain_IO_L1_out_wrapper_193__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_193__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_194__ap_start ap_done=C_drain_IO_L1_out_wrapper_194__ap_done ap_idle=C_drain_IO_L1_out_wrapper_194__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_194__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_195__ap_start ap_done=C_drain_IO_L1_out_wrapper_195__ap_done ap_idle=C_drain_IO_L1_out_wrapper_195__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_195__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_196__ap_start ap_done=C_drain_IO_L1_out_wrapper_196__ap_done ap_idle=C_drain_IO_L1_out_wrapper_196__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_196__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_197__ap_start ap_done=C_drain_IO_L1_out_wrapper_197__ap_done ap_idle=C_drain_IO_L1_out_wrapper_197__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_197__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_198__ap_start ap_done=C_drain_IO_L1_out_wrapper_198__ap_done ap_idle=C_drain_IO_L1_out_wrapper_198__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_198__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_199__ap_start ap_done=C_drain_IO_L1_out_wrapper_199__ap_done ap_idle=C_drain_IO_L1_out_wrapper_199__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_199__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_200__ap_start ap_done=C_drain_IO_L1_out_wrapper_200__ap_done ap_idle=C_drain_IO_L1_out_wrapper_200__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_200__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_201__ap_start ap_done=C_drain_IO_L1_out_wrapper_201__ap_done ap_idle=C_drain_IO_L1_out_wrapper_201__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_201__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_202__ap_start ap_done=C_drain_IO_L1_out_wrapper_202__ap_done ap_idle=C_drain_IO_L1_out_wrapper_202__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_202__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_203__ap_start ap_done=C_drain_IO_L1_out_wrapper_203__ap_done ap_idle=C_drain_IO_L1_out_wrapper_203__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_203__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_204__ap_start ap_done=C_drain_IO_L1_out_wrapper_204__ap_done ap_idle=C_drain_IO_L1_out_wrapper_204__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_204__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_205__ap_start ap_done=C_drain_IO_L1_out_wrapper_205__ap_done ap_idle=C_drain_IO_L1_out_wrapper_205__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_205__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_206__ap_start ap_done=C_drain_IO_L1_out_wrapper_206__ap_done ap_idle=C_drain_IO_L1_out_wrapper_206__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_206__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_207__ap_start ap_done=C_drain_IO_L1_out_wrapper_207__ap_done ap_idle=C_drain_IO_L1_out_wrapper_207__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_207__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_208__ap_start ap_done=C_drain_IO_L1_out_wrapper_208__ap_done ap_idle=C_drain_IO_L1_out_wrapper_208__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_208__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_209__ap_start ap_done=C_drain_IO_L1_out_wrapper_209__ap_done ap_idle=C_drain_IO_L1_out_wrapper_209__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_209__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_210__ap_start ap_done=C_drain_IO_L1_out_wrapper_210__ap_done ap_idle=C_drain_IO_L1_out_wrapper_210__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_210__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_211__ap_start ap_done=C_drain_IO_L1_out_wrapper_211__ap_done ap_idle=C_drain_IO_L1_out_wrapper_211__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_211__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_212__ap_start ap_done=C_drain_IO_L1_out_wrapper_212__ap_done ap_idle=C_drain_IO_L1_out_wrapper_212__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_212__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_213__ap_start ap_done=C_drain_IO_L1_out_wrapper_213__ap_done ap_idle=C_drain_IO_L1_out_wrapper_213__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_213__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_214__ap_start ap_done=C_drain_IO_L1_out_wrapper_214__ap_done ap_idle=C_drain_IO_L1_out_wrapper_214__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_214__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_215__ap_start ap_done=C_drain_IO_L1_out_wrapper_215__ap_done ap_idle=C_drain_IO_L1_out_wrapper_215__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_215__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_216__ap_start ap_done=C_drain_IO_L1_out_wrapper_216__ap_done ap_idle=C_drain_IO_L1_out_wrapper_216__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_216__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_217__ap_start ap_done=C_drain_IO_L1_out_wrapper_217__ap_done ap_idle=C_drain_IO_L1_out_wrapper_217__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_217__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_218__ap_start ap_done=C_drain_IO_L1_out_wrapper_218__ap_done ap_idle=C_drain_IO_L1_out_wrapper_218__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_218__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_219__ap_start ap_done=C_drain_IO_L1_out_wrapper_219__ap_done ap_idle=C_drain_IO_L1_out_wrapper_219__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_219__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_220__ap_start ap_done=C_drain_IO_L1_out_wrapper_220__ap_done ap_idle=C_drain_IO_L1_out_wrapper_220__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_220__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_221__ap_start ap_done=C_drain_IO_L1_out_wrapper_221__ap_done ap_idle=C_drain_IO_L1_out_wrapper_221__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_221__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_222__ap_start ap_done=C_drain_IO_L1_out_wrapper_222__ap_done ap_idle=C_drain_IO_L1_out_wrapper_222__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_222__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_223__ap_start ap_done=C_drain_IO_L1_out_wrapper_223__ap_done ap_idle=C_drain_IO_L1_out_wrapper_223__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_223__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_224__ap_start ap_done=C_drain_IO_L1_out_wrapper_224__ap_done ap_idle=C_drain_IO_L1_out_wrapper_224__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_224__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_225__ap_start ap_done=C_drain_IO_L1_out_wrapper_225__ap_done ap_idle=C_drain_IO_L1_out_wrapper_225__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_225__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_226__ap_start ap_done=C_drain_IO_L1_out_wrapper_226__ap_done ap_idle=C_drain_IO_L1_out_wrapper_226__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_226__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_227__ap_start ap_done=C_drain_IO_L1_out_wrapper_227__ap_done ap_idle=C_drain_IO_L1_out_wrapper_227__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_227__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_228__ap_start ap_done=C_drain_IO_L1_out_wrapper_228__ap_done ap_idle=C_drain_IO_L1_out_wrapper_228__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_228__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_229__ap_start ap_done=C_drain_IO_L1_out_wrapper_229__ap_done ap_idle=C_drain_IO_L1_out_wrapper_229__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_229__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_230__ap_start ap_done=C_drain_IO_L1_out_wrapper_230__ap_done ap_idle=C_drain_IO_L1_out_wrapper_230__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_230__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_231__ap_start ap_done=C_drain_IO_L1_out_wrapper_231__ap_done ap_idle=C_drain_IO_L1_out_wrapper_231__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_231__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_232__ap_start ap_done=C_drain_IO_L1_out_wrapper_232__ap_done ap_idle=C_drain_IO_L1_out_wrapper_232__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_232__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_233__ap_start ap_done=C_drain_IO_L1_out_wrapper_233__ap_done ap_idle=C_drain_IO_L1_out_wrapper_233__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_233__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_234__ap_start ap_done=C_drain_IO_L1_out_wrapper_234__ap_done ap_idle=C_drain_IO_L1_out_wrapper_234__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_234__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_235__ap_start ap_done=C_drain_IO_L1_out_wrapper_235__ap_done ap_idle=C_drain_IO_L1_out_wrapper_235__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_235__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_236__ap_start ap_done=C_drain_IO_L1_out_wrapper_236__ap_done ap_idle=C_drain_IO_L1_out_wrapper_236__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_236__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_237__ap_start ap_done=C_drain_IO_L1_out_wrapper_237__ap_done ap_idle=C_drain_IO_L1_out_wrapper_237__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_237__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_238__ap_start ap_done=C_drain_IO_L1_out_wrapper_238__ap_done ap_idle=C_drain_IO_L1_out_wrapper_238__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_238__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_239__ap_start ap_done=C_drain_IO_L1_out_wrapper_239__ap_done ap_idle=C_drain_IO_L1_out_wrapper_239__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_239__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_240__ap_start ap_done=C_drain_IO_L1_out_wrapper_240__ap_done ap_idle=C_drain_IO_L1_out_wrapper_240__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_240__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_241__ap_start ap_done=C_drain_IO_L1_out_wrapper_241__ap_done ap_idle=C_drain_IO_L1_out_wrapper_241__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_241__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_242__ap_start ap_done=C_drain_IO_L1_out_wrapper_242__ap_done ap_idle=C_drain_IO_L1_out_wrapper_242__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_242__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_243__ap_start ap_done=C_drain_IO_L1_out_wrapper_243__ap_done ap_idle=C_drain_IO_L1_out_wrapper_243__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_243__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_244__ap_start ap_done=C_drain_IO_L1_out_wrapper_244__ap_done ap_idle=C_drain_IO_L1_out_wrapper_244__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_244__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_245__ap_start ap_done=C_drain_IO_L1_out_wrapper_245__ap_done ap_idle=C_drain_IO_L1_out_wrapper_245__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_245__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_246__ap_start ap_done=C_drain_IO_L1_out_wrapper_246__ap_done ap_idle=C_drain_IO_L1_out_wrapper_246__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_246__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_247__ap_start ap_done=C_drain_IO_L1_out_wrapper_247__ap_done ap_idle=C_drain_IO_L1_out_wrapper_247__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_247__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_248__ap_start ap_done=C_drain_IO_L1_out_wrapper_248__ap_done ap_idle=C_drain_IO_L1_out_wrapper_248__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_248__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_249__ap_start ap_done=C_drain_IO_L1_out_wrapper_249__ap_done ap_idle=C_drain_IO_L1_out_wrapper_249__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_249__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_250__ap_start ap_done=C_drain_IO_L1_out_wrapper_250__ap_done ap_idle=C_drain_IO_L1_out_wrapper_250__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_250__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_251__ap_start ap_done=C_drain_IO_L1_out_wrapper_251__ap_done ap_idle=C_drain_IO_L1_out_wrapper_251__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_251__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_252__ap_start ap_done=C_drain_IO_L1_out_wrapper_252__ap_done ap_idle=C_drain_IO_L1_out_wrapper_252__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_252__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_253__ap_start ap_done=C_drain_IO_L1_out_wrapper_253__ap_done ap_idle=C_drain_IO_L1_out_wrapper_253__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_253__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_254__ap_start ap_done=C_drain_IO_L1_out_wrapper_254__ap_done ap_idle=C_drain_IO_L1_out_wrapper_254__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_254__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_255__ap_start ap_done=C_drain_IO_L1_out_wrapper_255__ap_done ap_idle=C_drain_IO_L1_out_wrapper_255__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_255__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_256__ap_start ap_done=C_drain_IO_L1_out_wrapper_256__ap_done ap_idle=C_drain_IO_L1_out_wrapper_256__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_256__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_257__ap_start ap_done=C_drain_IO_L1_out_wrapper_257__ap_done ap_idle=C_drain_IO_L1_out_wrapper_257__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_257__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_258__ap_start ap_done=C_drain_IO_L1_out_wrapper_258__ap_done ap_idle=C_drain_IO_L1_out_wrapper_258__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_258__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_259__ap_start ap_done=C_drain_IO_L1_out_wrapper_259__ap_done ap_idle=C_drain_IO_L1_out_wrapper_259__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_259__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_260__ap_start ap_done=C_drain_IO_L1_out_wrapper_260__ap_done ap_idle=C_drain_IO_L1_out_wrapper_260__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_260__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_261__ap_start ap_done=C_drain_IO_L1_out_wrapper_261__ap_done ap_idle=C_drain_IO_L1_out_wrapper_261__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_261__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_262__ap_start ap_done=C_drain_IO_L1_out_wrapper_262__ap_done ap_idle=C_drain_IO_L1_out_wrapper_262__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_262__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_263__ap_start ap_done=C_drain_IO_L1_out_wrapper_263__ap_done ap_idle=C_drain_IO_L1_out_wrapper_263__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_263__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_264__ap_start ap_done=C_drain_IO_L1_out_wrapper_264__ap_done ap_idle=C_drain_IO_L1_out_wrapper_264__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_264__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_265__ap_start ap_done=C_drain_IO_L1_out_wrapper_265__ap_done ap_idle=C_drain_IO_L1_out_wrapper_265__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_265__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_266__ap_start ap_done=C_drain_IO_L1_out_wrapper_266__ap_done ap_idle=C_drain_IO_L1_out_wrapper_266__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_266__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_267__ap_start ap_done=C_drain_IO_L1_out_wrapper_267__ap_done ap_idle=C_drain_IO_L1_out_wrapper_267__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_267__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_268__ap_start ap_done=C_drain_IO_L1_out_wrapper_268__ap_done ap_idle=C_drain_IO_L1_out_wrapper_268__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_268__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_269__ap_start ap_done=C_drain_IO_L1_out_wrapper_269__ap_done ap_idle=C_drain_IO_L1_out_wrapper_269__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_269__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_270__ap_start ap_done=C_drain_IO_L1_out_wrapper_270__ap_done ap_idle=C_drain_IO_L1_out_wrapper_270__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_270__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_271__ap_start ap_done=C_drain_IO_L1_out_wrapper_271__ap_done ap_idle=C_drain_IO_L1_out_wrapper_271__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_271__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_272__ap_start ap_done=C_drain_IO_L1_out_wrapper_272__ap_done ap_idle=C_drain_IO_L1_out_wrapper_272__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_272__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_273__ap_start ap_done=C_drain_IO_L1_out_wrapper_273__ap_done ap_idle=C_drain_IO_L1_out_wrapper_273__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_273__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_274__ap_start ap_done=C_drain_IO_L1_out_wrapper_274__ap_done ap_idle=C_drain_IO_L1_out_wrapper_274__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_274__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_275__ap_start ap_done=C_drain_IO_L1_out_wrapper_275__ap_done ap_idle=C_drain_IO_L1_out_wrapper_275__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_275__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_276__ap_start ap_done=C_drain_IO_L1_out_wrapper_276__ap_done ap_idle=C_drain_IO_L1_out_wrapper_276__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_276__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_277__ap_start ap_done=C_drain_IO_L1_out_wrapper_277__ap_done ap_idle=C_drain_IO_L1_out_wrapper_277__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_277__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_278__ap_start ap_done=C_drain_IO_L1_out_wrapper_278__ap_done ap_idle=C_drain_IO_L1_out_wrapper_278__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_278__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_279__ap_start ap_done=C_drain_IO_L1_out_wrapper_279__ap_done ap_idle=C_drain_IO_L1_out_wrapper_279__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_279__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_280__ap_start ap_done=C_drain_IO_L1_out_wrapper_280__ap_done ap_idle=C_drain_IO_L1_out_wrapper_280__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_280__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_281__ap_start ap_done=C_drain_IO_L1_out_wrapper_281__ap_done ap_idle=C_drain_IO_L1_out_wrapper_281__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_281__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_282__ap_start ap_done=C_drain_IO_L1_out_wrapper_282__ap_done ap_idle=C_drain_IO_L1_out_wrapper_282__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_282__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_283__ap_start ap_done=C_drain_IO_L1_out_wrapper_283__ap_done ap_idle=C_drain_IO_L1_out_wrapper_283__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_283__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_284__ap_start ap_done=C_drain_IO_L1_out_wrapper_284__ap_done ap_idle=C_drain_IO_L1_out_wrapper_284__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_284__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_285__ap_start ap_done=C_drain_IO_L1_out_wrapper_285__ap_done ap_idle=C_drain_IO_L1_out_wrapper_285__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_285__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_286__ap_start ap_done=C_drain_IO_L1_out_wrapper_286__ap_done ap_idle=C_drain_IO_L1_out_wrapper_286__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_286__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_287__ap_start ap_done=C_drain_IO_L1_out_wrapper_287__ap_done ap_idle=C_drain_IO_L1_out_wrapper_287__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_287__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L1_out_wrapper_288__ap_start ap_done=C_drain_IO_L1_out_wrapper_288__ap_done ap_idle=C_drain_IO_L1_out_wrapper_288__ap_idle ap_ready=C_drain_IO_L1_out_wrapper_288__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L2_out_0__ap_start ap_done=C_drain_IO_L2_out_0__ap_done ap_idle=C_drain_IO_L2_out_0__ap_idle ap_ready=C_drain_IO_L2_out_0__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L2_out_1__ap_start ap_done=C_drain_IO_L2_out_1__ap_done ap_idle=C_drain_IO_L2_out_1__ap_idle ap_ready=C_drain_IO_L2_out_1__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L2_out_2__ap_start ap_done=C_drain_IO_L2_out_2__ap_done ap_idle=C_drain_IO_L2_out_2__ap_idle ap_ready=C_drain_IO_L2_out_2__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L2_out_3__ap_start ap_done=C_drain_IO_L2_out_3__ap_done ap_idle=C_drain_IO_L2_out_3__ap_idle ap_ready=C_drain_IO_L2_out_3__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L2_out_4__ap_start ap_done=C_drain_IO_L2_out_4__ap_done ap_idle=C_drain_IO_L2_out_4__ap_idle ap_ready=C_drain_IO_L2_out_4__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L2_out_5__ap_start ap_done=C_drain_IO_L2_out_5__ap_done ap_idle=C_drain_IO_L2_out_5__ap_idle ap_ready=C_drain_IO_L2_out_5__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L2_out_6__ap_start ap_done=C_drain_IO_L2_out_6__ap_done ap_idle=C_drain_IO_L2_out_6__ap_idle ap_ready=C_drain_IO_L2_out_6__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L2_out_7__ap_start ap_done=C_drain_IO_L2_out_7__ap_done ap_idle=C_drain_IO_L2_out_7__ap_idle ap_ready=C_drain_IO_L2_out_7__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L2_out_8__ap_start ap_done=C_drain_IO_L2_out_8__ap_done ap_idle=C_drain_IO_L2_out_8__ap_idle ap_ready=C_drain_IO_L2_out_8__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L2_out_9__ap_start ap_done=C_drain_IO_L2_out_9__ap_done ap_idle=C_drain_IO_L2_out_9__ap_idle ap_ready=C_drain_IO_L2_out_9__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L2_out_10__ap_start ap_done=C_drain_IO_L2_out_10__ap_done ap_idle=C_drain_IO_L2_out_10__ap_idle ap_ready=C_drain_IO_L2_out_10__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L2_out_11__ap_start ap_done=C_drain_IO_L2_out_11__ap_done ap_idle=C_drain_IO_L2_out_11__ap_idle ap_ready=C_drain_IO_L2_out_11__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L2_out_12__ap_start ap_done=C_drain_IO_L2_out_12__ap_done ap_idle=C_drain_IO_L2_out_12__ap_idle ap_ready=C_drain_IO_L2_out_12__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L2_out_13__ap_start ap_done=C_drain_IO_L2_out_13__ap_done ap_idle=C_drain_IO_L2_out_13__ap_idle ap_ready=C_drain_IO_L2_out_13__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L2_out_14__ap_start ap_done=C_drain_IO_L2_out_14__ap_done ap_idle=C_drain_IO_L2_out_14__ap_idle ap_ready=C_drain_IO_L2_out_14__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L2_out_15__ap_start ap_done=C_drain_IO_L2_out_15__ap_done ap_idle=C_drain_IO_L2_out_15__ap_idle ap_ready=C_drain_IO_L2_out_15__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L2_out_boundary_0__ap_start ap_done=C_drain_IO_L2_out_boundary_0__ap_done ap_idle=C_drain_IO_L2_out_boundary_0__ap_idle ap_ready=C_drain_IO_L2_out_boundary_0__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L3_out_0__ap_start ap_done=C_drain_IO_L3_out_0__ap_done ap_idle=C_drain_IO_L3_out_0__ap_idle ap_ready=C_drain_IO_L3_out_0__ap_ready
  // pragma RS ap-ctrl ap_start=C_drain_IO_L3_out_serialize_0__ap_start ap_done=C_drain_IO_L3_out_serialize_0__ap_done ap_idle=C_drain_IO_L3_out_serialize_0__ap_idle ap_ready=C_drain_IO_L3_out_serialize_0__ap_ready scalar=C_drain_IO_L3_out_serialize_0___.*
  // pragma RS ap-ctrl ap_start=PE_wrapper_0__ap_start ap_done=PE_wrapper_0__ap_done ap_idle=PE_wrapper_0__ap_idle ap_ready=PE_wrapper_0__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_1__ap_start ap_done=PE_wrapper_1__ap_done ap_idle=PE_wrapper_1__ap_idle ap_ready=PE_wrapper_1__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_2__ap_start ap_done=PE_wrapper_2__ap_done ap_idle=PE_wrapper_2__ap_idle ap_ready=PE_wrapper_2__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_3__ap_start ap_done=PE_wrapper_3__ap_done ap_idle=PE_wrapper_3__ap_idle ap_ready=PE_wrapper_3__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_4__ap_start ap_done=PE_wrapper_4__ap_done ap_idle=PE_wrapper_4__ap_idle ap_ready=PE_wrapper_4__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_5__ap_start ap_done=PE_wrapper_5__ap_done ap_idle=PE_wrapper_5__ap_idle ap_ready=PE_wrapper_5__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_6__ap_start ap_done=PE_wrapper_6__ap_done ap_idle=PE_wrapper_6__ap_idle ap_ready=PE_wrapper_6__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_7__ap_start ap_done=PE_wrapper_7__ap_done ap_idle=PE_wrapper_7__ap_idle ap_ready=PE_wrapper_7__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_8__ap_start ap_done=PE_wrapper_8__ap_done ap_idle=PE_wrapper_8__ap_idle ap_ready=PE_wrapper_8__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_9__ap_start ap_done=PE_wrapper_9__ap_done ap_idle=PE_wrapper_9__ap_idle ap_ready=PE_wrapper_9__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_10__ap_start ap_done=PE_wrapper_10__ap_done ap_idle=PE_wrapper_10__ap_idle ap_ready=PE_wrapper_10__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_11__ap_start ap_done=PE_wrapper_11__ap_done ap_idle=PE_wrapper_11__ap_idle ap_ready=PE_wrapper_11__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_12__ap_start ap_done=PE_wrapper_12__ap_done ap_idle=PE_wrapper_12__ap_idle ap_ready=PE_wrapper_12__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_13__ap_start ap_done=PE_wrapper_13__ap_done ap_idle=PE_wrapper_13__ap_idle ap_ready=PE_wrapper_13__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_14__ap_start ap_done=PE_wrapper_14__ap_done ap_idle=PE_wrapper_14__ap_idle ap_ready=PE_wrapper_14__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_15__ap_start ap_done=PE_wrapper_15__ap_done ap_idle=PE_wrapper_15__ap_idle ap_ready=PE_wrapper_15__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_16__ap_start ap_done=PE_wrapper_16__ap_done ap_idle=PE_wrapper_16__ap_idle ap_ready=PE_wrapper_16__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_17__ap_start ap_done=PE_wrapper_17__ap_done ap_idle=PE_wrapper_17__ap_idle ap_ready=PE_wrapper_17__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_18__ap_start ap_done=PE_wrapper_18__ap_done ap_idle=PE_wrapper_18__ap_idle ap_ready=PE_wrapper_18__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_19__ap_start ap_done=PE_wrapper_19__ap_done ap_idle=PE_wrapper_19__ap_idle ap_ready=PE_wrapper_19__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_20__ap_start ap_done=PE_wrapper_20__ap_done ap_idle=PE_wrapper_20__ap_idle ap_ready=PE_wrapper_20__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_21__ap_start ap_done=PE_wrapper_21__ap_done ap_idle=PE_wrapper_21__ap_idle ap_ready=PE_wrapper_21__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_22__ap_start ap_done=PE_wrapper_22__ap_done ap_idle=PE_wrapper_22__ap_idle ap_ready=PE_wrapper_22__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_23__ap_start ap_done=PE_wrapper_23__ap_done ap_idle=PE_wrapper_23__ap_idle ap_ready=PE_wrapper_23__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_24__ap_start ap_done=PE_wrapper_24__ap_done ap_idle=PE_wrapper_24__ap_idle ap_ready=PE_wrapper_24__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_25__ap_start ap_done=PE_wrapper_25__ap_done ap_idle=PE_wrapper_25__ap_idle ap_ready=PE_wrapper_25__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_26__ap_start ap_done=PE_wrapper_26__ap_done ap_idle=PE_wrapper_26__ap_idle ap_ready=PE_wrapper_26__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_27__ap_start ap_done=PE_wrapper_27__ap_done ap_idle=PE_wrapper_27__ap_idle ap_ready=PE_wrapper_27__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_28__ap_start ap_done=PE_wrapper_28__ap_done ap_idle=PE_wrapper_28__ap_idle ap_ready=PE_wrapper_28__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_29__ap_start ap_done=PE_wrapper_29__ap_done ap_idle=PE_wrapper_29__ap_idle ap_ready=PE_wrapper_29__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_30__ap_start ap_done=PE_wrapper_30__ap_done ap_idle=PE_wrapper_30__ap_idle ap_ready=PE_wrapper_30__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_31__ap_start ap_done=PE_wrapper_31__ap_done ap_idle=PE_wrapper_31__ap_idle ap_ready=PE_wrapper_31__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_32__ap_start ap_done=PE_wrapper_32__ap_done ap_idle=PE_wrapper_32__ap_idle ap_ready=PE_wrapper_32__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_33__ap_start ap_done=PE_wrapper_33__ap_done ap_idle=PE_wrapper_33__ap_idle ap_ready=PE_wrapper_33__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_34__ap_start ap_done=PE_wrapper_34__ap_done ap_idle=PE_wrapper_34__ap_idle ap_ready=PE_wrapper_34__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_35__ap_start ap_done=PE_wrapper_35__ap_done ap_idle=PE_wrapper_35__ap_idle ap_ready=PE_wrapper_35__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_36__ap_start ap_done=PE_wrapper_36__ap_done ap_idle=PE_wrapper_36__ap_idle ap_ready=PE_wrapper_36__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_37__ap_start ap_done=PE_wrapper_37__ap_done ap_idle=PE_wrapper_37__ap_idle ap_ready=PE_wrapper_37__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_38__ap_start ap_done=PE_wrapper_38__ap_done ap_idle=PE_wrapper_38__ap_idle ap_ready=PE_wrapper_38__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_39__ap_start ap_done=PE_wrapper_39__ap_done ap_idle=PE_wrapper_39__ap_idle ap_ready=PE_wrapper_39__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_40__ap_start ap_done=PE_wrapper_40__ap_done ap_idle=PE_wrapper_40__ap_idle ap_ready=PE_wrapper_40__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_41__ap_start ap_done=PE_wrapper_41__ap_done ap_idle=PE_wrapper_41__ap_idle ap_ready=PE_wrapper_41__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_42__ap_start ap_done=PE_wrapper_42__ap_done ap_idle=PE_wrapper_42__ap_idle ap_ready=PE_wrapper_42__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_43__ap_start ap_done=PE_wrapper_43__ap_done ap_idle=PE_wrapper_43__ap_idle ap_ready=PE_wrapper_43__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_44__ap_start ap_done=PE_wrapper_44__ap_done ap_idle=PE_wrapper_44__ap_idle ap_ready=PE_wrapper_44__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_45__ap_start ap_done=PE_wrapper_45__ap_done ap_idle=PE_wrapper_45__ap_idle ap_ready=PE_wrapper_45__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_46__ap_start ap_done=PE_wrapper_46__ap_done ap_idle=PE_wrapper_46__ap_idle ap_ready=PE_wrapper_46__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_47__ap_start ap_done=PE_wrapper_47__ap_done ap_idle=PE_wrapper_47__ap_idle ap_ready=PE_wrapper_47__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_48__ap_start ap_done=PE_wrapper_48__ap_done ap_idle=PE_wrapper_48__ap_idle ap_ready=PE_wrapper_48__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_49__ap_start ap_done=PE_wrapper_49__ap_done ap_idle=PE_wrapper_49__ap_idle ap_ready=PE_wrapper_49__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_50__ap_start ap_done=PE_wrapper_50__ap_done ap_idle=PE_wrapper_50__ap_idle ap_ready=PE_wrapper_50__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_51__ap_start ap_done=PE_wrapper_51__ap_done ap_idle=PE_wrapper_51__ap_idle ap_ready=PE_wrapper_51__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_52__ap_start ap_done=PE_wrapper_52__ap_done ap_idle=PE_wrapper_52__ap_idle ap_ready=PE_wrapper_52__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_53__ap_start ap_done=PE_wrapper_53__ap_done ap_idle=PE_wrapper_53__ap_idle ap_ready=PE_wrapper_53__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_54__ap_start ap_done=PE_wrapper_54__ap_done ap_idle=PE_wrapper_54__ap_idle ap_ready=PE_wrapper_54__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_55__ap_start ap_done=PE_wrapper_55__ap_done ap_idle=PE_wrapper_55__ap_idle ap_ready=PE_wrapper_55__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_56__ap_start ap_done=PE_wrapper_56__ap_done ap_idle=PE_wrapper_56__ap_idle ap_ready=PE_wrapper_56__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_57__ap_start ap_done=PE_wrapper_57__ap_done ap_idle=PE_wrapper_57__ap_idle ap_ready=PE_wrapper_57__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_58__ap_start ap_done=PE_wrapper_58__ap_done ap_idle=PE_wrapper_58__ap_idle ap_ready=PE_wrapper_58__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_59__ap_start ap_done=PE_wrapper_59__ap_done ap_idle=PE_wrapper_59__ap_idle ap_ready=PE_wrapper_59__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_60__ap_start ap_done=PE_wrapper_60__ap_done ap_idle=PE_wrapper_60__ap_idle ap_ready=PE_wrapper_60__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_61__ap_start ap_done=PE_wrapper_61__ap_done ap_idle=PE_wrapper_61__ap_idle ap_ready=PE_wrapper_61__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_62__ap_start ap_done=PE_wrapper_62__ap_done ap_idle=PE_wrapper_62__ap_idle ap_ready=PE_wrapper_62__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_63__ap_start ap_done=PE_wrapper_63__ap_done ap_idle=PE_wrapper_63__ap_idle ap_ready=PE_wrapper_63__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_64__ap_start ap_done=PE_wrapper_64__ap_done ap_idle=PE_wrapper_64__ap_idle ap_ready=PE_wrapper_64__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_65__ap_start ap_done=PE_wrapper_65__ap_done ap_idle=PE_wrapper_65__ap_idle ap_ready=PE_wrapper_65__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_66__ap_start ap_done=PE_wrapper_66__ap_done ap_idle=PE_wrapper_66__ap_idle ap_ready=PE_wrapper_66__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_67__ap_start ap_done=PE_wrapper_67__ap_done ap_idle=PE_wrapper_67__ap_idle ap_ready=PE_wrapper_67__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_68__ap_start ap_done=PE_wrapper_68__ap_done ap_idle=PE_wrapper_68__ap_idle ap_ready=PE_wrapper_68__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_69__ap_start ap_done=PE_wrapper_69__ap_done ap_idle=PE_wrapper_69__ap_idle ap_ready=PE_wrapper_69__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_70__ap_start ap_done=PE_wrapper_70__ap_done ap_idle=PE_wrapper_70__ap_idle ap_ready=PE_wrapper_70__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_71__ap_start ap_done=PE_wrapper_71__ap_done ap_idle=PE_wrapper_71__ap_idle ap_ready=PE_wrapper_71__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_72__ap_start ap_done=PE_wrapper_72__ap_done ap_idle=PE_wrapper_72__ap_idle ap_ready=PE_wrapper_72__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_73__ap_start ap_done=PE_wrapper_73__ap_done ap_idle=PE_wrapper_73__ap_idle ap_ready=PE_wrapper_73__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_74__ap_start ap_done=PE_wrapper_74__ap_done ap_idle=PE_wrapper_74__ap_idle ap_ready=PE_wrapper_74__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_75__ap_start ap_done=PE_wrapper_75__ap_done ap_idle=PE_wrapper_75__ap_idle ap_ready=PE_wrapper_75__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_76__ap_start ap_done=PE_wrapper_76__ap_done ap_idle=PE_wrapper_76__ap_idle ap_ready=PE_wrapper_76__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_77__ap_start ap_done=PE_wrapper_77__ap_done ap_idle=PE_wrapper_77__ap_idle ap_ready=PE_wrapper_77__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_78__ap_start ap_done=PE_wrapper_78__ap_done ap_idle=PE_wrapper_78__ap_idle ap_ready=PE_wrapper_78__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_79__ap_start ap_done=PE_wrapper_79__ap_done ap_idle=PE_wrapper_79__ap_idle ap_ready=PE_wrapper_79__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_80__ap_start ap_done=PE_wrapper_80__ap_done ap_idle=PE_wrapper_80__ap_idle ap_ready=PE_wrapper_80__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_81__ap_start ap_done=PE_wrapper_81__ap_done ap_idle=PE_wrapper_81__ap_idle ap_ready=PE_wrapper_81__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_82__ap_start ap_done=PE_wrapper_82__ap_done ap_idle=PE_wrapper_82__ap_idle ap_ready=PE_wrapper_82__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_83__ap_start ap_done=PE_wrapper_83__ap_done ap_idle=PE_wrapper_83__ap_idle ap_ready=PE_wrapper_83__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_84__ap_start ap_done=PE_wrapper_84__ap_done ap_idle=PE_wrapper_84__ap_idle ap_ready=PE_wrapper_84__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_85__ap_start ap_done=PE_wrapper_85__ap_done ap_idle=PE_wrapper_85__ap_idle ap_ready=PE_wrapper_85__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_86__ap_start ap_done=PE_wrapper_86__ap_done ap_idle=PE_wrapper_86__ap_idle ap_ready=PE_wrapper_86__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_87__ap_start ap_done=PE_wrapper_87__ap_done ap_idle=PE_wrapper_87__ap_idle ap_ready=PE_wrapper_87__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_88__ap_start ap_done=PE_wrapper_88__ap_done ap_idle=PE_wrapper_88__ap_idle ap_ready=PE_wrapper_88__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_89__ap_start ap_done=PE_wrapper_89__ap_done ap_idle=PE_wrapper_89__ap_idle ap_ready=PE_wrapper_89__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_90__ap_start ap_done=PE_wrapper_90__ap_done ap_idle=PE_wrapper_90__ap_idle ap_ready=PE_wrapper_90__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_91__ap_start ap_done=PE_wrapper_91__ap_done ap_idle=PE_wrapper_91__ap_idle ap_ready=PE_wrapper_91__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_92__ap_start ap_done=PE_wrapper_92__ap_done ap_idle=PE_wrapper_92__ap_idle ap_ready=PE_wrapper_92__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_93__ap_start ap_done=PE_wrapper_93__ap_done ap_idle=PE_wrapper_93__ap_idle ap_ready=PE_wrapper_93__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_94__ap_start ap_done=PE_wrapper_94__ap_done ap_idle=PE_wrapper_94__ap_idle ap_ready=PE_wrapper_94__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_95__ap_start ap_done=PE_wrapper_95__ap_done ap_idle=PE_wrapper_95__ap_idle ap_ready=PE_wrapper_95__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_96__ap_start ap_done=PE_wrapper_96__ap_done ap_idle=PE_wrapper_96__ap_idle ap_ready=PE_wrapper_96__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_97__ap_start ap_done=PE_wrapper_97__ap_done ap_idle=PE_wrapper_97__ap_idle ap_ready=PE_wrapper_97__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_98__ap_start ap_done=PE_wrapper_98__ap_done ap_idle=PE_wrapper_98__ap_idle ap_ready=PE_wrapper_98__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_99__ap_start ap_done=PE_wrapper_99__ap_done ap_idle=PE_wrapper_99__ap_idle ap_ready=PE_wrapper_99__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_100__ap_start ap_done=PE_wrapper_100__ap_done ap_idle=PE_wrapper_100__ap_idle ap_ready=PE_wrapper_100__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_101__ap_start ap_done=PE_wrapper_101__ap_done ap_idle=PE_wrapper_101__ap_idle ap_ready=PE_wrapper_101__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_102__ap_start ap_done=PE_wrapper_102__ap_done ap_idle=PE_wrapper_102__ap_idle ap_ready=PE_wrapper_102__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_103__ap_start ap_done=PE_wrapper_103__ap_done ap_idle=PE_wrapper_103__ap_idle ap_ready=PE_wrapper_103__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_104__ap_start ap_done=PE_wrapper_104__ap_done ap_idle=PE_wrapper_104__ap_idle ap_ready=PE_wrapper_104__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_105__ap_start ap_done=PE_wrapper_105__ap_done ap_idle=PE_wrapper_105__ap_idle ap_ready=PE_wrapper_105__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_106__ap_start ap_done=PE_wrapper_106__ap_done ap_idle=PE_wrapper_106__ap_idle ap_ready=PE_wrapper_106__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_107__ap_start ap_done=PE_wrapper_107__ap_done ap_idle=PE_wrapper_107__ap_idle ap_ready=PE_wrapper_107__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_108__ap_start ap_done=PE_wrapper_108__ap_done ap_idle=PE_wrapper_108__ap_idle ap_ready=PE_wrapper_108__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_109__ap_start ap_done=PE_wrapper_109__ap_done ap_idle=PE_wrapper_109__ap_idle ap_ready=PE_wrapper_109__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_110__ap_start ap_done=PE_wrapper_110__ap_done ap_idle=PE_wrapper_110__ap_idle ap_ready=PE_wrapper_110__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_111__ap_start ap_done=PE_wrapper_111__ap_done ap_idle=PE_wrapper_111__ap_idle ap_ready=PE_wrapper_111__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_112__ap_start ap_done=PE_wrapper_112__ap_done ap_idle=PE_wrapper_112__ap_idle ap_ready=PE_wrapper_112__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_113__ap_start ap_done=PE_wrapper_113__ap_done ap_idle=PE_wrapper_113__ap_idle ap_ready=PE_wrapper_113__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_114__ap_start ap_done=PE_wrapper_114__ap_done ap_idle=PE_wrapper_114__ap_idle ap_ready=PE_wrapper_114__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_115__ap_start ap_done=PE_wrapper_115__ap_done ap_idle=PE_wrapper_115__ap_idle ap_ready=PE_wrapper_115__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_116__ap_start ap_done=PE_wrapper_116__ap_done ap_idle=PE_wrapper_116__ap_idle ap_ready=PE_wrapper_116__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_117__ap_start ap_done=PE_wrapper_117__ap_done ap_idle=PE_wrapper_117__ap_idle ap_ready=PE_wrapper_117__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_118__ap_start ap_done=PE_wrapper_118__ap_done ap_idle=PE_wrapper_118__ap_idle ap_ready=PE_wrapper_118__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_119__ap_start ap_done=PE_wrapper_119__ap_done ap_idle=PE_wrapper_119__ap_idle ap_ready=PE_wrapper_119__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_120__ap_start ap_done=PE_wrapper_120__ap_done ap_idle=PE_wrapper_120__ap_idle ap_ready=PE_wrapper_120__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_121__ap_start ap_done=PE_wrapper_121__ap_done ap_idle=PE_wrapper_121__ap_idle ap_ready=PE_wrapper_121__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_122__ap_start ap_done=PE_wrapper_122__ap_done ap_idle=PE_wrapper_122__ap_idle ap_ready=PE_wrapper_122__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_123__ap_start ap_done=PE_wrapper_123__ap_done ap_idle=PE_wrapper_123__ap_idle ap_ready=PE_wrapper_123__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_124__ap_start ap_done=PE_wrapper_124__ap_done ap_idle=PE_wrapper_124__ap_idle ap_ready=PE_wrapper_124__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_125__ap_start ap_done=PE_wrapper_125__ap_done ap_idle=PE_wrapper_125__ap_idle ap_ready=PE_wrapper_125__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_126__ap_start ap_done=PE_wrapper_126__ap_done ap_idle=PE_wrapper_126__ap_idle ap_ready=PE_wrapper_126__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_127__ap_start ap_done=PE_wrapper_127__ap_done ap_idle=PE_wrapper_127__ap_idle ap_ready=PE_wrapper_127__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_128__ap_start ap_done=PE_wrapper_128__ap_done ap_idle=PE_wrapper_128__ap_idle ap_ready=PE_wrapper_128__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_129__ap_start ap_done=PE_wrapper_129__ap_done ap_idle=PE_wrapper_129__ap_idle ap_ready=PE_wrapper_129__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_130__ap_start ap_done=PE_wrapper_130__ap_done ap_idle=PE_wrapper_130__ap_idle ap_ready=PE_wrapper_130__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_131__ap_start ap_done=PE_wrapper_131__ap_done ap_idle=PE_wrapper_131__ap_idle ap_ready=PE_wrapper_131__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_132__ap_start ap_done=PE_wrapper_132__ap_done ap_idle=PE_wrapper_132__ap_idle ap_ready=PE_wrapper_132__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_133__ap_start ap_done=PE_wrapper_133__ap_done ap_idle=PE_wrapper_133__ap_idle ap_ready=PE_wrapper_133__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_134__ap_start ap_done=PE_wrapper_134__ap_done ap_idle=PE_wrapper_134__ap_idle ap_ready=PE_wrapper_134__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_135__ap_start ap_done=PE_wrapper_135__ap_done ap_idle=PE_wrapper_135__ap_idle ap_ready=PE_wrapper_135__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_136__ap_start ap_done=PE_wrapper_136__ap_done ap_idle=PE_wrapper_136__ap_idle ap_ready=PE_wrapper_136__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_137__ap_start ap_done=PE_wrapper_137__ap_done ap_idle=PE_wrapper_137__ap_idle ap_ready=PE_wrapper_137__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_138__ap_start ap_done=PE_wrapper_138__ap_done ap_idle=PE_wrapper_138__ap_idle ap_ready=PE_wrapper_138__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_139__ap_start ap_done=PE_wrapper_139__ap_done ap_idle=PE_wrapper_139__ap_idle ap_ready=PE_wrapper_139__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_140__ap_start ap_done=PE_wrapper_140__ap_done ap_idle=PE_wrapper_140__ap_idle ap_ready=PE_wrapper_140__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_141__ap_start ap_done=PE_wrapper_141__ap_done ap_idle=PE_wrapper_141__ap_idle ap_ready=PE_wrapper_141__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_142__ap_start ap_done=PE_wrapper_142__ap_done ap_idle=PE_wrapper_142__ap_idle ap_ready=PE_wrapper_142__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_143__ap_start ap_done=PE_wrapper_143__ap_done ap_idle=PE_wrapper_143__ap_idle ap_ready=PE_wrapper_143__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_144__ap_start ap_done=PE_wrapper_144__ap_done ap_idle=PE_wrapper_144__ap_idle ap_ready=PE_wrapper_144__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_145__ap_start ap_done=PE_wrapper_145__ap_done ap_idle=PE_wrapper_145__ap_idle ap_ready=PE_wrapper_145__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_146__ap_start ap_done=PE_wrapper_146__ap_done ap_idle=PE_wrapper_146__ap_idle ap_ready=PE_wrapper_146__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_147__ap_start ap_done=PE_wrapper_147__ap_done ap_idle=PE_wrapper_147__ap_idle ap_ready=PE_wrapper_147__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_148__ap_start ap_done=PE_wrapper_148__ap_done ap_idle=PE_wrapper_148__ap_idle ap_ready=PE_wrapper_148__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_149__ap_start ap_done=PE_wrapper_149__ap_done ap_idle=PE_wrapper_149__ap_idle ap_ready=PE_wrapper_149__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_150__ap_start ap_done=PE_wrapper_150__ap_done ap_idle=PE_wrapper_150__ap_idle ap_ready=PE_wrapper_150__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_151__ap_start ap_done=PE_wrapper_151__ap_done ap_idle=PE_wrapper_151__ap_idle ap_ready=PE_wrapper_151__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_152__ap_start ap_done=PE_wrapper_152__ap_done ap_idle=PE_wrapper_152__ap_idle ap_ready=PE_wrapper_152__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_153__ap_start ap_done=PE_wrapper_153__ap_done ap_idle=PE_wrapper_153__ap_idle ap_ready=PE_wrapper_153__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_154__ap_start ap_done=PE_wrapper_154__ap_done ap_idle=PE_wrapper_154__ap_idle ap_ready=PE_wrapper_154__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_155__ap_start ap_done=PE_wrapper_155__ap_done ap_idle=PE_wrapper_155__ap_idle ap_ready=PE_wrapper_155__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_156__ap_start ap_done=PE_wrapper_156__ap_done ap_idle=PE_wrapper_156__ap_idle ap_ready=PE_wrapper_156__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_157__ap_start ap_done=PE_wrapper_157__ap_done ap_idle=PE_wrapper_157__ap_idle ap_ready=PE_wrapper_157__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_158__ap_start ap_done=PE_wrapper_158__ap_done ap_idle=PE_wrapper_158__ap_idle ap_ready=PE_wrapper_158__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_159__ap_start ap_done=PE_wrapper_159__ap_done ap_idle=PE_wrapper_159__ap_idle ap_ready=PE_wrapper_159__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_160__ap_start ap_done=PE_wrapper_160__ap_done ap_idle=PE_wrapper_160__ap_idle ap_ready=PE_wrapper_160__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_161__ap_start ap_done=PE_wrapper_161__ap_done ap_idle=PE_wrapper_161__ap_idle ap_ready=PE_wrapper_161__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_162__ap_start ap_done=PE_wrapper_162__ap_done ap_idle=PE_wrapper_162__ap_idle ap_ready=PE_wrapper_162__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_163__ap_start ap_done=PE_wrapper_163__ap_done ap_idle=PE_wrapper_163__ap_idle ap_ready=PE_wrapper_163__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_164__ap_start ap_done=PE_wrapper_164__ap_done ap_idle=PE_wrapper_164__ap_idle ap_ready=PE_wrapper_164__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_165__ap_start ap_done=PE_wrapper_165__ap_done ap_idle=PE_wrapper_165__ap_idle ap_ready=PE_wrapper_165__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_166__ap_start ap_done=PE_wrapper_166__ap_done ap_idle=PE_wrapper_166__ap_idle ap_ready=PE_wrapper_166__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_167__ap_start ap_done=PE_wrapper_167__ap_done ap_idle=PE_wrapper_167__ap_idle ap_ready=PE_wrapper_167__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_168__ap_start ap_done=PE_wrapper_168__ap_done ap_idle=PE_wrapper_168__ap_idle ap_ready=PE_wrapper_168__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_169__ap_start ap_done=PE_wrapper_169__ap_done ap_idle=PE_wrapper_169__ap_idle ap_ready=PE_wrapper_169__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_170__ap_start ap_done=PE_wrapper_170__ap_done ap_idle=PE_wrapper_170__ap_idle ap_ready=PE_wrapper_170__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_171__ap_start ap_done=PE_wrapper_171__ap_done ap_idle=PE_wrapper_171__ap_idle ap_ready=PE_wrapper_171__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_172__ap_start ap_done=PE_wrapper_172__ap_done ap_idle=PE_wrapper_172__ap_idle ap_ready=PE_wrapper_172__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_173__ap_start ap_done=PE_wrapper_173__ap_done ap_idle=PE_wrapper_173__ap_idle ap_ready=PE_wrapper_173__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_174__ap_start ap_done=PE_wrapper_174__ap_done ap_idle=PE_wrapper_174__ap_idle ap_ready=PE_wrapper_174__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_175__ap_start ap_done=PE_wrapper_175__ap_done ap_idle=PE_wrapper_175__ap_idle ap_ready=PE_wrapper_175__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_176__ap_start ap_done=PE_wrapper_176__ap_done ap_idle=PE_wrapper_176__ap_idle ap_ready=PE_wrapper_176__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_177__ap_start ap_done=PE_wrapper_177__ap_done ap_idle=PE_wrapper_177__ap_idle ap_ready=PE_wrapper_177__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_178__ap_start ap_done=PE_wrapper_178__ap_done ap_idle=PE_wrapper_178__ap_idle ap_ready=PE_wrapper_178__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_179__ap_start ap_done=PE_wrapper_179__ap_done ap_idle=PE_wrapper_179__ap_idle ap_ready=PE_wrapper_179__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_180__ap_start ap_done=PE_wrapper_180__ap_done ap_idle=PE_wrapper_180__ap_idle ap_ready=PE_wrapper_180__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_181__ap_start ap_done=PE_wrapper_181__ap_done ap_idle=PE_wrapper_181__ap_idle ap_ready=PE_wrapper_181__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_182__ap_start ap_done=PE_wrapper_182__ap_done ap_idle=PE_wrapper_182__ap_idle ap_ready=PE_wrapper_182__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_183__ap_start ap_done=PE_wrapper_183__ap_done ap_idle=PE_wrapper_183__ap_idle ap_ready=PE_wrapper_183__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_184__ap_start ap_done=PE_wrapper_184__ap_done ap_idle=PE_wrapper_184__ap_idle ap_ready=PE_wrapper_184__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_185__ap_start ap_done=PE_wrapper_185__ap_done ap_idle=PE_wrapper_185__ap_idle ap_ready=PE_wrapper_185__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_186__ap_start ap_done=PE_wrapper_186__ap_done ap_idle=PE_wrapper_186__ap_idle ap_ready=PE_wrapper_186__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_187__ap_start ap_done=PE_wrapper_187__ap_done ap_idle=PE_wrapper_187__ap_idle ap_ready=PE_wrapper_187__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_188__ap_start ap_done=PE_wrapper_188__ap_done ap_idle=PE_wrapper_188__ap_idle ap_ready=PE_wrapper_188__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_189__ap_start ap_done=PE_wrapper_189__ap_done ap_idle=PE_wrapper_189__ap_idle ap_ready=PE_wrapper_189__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_190__ap_start ap_done=PE_wrapper_190__ap_done ap_idle=PE_wrapper_190__ap_idle ap_ready=PE_wrapper_190__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_191__ap_start ap_done=PE_wrapper_191__ap_done ap_idle=PE_wrapper_191__ap_idle ap_ready=PE_wrapper_191__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_192__ap_start ap_done=PE_wrapper_192__ap_done ap_idle=PE_wrapper_192__ap_idle ap_ready=PE_wrapper_192__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_193__ap_start ap_done=PE_wrapper_193__ap_done ap_idle=PE_wrapper_193__ap_idle ap_ready=PE_wrapper_193__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_194__ap_start ap_done=PE_wrapper_194__ap_done ap_idle=PE_wrapper_194__ap_idle ap_ready=PE_wrapper_194__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_195__ap_start ap_done=PE_wrapper_195__ap_done ap_idle=PE_wrapper_195__ap_idle ap_ready=PE_wrapper_195__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_196__ap_start ap_done=PE_wrapper_196__ap_done ap_idle=PE_wrapper_196__ap_idle ap_ready=PE_wrapper_196__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_197__ap_start ap_done=PE_wrapper_197__ap_done ap_idle=PE_wrapper_197__ap_idle ap_ready=PE_wrapper_197__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_198__ap_start ap_done=PE_wrapper_198__ap_done ap_idle=PE_wrapper_198__ap_idle ap_ready=PE_wrapper_198__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_199__ap_start ap_done=PE_wrapper_199__ap_done ap_idle=PE_wrapper_199__ap_idle ap_ready=PE_wrapper_199__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_200__ap_start ap_done=PE_wrapper_200__ap_done ap_idle=PE_wrapper_200__ap_idle ap_ready=PE_wrapper_200__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_201__ap_start ap_done=PE_wrapper_201__ap_done ap_idle=PE_wrapper_201__ap_idle ap_ready=PE_wrapper_201__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_202__ap_start ap_done=PE_wrapper_202__ap_done ap_idle=PE_wrapper_202__ap_idle ap_ready=PE_wrapper_202__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_203__ap_start ap_done=PE_wrapper_203__ap_done ap_idle=PE_wrapper_203__ap_idle ap_ready=PE_wrapper_203__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_204__ap_start ap_done=PE_wrapper_204__ap_done ap_idle=PE_wrapper_204__ap_idle ap_ready=PE_wrapper_204__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_205__ap_start ap_done=PE_wrapper_205__ap_done ap_idle=PE_wrapper_205__ap_idle ap_ready=PE_wrapper_205__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_206__ap_start ap_done=PE_wrapper_206__ap_done ap_idle=PE_wrapper_206__ap_idle ap_ready=PE_wrapper_206__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_207__ap_start ap_done=PE_wrapper_207__ap_done ap_idle=PE_wrapper_207__ap_idle ap_ready=PE_wrapper_207__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_208__ap_start ap_done=PE_wrapper_208__ap_done ap_idle=PE_wrapper_208__ap_idle ap_ready=PE_wrapper_208__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_209__ap_start ap_done=PE_wrapper_209__ap_done ap_idle=PE_wrapper_209__ap_idle ap_ready=PE_wrapper_209__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_210__ap_start ap_done=PE_wrapper_210__ap_done ap_idle=PE_wrapper_210__ap_idle ap_ready=PE_wrapper_210__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_211__ap_start ap_done=PE_wrapper_211__ap_done ap_idle=PE_wrapper_211__ap_idle ap_ready=PE_wrapper_211__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_212__ap_start ap_done=PE_wrapper_212__ap_done ap_idle=PE_wrapper_212__ap_idle ap_ready=PE_wrapper_212__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_213__ap_start ap_done=PE_wrapper_213__ap_done ap_idle=PE_wrapper_213__ap_idle ap_ready=PE_wrapper_213__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_214__ap_start ap_done=PE_wrapper_214__ap_done ap_idle=PE_wrapper_214__ap_idle ap_ready=PE_wrapper_214__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_215__ap_start ap_done=PE_wrapper_215__ap_done ap_idle=PE_wrapper_215__ap_idle ap_ready=PE_wrapper_215__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_216__ap_start ap_done=PE_wrapper_216__ap_done ap_idle=PE_wrapper_216__ap_idle ap_ready=PE_wrapper_216__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_217__ap_start ap_done=PE_wrapper_217__ap_done ap_idle=PE_wrapper_217__ap_idle ap_ready=PE_wrapper_217__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_218__ap_start ap_done=PE_wrapper_218__ap_done ap_idle=PE_wrapper_218__ap_idle ap_ready=PE_wrapper_218__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_219__ap_start ap_done=PE_wrapper_219__ap_done ap_idle=PE_wrapper_219__ap_idle ap_ready=PE_wrapper_219__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_220__ap_start ap_done=PE_wrapper_220__ap_done ap_idle=PE_wrapper_220__ap_idle ap_ready=PE_wrapper_220__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_221__ap_start ap_done=PE_wrapper_221__ap_done ap_idle=PE_wrapper_221__ap_idle ap_ready=PE_wrapper_221__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_222__ap_start ap_done=PE_wrapper_222__ap_done ap_idle=PE_wrapper_222__ap_idle ap_ready=PE_wrapper_222__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_223__ap_start ap_done=PE_wrapper_223__ap_done ap_idle=PE_wrapper_223__ap_idle ap_ready=PE_wrapper_223__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_224__ap_start ap_done=PE_wrapper_224__ap_done ap_idle=PE_wrapper_224__ap_idle ap_ready=PE_wrapper_224__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_225__ap_start ap_done=PE_wrapper_225__ap_done ap_idle=PE_wrapper_225__ap_idle ap_ready=PE_wrapper_225__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_226__ap_start ap_done=PE_wrapper_226__ap_done ap_idle=PE_wrapper_226__ap_idle ap_ready=PE_wrapper_226__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_227__ap_start ap_done=PE_wrapper_227__ap_done ap_idle=PE_wrapper_227__ap_idle ap_ready=PE_wrapper_227__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_228__ap_start ap_done=PE_wrapper_228__ap_done ap_idle=PE_wrapper_228__ap_idle ap_ready=PE_wrapper_228__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_229__ap_start ap_done=PE_wrapper_229__ap_done ap_idle=PE_wrapper_229__ap_idle ap_ready=PE_wrapper_229__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_230__ap_start ap_done=PE_wrapper_230__ap_done ap_idle=PE_wrapper_230__ap_idle ap_ready=PE_wrapper_230__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_231__ap_start ap_done=PE_wrapper_231__ap_done ap_idle=PE_wrapper_231__ap_idle ap_ready=PE_wrapper_231__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_232__ap_start ap_done=PE_wrapper_232__ap_done ap_idle=PE_wrapper_232__ap_idle ap_ready=PE_wrapper_232__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_233__ap_start ap_done=PE_wrapper_233__ap_done ap_idle=PE_wrapper_233__ap_idle ap_ready=PE_wrapper_233__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_234__ap_start ap_done=PE_wrapper_234__ap_done ap_idle=PE_wrapper_234__ap_idle ap_ready=PE_wrapper_234__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_235__ap_start ap_done=PE_wrapper_235__ap_done ap_idle=PE_wrapper_235__ap_idle ap_ready=PE_wrapper_235__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_236__ap_start ap_done=PE_wrapper_236__ap_done ap_idle=PE_wrapper_236__ap_idle ap_ready=PE_wrapper_236__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_237__ap_start ap_done=PE_wrapper_237__ap_done ap_idle=PE_wrapper_237__ap_idle ap_ready=PE_wrapper_237__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_238__ap_start ap_done=PE_wrapper_238__ap_done ap_idle=PE_wrapper_238__ap_idle ap_ready=PE_wrapper_238__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_239__ap_start ap_done=PE_wrapper_239__ap_done ap_idle=PE_wrapper_239__ap_idle ap_ready=PE_wrapper_239__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_240__ap_start ap_done=PE_wrapper_240__ap_done ap_idle=PE_wrapper_240__ap_idle ap_ready=PE_wrapper_240__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_241__ap_start ap_done=PE_wrapper_241__ap_done ap_idle=PE_wrapper_241__ap_idle ap_ready=PE_wrapper_241__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_242__ap_start ap_done=PE_wrapper_242__ap_done ap_idle=PE_wrapper_242__ap_idle ap_ready=PE_wrapper_242__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_243__ap_start ap_done=PE_wrapper_243__ap_done ap_idle=PE_wrapper_243__ap_idle ap_ready=PE_wrapper_243__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_244__ap_start ap_done=PE_wrapper_244__ap_done ap_idle=PE_wrapper_244__ap_idle ap_ready=PE_wrapper_244__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_245__ap_start ap_done=PE_wrapper_245__ap_done ap_idle=PE_wrapper_245__ap_idle ap_ready=PE_wrapper_245__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_246__ap_start ap_done=PE_wrapper_246__ap_done ap_idle=PE_wrapper_246__ap_idle ap_ready=PE_wrapper_246__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_247__ap_start ap_done=PE_wrapper_247__ap_done ap_idle=PE_wrapper_247__ap_idle ap_ready=PE_wrapper_247__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_248__ap_start ap_done=PE_wrapper_248__ap_done ap_idle=PE_wrapper_248__ap_idle ap_ready=PE_wrapper_248__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_249__ap_start ap_done=PE_wrapper_249__ap_done ap_idle=PE_wrapper_249__ap_idle ap_ready=PE_wrapper_249__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_250__ap_start ap_done=PE_wrapper_250__ap_done ap_idle=PE_wrapper_250__ap_idle ap_ready=PE_wrapper_250__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_251__ap_start ap_done=PE_wrapper_251__ap_done ap_idle=PE_wrapper_251__ap_idle ap_ready=PE_wrapper_251__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_252__ap_start ap_done=PE_wrapper_252__ap_done ap_idle=PE_wrapper_252__ap_idle ap_ready=PE_wrapper_252__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_253__ap_start ap_done=PE_wrapper_253__ap_done ap_idle=PE_wrapper_253__ap_idle ap_ready=PE_wrapper_253__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_254__ap_start ap_done=PE_wrapper_254__ap_done ap_idle=PE_wrapper_254__ap_idle ap_ready=PE_wrapper_254__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_255__ap_start ap_done=PE_wrapper_255__ap_done ap_idle=PE_wrapper_255__ap_idle ap_ready=PE_wrapper_255__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_256__ap_start ap_done=PE_wrapper_256__ap_done ap_idle=PE_wrapper_256__ap_idle ap_ready=PE_wrapper_256__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_257__ap_start ap_done=PE_wrapper_257__ap_done ap_idle=PE_wrapper_257__ap_idle ap_ready=PE_wrapper_257__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_258__ap_start ap_done=PE_wrapper_258__ap_done ap_idle=PE_wrapper_258__ap_idle ap_ready=PE_wrapper_258__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_259__ap_start ap_done=PE_wrapper_259__ap_done ap_idle=PE_wrapper_259__ap_idle ap_ready=PE_wrapper_259__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_260__ap_start ap_done=PE_wrapper_260__ap_done ap_idle=PE_wrapper_260__ap_idle ap_ready=PE_wrapper_260__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_261__ap_start ap_done=PE_wrapper_261__ap_done ap_idle=PE_wrapper_261__ap_idle ap_ready=PE_wrapper_261__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_262__ap_start ap_done=PE_wrapper_262__ap_done ap_idle=PE_wrapper_262__ap_idle ap_ready=PE_wrapper_262__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_263__ap_start ap_done=PE_wrapper_263__ap_done ap_idle=PE_wrapper_263__ap_idle ap_ready=PE_wrapper_263__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_264__ap_start ap_done=PE_wrapper_264__ap_done ap_idle=PE_wrapper_264__ap_idle ap_ready=PE_wrapper_264__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_265__ap_start ap_done=PE_wrapper_265__ap_done ap_idle=PE_wrapper_265__ap_idle ap_ready=PE_wrapper_265__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_266__ap_start ap_done=PE_wrapper_266__ap_done ap_idle=PE_wrapper_266__ap_idle ap_ready=PE_wrapper_266__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_267__ap_start ap_done=PE_wrapper_267__ap_done ap_idle=PE_wrapper_267__ap_idle ap_ready=PE_wrapper_267__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_268__ap_start ap_done=PE_wrapper_268__ap_done ap_idle=PE_wrapper_268__ap_idle ap_ready=PE_wrapper_268__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_269__ap_start ap_done=PE_wrapper_269__ap_done ap_idle=PE_wrapper_269__ap_idle ap_ready=PE_wrapper_269__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_270__ap_start ap_done=PE_wrapper_270__ap_done ap_idle=PE_wrapper_270__ap_idle ap_ready=PE_wrapper_270__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_271__ap_start ap_done=PE_wrapper_271__ap_done ap_idle=PE_wrapper_271__ap_idle ap_ready=PE_wrapper_271__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_272__ap_start ap_done=PE_wrapper_272__ap_done ap_idle=PE_wrapper_272__ap_idle ap_ready=PE_wrapper_272__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_273__ap_start ap_done=PE_wrapper_273__ap_done ap_idle=PE_wrapper_273__ap_idle ap_ready=PE_wrapper_273__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_274__ap_start ap_done=PE_wrapper_274__ap_done ap_idle=PE_wrapper_274__ap_idle ap_ready=PE_wrapper_274__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_275__ap_start ap_done=PE_wrapper_275__ap_done ap_idle=PE_wrapper_275__ap_idle ap_ready=PE_wrapper_275__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_276__ap_start ap_done=PE_wrapper_276__ap_done ap_idle=PE_wrapper_276__ap_idle ap_ready=PE_wrapper_276__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_277__ap_start ap_done=PE_wrapper_277__ap_done ap_idle=PE_wrapper_277__ap_idle ap_ready=PE_wrapper_277__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_278__ap_start ap_done=PE_wrapper_278__ap_done ap_idle=PE_wrapper_278__ap_idle ap_ready=PE_wrapper_278__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_279__ap_start ap_done=PE_wrapper_279__ap_done ap_idle=PE_wrapper_279__ap_idle ap_ready=PE_wrapper_279__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_280__ap_start ap_done=PE_wrapper_280__ap_done ap_idle=PE_wrapper_280__ap_idle ap_ready=PE_wrapper_280__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_281__ap_start ap_done=PE_wrapper_281__ap_done ap_idle=PE_wrapper_281__ap_idle ap_ready=PE_wrapper_281__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_282__ap_start ap_done=PE_wrapper_282__ap_done ap_idle=PE_wrapper_282__ap_idle ap_ready=PE_wrapper_282__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_283__ap_start ap_done=PE_wrapper_283__ap_done ap_idle=PE_wrapper_283__ap_idle ap_ready=PE_wrapper_283__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_284__ap_start ap_done=PE_wrapper_284__ap_done ap_idle=PE_wrapper_284__ap_idle ap_ready=PE_wrapper_284__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_285__ap_start ap_done=PE_wrapper_285__ap_done ap_idle=PE_wrapper_285__ap_idle ap_ready=PE_wrapper_285__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_286__ap_start ap_done=PE_wrapper_286__ap_done ap_idle=PE_wrapper_286__ap_idle ap_ready=PE_wrapper_286__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_287__ap_start ap_done=PE_wrapper_287__ap_done ap_idle=PE_wrapper_287__ap_idle ap_ready=PE_wrapper_287__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_288__ap_start ap_done=PE_wrapper_288__ap_done ap_idle=PE_wrapper_288__ap_idle ap_ready=PE_wrapper_288__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_289__ap_start ap_done=PE_wrapper_289__ap_done ap_idle=PE_wrapper_289__ap_idle ap_ready=PE_wrapper_289__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_290__ap_start ap_done=PE_wrapper_290__ap_done ap_idle=PE_wrapper_290__ap_idle ap_ready=PE_wrapper_290__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_291__ap_start ap_done=PE_wrapper_291__ap_done ap_idle=PE_wrapper_291__ap_idle ap_ready=PE_wrapper_291__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_292__ap_start ap_done=PE_wrapper_292__ap_done ap_idle=PE_wrapper_292__ap_idle ap_ready=PE_wrapper_292__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_293__ap_start ap_done=PE_wrapper_293__ap_done ap_idle=PE_wrapper_293__ap_idle ap_ready=PE_wrapper_293__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_294__ap_start ap_done=PE_wrapper_294__ap_done ap_idle=PE_wrapper_294__ap_idle ap_ready=PE_wrapper_294__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_295__ap_start ap_done=PE_wrapper_295__ap_done ap_idle=PE_wrapper_295__ap_idle ap_ready=PE_wrapper_295__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_296__ap_start ap_done=PE_wrapper_296__ap_done ap_idle=PE_wrapper_296__ap_idle ap_ready=PE_wrapper_296__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_297__ap_start ap_done=PE_wrapper_297__ap_done ap_idle=PE_wrapper_297__ap_idle ap_ready=PE_wrapper_297__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_298__ap_start ap_done=PE_wrapper_298__ap_done ap_idle=PE_wrapper_298__ap_idle ap_ready=PE_wrapper_298__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_299__ap_start ap_done=PE_wrapper_299__ap_done ap_idle=PE_wrapper_299__ap_idle ap_ready=PE_wrapper_299__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_300__ap_start ap_done=PE_wrapper_300__ap_done ap_idle=PE_wrapper_300__ap_idle ap_ready=PE_wrapper_300__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_301__ap_start ap_done=PE_wrapper_301__ap_done ap_idle=PE_wrapper_301__ap_idle ap_ready=PE_wrapper_301__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_302__ap_start ap_done=PE_wrapper_302__ap_done ap_idle=PE_wrapper_302__ap_idle ap_ready=PE_wrapper_302__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_303__ap_start ap_done=PE_wrapper_303__ap_done ap_idle=PE_wrapper_303__ap_idle ap_ready=PE_wrapper_303__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_304__ap_start ap_done=PE_wrapper_304__ap_done ap_idle=PE_wrapper_304__ap_idle ap_ready=PE_wrapper_304__ap_ready
  // pragma RS ap-ctrl ap_start=PE_wrapper_305__ap_start ap_done=PE_wrapper_305__ap_done ap_idle=PE_wrapper_305__ap_idle ap_ready=PE_wrapper_305__ap_ready

  input ap_clk;
  input ap_rst_n;
  input ap_start;
  output ap_ready;
  output ap_done;
  output ap_idle;
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  output A_IO_L2_in_0__ap_start;
  input A_IO_L2_in_0__ap_ready;
  input A_IO_L2_in_0__ap_done;
  input A_IO_L2_in_0__ap_idle;
  output A_IO_L2_in_1__ap_start;
  input A_IO_L2_in_1__ap_ready;
  input A_IO_L2_in_1__ap_done;
  input A_IO_L2_in_1__ap_idle;
  output A_IO_L2_in_2__ap_start;
  input A_IO_L2_in_2__ap_ready;
  input A_IO_L2_in_2__ap_done;
  input A_IO_L2_in_2__ap_idle;
  output A_IO_L2_in_3__ap_start;
  input A_IO_L2_in_3__ap_ready;
  input A_IO_L2_in_3__ap_done;
  input A_IO_L2_in_3__ap_idle;
  output A_IO_L2_in_4__ap_start;
  input A_IO_L2_in_4__ap_ready;
  input A_IO_L2_in_4__ap_done;
  input A_IO_L2_in_4__ap_idle;
  output A_IO_L2_in_5__ap_start;
  input A_IO_L2_in_5__ap_ready;
  input A_IO_L2_in_5__ap_done;
  input A_IO_L2_in_5__ap_idle;
  output A_IO_L2_in_6__ap_start;
  input A_IO_L2_in_6__ap_ready;
  input A_IO_L2_in_6__ap_done;
  input A_IO_L2_in_6__ap_idle;
  output A_IO_L2_in_7__ap_start;
  input A_IO_L2_in_7__ap_ready;
  input A_IO_L2_in_7__ap_done;
  input A_IO_L2_in_7__ap_idle;
  output A_IO_L2_in_8__ap_start;
  input A_IO_L2_in_8__ap_ready;
  input A_IO_L2_in_8__ap_done;
  input A_IO_L2_in_8__ap_idle;
  output A_IO_L2_in_9__ap_start;
  input A_IO_L2_in_9__ap_ready;
  input A_IO_L2_in_9__ap_done;
  input A_IO_L2_in_9__ap_idle;
  output A_IO_L2_in_10__ap_start;
  input A_IO_L2_in_10__ap_ready;
  input A_IO_L2_in_10__ap_done;
  input A_IO_L2_in_10__ap_idle;
  output A_IO_L2_in_11__ap_start;
  input A_IO_L2_in_11__ap_ready;
  input A_IO_L2_in_11__ap_done;
  input A_IO_L2_in_11__ap_idle;
  output A_IO_L2_in_12__ap_start;
  input A_IO_L2_in_12__ap_ready;
  input A_IO_L2_in_12__ap_done;
  input A_IO_L2_in_12__ap_idle;
  output A_IO_L2_in_13__ap_start;
  input A_IO_L2_in_13__ap_ready;
  input A_IO_L2_in_13__ap_done;
  input A_IO_L2_in_13__ap_idle;
  output A_IO_L2_in_14__ap_start;
  input A_IO_L2_in_14__ap_ready;
  input A_IO_L2_in_14__ap_done;
  input A_IO_L2_in_14__ap_idle;
  output A_IO_L2_in_15__ap_start;
  input A_IO_L2_in_15__ap_ready;
  input A_IO_L2_in_15__ap_done;
  input A_IO_L2_in_15__ap_idle;
  output A_IO_L2_in_16__ap_start;
  input A_IO_L2_in_16__ap_ready;
  input A_IO_L2_in_16__ap_done;
  input A_IO_L2_in_16__ap_idle;
  output A_IO_L2_in_boundary_0__ap_start;
  input A_IO_L2_in_boundary_0__ap_ready;
  input A_IO_L2_in_boundary_0__ap_done;
  input A_IO_L2_in_boundary_0__ap_idle;
  output A_IO_L3_in_0__ap_start;
  input A_IO_L3_in_0__ap_ready;
  input A_IO_L3_in_0__ap_done;
  input A_IO_L3_in_0__ap_idle;
  output [63:0] A_IO_L3_in_serialize_0___A__q0;
  output A_IO_L3_in_serialize_0__ap_start;
  input A_IO_L3_in_serialize_0__ap_ready;
  input A_IO_L3_in_serialize_0__ap_done;
  input A_IO_L3_in_serialize_0__ap_idle;
  output A_PE_dummy_in_0__ap_start;
  input A_PE_dummy_in_0__ap_ready;
  input A_PE_dummy_in_0__ap_done;
  input A_PE_dummy_in_0__ap_idle;
  output A_PE_dummy_in_1__ap_start;
  input A_PE_dummy_in_1__ap_ready;
  input A_PE_dummy_in_1__ap_done;
  input A_PE_dummy_in_1__ap_idle;
  output A_PE_dummy_in_2__ap_start;
  input A_PE_dummy_in_2__ap_ready;
  input A_PE_dummy_in_2__ap_done;
  input A_PE_dummy_in_2__ap_idle;
  output A_PE_dummy_in_3__ap_start;
  input A_PE_dummy_in_3__ap_ready;
  input A_PE_dummy_in_3__ap_done;
  input A_PE_dummy_in_3__ap_idle;
  output A_PE_dummy_in_4__ap_start;
  input A_PE_dummy_in_4__ap_ready;
  input A_PE_dummy_in_4__ap_done;
  input A_PE_dummy_in_4__ap_idle;
  output A_PE_dummy_in_5__ap_start;
  input A_PE_dummy_in_5__ap_ready;
  input A_PE_dummy_in_5__ap_done;
  input A_PE_dummy_in_5__ap_idle;
  output A_PE_dummy_in_6__ap_start;
  input A_PE_dummy_in_6__ap_ready;
  input A_PE_dummy_in_6__ap_done;
  input A_PE_dummy_in_6__ap_idle;
  output A_PE_dummy_in_7__ap_start;
  input A_PE_dummy_in_7__ap_ready;
  input A_PE_dummy_in_7__ap_done;
  input A_PE_dummy_in_7__ap_idle;
  output A_PE_dummy_in_8__ap_start;
  input A_PE_dummy_in_8__ap_ready;
  input A_PE_dummy_in_8__ap_done;
  input A_PE_dummy_in_8__ap_idle;
  output A_PE_dummy_in_9__ap_start;
  input A_PE_dummy_in_9__ap_ready;
  input A_PE_dummy_in_9__ap_done;
  input A_PE_dummy_in_9__ap_idle;
  output A_PE_dummy_in_10__ap_start;
  input A_PE_dummy_in_10__ap_ready;
  input A_PE_dummy_in_10__ap_done;
  input A_PE_dummy_in_10__ap_idle;
  output A_PE_dummy_in_11__ap_start;
  input A_PE_dummy_in_11__ap_ready;
  input A_PE_dummy_in_11__ap_done;
  input A_PE_dummy_in_11__ap_idle;
  output A_PE_dummy_in_12__ap_start;
  input A_PE_dummy_in_12__ap_ready;
  input A_PE_dummy_in_12__ap_done;
  input A_PE_dummy_in_12__ap_idle;
  output A_PE_dummy_in_13__ap_start;
  input A_PE_dummy_in_13__ap_ready;
  input A_PE_dummy_in_13__ap_done;
  input A_PE_dummy_in_13__ap_idle;
  output A_PE_dummy_in_14__ap_start;
  input A_PE_dummy_in_14__ap_ready;
  input A_PE_dummy_in_14__ap_done;
  input A_PE_dummy_in_14__ap_idle;
  output A_PE_dummy_in_15__ap_start;
  input A_PE_dummy_in_15__ap_ready;
  input A_PE_dummy_in_15__ap_done;
  input A_PE_dummy_in_15__ap_idle;
  output A_PE_dummy_in_16__ap_start;
  input A_PE_dummy_in_16__ap_ready;
  input A_PE_dummy_in_16__ap_done;
  input A_PE_dummy_in_16__ap_idle;
  output A_PE_dummy_in_17__ap_start;
  input A_PE_dummy_in_17__ap_ready;
  input A_PE_dummy_in_17__ap_done;
  input A_PE_dummy_in_17__ap_idle;
  output B_IO_L2_in_0__ap_start;
  input B_IO_L2_in_0__ap_ready;
  input B_IO_L2_in_0__ap_done;
  input B_IO_L2_in_0__ap_idle;
  output B_IO_L2_in_1__ap_start;
  input B_IO_L2_in_1__ap_ready;
  input B_IO_L2_in_1__ap_done;
  input B_IO_L2_in_1__ap_idle;
  output B_IO_L2_in_2__ap_start;
  input B_IO_L2_in_2__ap_ready;
  input B_IO_L2_in_2__ap_done;
  input B_IO_L2_in_2__ap_idle;
  output B_IO_L2_in_3__ap_start;
  input B_IO_L2_in_3__ap_ready;
  input B_IO_L2_in_3__ap_done;
  input B_IO_L2_in_3__ap_idle;
  output B_IO_L2_in_4__ap_start;
  input B_IO_L2_in_4__ap_ready;
  input B_IO_L2_in_4__ap_done;
  input B_IO_L2_in_4__ap_idle;
  output B_IO_L2_in_5__ap_start;
  input B_IO_L2_in_5__ap_ready;
  input B_IO_L2_in_5__ap_done;
  input B_IO_L2_in_5__ap_idle;
  output B_IO_L2_in_6__ap_start;
  input B_IO_L2_in_6__ap_ready;
  input B_IO_L2_in_6__ap_done;
  input B_IO_L2_in_6__ap_idle;
  output B_IO_L2_in_7__ap_start;
  input B_IO_L2_in_7__ap_ready;
  input B_IO_L2_in_7__ap_done;
  input B_IO_L2_in_7__ap_idle;
  output B_IO_L2_in_8__ap_start;
  input B_IO_L2_in_8__ap_ready;
  input B_IO_L2_in_8__ap_done;
  input B_IO_L2_in_8__ap_idle;
  output B_IO_L2_in_9__ap_start;
  input B_IO_L2_in_9__ap_ready;
  input B_IO_L2_in_9__ap_done;
  input B_IO_L2_in_9__ap_idle;
  output B_IO_L2_in_10__ap_start;
  input B_IO_L2_in_10__ap_ready;
  input B_IO_L2_in_10__ap_done;
  input B_IO_L2_in_10__ap_idle;
  output B_IO_L2_in_11__ap_start;
  input B_IO_L2_in_11__ap_ready;
  input B_IO_L2_in_11__ap_done;
  input B_IO_L2_in_11__ap_idle;
  output B_IO_L2_in_12__ap_start;
  input B_IO_L2_in_12__ap_ready;
  input B_IO_L2_in_12__ap_done;
  input B_IO_L2_in_12__ap_idle;
  output B_IO_L2_in_13__ap_start;
  input B_IO_L2_in_13__ap_ready;
  input B_IO_L2_in_13__ap_done;
  input B_IO_L2_in_13__ap_idle;
  output B_IO_L2_in_14__ap_start;
  input B_IO_L2_in_14__ap_ready;
  input B_IO_L2_in_14__ap_done;
  input B_IO_L2_in_14__ap_idle;
  output B_IO_L2_in_15__ap_start;
  input B_IO_L2_in_15__ap_ready;
  input B_IO_L2_in_15__ap_done;
  input B_IO_L2_in_15__ap_idle;
  output B_IO_L2_in_boundary_0__ap_start;
  input B_IO_L2_in_boundary_0__ap_ready;
  input B_IO_L2_in_boundary_0__ap_done;
  input B_IO_L2_in_boundary_0__ap_idle;
  output B_IO_L3_in_0__ap_start;
  input B_IO_L3_in_0__ap_ready;
  input B_IO_L3_in_0__ap_done;
  input B_IO_L3_in_0__ap_idle;
  output [63:0] B_IO_L3_in_serialize_0___B__q0;
  output B_IO_L3_in_serialize_0__ap_start;
  input B_IO_L3_in_serialize_0__ap_ready;
  input B_IO_L3_in_serialize_0__ap_done;
  input B_IO_L3_in_serialize_0__ap_idle;
  output B_PE_dummy_in_0__ap_start;
  input B_PE_dummy_in_0__ap_ready;
  input B_PE_dummy_in_0__ap_done;
  input B_PE_dummy_in_0__ap_idle;
  output B_PE_dummy_in_1__ap_start;
  input B_PE_dummy_in_1__ap_ready;
  input B_PE_dummy_in_1__ap_done;
  input B_PE_dummy_in_1__ap_idle;
  output B_PE_dummy_in_2__ap_start;
  input B_PE_dummy_in_2__ap_ready;
  input B_PE_dummy_in_2__ap_done;
  input B_PE_dummy_in_2__ap_idle;
  output B_PE_dummy_in_3__ap_start;
  input B_PE_dummy_in_3__ap_ready;
  input B_PE_dummy_in_3__ap_done;
  input B_PE_dummy_in_3__ap_idle;
  output B_PE_dummy_in_4__ap_start;
  input B_PE_dummy_in_4__ap_ready;
  input B_PE_dummy_in_4__ap_done;
  input B_PE_dummy_in_4__ap_idle;
  output B_PE_dummy_in_5__ap_start;
  input B_PE_dummy_in_5__ap_ready;
  input B_PE_dummy_in_5__ap_done;
  input B_PE_dummy_in_5__ap_idle;
  output B_PE_dummy_in_6__ap_start;
  input B_PE_dummy_in_6__ap_ready;
  input B_PE_dummy_in_6__ap_done;
  input B_PE_dummy_in_6__ap_idle;
  output B_PE_dummy_in_7__ap_start;
  input B_PE_dummy_in_7__ap_ready;
  input B_PE_dummy_in_7__ap_done;
  input B_PE_dummy_in_7__ap_idle;
  output B_PE_dummy_in_8__ap_start;
  input B_PE_dummy_in_8__ap_ready;
  input B_PE_dummy_in_8__ap_done;
  input B_PE_dummy_in_8__ap_idle;
  output B_PE_dummy_in_9__ap_start;
  input B_PE_dummy_in_9__ap_ready;
  input B_PE_dummy_in_9__ap_done;
  input B_PE_dummy_in_9__ap_idle;
  output B_PE_dummy_in_10__ap_start;
  input B_PE_dummy_in_10__ap_ready;
  input B_PE_dummy_in_10__ap_done;
  input B_PE_dummy_in_10__ap_idle;
  output B_PE_dummy_in_11__ap_start;
  input B_PE_dummy_in_11__ap_ready;
  input B_PE_dummy_in_11__ap_done;
  input B_PE_dummy_in_11__ap_idle;
  output B_PE_dummy_in_12__ap_start;
  input B_PE_dummy_in_12__ap_ready;
  input B_PE_dummy_in_12__ap_done;
  input B_PE_dummy_in_12__ap_idle;
  output B_PE_dummy_in_13__ap_start;
  input B_PE_dummy_in_13__ap_ready;
  input B_PE_dummy_in_13__ap_done;
  input B_PE_dummy_in_13__ap_idle;
  output B_PE_dummy_in_14__ap_start;
  input B_PE_dummy_in_14__ap_ready;
  input B_PE_dummy_in_14__ap_done;
  input B_PE_dummy_in_14__ap_idle;
  output B_PE_dummy_in_15__ap_start;
  input B_PE_dummy_in_15__ap_ready;
  input B_PE_dummy_in_15__ap_done;
  input B_PE_dummy_in_15__ap_idle;
  output B_PE_dummy_in_16__ap_start;
  input B_PE_dummy_in_16__ap_ready;
  input B_PE_dummy_in_16__ap_done;
  input B_PE_dummy_in_16__ap_idle;
  output C_drain_IO_L1_out_boundary_wrapper_0__ap_start;
  input C_drain_IO_L1_out_boundary_wrapper_0__ap_ready;
  input C_drain_IO_L1_out_boundary_wrapper_0__ap_done;
  input C_drain_IO_L1_out_boundary_wrapper_0__ap_idle;
  output C_drain_IO_L1_out_boundary_wrapper_1__ap_start;
  input C_drain_IO_L1_out_boundary_wrapper_1__ap_ready;
  input C_drain_IO_L1_out_boundary_wrapper_1__ap_done;
  input C_drain_IO_L1_out_boundary_wrapper_1__ap_idle;
  output C_drain_IO_L1_out_boundary_wrapper_2__ap_start;
  input C_drain_IO_L1_out_boundary_wrapper_2__ap_ready;
  input C_drain_IO_L1_out_boundary_wrapper_2__ap_done;
  input C_drain_IO_L1_out_boundary_wrapper_2__ap_idle;
  output C_drain_IO_L1_out_boundary_wrapper_3__ap_start;
  input C_drain_IO_L1_out_boundary_wrapper_3__ap_ready;
  input C_drain_IO_L1_out_boundary_wrapper_3__ap_done;
  input C_drain_IO_L1_out_boundary_wrapper_3__ap_idle;
  output C_drain_IO_L1_out_boundary_wrapper_4__ap_start;
  input C_drain_IO_L1_out_boundary_wrapper_4__ap_ready;
  input C_drain_IO_L1_out_boundary_wrapper_4__ap_done;
  input C_drain_IO_L1_out_boundary_wrapper_4__ap_idle;
  output C_drain_IO_L1_out_boundary_wrapper_5__ap_start;
  input C_drain_IO_L1_out_boundary_wrapper_5__ap_ready;
  input C_drain_IO_L1_out_boundary_wrapper_5__ap_done;
  input C_drain_IO_L1_out_boundary_wrapper_5__ap_idle;
  output C_drain_IO_L1_out_boundary_wrapper_6__ap_start;
  input C_drain_IO_L1_out_boundary_wrapper_6__ap_ready;
  input C_drain_IO_L1_out_boundary_wrapper_6__ap_done;
  input C_drain_IO_L1_out_boundary_wrapper_6__ap_idle;
  output C_drain_IO_L1_out_boundary_wrapper_7__ap_start;
  input C_drain_IO_L1_out_boundary_wrapper_7__ap_ready;
  input C_drain_IO_L1_out_boundary_wrapper_7__ap_done;
  input C_drain_IO_L1_out_boundary_wrapper_7__ap_idle;
  output C_drain_IO_L1_out_boundary_wrapper_8__ap_start;
  input C_drain_IO_L1_out_boundary_wrapper_8__ap_ready;
  input C_drain_IO_L1_out_boundary_wrapper_8__ap_done;
  input C_drain_IO_L1_out_boundary_wrapper_8__ap_idle;
  output C_drain_IO_L1_out_boundary_wrapper_9__ap_start;
  input C_drain_IO_L1_out_boundary_wrapper_9__ap_ready;
  input C_drain_IO_L1_out_boundary_wrapper_9__ap_done;
  input C_drain_IO_L1_out_boundary_wrapper_9__ap_idle;
  output C_drain_IO_L1_out_boundary_wrapper_10__ap_start;
  input C_drain_IO_L1_out_boundary_wrapper_10__ap_ready;
  input C_drain_IO_L1_out_boundary_wrapper_10__ap_done;
  input C_drain_IO_L1_out_boundary_wrapper_10__ap_idle;
  output C_drain_IO_L1_out_boundary_wrapper_11__ap_start;
  input C_drain_IO_L1_out_boundary_wrapper_11__ap_ready;
  input C_drain_IO_L1_out_boundary_wrapper_11__ap_done;
  input C_drain_IO_L1_out_boundary_wrapper_11__ap_idle;
  output C_drain_IO_L1_out_boundary_wrapper_12__ap_start;
  input C_drain_IO_L1_out_boundary_wrapper_12__ap_ready;
  input C_drain_IO_L1_out_boundary_wrapper_12__ap_done;
  input C_drain_IO_L1_out_boundary_wrapper_12__ap_idle;
  output C_drain_IO_L1_out_boundary_wrapper_13__ap_start;
  input C_drain_IO_L1_out_boundary_wrapper_13__ap_ready;
  input C_drain_IO_L1_out_boundary_wrapper_13__ap_done;
  input C_drain_IO_L1_out_boundary_wrapper_13__ap_idle;
  output C_drain_IO_L1_out_boundary_wrapper_14__ap_start;
  input C_drain_IO_L1_out_boundary_wrapper_14__ap_ready;
  input C_drain_IO_L1_out_boundary_wrapper_14__ap_done;
  input C_drain_IO_L1_out_boundary_wrapper_14__ap_idle;
  output C_drain_IO_L1_out_boundary_wrapper_15__ap_start;
  input C_drain_IO_L1_out_boundary_wrapper_15__ap_ready;
  input C_drain_IO_L1_out_boundary_wrapper_15__ap_done;
  input C_drain_IO_L1_out_boundary_wrapper_15__ap_idle;
  output C_drain_IO_L1_out_boundary_wrapper_16__ap_start;
  input C_drain_IO_L1_out_boundary_wrapper_16__ap_ready;
  input C_drain_IO_L1_out_boundary_wrapper_16__ap_done;
  input C_drain_IO_L1_out_boundary_wrapper_16__ap_idle;
  output C_drain_IO_L1_out_wrapper_0__ap_start;
  input C_drain_IO_L1_out_wrapper_0__ap_ready;
  input C_drain_IO_L1_out_wrapper_0__ap_done;
  input C_drain_IO_L1_out_wrapper_0__ap_idle;
  output C_drain_IO_L1_out_wrapper_1__ap_start;
  input C_drain_IO_L1_out_wrapper_1__ap_ready;
  input C_drain_IO_L1_out_wrapper_1__ap_done;
  input C_drain_IO_L1_out_wrapper_1__ap_idle;
  output C_drain_IO_L1_out_wrapper_2__ap_start;
  input C_drain_IO_L1_out_wrapper_2__ap_ready;
  input C_drain_IO_L1_out_wrapper_2__ap_done;
  input C_drain_IO_L1_out_wrapper_2__ap_idle;
  output C_drain_IO_L1_out_wrapper_3__ap_start;
  input C_drain_IO_L1_out_wrapper_3__ap_ready;
  input C_drain_IO_L1_out_wrapper_3__ap_done;
  input C_drain_IO_L1_out_wrapper_3__ap_idle;
  output C_drain_IO_L1_out_wrapper_4__ap_start;
  input C_drain_IO_L1_out_wrapper_4__ap_ready;
  input C_drain_IO_L1_out_wrapper_4__ap_done;
  input C_drain_IO_L1_out_wrapper_4__ap_idle;
  output C_drain_IO_L1_out_wrapper_5__ap_start;
  input C_drain_IO_L1_out_wrapper_5__ap_ready;
  input C_drain_IO_L1_out_wrapper_5__ap_done;
  input C_drain_IO_L1_out_wrapper_5__ap_idle;
  output C_drain_IO_L1_out_wrapper_6__ap_start;
  input C_drain_IO_L1_out_wrapper_6__ap_ready;
  input C_drain_IO_L1_out_wrapper_6__ap_done;
  input C_drain_IO_L1_out_wrapper_6__ap_idle;
  output C_drain_IO_L1_out_wrapper_7__ap_start;
  input C_drain_IO_L1_out_wrapper_7__ap_ready;
  input C_drain_IO_L1_out_wrapper_7__ap_done;
  input C_drain_IO_L1_out_wrapper_7__ap_idle;
  output C_drain_IO_L1_out_wrapper_8__ap_start;
  input C_drain_IO_L1_out_wrapper_8__ap_ready;
  input C_drain_IO_L1_out_wrapper_8__ap_done;
  input C_drain_IO_L1_out_wrapper_8__ap_idle;
  output C_drain_IO_L1_out_wrapper_9__ap_start;
  input C_drain_IO_L1_out_wrapper_9__ap_ready;
  input C_drain_IO_L1_out_wrapper_9__ap_done;
  input C_drain_IO_L1_out_wrapper_9__ap_idle;
  output C_drain_IO_L1_out_wrapper_10__ap_start;
  input C_drain_IO_L1_out_wrapper_10__ap_ready;
  input C_drain_IO_L1_out_wrapper_10__ap_done;
  input C_drain_IO_L1_out_wrapper_10__ap_idle;
  output C_drain_IO_L1_out_wrapper_11__ap_start;
  input C_drain_IO_L1_out_wrapper_11__ap_ready;
  input C_drain_IO_L1_out_wrapper_11__ap_done;
  input C_drain_IO_L1_out_wrapper_11__ap_idle;
  output C_drain_IO_L1_out_wrapper_12__ap_start;
  input C_drain_IO_L1_out_wrapper_12__ap_ready;
  input C_drain_IO_L1_out_wrapper_12__ap_done;
  input C_drain_IO_L1_out_wrapper_12__ap_idle;
  output C_drain_IO_L1_out_wrapper_13__ap_start;
  input C_drain_IO_L1_out_wrapper_13__ap_ready;
  input C_drain_IO_L1_out_wrapper_13__ap_done;
  input C_drain_IO_L1_out_wrapper_13__ap_idle;
  output C_drain_IO_L1_out_wrapper_14__ap_start;
  input C_drain_IO_L1_out_wrapper_14__ap_ready;
  input C_drain_IO_L1_out_wrapper_14__ap_done;
  input C_drain_IO_L1_out_wrapper_14__ap_idle;
  output C_drain_IO_L1_out_wrapper_15__ap_start;
  input C_drain_IO_L1_out_wrapper_15__ap_ready;
  input C_drain_IO_L1_out_wrapper_15__ap_done;
  input C_drain_IO_L1_out_wrapper_15__ap_idle;
  output C_drain_IO_L1_out_wrapper_16__ap_start;
  input C_drain_IO_L1_out_wrapper_16__ap_ready;
  input C_drain_IO_L1_out_wrapper_16__ap_done;
  input C_drain_IO_L1_out_wrapper_16__ap_idle;
  output C_drain_IO_L1_out_wrapper_17__ap_start;
  input C_drain_IO_L1_out_wrapper_17__ap_ready;
  input C_drain_IO_L1_out_wrapper_17__ap_done;
  input C_drain_IO_L1_out_wrapper_17__ap_idle;
  output C_drain_IO_L1_out_wrapper_18__ap_start;
  input C_drain_IO_L1_out_wrapper_18__ap_ready;
  input C_drain_IO_L1_out_wrapper_18__ap_done;
  input C_drain_IO_L1_out_wrapper_18__ap_idle;
  output C_drain_IO_L1_out_wrapper_19__ap_start;
  input C_drain_IO_L1_out_wrapper_19__ap_ready;
  input C_drain_IO_L1_out_wrapper_19__ap_done;
  input C_drain_IO_L1_out_wrapper_19__ap_idle;
  output C_drain_IO_L1_out_wrapper_20__ap_start;
  input C_drain_IO_L1_out_wrapper_20__ap_ready;
  input C_drain_IO_L1_out_wrapper_20__ap_done;
  input C_drain_IO_L1_out_wrapper_20__ap_idle;
  output C_drain_IO_L1_out_wrapper_21__ap_start;
  input C_drain_IO_L1_out_wrapper_21__ap_ready;
  input C_drain_IO_L1_out_wrapper_21__ap_done;
  input C_drain_IO_L1_out_wrapper_21__ap_idle;
  output C_drain_IO_L1_out_wrapper_22__ap_start;
  input C_drain_IO_L1_out_wrapper_22__ap_ready;
  input C_drain_IO_L1_out_wrapper_22__ap_done;
  input C_drain_IO_L1_out_wrapper_22__ap_idle;
  output C_drain_IO_L1_out_wrapper_23__ap_start;
  input C_drain_IO_L1_out_wrapper_23__ap_ready;
  input C_drain_IO_L1_out_wrapper_23__ap_done;
  input C_drain_IO_L1_out_wrapper_23__ap_idle;
  output C_drain_IO_L1_out_wrapper_24__ap_start;
  input C_drain_IO_L1_out_wrapper_24__ap_ready;
  input C_drain_IO_L1_out_wrapper_24__ap_done;
  input C_drain_IO_L1_out_wrapper_24__ap_idle;
  output C_drain_IO_L1_out_wrapper_25__ap_start;
  input C_drain_IO_L1_out_wrapper_25__ap_ready;
  input C_drain_IO_L1_out_wrapper_25__ap_done;
  input C_drain_IO_L1_out_wrapper_25__ap_idle;
  output C_drain_IO_L1_out_wrapper_26__ap_start;
  input C_drain_IO_L1_out_wrapper_26__ap_ready;
  input C_drain_IO_L1_out_wrapper_26__ap_done;
  input C_drain_IO_L1_out_wrapper_26__ap_idle;
  output C_drain_IO_L1_out_wrapper_27__ap_start;
  input C_drain_IO_L1_out_wrapper_27__ap_ready;
  input C_drain_IO_L1_out_wrapper_27__ap_done;
  input C_drain_IO_L1_out_wrapper_27__ap_idle;
  output C_drain_IO_L1_out_wrapper_28__ap_start;
  input C_drain_IO_L1_out_wrapper_28__ap_ready;
  input C_drain_IO_L1_out_wrapper_28__ap_done;
  input C_drain_IO_L1_out_wrapper_28__ap_idle;
  output C_drain_IO_L1_out_wrapper_29__ap_start;
  input C_drain_IO_L1_out_wrapper_29__ap_ready;
  input C_drain_IO_L1_out_wrapper_29__ap_done;
  input C_drain_IO_L1_out_wrapper_29__ap_idle;
  output C_drain_IO_L1_out_wrapper_30__ap_start;
  input C_drain_IO_L1_out_wrapper_30__ap_ready;
  input C_drain_IO_L1_out_wrapper_30__ap_done;
  input C_drain_IO_L1_out_wrapper_30__ap_idle;
  output C_drain_IO_L1_out_wrapper_31__ap_start;
  input C_drain_IO_L1_out_wrapper_31__ap_ready;
  input C_drain_IO_L1_out_wrapper_31__ap_done;
  input C_drain_IO_L1_out_wrapper_31__ap_idle;
  output C_drain_IO_L1_out_wrapper_32__ap_start;
  input C_drain_IO_L1_out_wrapper_32__ap_ready;
  input C_drain_IO_L1_out_wrapper_32__ap_done;
  input C_drain_IO_L1_out_wrapper_32__ap_idle;
  output C_drain_IO_L1_out_wrapper_33__ap_start;
  input C_drain_IO_L1_out_wrapper_33__ap_ready;
  input C_drain_IO_L1_out_wrapper_33__ap_done;
  input C_drain_IO_L1_out_wrapper_33__ap_idle;
  output C_drain_IO_L1_out_wrapper_34__ap_start;
  input C_drain_IO_L1_out_wrapper_34__ap_ready;
  input C_drain_IO_L1_out_wrapper_34__ap_done;
  input C_drain_IO_L1_out_wrapper_34__ap_idle;
  output C_drain_IO_L1_out_wrapper_35__ap_start;
  input C_drain_IO_L1_out_wrapper_35__ap_ready;
  input C_drain_IO_L1_out_wrapper_35__ap_done;
  input C_drain_IO_L1_out_wrapper_35__ap_idle;
  output C_drain_IO_L1_out_wrapper_36__ap_start;
  input C_drain_IO_L1_out_wrapper_36__ap_ready;
  input C_drain_IO_L1_out_wrapper_36__ap_done;
  input C_drain_IO_L1_out_wrapper_36__ap_idle;
  output C_drain_IO_L1_out_wrapper_37__ap_start;
  input C_drain_IO_L1_out_wrapper_37__ap_ready;
  input C_drain_IO_L1_out_wrapper_37__ap_done;
  input C_drain_IO_L1_out_wrapper_37__ap_idle;
  output C_drain_IO_L1_out_wrapper_38__ap_start;
  input C_drain_IO_L1_out_wrapper_38__ap_ready;
  input C_drain_IO_L1_out_wrapper_38__ap_done;
  input C_drain_IO_L1_out_wrapper_38__ap_idle;
  output C_drain_IO_L1_out_wrapper_39__ap_start;
  input C_drain_IO_L1_out_wrapper_39__ap_ready;
  input C_drain_IO_L1_out_wrapper_39__ap_done;
  input C_drain_IO_L1_out_wrapper_39__ap_idle;
  output C_drain_IO_L1_out_wrapper_40__ap_start;
  input C_drain_IO_L1_out_wrapper_40__ap_ready;
  input C_drain_IO_L1_out_wrapper_40__ap_done;
  input C_drain_IO_L1_out_wrapper_40__ap_idle;
  output C_drain_IO_L1_out_wrapper_41__ap_start;
  input C_drain_IO_L1_out_wrapper_41__ap_ready;
  input C_drain_IO_L1_out_wrapper_41__ap_done;
  input C_drain_IO_L1_out_wrapper_41__ap_idle;
  output C_drain_IO_L1_out_wrapper_42__ap_start;
  input C_drain_IO_L1_out_wrapper_42__ap_ready;
  input C_drain_IO_L1_out_wrapper_42__ap_done;
  input C_drain_IO_L1_out_wrapper_42__ap_idle;
  output C_drain_IO_L1_out_wrapper_43__ap_start;
  input C_drain_IO_L1_out_wrapper_43__ap_ready;
  input C_drain_IO_L1_out_wrapper_43__ap_done;
  input C_drain_IO_L1_out_wrapper_43__ap_idle;
  output C_drain_IO_L1_out_wrapper_44__ap_start;
  input C_drain_IO_L1_out_wrapper_44__ap_ready;
  input C_drain_IO_L1_out_wrapper_44__ap_done;
  input C_drain_IO_L1_out_wrapper_44__ap_idle;
  output C_drain_IO_L1_out_wrapper_45__ap_start;
  input C_drain_IO_L1_out_wrapper_45__ap_ready;
  input C_drain_IO_L1_out_wrapper_45__ap_done;
  input C_drain_IO_L1_out_wrapper_45__ap_idle;
  output C_drain_IO_L1_out_wrapper_46__ap_start;
  input C_drain_IO_L1_out_wrapper_46__ap_ready;
  input C_drain_IO_L1_out_wrapper_46__ap_done;
  input C_drain_IO_L1_out_wrapper_46__ap_idle;
  output C_drain_IO_L1_out_wrapper_47__ap_start;
  input C_drain_IO_L1_out_wrapper_47__ap_ready;
  input C_drain_IO_L1_out_wrapper_47__ap_done;
  input C_drain_IO_L1_out_wrapper_47__ap_idle;
  output C_drain_IO_L1_out_wrapper_48__ap_start;
  input C_drain_IO_L1_out_wrapper_48__ap_ready;
  input C_drain_IO_L1_out_wrapper_48__ap_done;
  input C_drain_IO_L1_out_wrapper_48__ap_idle;
  output C_drain_IO_L1_out_wrapper_49__ap_start;
  input C_drain_IO_L1_out_wrapper_49__ap_ready;
  input C_drain_IO_L1_out_wrapper_49__ap_done;
  input C_drain_IO_L1_out_wrapper_49__ap_idle;
  output C_drain_IO_L1_out_wrapper_50__ap_start;
  input C_drain_IO_L1_out_wrapper_50__ap_ready;
  input C_drain_IO_L1_out_wrapper_50__ap_done;
  input C_drain_IO_L1_out_wrapper_50__ap_idle;
  output C_drain_IO_L1_out_wrapper_51__ap_start;
  input C_drain_IO_L1_out_wrapper_51__ap_ready;
  input C_drain_IO_L1_out_wrapper_51__ap_done;
  input C_drain_IO_L1_out_wrapper_51__ap_idle;
  output C_drain_IO_L1_out_wrapper_52__ap_start;
  input C_drain_IO_L1_out_wrapper_52__ap_ready;
  input C_drain_IO_L1_out_wrapper_52__ap_done;
  input C_drain_IO_L1_out_wrapper_52__ap_idle;
  output C_drain_IO_L1_out_wrapper_53__ap_start;
  input C_drain_IO_L1_out_wrapper_53__ap_ready;
  input C_drain_IO_L1_out_wrapper_53__ap_done;
  input C_drain_IO_L1_out_wrapper_53__ap_idle;
  output C_drain_IO_L1_out_wrapper_54__ap_start;
  input C_drain_IO_L1_out_wrapper_54__ap_ready;
  input C_drain_IO_L1_out_wrapper_54__ap_done;
  input C_drain_IO_L1_out_wrapper_54__ap_idle;
  output C_drain_IO_L1_out_wrapper_55__ap_start;
  input C_drain_IO_L1_out_wrapper_55__ap_ready;
  input C_drain_IO_L1_out_wrapper_55__ap_done;
  input C_drain_IO_L1_out_wrapper_55__ap_idle;
  output C_drain_IO_L1_out_wrapper_56__ap_start;
  input C_drain_IO_L1_out_wrapper_56__ap_ready;
  input C_drain_IO_L1_out_wrapper_56__ap_done;
  input C_drain_IO_L1_out_wrapper_56__ap_idle;
  output C_drain_IO_L1_out_wrapper_57__ap_start;
  input C_drain_IO_L1_out_wrapper_57__ap_ready;
  input C_drain_IO_L1_out_wrapper_57__ap_done;
  input C_drain_IO_L1_out_wrapper_57__ap_idle;
  output C_drain_IO_L1_out_wrapper_58__ap_start;
  input C_drain_IO_L1_out_wrapper_58__ap_ready;
  input C_drain_IO_L1_out_wrapper_58__ap_done;
  input C_drain_IO_L1_out_wrapper_58__ap_idle;
  output C_drain_IO_L1_out_wrapper_59__ap_start;
  input C_drain_IO_L1_out_wrapper_59__ap_ready;
  input C_drain_IO_L1_out_wrapper_59__ap_done;
  input C_drain_IO_L1_out_wrapper_59__ap_idle;
  output C_drain_IO_L1_out_wrapper_60__ap_start;
  input C_drain_IO_L1_out_wrapper_60__ap_ready;
  input C_drain_IO_L1_out_wrapper_60__ap_done;
  input C_drain_IO_L1_out_wrapper_60__ap_idle;
  output C_drain_IO_L1_out_wrapper_61__ap_start;
  input C_drain_IO_L1_out_wrapper_61__ap_ready;
  input C_drain_IO_L1_out_wrapper_61__ap_done;
  input C_drain_IO_L1_out_wrapper_61__ap_idle;
  output C_drain_IO_L1_out_wrapper_62__ap_start;
  input C_drain_IO_L1_out_wrapper_62__ap_ready;
  input C_drain_IO_L1_out_wrapper_62__ap_done;
  input C_drain_IO_L1_out_wrapper_62__ap_idle;
  output C_drain_IO_L1_out_wrapper_63__ap_start;
  input C_drain_IO_L1_out_wrapper_63__ap_ready;
  input C_drain_IO_L1_out_wrapper_63__ap_done;
  input C_drain_IO_L1_out_wrapper_63__ap_idle;
  output C_drain_IO_L1_out_wrapper_64__ap_start;
  input C_drain_IO_L1_out_wrapper_64__ap_ready;
  input C_drain_IO_L1_out_wrapper_64__ap_done;
  input C_drain_IO_L1_out_wrapper_64__ap_idle;
  output C_drain_IO_L1_out_wrapper_65__ap_start;
  input C_drain_IO_L1_out_wrapper_65__ap_ready;
  input C_drain_IO_L1_out_wrapper_65__ap_done;
  input C_drain_IO_L1_out_wrapper_65__ap_idle;
  output C_drain_IO_L1_out_wrapper_66__ap_start;
  input C_drain_IO_L1_out_wrapper_66__ap_ready;
  input C_drain_IO_L1_out_wrapper_66__ap_done;
  input C_drain_IO_L1_out_wrapper_66__ap_idle;
  output C_drain_IO_L1_out_wrapper_67__ap_start;
  input C_drain_IO_L1_out_wrapper_67__ap_ready;
  input C_drain_IO_L1_out_wrapper_67__ap_done;
  input C_drain_IO_L1_out_wrapper_67__ap_idle;
  output C_drain_IO_L1_out_wrapper_68__ap_start;
  input C_drain_IO_L1_out_wrapper_68__ap_ready;
  input C_drain_IO_L1_out_wrapper_68__ap_done;
  input C_drain_IO_L1_out_wrapper_68__ap_idle;
  output C_drain_IO_L1_out_wrapper_69__ap_start;
  input C_drain_IO_L1_out_wrapper_69__ap_ready;
  input C_drain_IO_L1_out_wrapper_69__ap_done;
  input C_drain_IO_L1_out_wrapper_69__ap_idle;
  output C_drain_IO_L1_out_wrapper_70__ap_start;
  input C_drain_IO_L1_out_wrapper_70__ap_ready;
  input C_drain_IO_L1_out_wrapper_70__ap_done;
  input C_drain_IO_L1_out_wrapper_70__ap_idle;
  output C_drain_IO_L1_out_wrapper_71__ap_start;
  input C_drain_IO_L1_out_wrapper_71__ap_ready;
  input C_drain_IO_L1_out_wrapper_71__ap_done;
  input C_drain_IO_L1_out_wrapper_71__ap_idle;
  output C_drain_IO_L1_out_wrapper_72__ap_start;
  input C_drain_IO_L1_out_wrapper_72__ap_ready;
  input C_drain_IO_L1_out_wrapper_72__ap_done;
  input C_drain_IO_L1_out_wrapper_72__ap_idle;
  output C_drain_IO_L1_out_wrapper_73__ap_start;
  input C_drain_IO_L1_out_wrapper_73__ap_ready;
  input C_drain_IO_L1_out_wrapper_73__ap_done;
  input C_drain_IO_L1_out_wrapper_73__ap_idle;
  output C_drain_IO_L1_out_wrapper_74__ap_start;
  input C_drain_IO_L1_out_wrapper_74__ap_ready;
  input C_drain_IO_L1_out_wrapper_74__ap_done;
  input C_drain_IO_L1_out_wrapper_74__ap_idle;
  output C_drain_IO_L1_out_wrapper_75__ap_start;
  input C_drain_IO_L1_out_wrapper_75__ap_ready;
  input C_drain_IO_L1_out_wrapper_75__ap_done;
  input C_drain_IO_L1_out_wrapper_75__ap_idle;
  output C_drain_IO_L1_out_wrapper_76__ap_start;
  input C_drain_IO_L1_out_wrapper_76__ap_ready;
  input C_drain_IO_L1_out_wrapper_76__ap_done;
  input C_drain_IO_L1_out_wrapper_76__ap_idle;
  output C_drain_IO_L1_out_wrapper_77__ap_start;
  input C_drain_IO_L1_out_wrapper_77__ap_ready;
  input C_drain_IO_L1_out_wrapper_77__ap_done;
  input C_drain_IO_L1_out_wrapper_77__ap_idle;
  output C_drain_IO_L1_out_wrapper_78__ap_start;
  input C_drain_IO_L1_out_wrapper_78__ap_ready;
  input C_drain_IO_L1_out_wrapper_78__ap_done;
  input C_drain_IO_L1_out_wrapper_78__ap_idle;
  output C_drain_IO_L1_out_wrapper_79__ap_start;
  input C_drain_IO_L1_out_wrapper_79__ap_ready;
  input C_drain_IO_L1_out_wrapper_79__ap_done;
  input C_drain_IO_L1_out_wrapper_79__ap_idle;
  output C_drain_IO_L1_out_wrapper_80__ap_start;
  input C_drain_IO_L1_out_wrapper_80__ap_ready;
  input C_drain_IO_L1_out_wrapper_80__ap_done;
  input C_drain_IO_L1_out_wrapper_80__ap_idle;
  output C_drain_IO_L1_out_wrapper_81__ap_start;
  input C_drain_IO_L1_out_wrapper_81__ap_ready;
  input C_drain_IO_L1_out_wrapper_81__ap_done;
  input C_drain_IO_L1_out_wrapper_81__ap_idle;
  output C_drain_IO_L1_out_wrapper_82__ap_start;
  input C_drain_IO_L1_out_wrapper_82__ap_ready;
  input C_drain_IO_L1_out_wrapper_82__ap_done;
  input C_drain_IO_L1_out_wrapper_82__ap_idle;
  output C_drain_IO_L1_out_wrapper_83__ap_start;
  input C_drain_IO_L1_out_wrapper_83__ap_ready;
  input C_drain_IO_L1_out_wrapper_83__ap_done;
  input C_drain_IO_L1_out_wrapper_83__ap_idle;
  output C_drain_IO_L1_out_wrapper_84__ap_start;
  input C_drain_IO_L1_out_wrapper_84__ap_ready;
  input C_drain_IO_L1_out_wrapper_84__ap_done;
  input C_drain_IO_L1_out_wrapper_84__ap_idle;
  output C_drain_IO_L1_out_wrapper_85__ap_start;
  input C_drain_IO_L1_out_wrapper_85__ap_ready;
  input C_drain_IO_L1_out_wrapper_85__ap_done;
  input C_drain_IO_L1_out_wrapper_85__ap_idle;
  output C_drain_IO_L1_out_wrapper_86__ap_start;
  input C_drain_IO_L1_out_wrapper_86__ap_ready;
  input C_drain_IO_L1_out_wrapper_86__ap_done;
  input C_drain_IO_L1_out_wrapper_86__ap_idle;
  output C_drain_IO_L1_out_wrapper_87__ap_start;
  input C_drain_IO_L1_out_wrapper_87__ap_ready;
  input C_drain_IO_L1_out_wrapper_87__ap_done;
  input C_drain_IO_L1_out_wrapper_87__ap_idle;
  output C_drain_IO_L1_out_wrapper_88__ap_start;
  input C_drain_IO_L1_out_wrapper_88__ap_ready;
  input C_drain_IO_L1_out_wrapper_88__ap_done;
  input C_drain_IO_L1_out_wrapper_88__ap_idle;
  output C_drain_IO_L1_out_wrapper_89__ap_start;
  input C_drain_IO_L1_out_wrapper_89__ap_ready;
  input C_drain_IO_L1_out_wrapper_89__ap_done;
  input C_drain_IO_L1_out_wrapper_89__ap_idle;
  output C_drain_IO_L1_out_wrapper_90__ap_start;
  input C_drain_IO_L1_out_wrapper_90__ap_ready;
  input C_drain_IO_L1_out_wrapper_90__ap_done;
  input C_drain_IO_L1_out_wrapper_90__ap_idle;
  output C_drain_IO_L1_out_wrapper_91__ap_start;
  input C_drain_IO_L1_out_wrapper_91__ap_ready;
  input C_drain_IO_L1_out_wrapper_91__ap_done;
  input C_drain_IO_L1_out_wrapper_91__ap_idle;
  output C_drain_IO_L1_out_wrapper_92__ap_start;
  input C_drain_IO_L1_out_wrapper_92__ap_ready;
  input C_drain_IO_L1_out_wrapper_92__ap_done;
  input C_drain_IO_L1_out_wrapper_92__ap_idle;
  output C_drain_IO_L1_out_wrapper_93__ap_start;
  input C_drain_IO_L1_out_wrapper_93__ap_ready;
  input C_drain_IO_L1_out_wrapper_93__ap_done;
  input C_drain_IO_L1_out_wrapper_93__ap_idle;
  output C_drain_IO_L1_out_wrapper_94__ap_start;
  input C_drain_IO_L1_out_wrapper_94__ap_ready;
  input C_drain_IO_L1_out_wrapper_94__ap_done;
  input C_drain_IO_L1_out_wrapper_94__ap_idle;
  output C_drain_IO_L1_out_wrapper_95__ap_start;
  input C_drain_IO_L1_out_wrapper_95__ap_ready;
  input C_drain_IO_L1_out_wrapper_95__ap_done;
  input C_drain_IO_L1_out_wrapper_95__ap_idle;
  output C_drain_IO_L1_out_wrapper_96__ap_start;
  input C_drain_IO_L1_out_wrapper_96__ap_ready;
  input C_drain_IO_L1_out_wrapper_96__ap_done;
  input C_drain_IO_L1_out_wrapper_96__ap_idle;
  output C_drain_IO_L1_out_wrapper_97__ap_start;
  input C_drain_IO_L1_out_wrapper_97__ap_ready;
  input C_drain_IO_L1_out_wrapper_97__ap_done;
  input C_drain_IO_L1_out_wrapper_97__ap_idle;
  output C_drain_IO_L1_out_wrapper_98__ap_start;
  input C_drain_IO_L1_out_wrapper_98__ap_ready;
  input C_drain_IO_L1_out_wrapper_98__ap_done;
  input C_drain_IO_L1_out_wrapper_98__ap_idle;
  output C_drain_IO_L1_out_wrapper_99__ap_start;
  input C_drain_IO_L1_out_wrapper_99__ap_ready;
  input C_drain_IO_L1_out_wrapper_99__ap_done;
  input C_drain_IO_L1_out_wrapper_99__ap_idle;
  output C_drain_IO_L1_out_wrapper_100__ap_start;
  input C_drain_IO_L1_out_wrapper_100__ap_ready;
  input C_drain_IO_L1_out_wrapper_100__ap_done;
  input C_drain_IO_L1_out_wrapper_100__ap_idle;
  output C_drain_IO_L1_out_wrapper_101__ap_start;
  input C_drain_IO_L1_out_wrapper_101__ap_ready;
  input C_drain_IO_L1_out_wrapper_101__ap_done;
  input C_drain_IO_L1_out_wrapper_101__ap_idle;
  output C_drain_IO_L1_out_wrapper_102__ap_start;
  input C_drain_IO_L1_out_wrapper_102__ap_ready;
  input C_drain_IO_L1_out_wrapper_102__ap_done;
  input C_drain_IO_L1_out_wrapper_102__ap_idle;
  output C_drain_IO_L1_out_wrapper_103__ap_start;
  input C_drain_IO_L1_out_wrapper_103__ap_ready;
  input C_drain_IO_L1_out_wrapper_103__ap_done;
  input C_drain_IO_L1_out_wrapper_103__ap_idle;
  output C_drain_IO_L1_out_wrapper_104__ap_start;
  input C_drain_IO_L1_out_wrapper_104__ap_ready;
  input C_drain_IO_L1_out_wrapper_104__ap_done;
  input C_drain_IO_L1_out_wrapper_104__ap_idle;
  output C_drain_IO_L1_out_wrapper_105__ap_start;
  input C_drain_IO_L1_out_wrapper_105__ap_ready;
  input C_drain_IO_L1_out_wrapper_105__ap_done;
  input C_drain_IO_L1_out_wrapper_105__ap_idle;
  output C_drain_IO_L1_out_wrapper_106__ap_start;
  input C_drain_IO_L1_out_wrapper_106__ap_ready;
  input C_drain_IO_L1_out_wrapper_106__ap_done;
  input C_drain_IO_L1_out_wrapper_106__ap_idle;
  output C_drain_IO_L1_out_wrapper_107__ap_start;
  input C_drain_IO_L1_out_wrapper_107__ap_ready;
  input C_drain_IO_L1_out_wrapper_107__ap_done;
  input C_drain_IO_L1_out_wrapper_107__ap_idle;
  output C_drain_IO_L1_out_wrapper_108__ap_start;
  input C_drain_IO_L1_out_wrapper_108__ap_ready;
  input C_drain_IO_L1_out_wrapper_108__ap_done;
  input C_drain_IO_L1_out_wrapper_108__ap_idle;
  output C_drain_IO_L1_out_wrapper_109__ap_start;
  input C_drain_IO_L1_out_wrapper_109__ap_ready;
  input C_drain_IO_L1_out_wrapper_109__ap_done;
  input C_drain_IO_L1_out_wrapper_109__ap_idle;
  output C_drain_IO_L1_out_wrapper_110__ap_start;
  input C_drain_IO_L1_out_wrapper_110__ap_ready;
  input C_drain_IO_L1_out_wrapper_110__ap_done;
  input C_drain_IO_L1_out_wrapper_110__ap_idle;
  output C_drain_IO_L1_out_wrapper_111__ap_start;
  input C_drain_IO_L1_out_wrapper_111__ap_ready;
  input C_drain_IO_L1_out_wrapper_111__ap_done;
  input C_drain_IO_L1_out_wrapper_111__ap_idle;
  output C_drain_IO_L1_out_wrapper_112__ap_start;
  input C_drain_IO_L1_out_wrapper_112__ap_ready;
  input C_drain_IO_L1_out_wrapper_112__ap_done;
  input C_drain_IO_L1_out_wrapper_112__ap_idle;
  output C_drain_IO_L1_out_wrapper_113__ap_start;
  input C_drain_IO_L1_out_wrapper_113__ap_ready;
  input C_drain_IO_L1_out_wrapper_113__ap_done;
  input C_drain_IO_L1_out_wrapper_113__ap_idle;
  output C_drain_IO_L1_out_wrapper_114__ap_start;
  input C_drain_IO_L1_out_wrapper_114__ap_ready;
  input C_drain_IO_L1_out_wrapper_114__ap_done;
  input C_drain_IO_L1_out_wrapper_114__ap_idle;
  output C_drain_IO_L1_out_wrapper_115__ap_start;
  input C_drain_IO_L1_out_wrapper_115__ap_ready;
  input C_drain_IO_L1_out_wrapper_115__ap_done;
  input C_drain_IO_L1_out_wrapper_115__ap_idle;
  output C_drain_IO_L1_out_wrapper_116__ap_start;
  input C_drain_IO_L1_out_wrapper_116__ap_ready;
  input C_drain_IO_L1_out_wrapper_116__ap_done;
  input C_drain_IO_L1_out_wrapper_116__ap_idle;
  output C_drain_IO_L1_out_wrapper_117__ap_start;
  input C_drain_IO_L1_out_wrapper_117__ap_ready;
  input C_drain_IO_L1_out_wrapper_117__ap_done;
  input C_drain_IO_L1_out_wrapper_117__ap_idle;
  output C_drain_IO_L1_out_wrapper_118__ap_start;
  input C_drain_IO_L1_out_wrapper_118__ap_ready;
  input C_drain_IO_L1_out_wrapper_118__ap_done;
  input C_drain_IO_L1_out_wrapper_118__ap_idle;
  output C_drain_IO_L1_out_wrapper_119__ap_start;
  input C_drain_IO_L1_out_wrapper_119__ap_ready;
  input C_drain_IO_L1_out_wrapper_119__ap_done;
  input C_drain_IO_L1_out_wrapper_119__ap_idle;
  output C_drain_IO_L1_out_wrapper_120__ap_start;
  input C_drain_IO_L1_out_wrapper_120__ap_ready;
  input C_drain_IO_L1_out_wrapper_120__ap_done;
  input C_drain_IO_L1_out_wrapper_120__ap_idle;
  output C_drain_IO_L1_out_wrapper_121__ap_start;
  input C_drain_IO_L1_out_wrapper_121__ap_ready;
  input C_drain_IO_L1_out_wrapper_121__ap_done;
  input C_drain_IO_L1_out_wrapper_121__ap_idle;
  output C_drain_IO_L1_out_wrapper_122__ap_start;
  input C_drain_IO_L1_out_wrapper_122__ap_ready;
  input C_drain_IO_L1_out_wrapper_122__ap_done;
  input C_drain_IO_L1_out_wrapper_122__ap_idle;
  output C_drain_IO_L1_out_wrapper_123__ap_start;
  input C_drain_IO_L1_out_wrapper_123__ap_ready;
  input C_drain_IO_L1_out_wrapper_123__ap_done;
  input C_drain_IO_L1_out_wrapper_123__ap_idle;
  output C_drain_IO_L1_out_wrapper_124__ap_start;
  input C_drain_IO_L1_out_wrapper_124__ap_ready;
  input C_drain_IO_L1_out_wrapper_124__ap_done;
  input C_drain_IO_L1_out_wrapper_124__ap_idle;
  output C_drain_IO_L1_out_wrapper_125__ap_start;
  input C_drain_IO_L1_out_wrapper_125__ap_ready;
  input C_drain_IO_L1_out_wrapper_125__ap_done;
  input C_drain_IO_L1_out_wrapper_125__ap_idle;
  output C_drain_IO_L1_out_wrapper_126__ap_start;
  input C_drain_IO_L1_out_wrapper_126__ap_ready;
  input C_drain_IO_L1_out_wrapper_126__ap_done;
  input C_drain_IO_L1_out_wrapper_126__ap_idle;
  output C_drain_IO_L1_out_wrapper_127__ap_start;
  input C_drain_IO_L1_out_wrapper_127__ap_ready;
  input C_drain_IO_L1_out_wrapper_127__ap_done;
  input C_drain_IO_L1_out_wrapper_127__ap_idle;
  output C_drain_IO_L1_out_wrapper_128__ap_start;
  input C_drain_IO_L1_out_wrapper_128__ap_ready;
  input C_drain_IO_L1_out_wrapper_128__ap_done;
  input C_drain_IO_L1_out_wrapper_128__ap_idle;
  output C_drain_IO_L1_out_wrapper_129__ap_start;
  input C_drain_IO_L1_out_wrapper_129__ap_ready;
  input C_drain_IO_L1_out_wrapper_129__ap_done;
  input C_drain_IO_L1_out_wrapper_129__ap_idle;
  output C_drain_IO_L1_out_wrapper_130__ap_start;
  input C_drain_IO_L1_out_wrapper_130__ap_ready;
  input C_drain_IO_L1_out_wrapper_130__ap_done;
  input C_drain_IO_L1_out_wrapper_130__ap_idle;
  output C_drain_IO_L1_out_wrapper_131__ap_start;
  input C_drain_IO_L1_out_wrapper_131__ap_ready;
  input C_drain_IO_L1_out_wrapper_131__ap_done;
  input C_drain_IO_L1_out_wrapper_131__ap_idle;
  output C_drain_IO_L1_out_wrapper_132__ap_start;
  input C_drain_IO_L1_out_wrapper_132__ap_ready;
  input C_drain_IO_L1_out_wrapper_132__ap_done;
  input C_drain_IO_L1_out_wrapper_132__ap_idle;
  output C_drain_IO_L1_out_wrapper_133__ap_start;
  input C_drain_IO_L1_out_wrapper_133__ap_ready;
  input C_drain_IO_L1_out_wrapper_133__ap_done;
  input C_drain_IO_L1_out_wrapper_133__ap_idle;
  output C_drain_IO_L1_out_wrapper_134__ap_start;
  input C_drain_IO_L1_out_wrapper_134__ap_ready;
  input C_drain_IO_L1_out_wrapper_134__ap_done;
  input C_drain_IO_L1_out_wrapper_134__ap_idle;
  output C_drain_IO_L1_out_wrapper_135__ap_start;
  input C_drain_IO_L1_out_wrapper_135__ap_ready;
  input C_drain_IO_L1_out_wrapper_135__ap_done;
  input C_drain_IO_L1_out_wrapper_135__ap_idle;
  output C_drain_IO_L1_out_wrapper_136__ap_start;
  input C_drain_IO_L1_out_wrapper_136__ap_ready;
  input C_drain_IO_L1_out_wrapper_136__ap_done;
  input C_drain_IO_L1_out_wrapper_136__ap_idle;
  output C_drain_IO_L1_out_wrapper_137__ap_start;
  input C_drain_IO_L1_out_wrapper_137__ap_ready;
  input C_drain_IO_L1_out_wrapper_137__ap_done;
  input C_drain_IO_L1_out_wrapper_137__ap_idle;
  output C_drain_IO_L1_out_wrapper_138__ap_start;
  input C_drain_IO_L1_out_wrapper_138__ap_ready;
  input C_drain_IO_L1_out_wrapper_138__ap_done;
  input C_drain_IO_L1_out_wrapper_138__ap_idle;
  output C_drain_IO_L1_out_wrapper_139__ap_start;
  input C_drain_IO_L1_out_wrapper_139__ap_ready;
  input C_drain_IO_L1_out_wrapper_139__ap_done;
  input C_drain_IO_L1_out_wrapper_139__ap_idle;
  output C_drain_IO_L1_out_wrapper_140__ap_start;
  input C_drain_IO_L1_out_wrapper_140__ap_ready;
  input C_drain_IO_L1_out_wrapper_140__ap_done;
  input C_drain_IO_L1_out_wrapper_140__ap_idle;
  output C_drain_IO_L1_out_wrapper_141__ap_start;
  input C_drain_IO_L1_out_wrapper_141__ap_ready;
  input C_drain_IO_L1_out_wrapper_141__ap_done;
  input C_drain_IO_L1_out_wrapper_141__ap_idle;
  output C_drain_IO_L1_out_wrapper_142__ap_start;
  input C_drain_IO_L1_out_wrapper_142__ap_ready;
  input C_drain_IO_L1_out_wrapper_142__ap_done;
  input C_drain_IO_L1_out_wrapper_142__ap_idle;
  output C_drain_IO_L1_out_wrapper_143__ap_start;
  input C_drain_IO_L1_out_wrapper_143__ap_ready;
  input C_drain_IO_L1_out_wrapper_143__ap_done;
  input C_drain_IO_L1_out_wrapper_143__ap_idle;
  output C_drain_IO_L1_out_wrapper_144__ap_start;
  input C_drain_IO_L1_out_wrapper_144__ap_ready;
  input C_drain_IO_L1_out_wrapper_144__ap_done;
  input C_drain_IO_L1_out_wrapper_144__ap_idle;
  output C_drain_IO_L1_out_wrapper_145__ap_start;
  input C_drain_IO_L1_out_wrapper_145__ap_ready;
  input C_drain_IO_L1_out_wrapper_145__ap_done;
  input C_drain_IO_L1_out_wrapper_145__ap_idle;
  output C_drain_IO_L1_out_wrapper_146__ap_start;
  input C_drain_IO_L1_out_wrapper_146__ap_ready;
  input C_drain_IO_L1_out_wrapper_146__ap_done;
  input C_drain_IO_L1_out_wrapper_146__ap_idle;
  output C_drain_IO_L1_out_wrapper_147__ap_start;
  input C_drain_IO_L1_out_wrapper_147__ap_ready;
  input C_drain_IO_L1_out_wrapper_147__ap_done;
  input C_drain_IO_L1_out_wrapper_147__ap_idle;
  output C_drain_IO_L1_out_wrapper_148__ap_start;
  input C_drain_IO_L1_out_wrapper_148__ap_ready;
  input C_drain_IO_L1_out_wrapper_148__ap_done;
  input C_drain_IO_L1_out_wrapper_148__ap_idle;
  output C_drain_IO_L1_out_wrapper_149__ap_start;
  input C_drain_IO_L1_out_wrapper_149__ap_ready;
  input C_drain_IO_L1_out_wrapper_149__ap_done;
  input C_drain_IO_L1_out_wrapper_149__ap_idle;
  output C_drain_IO_L1_out_wrapper_150__ap_start;
  input C_drain_IO_L1_out_wrapper_150__ap_ready;
  input C_drain_IO_L1_out_wrapper_150__ap_done;
  input C_drain_IO_L1_out_wrapper_150__ap_idle;
  output C_drain_IO_L1_out_wrapper_151__ap_start;
  input C_drain_IO_L1_out_wrapper_151__ap_ready;
  input C_drain_IO_L1_out_wrapper_151__ap_done;
  input C_drain_IO_L1_out_wrapper_151__ap_idle;
  output C_drain_IO_L1_out_wrapper_152__ap_start;
  input C_drain_IO_L1_out_wrapper_152__ap_ready;
  input C_drain_IO_L1_out_wrapper_152__ap_done;
  input C_drain_IO_L1_out_wrapper_152__ap_idle;
  output C_drain_IO_L1_out_wrapper_153__ap_start;
  input C_drain_IO_L1_out_wrapper_153__ap_ready;
  input C_drain_IO_L1_out_wrapper_153__ap_done;
  input C_drain_IO_L1_out_wrapper_153__ap_idle;
  output C_drain_IO_L1_out_wrapper_154__ap_start;
  input C_drain_IO_L1_out_wrapper_154__ap_ready;
  input C_drain_IO_L1_out_wrapper_154__ap_done;
  input C_drain_IO_L1_out_wrapper_154__ap_idle;
  output C_drain_IO_L1_out_wrapper_155__ap_start;
  input C_drain_IO_L1_out_wrapper_155__ap_ready;
  input C_drain_IO_L1_out_wrapper_155__ap_done;
  input C_drain_IO_L1_out_wrapper_155__ap_idle;
  output C_drain_IO_L1_out_wrapper_156__ap_start;
  input C_drain_IO_L1_out_wrapper_156__ap_ready;
  input C_drain_IO_L1_out_wrapper_156__ap_done;
  input C_drain_IO_L1_out_wrapper_156__ap_idle;
  output C_drain_IO_L1_out_wrapper_157__ap_start;
  input C_drain_IO_L1_out_wrapper_157__ap_ready;
  input C_drain_IO_L1_out_wrapper_157__ap_done;
  input C_drain_IO_L1_out_wrapper_157__ap_idle;
  output C_drain_IO_L1_out_wrapper_158__ap_start;
  input C_drain_IO_L1_out_wrapper_158__ap_ready;
  input C_drain_IO_L1_out_wrapper_158__ap_done;
  input C_drain_IO_L1_out_wrapper_158__ap_idle;
  output C_drain_IO_L1_out_wrapper_159__ap_start;
  input C_drain_IO_L1_out_wrapper_159__ap_ready;
  input C_drain_IO_L1_out_wrapper_159__ap_done;
  input C_drain_IO_L1_out_wrapper_159__ap_idle;
  output C_drain_IO_L1_out_wrapper_160__ap_start;
  input C_drain_IO_L1_out_wrapper_160__ap_ready;
  input C_drain_IO_L1_out_wrapper_160__ap_done;
  input C_drain_IO_L1_out_wrapper_160__ap_idle;
  output C_drain_IO_L1_out_wrapper_161__ap_start;
  input C_drain_IO_L1_out_wrapper_161__ap_ready;
  input C_drain_IO_L1_out_wrapper_161__ap_done;
  input C_drain_IO_L1_out_wrapper_161__ap_idle;
  output C_drain_IO_L1_out_wrapper_162__ap_start;
  input C_drain_IO_L1_out_wrapper_162__ap_ready;
  input C_drain_IO_L1_out_wrapper_162__ap_done;
  input C_drain_IO_L1_out_wrapper_162__ap_idle;
  output C_drain_IO_L1_out_wrapper_163__ap_start;
  input C_drain_IO_L1_out_wrapper_163__ap_ready;
  input C_drain_IO_L1_out_wrapper_163__ap_done;
  input C_drain_IO_L1_out_wrapper_163__ap_idle;
  output C_drain_IO_L1_out_wrapper_164__ap_start;
  input C_drain_IO_L1_out_wrapper_164__ap_ready;
  input C_drain_IO_L1_out_wrapper_164__ap_done;
  input C_drain_IO_L1_out_wrapper_164__ap_idle;
  output C_drain_IO_L1_out_wrapper_165__ap_start;
  input C_drain_IO_L1_out_wrapper_165__ap_ready;
  input C_drain_IO_L1_out_wrapper_165__ap_done;
  input C_drain_IO_L1_out_wrapper_165__ap_idle;
  output C_drain_IO_L1_out_wrapper_166__ap_start;
  input C_drain_IO_L1_out_wrapper_166__ap_ready;
  input C_drain_IO_L1_out_wrapper_166__ap_done;
  input C_drain_IO_L1_out_wrapper_166__ap_idle;
  output C_drain_IO_L1_out_wrapper_167__ap_start;
  input C_drain_IO_L1_out_wrapper_167__ap_ready;
  input C_drain_IO_L1_out_wrapper_167__ap_done;
  input C_drain_IO_L1_out_wrapper_167__ap_idle;
  output C_drain_IO_L1_out_wrapper_168__ap_start;
  input C_drain_IO_L1_out_wrapper_168__ap_ready;
  input C_drain_IO_L1_out_wrapper_168__ap_done;
  input C_drain_IO_L1_out_wrapper_168__ap_idle;
  output C_drain_IO_L1_out_wrapper_169__ap_start;
  input C_drain_IO_L1_out_wrapper_169__ap_ready;
  input C_drain_IO_L1_out_wrapper_169__ap_done;
  input C_drain_IO_L1_out_wrapper_169__ap_idle;
  output C_drain_IO_L1_out_wrapper_170__ap_start;
  input C_drain_IO_L1_out_wrapper_170__ap_ready;
  input C_drain_IO_L1_out_wrapper_170__ap_done;
  input C_drain_IO_L1_out_wrapper_170__ap_idle;
  output C_drain_IO_L1_out_wrapper_171__ap_start;
  input C_drain_IO_L1_out_wrapper_171__ap_ready;
  input C_drain_IO_L1_out_wrapper_171__ap_done;
  input C_drain_IO_L1_out_wrapper_171__ap_idle;
  output C_drain_IO_L1_out_wrapper_172__ap_start;
  input C_drain_IO_L1_out_wrapper_172__ap_ready;
  input C_drain_IO_L1_out_wrapper_172__ap_done;
  input C_drain_IO_L1_out_wrapper_172__ap_idle;
  output C_drain_IO_L1_out_wrapper_173__ap_start;
  input C_drain_IO_L1_out_wrapper_173__ap_ready;
  input C_drain_IO_L1_out_wrapper_173__ap_done;
  input C_drain_IO_L1_out_wrapper_173__ap_idle;
  output C_drain_IO_L1_out_wrapper_174__ap_start;
  input C_drain_IO_L1_out_wrapper_174__ap_ready;
  input C_drain_IO_L1_out_wrapper_174__ap_done;
  input C_drain_IO_L1_out_wrapper_174__ap_idle;
  output C_drain_IO_L1_out_wrapper_175__ap_start;
  input C_drain_IO_L1_out_wrapper_175__ap_ready;
  input C_drain_IO_L1_out_wrapper_175__ap_done;
  input C_drain_IO_L1_out_wrapper_175__ap_idle;
  output C_drain_IO_L1_out_wrapper_176__ap_start;
  input C_drain_IO_L1_out_wrapper_176__ap_ready;
  input C_drain_IO_L1_out_wrapper_176__ap_done;
  input C_drain_IO_L1_out_wrapper_176__ap_idle;
  output C_drain_IO_L1_out_wrapper_177__ap_start;
  input C_drain_IO_L1_out_wrapper_177__ap_ready;
  input C_drain_IO_L1_out_wrapper_177__ap_done;
  input C_drain_IO_L1_out_wrapper_177__ap_idle;
  output C_drain_IO_L1_out_wrapper_178__ap_start;
  input C_drain_IO_L1_out_wrapper_178__ap_ready;
  input C_drain_IO_L1_out_wrapper_178__ap_done;
  input C_drain_IO_L1_out_wrapper_178__ap_idle;
  output C_drain_IO_L1_out_wrapper_179__ap_start;
  input C_drain_IO_L1_out_wrapper_179__ap_ready;
  input C_drain_IO_L1_out_wrapper_179__ap_done;
  input C_drain_IO_L1_out_wrapper_179__ap_idle;
  output C_drain_IO_L1_out_wrapper_180__ap_start;
  input C_drain_IO_L1_out_wrapper_180__ap_ready;
  input C_drain_IO_L1_out_wrapper_180__ap_done;
  input C_drain_IO_L1_out_wrapper_180__ap_idle;
  output C_drain_IO_L1_out_wrapper_181__ap_start;
  input C_drain_IO_L1_out_wrapper_181__ap_ready;
  input C_drain_IO_L1_out_wrapper_181__ap_done;
  input C_drain_IO_L1_out_wrapper_181__ap_idle;
  output C_drain_IO_L1_out_wrapper_182__ap_start;
  input C_drain_IO_L1_out_wrapper_182__ap_ready;
  input C_drain_IO_L1_out_wrapper_182__ap_done;
  input C_drain_IO_L1_out_wrapper_182__ap_idle;
  output C_drain_IO_L1_out_wrapper_183__ap_start;
  input C_drain_IO_L1_out_wrapper_183__ap_ready;
  input C_drain_IO_L1_out_wrapper_183__ap_done;
  input C_drain_IO_L1_out_wrapper_183__ap_idle;
  output C_drain_IO_L1_out_wrapper_184__ap_start;
  input C_drain_IO_L1_out_wrapper_184__ap_ready;
  input C_drain_IO_L1_out_wrapper_184__ap_done;
  input C_drain_IO_L1_out_wrapper_184__ap_idle;
  output C_drain_IO_L1_out_wrapper_185__ap_start;
  input C_drain_IO_L1_out_wrapper_185__ap_ready;
  input C_drain_IO_L1_out_wrapper_185__ap_done;
  input C_drain_IO_L1_out_wrapper_185__ap_idle;
  output C_drain_IO_L1_out_wrapper_186__ap_start;
  input C_drain_IO_L1_out_wrapper_186__ap_ready;
  input C_drain_IO_L1_out_wrapper_186__ap_done;
  input C_drain_IO_L1_out_wrapper_186__ap_idle;
  output C_drain_IO_L1_out_wrapper_187__ap_start;
  input C_drain_IO_L1_out_wrapper_187__ap_ready;
  input C_drain_IO_L1_out_wrapper_187__ap_done;
  input C_drain_IO_L1_out_wrapper_187__ap_idle;
  output C_drain_IO_L1_out_wrapper_188__ap_start;
  input C_drain_IO_L1_out_wrapper_188__ap_ready;
  input C_drain_IO_L1_out_wrapper_188__ap_done;
  input C_drain_IO_L1_out_wrapper_188__ap_idle;
  output C_drain_IO_L1_out_wrapper_189__ap_start;
  input C_drain_IO_L1_out_wrapper_189__ap_ready;
  input C_drain_IO_L1_out_wrapper_189__ap_done;
  input C_drain_IO_L1_out_wrapper_189__ap_idle;
  output C_drain_IO_L1_out_wrapper_190__ap_start;
  input C_drain_IO_L1_out_wrapper_190__ap_ready;
  input C_drain_IO_L1_out_wrapper_190__ap_done;
  input C_drain_IO_L1_out_wrapper_190__ap_idle;
  output C_drain_IO_L1_out_wrapper_191__ap_start;
  input C_drain_IO_L1_out_wrapper_191__ap_ready;
  input C_drain_IO_L1_out_wrapper_191__ap_done;
  input C_drain_IO_L1_out_wrapper_191__ap_idle;
  output C_drain_IO_L1_out_wrapper_192__ap_start;
  input C_drain_IO_L1_out_wrapper_192__ap_ready;
  input C_drain_IO_L1_out_wrapper_192__ap_done;
  input C_drain_IO_L1_out_wrapper_192__ap_idle;
  output C_drain_IO_L1_out_wrapper_193__ap_start;
  input C_drain_IO_L1_out_wrapper_193__ap_ready;
  input C_drain_IO_L1_out_wrapper_193__ap_done;
  input C_drain_IO_L1_out_wrapper_193__ap_idle;
  output C_drain_IO_L1_out_wrapper_194__ap_start;
  input C_drain_IO_L1_out_wrapper_194__ap_ready;
  input C_drain_IO_L1_out_wrapper_194__ap_done;
  input C_drain_IO_L1_out_wrapper_194__ap_idle;
  output C_drain_IO_L1_out_wrapper_195__ap_start;
  input C_drain_IO_L1_out_wrapper_195__ap_ready;
  input C_drain_IO_L1_out_wrapper_195__ap_done;
  input C_drain_IO_L1_out_wrapper_195__ap_idle;
  output C_drain_IO_L1_out_wrapper_196__ap_start;
  input C_drain_IO_L1_out_wrapper_196__ap_ready;
  input C_drain_IO_L1_out_wrapper_196__ap_done;
  input C_drain_IO_L1_out_wrapper_196__ap_idle;
  output C_drain_IO_L1_out_wrapper_197__ap_start;
  input C_drain_IO_L1_out_wrapper_197__ap_ready;
  input C_drain_IO_L1_out_wrapper_197__ap_done;
  input C_drain_IO_L1_out_wrapper_197__ap_idle;
  output C_drain_IO_L1_out_wrapper_198__ap_start;
  input C_drain_IO_L1_out_wrapper_198__ap_ready;
  input C_drain_IO_L1_out_wrapper_198__ap_done;
  input C_drain_IO_L1_out_wrapper_198__ap_idle;
  output C_drain_IO_L1_out_wrapper_199__ap_start;
  input C_drain_IO_L1_out_wrapper_199__ap_ready;
  input C_drain_IO_L1_out_wrapper_199__ap_done;
  input C_drain_IO_L1_out_wrapper_199__ap_idle;
  output C_drain_IO_L1_out_wrapper_200__ap_start;
  input C_drain_IO_L1_out_wrapper_200__ap_ready;
  input C_drain_IO_L1_out_wrapper_200__ap_done;
  input C_drain_IO_L1_out_wrapper_200__ap_idle;
  output C_drain_IO_L1_out_wrapper_201__ap_start;
  input C_drain_IO_L1_out_wrapper_201__ap_ready;
  input C_drain_IO_L1_out_wrapper_201__ap_done;
  input C_drain_IO_L1_out_wrapper_201__ap_idle;
  output C_drain_IO_L1_out_wrapper_202__ap_start;
  input C_drain_IO_L1_out_wrapper_202__ap_ready;
  input C_drain_IO_L1_out_wrapper_202__ap_done;
  input C_drain_IO_L1_out_wrapper_202__ap_idle;
  output C_drain_IO_L1_out_wrapper_203__ap_start;
  input C_drain_IO_L1_out_wrapper_203__ap_ready;
  input C_drain_IO_L1_out_wrapper_203__ap_done;
  input C_drain_IO_L1_out_wrapper_203__ap_idle;
  output C_drain_IO_L1_out_wrapper_204__ap_start;
  input C_drain_IO_L1_out_wrapper_204__ap_ready;
  input C_drain_IO_L1_out_wrapper_204__ap_done;
  input C_drain_IO_L1_out_wrapper_204__ap_idle;
  output C_drain_IO_L1_out_wrapper_205__ap_start;
  input C_drain_IO_L1_out_wrapper_205__ap_ready;
  input C_drain_IO_L1_out_wrapper_205__ap_done;
  input C_drain_IO_L1_out_wrapper_205__ap_idle;
  output C_drain_IO_L1_out_wrapper_206__ap_start;
  input C_drain_IO_L1_out_wrapper_206__ap_ready;
  input C_drain_IO_L1_out_wrapper_206__ap_done;
  input C_drain_IO_L1_out_wrapper_206__ap_idle;
  output C_drain_IO_L1_out_wrapper_207__ap_start;
  input C_drain_IO_L1_out_wrapper_207__ap_ready;
  input C_drain_IO_L1_out_wrapper_207__ap_done;
  input C_drain_IO_L1_out_wrapper_207__ap_idle;
  output C_drain_IO_L1_out_wrapper_208__ap_start;
  input C_drain_IO_L1_out_wrapper_208__ap_ready;
  input C_drain_IO_L1_out_wrapper_208__ap_done;
  input C_drain_IO_L1_out_wrapper_208__ap_idle;
  output C_drain_IO_L1_out_wrapper_209__ap_start;
  input C_drain_IO_L1_out_wrapper_209__ap_ready;
  input C_drain_IO_L1_out_wrapper_209__ap_done;
  input C_drain_IO_L1_out_wrapper_209__ap_idle;
  output C_drain_IO_L1_out_wrapper_210__ap_start;
  input C_drain_IO_L1_out_wrapper_210__ap_ready;
  input C_drain_IO_L1_out_wrapper_210__ap_done;
  input C_drain_IO_L1_out_wrapper_210__ap_idle;
  output C_drain_IO_L1_out_wrapper_211__ap_start;
  input C_drain_IO_L1_out_wrapper_211__ap_ready;
  input C_drain_IO_L1_out_wrapper_211__ap_done;
  input C_drain_IO_L1_out_wrapper_211__ap_idle;
  output C_drain_IO_L1_out_wrapper_212__ap_start;
  input C_drain_IO_L1_out_wrapper_212__ap_ready;
  input C_drain_IO_L1_out_wrapper_212__ap_done;
  input C_drain_IO_L1_out_wrapper_212__ap_idle;
  output C_drain_IO_L1_out_wrapper_213__ap_start;
  input C_drain_IO_L1_out_wrapper_213__ap_ready;
  input C_drain_IO_L1_out_wrapper_213__ap_done;
  input C_drain_IO_L1_out_wrapper_213__ap_idle;
  output C_drain_IO_L1_out_wrapper_214__ap_start;
  input C_drain_IO_L1_out_wrapper_214__ap_ready;
  input C_drain_IO_L1_out_wrapper_214__ap_done;
  input C_drain_IO_L1_out_wrapper_214__ap_idle;
  output C_drain_IO_L1_out_wrapper_215__ap_start;
  input C_drain_IO_L1_out_wrapper_215__ap_ready;
  input C_drain_IO_L1_out_wrapper_215__ap_done;
  input C_drain_IO_L1_out_wrapper_215__ap_idle;
  output C_drain_IO_L1_out_wrapper_216__ap_start;
  input C_drain_IO_L1_out_wrapper_216__ap_ready;
  input C_drain_IO_L1_out_wrapper_216__ap_done;
  input C_drain_IO_L1_out_wrapper_216__ap_idle;
  output C_drain_IO_L1_out_wrapper_217__ap_start;
  input C_drain_IO_L1_out_wrapper_217__ap_ready;
  input C_drain_IO_L1_out_wrapper_217__ap_done;
  input C_drain_IO_L1_out_wrapper_217__ap_idle;
  output C_drain_IO_L1_out_wrapper_218__ap_start;
  input C_drain_IO_L1_out_wrapper_218__ap_ready;
  input C_drain_IO_L1_out_wrapper_218__ap_done;
  input C_drain_IO_L1_out_wrapper_218__ap_idle;
  output C_drain_IO_L1_out_wrapper_219__ap_start;
  input C_drain_IO_L1_out_wrapper_219__ap_ready;
  input C_drain_IO_L1_out_wrapper_219__ap_done;
  input C_drain_IO_L1_out_wrapper_219__ap_idle;
  output C_drain_IO_L1_out_wrapper_220__ap_start;
  input C_drain_IO_L1_out_wrapper_220__ap_ready;
  input C_drain_IO_L1_out_wrapper_220__ap_done;
  input C_drain_IO_L1_out_wrapper_220__ap_idle;
  output C_drain_IO_L1_out_wrapper_221__ap_start;
  input C_drain_IO_L1_out_wrapper_221__ap_ready;
  input C_drain_IO_L1_out_wrapper_221__ap_done;
  input C_drain_IO_L1_out_wrapper_221__ap_idle;
  output C_drain_IO_L1_out_wrapper_222__ap_start;
  input C_drain_IO_L1_out_wrapper_222__ap_ready;
  input C_drain_IO_L1_out_wrapper_222__ap_done;
  input C_drain_IO_L1_out_wrapper_222__ap_idle;
  output C_drain_IO_L1_out_wrapper_223__ap_start;
  input C_drain_IO_L1_out_wrapper_223__ap_ready;
  input C_drain_IO_L1_out_wrapper_223__ap_done;
  input C_drain_IO_L1_out_wrapper_223__ap_idle;
  output C_drain_IO_L1_out_wrapper_224__ap_start;
  input C_drain_IO_L1_out_wrapper_224__ap_ready;
  input C_drain_IO_L1_out_wrapper_224__ap_done;
  input C_drain_IO_L1_out_wrapper_224__ap_idle;
  output C_drain_IO_L1_out_wrapper_225__ap_start;
  input C_drain_IO_L1_out_wrapper_225__ap_ready;
  input C_drain_IO_L1_out_wrapper_225__ap_done;
  input C_drain_IO_L1_out_wrapper_225__ap_idle;
  output C_drain_IO_L1_out_wrapper_226__ap_start;
  input C_drain_IO_L1_out_wrapper_226__ap_ready;
  input C_drain_IO_L1_out_wrapper_226__ap_done;
  input C_drain_IO_L1_out_wrapper_226__ap_idle;
  output C_drain_IO_L1_out_wrapper_227__ap_start;
  input C_drain_IO_L1_out_wrapper_227__ap_ready;
  input C_drain_IO_L1_out_wrapper_227__ap_done;
  input C_drain_IO_L1_out_wrapper_227__ap_idle;
  output C_drain_IO_L1_out_wrapper_228__ap_start;
  input C_drain_IO_L1_out_wrapper_228__ap_ready;
  input C_drain_IO_L1_out_wrapper_228__ap_done;
  input C_drain_IO_L1_out_wrapper_228__ap_idle;
  output C_drain_IO_L1_out_wrapper_229__ap_start;
  input C_drain_IO_L1_out_wrapper_229__ap_ready;
  input C_drain_IO_L1_out_wrapper_229__ap_done;
  input C_drain_IO_L1_out_wrapper_229__ap_idle;
  output C_drain_IO_L1_out_wrapper_230__ap_start;
  input C_drain_IO_L1_out_wrapper_230__ap_ready;
  input C_drain_IO_L1_out_wrapper_230__ap_done;
  input C_drain_IO_L1_out_wrapper_230__ap_idle;
  output C_drain_IO_L1_out_wrapper_231__ap_start;
  input C_drain_IO_L1_out_wrapper_231__ap_ready;
  input C_drain_IO_L1_out_wrapper_231__ap_done;
  input C_drain_IO_L1_out_wrapper_231__ap_idle;
  output C_drain_IO_L1_out_wrapper_232__ap_start;
  input C_drain_IO_L1_out_wrapper_232__ap_ready;
  input C_drain_IO_L1_out_wrapper_232__ap_done;
  input C_drain_IO_L1_out_wrapper_232__ap_idle;
  output C_drain_IO_L1_out_wrapper_233__ap_start;
  input C_drain_IO_L1_out_wrapper_233__ap_ready;
  input C_drain_IO_L1_out_wrapper_233__ap_done;
  input C_drain_IO_L1_out_wrapper_233__ap_idle;
  output C_drain_IO_L1_out_wrapper_234__ap_start;
  input C_drain_IO_L1_out_wrapper_234__ap_ready;
  input C_drain_IO_L1_out_wrapper_234__ap_done;
  input C_drain_IO_L1_out_wrapper_234__ap_idle;
  output C_drain_IO_L1_out_wrapper_235__ap_start;
  input C_drain_IO_L1_out_wrapper_235__ap_ready;
  input C_drain_IO_L1_out_wrapper_235__ap_done;
  input C_drain_IO_L1_out_wrapper_235__ap_idle;
  output C_drain_IO_L1_out_wrapper_236__ap_start;
  input C_drain_IO_L1_out_wrapper_236__ap_ready;
  input C_drain_IO_L1_out_wrapper_236__ap_done;
  input C_drain_IO_L1_out_wrapper_236__ap_idle;
  output C_drain_IO_L1_out_wrapper_237__ap_start;
  input C_drain_IO_L1_out_wrapper_237__ap_ready;
  input C_drain_IO_L1_out_wrapper_237__ap_done;
  input C_drain_IO_L1_out_wrapper_237__ap_idle;
  output C_drain_IO_L1_out_wrapper_238__ap_start;
  input C_drain_IO_L1_out_wrapper_238__ap_ready;
  input C_drain_IO_L1_out_wrapper_238__ap_done;
  input C_drain_IO_L1_out_wrapper_238__ap_idle;
  output C_drain_IO_L1_out_wrapper_239__ap_start;
  input C_drain_IO_L1_out_wrapper_239__ap_ready;
  input C_drain_IO_L1_out_wrapper_239__ap_done;
  input C_drain_IO_L1_out_wrapper_239__ap_idle;
  output C_drain_IO_L1_out_wrapper_240__ap_start;
  input C_drain_IO_L1_out_wrapper_240__ap_ready;
  input C_drain_IO_L1_out_wrapper_240__ap_done;
  input C_drain_IO_L1_out_wrapper_240__ap_idle;
  output C_drain_IO_L1_out_wrapper_241__ap_start;
  input C_drain_IO_L1_out_wrapper_241__ap_ready;
  input C_drain_IO_L1_out_wrapper_241__ap_done;
  input C_drain_IO_L1_out_wrapper_241__ap_idle;
  output C_drain_IO_L1_out_wrapper_242__ap_start;
  input C_drain_IO_L1_out_wrapper_242__ap_ready;
  input C_drain_IO_L1_out_wrapper_242__ap_done;
  input C_drain_IO_L1_out_wrapper_242__ap_idle;
  output C_drain_IO_L1_out_wrapper_243__ap_start;
  input C_drain_IO_L1_out_wrapper_243__ap_ready;
  input C_drain_IO_L1_out_wrapper_243__ap_done;
  input C_drain_IO_L1_out_wrapper_243__ap_idle;
  output C_drain_IO_L1_out_wrapper_244__ap_start;
  input C_drain_IO_L1_out_wrapper_244__ap_ready;
  input C_drain_IO_L1_out_wrapper_244__ap_done;
  input C_drain_IO_L1_out_wrapper_244__ap_idle;
  output C_drain_IO_L1_out_wrapper_245__ap_start;
  input C_drain_IO_L1_out_wrapper_245__ap_ready;
  input C_drain_IO_L1_out_wrapper_245__ap_done;
  input C_drain_IO_L1_out_wrapper_245__ap_idle;
  output C_drain_IO_L1_out_wrapper_246__ap_start;
  input C_drain_IO_L1_out_wrapper_246__ap_ready;
  input C_drain_IO_L1_out_wrapper_246__ap_done;
  input C_drain_IO_L1_out_wrapper_246__ap_idle;
  output C_drain_IO_L1_out_wrapper_247__ap_start;
  input C_drain_IO_L1_out_wrapper_247__ap_ready;
  input C_drain_IO_L1_out_wrapper_247__ap_done;
  input C_drain_IO_L1_out_wrapper_247__ap_idle;
  output C_drain_IO_L1_out_wrapper_248__ap_start;
  input C_drain_IO_L1_out_wrapper_248__ap_ready;
  input C_drain_IO_L1_out_wrapper_248__ap_done;
  input C_drain_IO_L1_out_wrapper_248__ap_idle;
  output C_drain_IO_L1_out_wrapper_249__ap_start;
  input C_drain_IO_L1_out_wrapper_249__ap_ready;
  input C_drain_IO_L1_out_wrapper_249__ap_done;
  input C_drain_IO_L1_out_wrapper_249__ap_idle;
  output C_drain_IO_L1_out_wrapper_250__ap_start;
  input C_drain_IO_L1_out_wrapper_250__ap_ready;
  input C_drain_IO_L1_out_wrapper_250__ap_done;
  input C_drain_IO_L1_out_wrapper_250__ap_idle;
  output C_drain_IO_L1_out_wrapper_251__ap_start;
  input C_drain_IO_L1_out_wrapper_251__ap_ready;
  input C_drain_IO_L1_out_wrapper_251__ap_done;
  input C_drain_IO_L1_out_wrapper_251__ap_idle;
  output C_drain_IO_L1_out_wrapper_252__ap_start;
  input C_drain_IO_L1_out_wrapper_252__ap_ready;
  input C_drain_IO_L1_out_wrapper_252__ap_done;
  input C_drain_IO_L1_out_wrapper_252__ap_idle;
  output C_drain_IO_L1_out_wrapper_253__ap_start;
  input C_drain_IO_L1_out_wrapper_253__ap_ready;
  input C_drain_IO_L1_out_wrapper_253__ap_done;
  input C_drain_IO_L1_out_wrapper_253__ap_idle;
  output C_drain_IO_L1_out_wrapper_254__ap_start;
  input C_drain_IO_L1_out_wrapper_254__ap_ready;
  input C_drain_IO_L1_out_wrapper_254__ap_done;
  input C_drain_IO_L1_out_wrapper_254__ap_idle;
  output C_drain_IO_L1_out_wrapper_255__ap_start;
  input C_drain_IO_L1_out_wrapper_255__ap_ready;
  input C_drain_IO_L1_out_wrapper_255__ap_done;
  input C_drain_IO_L1_out_wrapper_255__ap_idle;
  output C_drain_IO_L1_out_wrapper_256__ap_start;
  input C_drain_IO_L1_out_wrapper_256__ap_ready;
  input C_drain_IO_L1_out_wrapper_256__ap_done;
  input C_drain_IO_L1_out_wrapper_256__ap_idle;
  output C_drain_IO_L1_out_wrapper_257__ap_start;
  input C_drain_IO_L1_out_wrapper_257__ap_ready;
  input C_drain_IO_L1_out_wrapper_257__ap_done;
  input C_drain_IO_L1_out_wrapper_257__ap_idle;
  output C_drain_IO_L1_out_wrapper_258__ap_start;
  input C_drain_IO_L1_out_wrapper_258__ap_ready;
  input C_drain_IO_L1_out_wrapper_258__ap_done;
  input C_drain_IO_L1_out_wrapper_258__ap_idle;
  output C_drain_IO_L1_out_wrapper_259__ap_start;
  input C_drain_IO_L1_out_wrapper_259__ap_ready;
  input C_drain_IO_L1_out_wrapper_259__ap_done;
  input C_drain_IO_L1_out_wrapper_259__ap_idle;
  output C_drain_IO_L1_out_wrapper_260__ap_start;
  input C_drain_IO_L1_out_wrapper_260__ap_ready;
  input C_drain_IO_L1_out_wrapper_260__ap_done;
  input C_drain_IO_L1_out_wrapper_260__ap_idle;
  output C_drain_IO_L1_out_wrapper_261__ap_start;
  input C_drain_IO_L1_out_wrapper_261__ap_ready;
  input C_drain_IO_L1_out_wrapper_261__ap_done;
  input C_drain_IO_L1_out_wrapper_261__ap_idle;
  output C_drain_IO_L1_out_wrapper_262__ap_start;
  input C_drain_IO_L1_out_wrapper_262__ap_ready;
  input C_drain_IO_L1_out_wrapper_262__ap_done;
  input C_drain_IO_L1_out_wrapper_262__ap_idle;
  output C_drain_IO_L1_out_wrapper_263__ap_start;
  input C_drain_IO_L1_out_wrapper_263__ap_ready;
  input C_drain_IO_L1_out_wrapper_263__ap_done;
  input C_drain_IO_L1_out_wrapper_263__ap_idle;
  output C_drain_IO_L1_out_wrapper_264__ap_start;
  input C_drain_IO_L1_out_wrapper_264__ap_ready;
  input C_drain_IO_L1_out_wrapper_264__ap_done;
  input C_drain_IO_L1_out_wrapper_264__ap_idle;
  output C_drain_IO_L1_out_wrapper_265__ap_start;
  input C_drain_IO_L1_out_wrapper_265__ap_ready;
  input C_drain_IO_L1_out_wrapper_265__ap_done;
  input C_drain_IO_L1_out_wrapper_265__ap_idle;
  output C_drain_IO_L1_out_wrapper_266__ap_start;
  input C_drain_IO_L1_out_wrapper_266__ap_ready;
  input C_drain_IO_L1_out_wrapper_266__ap_done;
  input C_drain_IO_L1_out_wrapper_266__ap_idle;
  output C_drain_IO_L1_out_wrapper_267__ap_start;
  input C_drain_IO_L1_out_wrapper_267__ap_ready;
  input C_drain_IO_L1_out_wrapper_267__ap_done;
  input C_drain_IO_L1_out_wrapper_267__ap_idle;
  output C_drain_IO_L1_out_wrapper_268__ap_start;
  input C_drain_IO_L1_out_wrapper_268__ap_ready;
  input C_drain_IO_L1_out_wrapper_268__ap_done;
  input C_drain_IO_L1_out_wrapper_268__ap_idle;
  output C_drain_IO_L1_out_wrapper_269__ap_start;
  input C_drain_IO_L1_out_wrapper_269__ap_ready;
  input C_drain_IO_L1_out_wrapper_269__ap_done;
  input C_drain_IO_L1_out_wrapper_269__ap_idle;
  output C_drain_IO_L1_out_wrapper_270__ap_start;
  input C_drain_IO_L1_out_wrapper_270__ap_ready;
  input C_drain_IO_L1_out_wrapper_270__ap_done;
  input C_drain_IO_L1_out_wrapper_270__ap_idle;
  output C_drain_IO_L1_out_wrapper_271__ap_start;
  input C_drain_IO_L1_out_wrapper_271__ap_ready;
  input C_drain_IO_L1_out_wrapper_271__ap_done;
  input C_drain_IO_L1_out_wrapper_271__ap_idle;
  output C_drain_IO_L1_out_wrapper_272__ap_start;
  input C_drain_IO_L1_out_wrapper_272__ap_ready;
  input C_drain_IO_L1_out_wrapper_272__ap_done;
  input C_drain_IO_L1_out_wrapper_272__ap_idle;
  output C_drain_IO_L1_out_wrapper_273__ap_start;
  input C_drain_IO_L1_out_wrapper_273__ap_ready;
  input C_drain_IO_L1_out_wrapper_273__ap_done;
  input C_drain_IO_L1_out_wrapper_273__ap_idle;
  output C_drain_IO_L1_out_wrapper_274__ap_start;
  input C_drain_IO_L1_out_wrapper_274__ap_ready;
  input C_drain_IO_L1_out_wrapper_274__ap_done;
  input C_drain_IO_L1_out_wrapper_274__ap_idle;
  output C_drain_IO_L1_out_wrapper_275__ap_start;
  input C_drain_IO_L1_out_wrapper_275__ap_ready;
  input C_drain_IO_L1_out_wrapper_275__ap_done;
  input C_drain_IO_L1_out_wrapper_275__ap_idle;
  output C_drain_IO_L1_out_wrapper_276__ap_start;
  input C_drain_IO_L1_out_wrapper_276__ap_ready;
  input C_drain_IO_L1_out_wrapper_276__ap_done;
  input C_drain_IO_L1_out_wrapper_276__ap_idle;
  output C_drain_IO_L1_out_wrapper_277__ap_start;
  input C_drain_IO_L1_out_wrapper_277__ap_ready;
  input C_drain_IO_L1_out_wrapper_277__ap_done;
  input C_drain_IO_L1_out_wrapper_277__ap_idle;
  output C_drain_IO_L1_out_wrapper_278__ap_start;
  input C_drain_IO_L1_out_wrapper_278__ap_ready;
  input C_drain_IO_L1_out_wrapper_278__ap_done;
  input C_drain_IO_L1_out_wrapper_278__ap_idle;
  output C_drain_IO_L1_out_wrapper_279__ap_start;
  input C_drain_IO_L1_out_wrapper_279__ap_ready;
  input C_drain_IO_L1_out_wrapper_279__ap_done;
  input C_drain_IO_L1_out_wrapper_279__ap_idle;
  output C_drain_IO_L1_out_wrapper_280__ap_start;
  input C_drain_IO_L1_out_wrapper_280__ap_ready;
  input C_drain_IO_L1_out_wrapper_280__ap_done;
  input C_drain_IO_L1_out_wrapper_280__ap_idle;
  output C_drain_IO_L1_out_wrapper_281__ap_start;
  input C_drain_IO_L1_out_wrapper_281__ap_ready;
  input C_drain_IO_L1_out_wrapper_281__ap_done;
  input C_drain_IO_L1_out_wrapper_281__ap_idle;
  output C_drain_IO_L1_out_wrapper_282__ap_start;
  input C_drain_IO_L1_out_wrapper_282__ap_ready;
  input C_drain_IO_L1_out_wrapper_282__ap_done;
  input C_drain_IO_L1_out_wrapper_282__ap_idle;
  output C_drain_IO_L1_out_wrapper_283__ap_start;
  input C_drain_IO_L1_out_wrapper_283__ap_ready;
  input C_drain_IO_L1_out_wrapper_283__ap_done;
  input C_drain_IO_L1_out_wrapper_283__ap_idle;
  output C_drain_IO_L1_out_wrapper_284__ap_start;
  input C_drain_IO_L1_out_wrapper_284__ap_ready;
  input C_drain_IO_L1_out_wrapper_284__ap_done;
  input C_drain_IO_L1_out_wrapper_284__ap_idle;
  output C_drain_IO_L1_out_wrapper_285__ap_start;
  input C_drain_IO_L1_out_wrapper_285__ap_ready;
  input C_drain_IO_L1_out_wrapper_285__ap_done;
  input C_drain_IO_L1_out_wrapper_285__ap_idle;
  output C_drain_IO_L1_out_wrapper_286__ap_start;
  input C_drain_IO_L1_out_wrapper_286__ap_ready;
  input C_drain_IO_L1_out_wrapper_286__ap_done;
  input C_drain_IO_L1_out_wrapper_286__ap_idle;
  output C_drain_IO_L1_out_wrapper_287__ap_start;
  input C_drain_IO_L1_out_wrapper_287__ap_ready;
  input C_drain_IO_L1_out_wrapper_287__ap_done;
  input C_drain_IO_L1_out_wrapper_287__ap_idle;
  output C_drain_IO_L1_out_wrapper_288__ap_start;
  input C_drain_IO_L1_out_wrapper_288__ap_ready;
  input C_drain_IO_L1_out_wrapper_288__ap_done;
  input C_drain_IO_L1_out_wrapper_288__ap_idle;
  output C_drain_IO_L2_out_0__ap_start;
  input C_drain_IO_L2_out_0__ap_ready;
  input C_drain_IO_L2_out_0__ap_done;
  input C_drain_IO_L2_out_0__ap_idle;
  output C_drain_IO_L2_out_1__ap_start;
  input C_drain_IO_L2_out_1__ap_ready;
  input C_drain_IO_L2_out_1__ap_done;
  input C_drain_IO_L2_out_1__ap_idle;
  output C_drain_IO_L2_out_2__ap_start;
  input C_drain_IO_L2_out_2__ap_ready;
  input C_drain_IO_L2_out_2__ap_done;
  input C_drain_IO_L2_out_2__ap_idle;
  output C_drain_IO_L2_out_3__ap_start;
  input C_drain_IO_L2_out_3__ap_ready;
  input C_drain_IO_L2_out_3__ap_done;
  input C_drain_IO_L2_out_3__ap_idle;
  output C_drain_IO_L2_out_4__ap_start;
  input C_drain_IO_L2_out_4__ap_ready;
  input C_drain_IO_L2_out_4__ap_done;
  input C_drain_IO_L2_out_4__ap_idle;
  output C_drain_IO_L2_out_5__ap_start;
  input C_drain_IO_L2_out_5__ap_ready;
  input C_drain_IO_L2_out_5__ap_done;
  input C_drain_IO_L2_out_5__ap_idle;
  output C_drain_IO_L2_out_6__ap_start;
  input C_drain_IO_L2_out_6__ap_ready;
  input C_drain_IO_L2_out_6__ap_done;
  input C_drain_IO_L2_out_6__ap_idle;
  output C_drain_IO_L2_out_7__ap_start;
  input C_drain_IO_L2_out_7__ap_ready;
  input C_drain_IO_L2_out_7__ap_done;
  input C_drain_IO_L2_out_7__ap_idle;
  output C_drain_IO_L2_out_8__ap_start;
  input C_drain_IO_L2_out_8__ap_ready;
  input C_drain_IO_L2_out_8__ap_done;
  input C_drain_IO_L2_out_8__ap_idle;
  output C_drain_IO_L2_out_9__ap_start;
  input C_drain_IO_L2_out_9__ap_ready;
  input C_drain_IO_L2_out_9__ap_done;
  input C_drain_IO_L2_out_9__ap_idle;
  output C_drain_IO_L2_out_10__ap_start;
  input C_drain_IO_L2_out_10__ap_ready;
  input C_drain_IO_L2_out_10__ap_done;
  input C_drain_IO_L2_out_10__ap_idle;
  output C_drain_IO_L2_out_11__ap_start;
  input C_drain_IO_L2_out_11__ap_ready;
  input C_drain_IO_L2_out_11__ap_done;
  input C_drain_IO_L2_out_11__ap_idle;
  output C_drain_IO_L2_out_12__ap_start;
  input C_drain_IO_L2_out_12__ap_ready;
  input C_drain_IO_L2_out_12__ap_done;
  input C_drain_IO_L2_out_12__ap_idle;
  output C_drain_IO_L2_out_13__ap_start;
  input C_drain_IO_L2_out_13__ap_ready;
  input C_drain_IO_L2_out_13__ap_done;
  input C_drain_IO_L2_out_13__ap_idle;
  output C_drain_IO_L2_out_14__ap_start;
  input C_drain_IO_L2_out_14__ap_ready;
  input C_drain_IO_L2_out_14__ap_done;
  input C_drain_IO_L2_out_14__ap_idle;
  output C_drain_IO_L2_out_15__ap_start;
  input C_drain_IO_L2_out_15__ap_ready;
  input C_drain_IO_L2_out_15__ap_done;
  input C_drain_IO_L2_out_15__ap_idle;
  output C_drain_IO_L2_out_boundary_0__ap_start;
  input C_drain_IO_L2_out_boundary_0__ap_ready;
  input C_drain_IO_L2_out_boundary_0__ap_done;
  input C_drain_IO_L2_out_boundary_0__ap_idle;
  output C_drain_IO_L3_out_0__ap_start;
  input C_drain_IO_L3_out_0__ap_ready;
  input C_drain_IO_L3_out_0__ap_done;
  input C_drain_IO_L3_out_0__ap_idle;
  output [63:0] C_drain_IO_L3_out_serialize_0___C__q0;
  output C_drain_IO_L3_out_serialize_0__ap_start;
  input C_drain_IO_L3_out_serialize_0__ap_ready;
  input C_drain_IO_L3_out_serialize_0__ap_done;
  input C_drain_IO_L3_out_serialize_0__ap_idle;
  output PE_wrapper_0__ap_start;
  input PE_wrapper_0__ap_ready;
  input PE_wrapper_0__ap_done;
  input PE_wrapper_0__ap_idle;
  output PE_wrapper_1__ap_start;
  input PE_wrapper_1__ap_ready;
  input PE_wrapper_1__ap_done;
  input PE_wrapper_1__ap_idle;
  output PE_wrapper_2__ap_start;
  input PE_wrapper_2__ap_ready;
  input PE_wrapper_2__ap_done;
  input PE_wrapper_2__ap_idle;
  output PE_wrapper_3__ap_start;
  input PE_wrapper_3__ap_ready;
  input PE_wrapper_3__ap_done;
  input PE_wrapper_3__ap_idle;
  output PE_wrapper_4__ap_start;
  input PE_wrapper_4__ap_ready;
  input PE_wrapper_4__ap_done;
  input PE_wrapper_4__ap_idle;
  output PE_wrapper_5__ap_start;
  input PE_wrapper_5__ap_ready;
  input PE_wrapper_5__ap_done;
  input PE_wrapper_5__ap_idle;
  output PE_wrapper_6__ap_start;
  input PE_wrapper_6__ap_ready;
  input PE_wrapper_6__ap_done;
  input PE_wrapper_6__ap_idle;
  output PE_wrapper_7__ap_start;
  input PE_wrapper_7__ap_ready;
  input PE_wrapper_7__ap_done;
  input PE_wrapper_7__ap_idle;
  output PE_wrapper_8__ap_start;
  input PE_wrapper_8__ap_ready;
  input PE_wrapper_8__ap_done;
  input PE_wrapper_8__ap_idle;
  output PE_wrapper_9__ap_start;
  input PE_wrapper_9__ap_ready;
  input PE_wrapper_9__ap_done;
  input PE_wrapper_9__ap_idle;
  output PE_wrapper_10__ap_start;
  input PE_wrapper_10__ap_ready;
  input PE_wrapper_10__ap_done;
  input PE_wrapper_10__ap_idle;
  output PE_wrapper_11__ap_start;
  input PE_wrapper_11__ap_ready;
  input PE_wrapper_11__ap_done;
  input PE_wrapper_11__ap_idle;
  output PE_wrapper_12__ap_start;
  input PE_wrapper_12__ap_ready;
  input PE_wrapper_12__ap_done;
  input PE_wrapper_12__ap_idle;
  output PE_wrapper_13__ap_start;
  input PE_wrapper_13__ap_ready;
  input PE_wrapper_13__ap_done;
  input PE_wrapper_13__ap_idle;
  output PE_wrapper_14__ap_start;
  input PE_wrapper_14__ap_ready;
  input PE_wrapper_14__ap_done;
  input PE_wrapper_14__ap_idle;
  output PE_wrapper_15__ap_start;
  input PE_wrapper_15__ap_ready;
  input PE_wrapper_15__ap_done;
  input PE_wrapper_15__ap_idle;
  output PE_wrapper_16__ap_start;
  input PE_wrapper_16__ap_ready;
  input PE_wrapper_16__ap_done;
  input PE_wrapper_16__ap_idle;
  output PE_wrapper_17__ap_start;
  input PE_wrapper_17__ap_ready;
  input PE_wrapper_17__ap_done;
  input PE_wrapper_17__ap_idle;
  output PE_wrapper_18__ap_start;
  input PE_wrapper_18__ap_ready;
  input PE_wrapper_18__ap_done;
  input PE_wrapper_18__ap_idle;
  output PE_wrapper_19__ap_start;
  input PE_wrapper_19__ap_ready;
  input PE_wrapper_19__ap_done;
  input PE_wrapper_19__ap_idle;
  output PE_wrapper_20__ap_start;
  input PE_wrapper_20__ap_ready;
  input PE_wrapper_20__ap_done;
  input PE_wrapper_20__ap_idle;
  output PE_wrapper_21__ap_start;
  input PE_wrapper_21__ap_ready;
  input PE_wrapper_21__ap_done;
  input PE_wrapper_21__ap_idle;
  output PE_wrapper_22__ap_start;
  input PE_wrapper_22__ap_ready;
  input PE_wrapper_22__ap_done;
  input PE_wrapper_22__ap_idle;
  output PE_wrapper_23__ap_start;
  input PE_wrapper_23__ap_ready;
  input PE_wrapper_23__ap_done;
  input PE_wrapper_23__ap_idle;
  output PE_wrapper_24__ap_start;
  input PE_wrapper_24__ap_ready;
  input PE_wrapper_24__ap_done;
  input PE_wrapper_24__ap_idle;
  output PE_wrapper_25__ap_start;
  input PE_wrapper_25__ap_ready;
  input PE_wrapper_25__ap_done;
  input PE_wrapper_25__ap_idle;
  output PE_wrapper_26__ap_start;
  input PE_wrapper_26__ap_ready;
  input PE_wrapper_26__ap_done;
  input PE_wrapper_26__ap_idle;
  output PE_wrapper_27__ap_start;
  input PE_wrapper_27__ap_ready;
  input PE_wrapper_27__ap_done;
  input PE_wrapper_27__ap_idle;
  output PE_wrapper_28__ap_start;
  input PE_wrapper_28__ap_ready;
  input PE_wrapper_28__ap_done;
  input PE_wrapper_28__ap_idle;
  output PE_wrapper_29__ap_start;
  input PE_wrapper_29__ap_ready;
  input PE_wrapper_29__ap_done;
  input PE_wrapper_29__ap_idle;
  output PE_wrapper_30__ap_start;
  input PE_wrapper_30__ap_ready;
  input PE_wrapper_30__ap_done;
  input PE_wrapper_30__ap_idle;
  output PE_wrapper_31__ap_start;
  input PE_wrapper_31__ap_ready;
  input PE_wrapper_31__ap_done;
  input PE_wrapper_31__ap_idle;
  output PE_wrapper_32__ap_start;
  input PE_wrapper_32__ap_ready;
  input PE_wrapper_32__ap_done;
  input PE_wrapper_32__ap_idle;
  output PE_wrapper_33__ap_start;
  input PE_wrapper_33__ap_ready;
  input PE_wrapper_33__ap_done;
  input PE_wrapper_33__ap_idle;
  output PE_wrapper_34__ap_start;
  input PE_wrapper_34__ap_ready;
  input PE_wrapper_34__ap_done;
  input PE_wrapper_34__ap_idle;
  output PE_wrapper_35__ap_start;
  input PE_wrapper_35__ap_ready;
  input PE_wrapper_35__ap_done;
  input PE_wrapper_35__ap_idle;
  output PE_wrapper_36__ap_start;
  input PE_wrapper_36__ap_ready;
  input PE_wrapper_36__ap_done;
  input PE_wrapper_36__ap_idle;
  output PE_wrapper_37__ap_start;
  input PE_wrapper_37__ap_ready;
  input PE_wrapper_37__ap_done;
  input PE_wrapper_37__ap_idle;
  output PE_wrapper_38__ap_start;
  input PE_wrapper_38__ap_ready;
  input PE_wrapper_38__ap_done;
  input PE_wrapper_38__ap_idle;
  output PE_wrapper_39__ap_start;
  input PE_wrapper_39__ap_ready;
  input PE_wrapper_39__ap_done;
  input PE_wrapper_39__ap_idle;
  output PE_wrapper_40__ap_start;
  input PE_wrapper_40__ap_ready;
  input PE_wrapper_40__ap_done;
  input PE_wrapper_40__ap_idle;
  output PE_wrapper_41__ap_start;
  input PE_wrapper_41__ap_ready;
  input PE_wrapper_41__ap_done;
  input PE_wrapper_41__ap_idle;
  output PE_wrapper_42__ap_start;
  input PE_wrapper_42__ap_ready;
  input PE_wrapper_42__ap_done;
  input PE_wrapper_42__ap_idle;
  output PE_wrapper_43__ap_start;
  input PE_wrapper_43__ap_ready;
  input PE_wrapper_43__ap_done;
  input PE_wrapper_43__ap_idle;
  output PE_wrapper_44__ap_start;
  input PE_wrapper_44__ap_ready;
  input PE_wrapper_44__ap_done;
  input PE_wrapper_44__ap_idle;
  output PE_wrapper_45__ap_start;
  input PE_wrapper_45__ap_ready;
  input PE_wrapper_45__ap_done;
  input PE_wrapper_45__ap_idle;
  output PE_wrapper_46__ap_start;
  input PE_wrapper_46__ap_ready;
  input PE_wrapper_46__ap_done;
  input PE_wrapper_46__ap_idle;
  output PE_wrapper_47__ap_start;
  input PE_wrapper_47__ap_ready;
  input PE_wrapper_47__ap_done;
  input PE_wrapper_47__ap_idle;
  output PE_wrapper_48__ap_start;
  input PE_wrapper_48__ap_ready;
  input PE_wrapper_48__ap_done;
  input PE_wrapper_48__ap_idle;
  output PE_wrapper_49__ap_start;
  input PE_wrapper_49__ap_ready;
  input PE_wrapper_49__ap_done;
  input PE_wrapper_49__ap_idle;
  output PE_wrapper_50__ap_start;
  input PE_wrapper_50__ap_ready;
  input PE_wrapper_50__ap_done;
  input PE_wrapper_50__ap_idle;
  output PE_wrapper_51__ap_start;
  input PE_wrapper_51__ap_ready;
  input PE_wrapper_51__ap_done;
  input PE_wrapper_51__ap_idle;
  output PE_wrapper_52__ap_start;
  input PE_wrapper_52__ap_ready;
  input PE_wrapper_52__ap_done;
  input PE_wrapper_52__ap_idle;
  output PE_wrapper_53__ap_start;
  input PE_wrapper_53__ap_ready;
  input PE_wrapper_53__ap_done;
  input PE_wrapper_53__ap_idle;
  output PE_wrapper_54__ap_start;
  input PE_wrapper_54__ap_ready;
  input PE_wrapper_54__ap_done;
  input PE_wrapper_54__ap_idle;
  output PE_wrapper_55__ap_start;
  input PE_wrapper_55__ap_ready;
  input PE_wrapper_55__ap_done;
  input PE_wrapper_55__ap_idle;
  output PE_wrapper_56__ap_start;
  input PE_wrapper_56__ap_ready;
  input PE_wrapper_56__ap_done;
  input PE_wrapper_56__ap_idle;
  output PE_wrapper_57__ap_start;
  input PE_wrapper_57__ap_ready;
  input PE_wrapper_57__ap_done;
  input PE_wrapper_57__ap_idle;
  output PE_wrapper_58__ap_start;
  input PE_wrapper_58__ap_ready;
  input PE_wrapper_58__ap_done;
  input PE_wrapper_58__ap_idle;
  output PE_wrapper_59__ap_start;
  input PE_wrapper_59__ap_ready;
  input PE_wrapper_59__ap_done;
  input PE_wrapper_59__ap_idle;
  output PE_wrapper_60__ap_start;
  input PE_wrapper_60__ap_ready;
  input PE_wrapper_60__ap_done;
  input PE_wrapper_60__ap_idle;
  output PE_wrapper_61__ap_start;
  input PE_wrapper_61__ap_ready;
  input PE_wrapper_61__ap_done;
  input PE_wrapper_61__ap_idle;
  output PE_wrapper_62__ap_start;
  input PE_wrapper_62__ap_ready;
  input PE_wrapper_62__ap_done;
  input PE_wrapper_62__ap_idle;
  output PE_wrapper_63__ap_start;
  input PE_wrapper_63__ap_ready;
  input PE_wrapper_63__ap_done;
  input PE_wrapper_63__ap_idle;
  output PE_wrapper_64__ap_start;
  input PE_wrapper_64__ap_ready;
  input PE_wrapper_64__ap_done;
  input PE_wrapper_64__ap_idle;
  output PE_wrapper_65__ap_start;
  input PE_wrapper_65__ap_ready;
  input PE_wrapper_65__ap_done;
  input PE_wrapper_65__ap_idle;
  output PE_wrapper_66__ap_start;
  input PE_wrapper_66__ap_ready;
  input PE_wrapper_66__ap_done;
  input PE_wrapper_66__ap_idle;
  output PE_wrapper_67__ap_start;
  input PE_wrapper_67__ap_ready;
  input PE_wrapper_67__ap_done;
  input PE_wrapper_67__ap_idle;
  output PE_wrapper_68__ap_start;
  input PE_wrapper_68__ap_ready;
  input PE_wrapper_68__ap_done;
  input PE_wrapper_68__ap_idle;
  output PE_wrapper_69__ap_start;
  input PE_wrapper_69__ap_ready;
  input PE_wrapper_69__ap_done;
  input PE_wrapper_69__ap_idle;
  output PE_wrapper_70__ap_start;
  input PE_wrapper_70__ap_ready;
  input PE_wrapper_70__ap_done;
  input PE_wrapper_70__ap_idle;
  output PE_wrapper_71__ap_start;
  input PE_wrapper_71__ap_ready;
  input PE_wrapper_71__ap_done;
  input PE_wrapper_71__ap_idle;
  output PE_wrapper_72__ap_start;
  input PE_wrapper_72__ap_ready;
  input PE_wrapper_72__ap_done;
  input PE_wrapper_72__ap_idle;
  output PE_wrapper_73__ap_start;
  input PE_wrapper_73__ap_ready;
  input PE_wrapper_73__ap_done;
  input PE_wrapper_73__ap_idle;
  output PE_wrapper_74__ap_start;
  input PE_wrapper_74__ap_ready;
  input PE_wrapper_74__ap_done;
  input PE_wrapper_74__ap_idle;
  output PE_wrapper_75__ap_start;
  input PE_wrapper_75__ap_ready;
  input PE_wrapper_75__ap_done;
  input PE_wrapper_75__ap_idle;
  output PE_wrapper_76__ap_start;
  input PE_wrapper_76__ap_ready;
  input PE_wrapper_76__ap_done;
  input PE_wrapper_76__ap_idle;
  output PE_wrapper_77__ap_start;
  input PE_wrapper_77__ap_ready;
  input PE_wrapper_77__ap_done;
  input PE_wrapper_77__ap_idle;
  output PE_wrapper_78__ap_start;
  input PE_wrapper_78__ap_ready;
  input PE_wrapper_78__ap_done;
  input PE_wrapper_78__ap_idle;
  output PE_wrapper_79__ap_start;
  input PE_wrapper_79__ap_ready;
  input PE_wrapper_79__ap_done;
  input PE_wrapper_79__ap_idle;
  output PE_wrapper_80__ap_start;
  input PE_wrapper_80__ap_ready;
  input PE_wrapper_80__ap_done;
  input PE_wrapper_80__ap_idle;
  output PE_wrapper_81__ap_start;
  input PE_wrapper_81__ap_ready;
  input PE_wrapper_81__ap_done;
  input PE_wrapper_81__ap_idle;
  output PE_wrapper_82__ap_start;
  input PE_wrapper_82__ap_ready;
  input PE_wrapper_82__ap_done;
  input PE_wrapper_82__ap_idle;
  output PE_wrapper_83__ap_start;
  input PE_wrapper_83__ap_ready;
  input PE_wrapper_83__ap_done;
  input PE_wrapper_83__ap_idle;
  output PE_wrapper_84__ap_start;
  input PE_wrapper_84__ap_ready;
  input PE_wrapper_84__ap_done;
  input PE_wrapper_84__ap_idle;
  output PE_wrapper_85__ap_start;
  input PE_wrapper_85__ap_ready;
  input PE_wrapper_85__ap_done;
  input PE_wrapper_85__ap_idle;
  output PE_wrapper_86__ap_start;
  input PE_wrapper_86__ap_ready;
  input PE_wrapper_86__ap_done;
  input PE_wrapper_86__ap_idle;
  output PE_wrapper_87__ap_start;
  input PE_wrapper_87__ap_ready;
  input PE_wrapper_87__ap_done;
  input PE_wrapper_87__ap_idle;
  output PE_wrapper_88__ap_start;
  input PE_wrapper_88__ap_ready;
  input PE_wrapper_88__ap_done;
  input PE_wrapper_88__ap_idle;
  output PE_wrapper_89__ap_start;
  input PE_wrapper_89__ap_ready;
  input PE_wrapper_89__ap_done;
  input PE_wrapper_89__ap_idle;
  output PE_wrapper_90__ap_start;
  input PE_wrapper_90__ap_ready;
  input PE_wrapper_90__ap_done;
  input PE_wrapper_90__ap_idle;
  output PE_wrapper_91__ap_start;
  input PE_wrapper_91__ap_ready;
  input PE_wrapper_91__ap_done;
  input PE_wrapper_91__ap_idle;
  output PE_wrapper_92__ap_start;
  input PE_wrapper_92__ap_ready;
  input PE_wrapper_92__ap_done;
  input PE_wrapper_92__ap_idle;
  output PE_wrapper_93__ap_start;
  input PE_wrapper_93__ap_ready;
  input PE_wrapper_93__ap_done;
  input PE_wrapper_93__ap_idle;
  output PE_wrapper_94__ap_start;
  input PE_wrapper_94__ap_ready;
  input PE_wrapper_94__ap_done;
  input PE_wrapper_94__ap_idle;
  output PE_wrapper_95__ap_start;
  input PE_wrapper_95__ap_ready;
  input PE_wrapper_95__ap_done;
  input PE_wrapper_95__ap_idle;
  output PE_wrapper_96__ap_start;
  input PE_wrapper_96__ap_ready;
  input PE_wrapper_96__ap_done;
  input PE_wrapper_96__ap_idle;
  output PE_wrapper_97__ap_start;
  input PE_wrapper_97__ap_ready;
  input PE_wrapper_97__ap_done;
  input PE_wrapper_97__ap_idle;
  output PE_wrapper_98__ap_start;
  input PE_wrapper_98__ap_ready;
  input PE_wrapper_98__ap_done;
  input PE_wrapper_98__ap_idle;
  output PE_wrapper_99__ap_start;
  input PE_wrapper_99__ap_ready;
  input PE_wrapper_99__ap_done;
  input PE_wrapper_99__ap_idle;
  output PE_wrapper_100__ap_start;
  input PE_wrapper_100__ap_ready;
  input PE_wrapper_100__ap_done;
  input PE_wrapper_100__ap_idle;
  output PE_wrapper_101__ap_start;
  input PE_wrapper_101__ap_ready;
  input PE_wrapper_101__ap_done;
  input PE_wrapper_101__ap_idle;
  output PE_wrapper_102__ap_start;
  input PE_wrapper_102__ap_ready;
  input PE_wrapper_102__ap_done;
  input PE_wrapper_102__ap_idle;
  output PE_wrapper_103__ap_start;
  input PE_wrapper_103__ap_ready;
  input PE_wrapper_103__ap_done;
  input PE_wrapper_103__ap_idle;
  output PE_wrapper_104__ap_start;
  input PE_wrapper_104__ap_ready;
  input PE_wrapper_104__ap_done;
  input PE_wrapper_104__ap_idle;
  output PE_wrapper_105__ap_start;
  input PE_wrapper_105__ap_ready;
  input PE_wrapper_105__ap_done;
  input PE_wrapper_105__ap_idle;
  output PE_wrapper_106__ap_start;
  input PE_wrapper_106__ap_ready;
  input PE_wrapper_106__ap_done;
  input PE_wrapper_106__ap_idle;
  output PE_wrapper_107__ap_start;
  input PE_wrapper_107__ap_ready;
  input PE_wrapper_107__ap_done;
  input PE_wrapper_107__ap_idle;
  output PE_wrapper_108__ap_start;
  input PE_wrapper_108__ap_ready;
  input PE_wrapper_108__ap_done;
  input PE_wrapper_108__ap_idle;
  output PE_wrapper_109__ap_start;
  input PE_wrapper_109__ap_ready;
  input PE_wrapper_109__ap_done;
  input PE_wrapper_109__ap_idle;
  output PE_wrapper_110__ap_start;
  input PE_wrapper_110__ap_ready;
  input PE_wrapper_110__ap_done;
  input PE_wrapper_110__ap_idle;
  output PE_wrapper_111__ap_start;
  input PE_wrapper_111__ap_ready;
  input PE_wrapper_111__ap_done;
  input PE_wrapper_111__ap_idle;
  output PE_wrapper_112__ap_start;
  input PE_wrapper_112__ap_ready;
  input PE_wrapper_112__ap_done;
  input PE_wrapper_112__ap_idle;
  output PE_wrapper_113__ap_start;
  input PE_wrapper_113__ap_ready;
  input PE_wrapper_113__ap_done;
  input PE_wrapper_113__ap_idle;
  output PE_wrapper_114__ap_start;
  input PE_wrapper_114__ap_ready;
  input PE_wrapper_114__ap_done;
  input PE_wrapper_114__ap_idle;
  output PE_wrapper_115__ap_start;
  input PE_wrapper_115__ap_ready;
  input PE_wrapper_115__ap_done;
  input PE_wrapper_115__ap_idle;
  output PE_wrapper_116__ap_start;
  input PE_wrapper_116__ap_ready;
  input PE_wrapper_116__ap_done;
  input PE_wrapper_116__ap_idle;
  output PE_wrapper_117__ap_start;
  input PE_wrapper_117__ap_ready;
  input PE_wrapper_117__ap_done;
  input PE_wrapper_117__ap_idle;
  output PE_wrapper_118__ap_start;
  input PE_wrapper_118__ap_ready;
  input PE_wrapper_118__ap_done;
  input PE_wrapper_118__ap_idle;
  output PE_wrapper_119__ap_start;
  input PE_wrapper_119__ap_ready;
  input PE_wrapper_119__ap_done;
  input PE_wrapper_119__ap_idle;
  output PE_wrapper_120__ap_start;
  input PE_wrapper_120__ap_ready;
  input PE_wrapper_120__ap_done;
  input PE_wrapper_120__ap_idle;
  output PE_wrapper_121__ap_start;
  input PE_wrapper_121__ap_ready;
  input PE_wrapper_121__ap_done;
  input PE_wrapper_121__ap_idle;
  output PE_wrapper_122__ap_start;
  input PE_wrapper_122__ap_ready;
  input PE_wrapper_122__ap_done;
  input PE_wrapper_122__ap_idle;
  output PE_wrapper_123__ap_start;
  input PE_wrapper_123__ap_ready;
  input PE_wrapper_123__ap_done;
  input PE_wrapper_123__ap_idle;
  output PE_wrapper_124__ap_start;
  input PE_wrapper_124__ap_ready;
  input PE_wrapper_124__ap_done;
  input PE_wrapper_124__ap_idle;
  output PE_wrapper_125__ap_start;
  input PE_wrapper_125__ap_ready;
  input PE_wrapper_125__ap_done;
  input PE_wrapper_125__ap_idle;
  output PE_wrapper_126__ap_start;
  input PE_wrapper_126__ap_ready;
  input PE_wrapper_126__ap_done;
  input PE_wrapper_126__ap_idle;
  output PE_wrapper_127__ap_start;
  input PE_wrapper_127__ap_ready;
  input PE_wrapper_127__ap_done;
  input PE_wrapper_127__ap_idle;
  output PE_wrapper_128__ap_start;
  input PE_wrapper_128__ap_ready;
  input PE_wrapper_128__ap_done;
  input PE_wrapper_128__ap_idle;
  output PE_wrapper_129__ap_start;
  input PE_wrapper_129__ap_ready;
  input PE_wrapper_129__ap_done;
  input PE_wrapper_129__ap_idle;
  output PE_wrapper_130__ap_start;
  input PE_wrapper_130__ap_ready;
  input PE_wrapper_130__ap_done;
  input PE_wrapper_130__ap_idle;
  output PE_wrapper_131__ap_start;
  input PE_wrapper_131__ap_ready;
  input PE_wrapper_131__ap_done;
  input PE_wrapper_131__ap_idle;
  output PE_wrapper_132__ap_start;
  input PE_wrapper_132__ap_ready;
  input PE_wrapper_132__ap_done;
  input PE_wrapper_132__ap_idle;
  output PE_wrapper_133__ap_start;
  input PE_wrapper_133__ap_ready;
  input PE_wrapper_133__ap_done;
  input PE_wrapper_133__ap_idle;
  output PE_wrapper_134__ap_start;
  input PE_wrapper_134__ap_ready;
  input PE_wrapper_134__ap_done;
  input PE_wrapper_134__ap_idle;
  output PE_wrapper_135__ap_start;
  input PE_wrapper_135__ap_ready;
  input PE_wrapper_135__ap_done;
  input PE_wrapper_135__ap_idle;
  output PE_wrapper_136__ap_start;
  input PE_wrapper_136__ap_ready;
  input PE_wrapper_136__ap_done;
  input PE_wrapper_136__ap_idle;
  output PE_wrapper_137__ap_start;
  input PE_wrapper_137__ap_ready;
  input PE_wrapper_137__ap_done;
  input PE_wrapper_137__ap_idle;
  output PE_wrapper_138__ap_start;
  input PE_wrapper_138__ap_ready;
  input PE_wrapper_138__ap_done;
  input PE_wrapper_138__ap_idle;
  output PE_wrapper_139__ap_start;
  input PE_wrapper_139__ap_ready;
  input PE_wrapper_139__ap_done;
  input PE_wrapper_139__ap_idle;
  output PE_wrapper_140__ap_start;
  input PE_wrapper_140__ap_ready;
  input PE_wrapper_140__ap_done;
  input PE_wrapper_140__ap_idle;
  output PE_wrapper_141__ap_start;
  input PE_wrapper_141__ap_ready;
  input PE_wrapper_141__ap_done;
  input PE_wrapper_141__ap_idle;
  output PE_wrapper_142__ap_start;
  input PE_wrapper_142__ap_ready;
  input PE_wrapper_142__ap_done;
  input PE_wrapper_142__ap_idle;
  output PE_wrapper_143__ap_start;
  input PE_wrapper_143__ap_ready;
  input PE_wrapper_143__ap_done;
  input PE_wrapper_143__ap_idle;
  output PE_wrapper_144__ap_start;
  input PE_wrapper_144__ap_ready;
  input PE_wrapper_144__ap_done;
  input PE_wrapper_144__ap_idle;
  output PE_wrapper_145__ap_start;
  input PE_wrapper_145__ap_ready;
  input PE_wrapper_145__ap_done;
  input PE_wrapper_145__ap_idle;
  output PE_wrapper_146__ap_start;
  input PE_wrapper_146__ap_ready;
  input PE_wrapper_146__ap_done;
  input PE_wrapper_146__ap_idle;
  output PE_wrapper_147__ap_start;
  input PE_wrapper_147__ap_ready;
  input PE_wrapper_147__ap_done;
  input PE_wrapper_147__ap_idle;
  output PE_wrapper_148__ap_start;
  input PE_wrapper_148__ap_ready;
  input PE_wrapper_148__ap_done;
  input PE_wrapper_148__ap_idle;
  output PE_wrapper_149__ap_start;
  input PE_wrapper_149__ap_ready;
  input PE_wrapper_149__ap_done;
  input PE_wrapper_149__ap_idle;
  output PE_wrapper_150__ap_start;
  input PE_wrapper_150__ap_ready;
  input PE_wrapper_150__ap_done;
  input PE_wrapper_150__ap_idle;
  output PE_wrapper_151__ap_start;
  input PE_wrapper_151__ap_ready;
  input PE_wrapper_151__ap_done;
  input PE_wrapper_151__ap_idle;
  output PE_wrapper_152__ap_start;
  input PE_wrapper_152__ap_ready;
  input PE_wrapper_152__ap_done;
  input PE_wrapper_152__ap_idle;
  output PE_wrapper_153__ap_start;
  input PE_wrapper_153__ap_ready;
  input PE_wrapper_153__ap_done;
  input PE_wrapper_153__ap_idle;
  output PE_wrapper_154__ap_start;
  input PE_wrapper_154__ap_ready;
  input PE_wrapper_154__ap_done;
  input PE_wrapper_154__ap_idle;
  output PE_wrapper_155__ap_start;
  input PE_wrapper_155__ap_ready;
  input PE_wrapper_155__ap_done;
  input PE_wrapper_155__ap_idle;
  output PE_wrapper_156__ap_start;
  input PE_wrapper_156__ap_ready;
  input PE_wrapper_156__ap_done;
  input PE_wrapper_156__ap_idle;
  output PE_wrapper_157__ap_start;
  input PE_wrapper_157__ap_ready;
  input PE_wrapper_157__ap_done;
  input PE_wrapper_157__ap_idle;
  output PE_wrapper_158__ap_start;
  input PE_wrapper_158__ap_ready;
  input PE_wrapper_158__ap_done;
  input PE_wrapper_158__ap_idle;
  output PE_wrapper_159__ap_start;
  input PE_wrapper_159__ap_ready;
  input PE_wrapper_159__ap_done;
  input PE_wrapper_159__ap_idle;
  output PE_wrapper_160__ap_start;
  input PE_wrapper_160__ap_ready;
  input PE_wrapper_160__ap_done;
  input PE_wrapper_160__ap_idle;
  output PE_wrapper_161__ap_start;
  input PE_wrapper_161__ap_ready;
  input PE_wrapper_161__ap_done;
  input PE_wrapper_161__ap_idle;
  output PE_wrapper_162__ap_start;
  input PE_wrapper_162__ap_ready;
  input PE_wrapper_162__ap_done;
  input PE_wrapper_162__ap_idle;
  output PE_wrapper_163__ap_start;
  input PE_wrapper_163__ap_ready;
  input PE_wrapper_163__ap_done;
  input PE_wrapper_163__ap_idle;
  output PE_wrapper_164__ap_start;
  input PE_wrapper_164__ap_ready;
  input PE_wrapper_164__ap_done;
  input PE_wrapper_164__ap_idle;
  output PE_wrapper_165__ap_start;
  input PE_wrapper_165__ap_ready;
  input PE_wrapper_165__ap_done;
  input PE_wrapper_165__ap_idle;
  output PE_wrapper_166__ap_start;
  input PE_wrapper_166__ap_ready;
  input PE_wrapper_166__ap_done;
  input PE_wrapper_166__ap_idle;
  output PE_wrapper_167__ap_start;
  input PE_wrapper_167__ap_ready;
  input PE_wrapper_167__ap_done;
  input PE_wrapper_167__ap_idle;
  output PE_wrapper_168__ap_start;
  input PE_wrapper_168__ap_ready;
  input PE_wrapper_168__ap_done;
  input PE_wrapper_168__ap_idle;
  output PE_wrapper_169__ap_start;
  input PE_wrapper_169__ap_ready;
  input PE_wrapper_169__ap_done;
  input PE_wrapper_169__ap_idle;
  output PE_wrapper_170__ap_start;
  input PE_wrapper_170__ap_ready;
  input PE_wrapper_170__ap_done;
  input PE_wrapper_170__ap_idle;
  output PE_wrapper_171__ap_start;
  input PE_wrapper_171__ap_ready;
  input PE_wrapper_171__ap_done;
  input PE_wrapper_171__ap_idle;
  output PE_wrapper_172__ap_start;
  input PE_wrapper_172__ap_ready;
  input PE_wrapper_172__ap_done;
  input PE_wrapper_172__ap_idle;
  output PE_wrapper_173__ap_start;
  input PE_wrapper_173__ap_ready;
  input PE_wrapper_173__ap_done;
  input PE_wrapper_173__ap_idle;
  output PE_wrapper_174__ap_start;
  input PE_wrapper_174__ap_ready;
  input PE_wrapper_174__ap_done;
  input PE_wrapper_174__ap_idle;
  output PE_wrapper_175__ap_start;
  input PE_wrapper_175__ap_ready;
  input PE_wrapper_175__ap_done;
  input PE_wrapper_175__ap_idle;
  output PE_wrapper_176__ap_start;
  input PE_wrapper_176__ap_ready;
  input PE_wrapper_176__ap_done;
  input PE_wrapper_176__ap_idle;
  output PE_wrapper_177__ap_start;
  input PE_wrapper_177__ap_ready;
  input PE_wrapper_177__ap_done;
  input PE_wrapper_177__ap_idle;
  output PE_wrapper_178__ap_start;
  input PE_wrapper_178__ap_ready;
  input PE_wrapper_178__ap_done;
  input PE_wrapper_178__ap_idle;
  output PE_wrapper_179__ap_start;
  input PE_wrapper_179__ap_ready;
  input PE_wrapper_179__ap_done;
  input PE_wrapper_179__ap_idle;
  output PE_wrapper_180__ap_start;
  input PE_wrapper_180__ap_ready;
  input PE_wrapper_180__ap_done;
  input PE_wrapper_180__ap_idle;
  output PE_wrapper_181__ap_start;
  input PE_wrapper_181__ap_ready;
  input PE_wrapper_181__ap_done;
  input PE_wrapper_181__ap_idle;
  output PE_wrapper_182__ap_start;
  input PE_wrapper_182__ap_ready;
  input PE_wrapper_182__ap_done;
  input PE_wrapper_182__ap_idle;
  output PE_wrapper_183__ap_start;
  input PE_wrapper_183__ap_ready;
  input PE_wrapper_183__ap_done;
  input PE_wrapper_183__ap_idle;
  output PE_wrapper_184__ap_start;
  input PE_wrapper_184__ap_ready;
  input PE_wrapper_184__ap_done;
  input PE_wrapper_184__ap_idle;
  output PE_wrapper_185__ap_start;
  input PE_wrapper_185__ap_ready;
  input PE_wrapper_185__ap_done;
  input PE_wrapper_185__ap_idle;
  output PE_wrapper_186__ap_start;
  input PE_wrapper_186__ap_ready;
  input PE_wrapper_186__ap_done;
  input PE_wrapper_186__ap_idle;
  output PE_wrapper_187__ap_start;
  input PE_wrapper_187__ap_ready;
  input PE_wrapper_187__ap_done;
  input PE_wrapper_187__ap_idle;
  output PE_wrapper_188__ap_start;
  input PE_wrapper_188__ap_ready;
  input PE_wrapper_188__ap_done;
  input PE_wrapper_188__ap_idle;
  output PE_wrapper_189__ap_start;
  input PE_wrapper_189__ap_ready;
  input PE_wrapper_189__ap_done;
  input PE_wrapper_189__ap_idle;
  output PE_wrapper_190__ap_start;
  input PE_wrapper_190__ap_ready;
  input PE_wrapper_190__ap_done;
  input PE_wrapper_190__ap_idle;
  output PE_wrapper_191__ap_start;
  input PE_wrapper_191__ap_ready;
  input PE_wrapper_191__ap_done;
  input PE_wrapper_191__ap_idle;
  output PE_wrapper_192__ap_start;
  input PE_wrapper_192__ap_ready;
  input PE_wrapper_192__ap_done;
  input PE_wrapper_192__ap_idle;
  output PE_wrapper_193__ap_start;
  input PE_wrapper_193__ap_ready;
  input PE_wrapper_193__ap_done;
  input PE_wrapper_193__ap_idle;
  output PE_wrapper_194__ap_start;
  input PE_wrapper_194__ap_ready;
  input PE_wrapper_194__ap_done;
  input PE_wrapper_194__ap_idle;
  output PE_wrapper_195__ap_start;
  input PE_wrapper_195__ap_ready;
  input PE_wrapper_195__ap_done;
  input PE_wrapper_195__ap_idle;
  output PE_wrapper_196__ap_start;
  input PE_wrapper_196__ap_ready;
  input PE_wrapper_196__ap_done;
  input PE_wrapper_196__ap_idle;
  output PE_wrapper_197__ap_start;
  input PE_wrapper_197__ap_ready;
  input PE_wrapper_197__ap_done;
  input PE_wrapper_197__ap_idle;
  output PE_wrapper_198__ap_start;
  input PE_wrapper_198__ap_ready;
  input PE_wrapper_198__ap_done;
  input PE_wrapper_198__ap_idle;
  output PE_wrapper_199__ap_start;
  input PE_wrapper_199__ap_ready;
  input PE_wrapper_199__ap_done;
  input PE_wrapper_199__ap_idle;
  output PE_wrapper_200__ap_start;
  input PE_wrapper_200__ap_ready;
  input PE_wrapper_200__ap_done;
  input PE_wrapper_200__ap_idle;
  output PE_wrapper_201__ap_start;
  input PE_wrapper_201__ap_ready;
  input PE_wrapper_201__ap_done;
  input PE_wrapper_201__ap_idle;
  output PE_wrapper_202__ap_start;
  input PE_wrapper_202__ap_ready;
  input PE_wrapper_202__ap_done;
  input PE_wrapper_202__ap_idle;
  output PE_wrapper_203__ap_start;
  input PE_wrapper_203__ap_ready;
  input PE_wrapper_203__ap_done;
  input PE_wrapper_203__ap_idle;
  output PE_wrapper_204__ap_start;
  input PE_wrapper_204__ap_ready;
  input PE_wrapper_204__ap_done;
  input PE_wrapper_204__ap_idle;
  output PE_wrapper_205__ap_start;
  input PE_wrapper_205__ap_ready;
  input PE_wrapper_205__ap_done;
  input PE_wrapper_205__ap_idle;
  output PE_wrapper_206__ap_start;
  input PE_wrapper_206__ap_ready;
  input PE_wrapper_206__ap_done;
  input PE_wrapper_206__ap_idle;
  output PE_wrapper_207__ap_start;
  input PE_wrapper_207__ap_ready;
  input PE_wrapper_207__ap_done;
  input PE_wrapper_207__ap_idle;
  output PE_wrapper_208__ap_start;
  input PE_wrapper_208__ap_ready;
  input PE_wrapper_208__ap_done;
  input PE_wrapper_208__ap_idle;
  output PE_wrapper_209__ap_start;
  input PE_wrapper_209__ap_ready;
  input PE_wrapper_209__ap_done;
  input PE_wrapper_209__ap_idle;
  output PE_wrapper_210__ap_start;
  input PE_wrapper_210__ap_ready;
  input PE_wrapper_210__ap_done;
  input PE_wrapper_210__ap_idle;
  output PE_wrapper_211__ap_start;
  input PE_wrapper_211__ap_ready;
  input PE_wrapper_211__ap_done;
  input PE_wrapper_211__ap_idle;
  output PE_wrapper_212__ap_start;
  input PE_wrapper_212__ap_ready;
  input PE_wrapper_212__ap_done;
  input PE_wrapper_212__ap_idle;
  output PE_wrapper_213__ap_start;
  input PE_wrapper_213__ap_ready;
  input PE_wrapper_213__ap_done;
  input PE_wrapper_213__ap_idle;
  output PE_wrapper_214__ap_start;
  input PE_wrapper_214__ap_ready;
  input PE_wrapper_214__ap_done;
  input PE_wrapper_214__ap_idle;
  output PE_wrapper_215__ap_start;
  input PE_wrapper_215__ap_ready;
  input PE_wrapper_215__ap_done;
  input PE_wrapper_215__ap_idle;
  output PE_wrapper_216__ap_start;
  input PE_wrapper_216__ap_ready;
  input PE_wrapper_216__ap_done;
  input PE_wrapper_216__ap_idle;
  output PE_wrapper_217__ap_start;
  input PE_wrapper_217__ap_ready;
  input PE_wrapper_217__ap_done;
  input PE_wrapper_217__ap_idle;
  output PE_wrapper_218__ap_start;
  input PE_wrapper_218__ap_ready;
  input PE_wrapper_218__ap_done;
  input PE_wrapper_218__ap_idle;
  output PE_wrapper_219__ap_start;
  input PE_wrapper_219__ap_ready;
  input PE_wrapper_219__ap_done;
  input PE_wrapper_219__ap_idle;
  output PE_wrapper_220__ap_start;
  input PE_wrapper_220__ap_ready;
  input PE_wrapper_220__ap_done;
  input PE_wrapper_220__ap_idle;
  output PE_wrapper_221__ap_start;
  input PE_wrapper_221__ap_ready;
  input PE_wrapper_221__ap_done;
  input PE_wrapper_221__ap_idle;
  output PE_wrapper_222__ap_start;
  input PE_wrapper_222__ap_ready;
  input PE_wrapper_222__ap_done;
  input PE_wrapper_222__ap_idle;
  output PE_wrapper_223__ap_start;
  input PE_wrapper_223__ap_ready;
  input PE_wrapper_223__ap_done;
  input PE_wrapper_223__ap_idle;
  output PE_wrapper_224__ap_start;
  input PE_wrapper_224__ap_ready;
  input PE_wrapper_224__ap_done;
  input PE_wrapper_224__ap_idle;
  output PE_wrapper_225__ap_start;
  input PE_wrapper_225__ap_ready;
  input PE_wrapper_225__ap_done;
  input PE_wrapper_225__ap_idle;
  output PE_wrapper_226__ap_start;
  input PE_wrapper_226__ap_ready;
  input PE_wrapper_226__ap_done;
  input PE_wrapper_226__ap_idle;
  output PE_wrapper_227__ap_start;
  input PE_wrapper_227__ap_ready;
  input PE_wrapper_227__ap_done;
  input PE_wrapper_227__ap_idle;
  output PE_wrapper_228__ap_start;
  input PE_wrapper_228__ap_ready;
  input PE_wrapper_228__ap_done;
  input PE_wrapper_228__ap_idle;
  output PE_wrapper_229__ap_start;
  input PE_wrapper_229__ap_ready;
  input PE_wrapper_229__ap_done;
  input PE_wrapper_229__ap_idle;
  output PE_wrapper_230__ap_start;
  input PE_wrapper_230__ap_ready;
  input PE_wrapper_230__ap_done;
  input PE_wrapper_230__ap_idle;
  output PE_wrapper_231__ap_start;
  input PE_wrapper_231__ap_ready;
  input PE_wrapper_231__ap_done;
  input PE_wrapper_231__ap_idle;
  output PE_wrapper_232__ap_start;
  input PE_wrapper_232__ap_ready;
  input PE_wrapper_232__ap_done;
  input PE_wrapper_232__ap_idle;
  output PE_wrapper_233__ap_start;
  input PE_wrapper_233__ap_ready;
  input PE_wrapper_233__ap_done;
  input PE_wrapper_233__ap_idle;
  output PE_wrapper_234__ap_start;
  input PE_wrapper_234__ap_ready;
  input PE_wrapper_234__ap_done;
  input PE_wrapper_234__ap_idle;
  output PE_wrapper_235__ap_start;
  input PE_wrapper_235__ap_ready;
  input PE_wrapper_235__ap_done;
  input PE_wrapper_235__ap_idle;
  output PE_wrapper_236__ap_start;
  input PE_wrapper_236__ap_ready;
  input PE_wrapper_236__ap_done;
  input PE_wrapper_236__ap_idle;
  output PE_wrapper_237__ap_start;
  input PE_wrapper_237__ap_ready;
  input PE_wrapper_237__ap_done;
  input PE_wrapper_237__ap_idle;
  output PE_wrapper_238__ap_start;
  input PE_wrapper_238__ap_ready;
  input PE_wrapper_238__ap_done;
  input PE_wrapper_238__ap_idle;
  output PE_wrapper_239__ap_start;
  input PE_wrapper_239__ap_ready;
  input PE_wrapper_239__ap_done;
  input PE_wrapper_239__ap_idle;
  output PE_wrapper_240__ap_start;
  input PE_wrapper_240__ap_ready;
  input PE_wrapper_240__ap_done;
  input PE_wrapper_240__ap_idle;
  output PE_wrapper_241__ap_start;
  input PE_wrapper_241__ap_ready;
  input PE_wrapper_241__ap_done;
  input PE_wrapper_241__ap_idle;
  output PE_wrapper_242__ap_start;
  input PE_wrapper_242__ap_ready;
  input PE_wrapper_242__ap_done;
  input PE_wrapper_242__ap_idle;
  output PE_wrapper_243__ap_start;
  input PE_wrapper_243__ap_ready;
  input PE_wrapper_243__ap_done;
  input PE_wrapper_243__ap_idle;
  output PE_wrapper_244__ap_start;
  input PE_wrapper_244__ap_ready;
  input PE_wrapper_244__ap_done;
  input PE_wrapper_244__ap_idle;
  output PE_wrapper_245__ap_start;
  input PE_wrapper_245__ap_ready;
  input PE_wrapper_245__ap_done;
  input PE_wrapper_245__ap_idle;
  output PE_wrapper_246__ap_start;
  input PE_wrapper_246__ap_ready;
  input PE_wrapper_246__ap_done;
  input PE_wrapper_246__ap_idle;
  output PE_wrapper_247__ap_start;
  input PE_wrapper_247__ap_ready;
  input PE_wrapper_247__ap_done;
  input PE_wrapper_247__ap_idle;
  output PE_wrapper_248__ap_start;
  input PE_wrapper_248__ap_ready;
  input PE_wrapper_248__ap_done;
  input PE_wrapper_248__ap_idle;
  output PE_wrapper_249__ap_start;
  input PE_wrapper_249__ap_ready;
  input PE_wrapper_249__ap_done;
  input PE_wrapper_249__ap_idle;
  output PE_wrapper_250__ap_start;
  input PE_wrapper_250__ap_ready;
  input PE_wrapper_250__ap_done;
  input PE_wrapper_250__ap_idle;
  output PE_wrapper_251__ap_start;
  input PE_wrapper_251__ap_ready;
  input PE_wrapper_251__ap_done;
  input PE_wrapper_251__ap_idle;
  output PE_wrapper_252__ap_start;
  input PE_wrapper_252__ap_ready;
  input PE_wrapper_252__ap_done;
  input PE_wrapper_252__ap_idle;
  output PE_wrapper_253__ap_start;
  input PE_wrapper_253__ap_ready;
  input PE_wrapper_253__ap_done;
  input PE_wrapper_253__ap_idle;
  output PE_wrapper_254__ap_start;
  input PE_wrapper_254__ap_ready;
  input PE_wrapper_254__ap_done;
  input PE_wrapper_254__ap_idle;
  output PE_wrapper_255__ap_start;
  input PE_wrapper_255__ap_ready;
  input PE_wrapper_255__ap_done;
  input PE_wrapper_255__ap_idle;
  output PE_wrapper_256__ap_start;
  input PE_wrapper_256__ap_ready;
  input PE_wrapper_256__ap_done;
  input PE_wrapper_256__ap_idle;
  output PE_wrapper_257__ap_start;
  input PE_wrapper_257__ap_ready;
  input PE_wrapper_257__ap_done;
  input PE_wrapper_257__ap_idle;
  output PE_wrapper_258__ap_start;
  input PE_wrapper_258__ap_ready;
  input PE_wrapper_258__ap_done;
  input PE_wrapper_258__ap_idle;
  output PE_wrapper_259__ap_start;
  input PE_wrapper_259__ap_ready;
  input PE_wrapper_259__ap_done;
  input PE_wrapper_259__ap_idle;
  output PE_wrapper_260__ap_start;
  input PE_wrapper_260__ap_ready;
  input PE_wrapper_260__ap_done;
  input PE_wrapper_260__ap_idle;
  output PE_wrapper_261__ap_start;
  input PE_wrapper_261__ap_ready;
  input PE_wrapper_261__ap_done;
  input PE_wrapper_261__ap_idle;
  output PE_wrapper_262__ap_start;
  input PE_wrapper_262__ap_ready;
  input PE_wrapper_262__ap_done;
  input PE_wrapper_262__ap_idle;
  output PE_wrapper_263__ap_start;
  input PE_wrapper_263__ap_ready;
  input PE_wrapper_263__ap_done;
  input PE_wrapper_263__ap_idle;
  output PE_wrapper_264__ap_start;
  input PE_wrapper_264__ap_ready;
  input PE_wrapper_264__ap_done;
  input PE_wrapper_264__ap_idle;
  output PE_wrapper_265__ap_start;
  input PE_wrapper_265__ap_ready;
  input PE_wrapper_265__ap_done;
  input PE_wrapper_265__ap_idle;
  output PE_wrapper_266__ap_start;
  input PE_wrapper_266__ap_ready;
  input PE_wrapper_266__ap_done;
  input PE_wrapper_266__ap_idle;
  output PE_wrapper_267__ap_start;
  input PE_wrapper_267__ap_ready;
  input PE_wrapper_267__ap_done;
  input PE_wrapper_267__ap_idle;
  output PE_wrapper_268__ap_start;
  input PE_wrapper_268__ap_ready;
  input PE_wrapper_268__ap_done;
  input PE_wrapper_268__ap_idle;
  output PE_wrapper_269__ap_start;
  input PE_wrapper_269__ap_ready;
  input PE_wrapper_269__ap_done;
  input PE_wrapper_269__ap_idle;
  output PE_wrapper_270__ap_start;
  input PE_wrapper_270__ap_ready;
  input PE_wrapper_270__ap_done;
  input PE_wrapper_270__ap_idle;
  output PE_wrapper_271__ap_start;
  input PE_wrapper_271__ap_ready;
  input PE_wrapper_271__ap_done;
  input PE_wrapper_271__ap_idle;
  output PE_wrapper_272__ap_start;
  input PE_wrapper_272__ap_ready;
  input PE_wrapper_272__ap_done;
  input PE_wrapper_272__ap_idle;
  output PE_wrapper_273__ap_start;
  input PE_wrapper_273__ap_ready;
  input PE_wrapper_273__ap_done;
  input PE_wrapper_273__ap_idle;
  output PE_wrapper_274__ap_start;
  input PE_wrapper_274__ap_ready;
  input PE_wrapper_274__ap_done;
  input PE_wrapper_274__ap_idle;
  output PE_wrapper_275__ap_start;
  input PE_wrapper_275__ap_ready;
  input PE_wrapper_275__ap_done;
  input PE_wrapper_275__ap_idle;
  output PE_wrapper_276__ap_start;
  input PE_wrapper_276__ap_ready;
  input PE_wrapper_276__ap_done;
  input PE_wrapper_276__ap_idle;
  output PE_wrapper_277__ap_start;
  input PE_wrapper_277__ap_ready;
  input PE_wrapper_277__ap_done;
  input PE_wrapper_277__ap_idle;
  output PE_wrapper_278__ap_start;
  input PE_wrapper_278__ap_ready;
  input PE_wrapper_278__ap_done;
  input PE_wrapper_278__ap_idle;
  output PE_wrapper_279__ap_start;
  input PE_wrapper_279__ap_ready;
  input PE_wrapper_279__ap_done;
  input PE_wrapper_279__ap_idle;
  output PE_wrapper_280__ap_start;
  input PE_wrapper_280__ap_ready;
  input PE_wrapper_280__ap_done;
  input PE_wrapper_280__ap_idle;
  output PE_wrapper_281__ap_start;
  input PE_wrapper_281__ap_ready;
  input PE_wrapper_281__ap_done;
  input PE_wrapper_281__ap_idle;
  output PE_wrapper_282__ap_start;
  input PE_wrapper_282__ap_ready;
  input PE_wrapper_282__ap_done;
  input PE_wrapper_282__ap_idle;
  output PE_wrapper_283__ap_start;
  input PE_wrapper_283__ap_ready;
  input PE_wrapper_283__ap_done;
  input PE_wrapper_283__ap_idle;
  output PE_wrapper_284__ap_start;
  input PE_wrapper_284__ap_ready;
  input PE_wrapper_284__ap_done;
  input PE_wrapper_284__ap_idle;
  output PE_wrapper_285__ap_start;
  input PE_wrapper_285__ap_ready;
  input PE_wrapper_285__ap_done;
  input PE_wrapper_285__ap_idle;
  output PE_wrapper_286__ap_start;
  input PE_wrapper_286__ap_ready;
  input PE_wrapper_286__ap_done;
  input PE_wrapper_286__ap_idle;
  output PE_wrapper_287__ap_start;
  input PE_wrapper_287__ap_ready;
  input PE_wrapper_287__ap_done;
  input PE_wrapper_287__ap_idle;
  output PE_wrapper_288__ap_start;
  input PE_wrapper_288__ap_ready;
  input PE_wrapper_288__ap_done;
  input PE_wrapper_288__ap_idle;
  output PE_wrapper_289__ap_start;
  input PE_wrapper_289__ap_ready;
  input PE_wrapper_289__ap_done;
  input PE_wrapper_289__ap_idle;
  output PE_wrapper_290__ap_start;
  input PE_wrapper_290__ap_ready;
  input PE_wrapper_290__ap_done;
  input PE_wrapper_290__ap_idle;
  output PE_wrapper_291__ap_start;
  input PE_wrapper_291__ap_ready;
  input PE_wrapper_291__ap_done;
  input PE_wrapper_291__ap_idle;
  output PE_wrapper_292__ap_start;
  input PE_wrapper_292__ap_ready;
  input PE_wrapper_292__ap_done;
  input PE_wrapper_292__ap_idle;
  output PE_wrapper_293__ap_start;
  input PE_wrapper_293__ap_ready;
  input PE_wrapper_293__ap_done;
  input PE_wrapper_293__ap_idle;
  output PE_wrapper_294__ap_start;
  input PE_wrapper_294__ap_ready;
  input PE_wrapper_294__ap_done;
  input PE_wrapper_294__ap_idle;
  output PE_wrapper_295__ap_start;
  input PE_wrapper_295__ap_ready;
  input PE_wrapper_295__ap_done;
  input PE_wrapper_295__ap_idle;
  output PE_wrapper_296__ap_start;
  input PE_wrapper_296__ap_ready;
  input PE_wrapper_296__ap_done;
  input PE_wrapper_296__ap_idle;
  output PE_wrapper_297__ap_start;
  input PE_wrapper_297__ap_ready;
  input PE_wrapper_297__ap_done;
  input PE_wrapper_297__ap_idle;
  output PE_wrapper_298__ap_start;
  input PE_wrapper_298__ap_ready;
  input PE_wrapper_298__ap_done;
  input PE_wrapper_298__ap_idle;
  output PE_wrapper_299__ap_start;
  input PE_wrapper_299__ap_ready;
  input PE_wrapper_299__ap_done;
  input PE_wrapper_299__ap_idle;
  output PE_wrapper_300__ap_start;
  input PE_wrapper_300__ap_ready;
  input PE_wrapper_300__ap_done;
  input PE_wrapper_300__ap_idle;
  output PE_wrapper_301__ap_start;
  input PE_wrapper_301__ap_ready;
  input PE_wrapper_301__ap_done;
  input PE_wrapper_301__ap_idle;
  output PE_wrapper_302__ap_start;
  input PE_wrapper_302__ap_ready;
  input PE_wrapper_302__ap_done;
  input PE_wrapper_302__ap_idle;
  output PE_wrapper_303__ap_start;
  input PE_wrapper_303__ap_ready;
  input PE_wrapper_303__ap_done;
  input PE_wrapper_303__ap_idle;
  output PE_wrapper_304__ap_start;
  input PE_wrapper_304__ap_ready;
  input PE_wrapper_304__ap_done;
  input PE_wrapper_304__ap_idle;
  output PE_wrapper_305__ap_start;
  input PE_wrapper_305__ap_ready;
  input PE_wrapper_305__ap_done;
  input PE_wrapper_305__ap_idle;
  wire A_IO_L2_in_0__ap_start_global__q0;
  wire A_IO_L2_in_0__is_done__q0;
  wire A_IO_L2_in_0__ap_done_global__q0;
  wire A_IO_L2_in_0__ap_start;
  wire A_IO_L2_in_0__ap_ready;
  wire A_IO_L2_in_0__ap_done;
  wire A_IO_L2_in_0__ap_idle;
  reg [1:0] A_IO_L2_in_0__state;
  wire A_IO_L2_in_1__ap_start_global__q0;
  wire A_IO_L2_in_1__is_done__q0;
  wire A_IO_L2_in_1__ap_done_global__q0;
  wire A_IO_L2_in_1__ap_start;
  wire A_IO_L2_in_1__ap_ready;
  wire A_IO_L2_in_1__ap_done;
  wire A_IO_L2_in_1__ap_idle;
  reg [1:0] A_IO_L2_in_1__state;
  wire A_IO_L2_in_2__ap_start_global__q0;
  wire A_IO_L2_in_2__is_done__q0;
  wire A_IO_L2_in_2__ap_done_global__q0;
  wire A_IO_L2_in_2__ap_start;
  wire A_IO_L2_in_2__ap_ready;
  wire A_IO_L2_in_2__ap_done;
  wire A_IO_L2_in_2__ap_idle;
  reg [1:0] A_IO_L2_in_2__state;
  wire A_IO_L2_in_3__ap_start_global__q0;
  wire A_IO_L2_in_3__is_done__q0;
  wire A_IO_L2_in_3__ap_done_global__q0;
  wire A_IO_L2_in_3__ap_start;
  wire A_IO_L2_in_3__ap_ready;
  wire A_IO_L2_in_3__ap_done;
  wire A_IO_L2_in_3__ap_idle;
  reg [1:0] A_IO_L2_in_3__state;
  wire A_IO_L2_in_4__ap_start_global__q0;
  wire A_IO_L2_in_4__is_done__q0;
  wire A_IO_L2_in_4__ap_done_global__q0;
  wire A_IO_L2_in_4__ap_start;
  wire A_IO_L2_in_4__ap_ready;
  wire A_IO_L2_in_4__ap_done;
  wire A_IO_L2_in_4__ap_idle;
  reg [1:0] A_IO_L2_in_4__state;
  wire A_IO_L2_in_5__ap_start_global__q0;
  wire A_IO_L2_in_5__is_done__q0;
  wire A_IO_L2_in_5__ap_done_global__q0;
  wire A_IO_L2_in_5__ap_start;
  wire A_IO_L2_in_5__ap_ready;
  wire A_IO_L2_in_5__ap_done;
  wire A_IO_L2_in_5__ap_idle;
  reg [1:0] A_IO_L2_in_5__state;
  wire A_IO_L2_in_6__ap_start_global__q0;
  wire A_IO_L2_in_6__is_done__q0;
  wire A_IO_L2_in_6__ap_done_global__q0;
  wire A_IO_L2_in_6__ap_start;
  wire A_IO_L2_in_6__ap_ready;
  wire A_IO_L2_in_6__ap_done;
  wire A_IO_L2_in_6__ap_idle;
  reg [1:0] A_IO_L2_in_6__state;
  wire A_IO_L2_in_7__ap_start_global__q0;
  wire A_IO_L2_in_7__is_done__q0;
  wire A_IO_L2_in_7__ap_done_global__q0;
  wire A_IO_L2_in_7__ap_start;
  wire A_IO_L2_in_7__ap_ready;
  wire A_IO_L2_in_7__ap_done;
  wire A_IO_L2_in_7__ap_idle;
  reg [1:0] A_IO_L2_in_7__state;
  wire A_IO_L2_in_8__ap_start_global__q0;
  wire A_IO_L2_in_8__is_done__q0;
  wire A_IO_L2_in_8__ap_done_global__q0;
  wire A_IO_L2_in_8__ap_start;
  wire A_IO_L2_in_8__ap_ready;
  wire A_IO_L2_in_8__ap_done;
  wire A_IO_L2_in_8__ap_idle;
  reg [1:0] A_IO_L2_in_8__state;
  wire A_IO_L2_in_9__ap_start_global__q0;
  wire A_IO_L2_in_9__is_done__q0;
  wire A_IO_L2_in_9__ap_done_global__q0;
  wire A_IO_L2_in_9__ap_start;
  wire A_IO_L2_in_9__ap_ready;
  wire A_IO_L2_in_9__ap_done;
  wire A_IO_L2_in_9__ap_idle;
  reg [1:0] A_IO_L2_in_9__state;
  wire A_IO_L2_in_10__ap_start_global__q0;
  wire A_IO_L2_in_10__is_done__q0;
  wire A_IO_L2_in_10__ap_done_global__q0;
  wire A_IO_L2_in_10__ap_start;
  wire A_IO_L2_in_10__ap_ready;
  wire A_IO_L2_in_10__ap_done;
  wire A_IO_L2_in_10__ap_idle;
  reg [1:0] A_IO_L2_in_10__state;
  wire A_IO_L2_in_11__ap_start_global__q0;
  wire A_IO_L2_in_11__is_done__q0;
  wire A_IO_L2_in_11__ap_done_global__q0;
  wire A_IO_L2_in_11__ap_start;
  wire A_IO_L2_in_11__ap_ready;
  wire A_IO_L2_in_11__ap_done;
  wire A_IO_L2_in_11__ap_idle;
  reg [1:0] A_IO_L2_in_11__state;
  wire A_IO_L2_in_12__ap_start_global__q0;
  wire A_IO_L2_in_12__is_done__q0;
  wire A_IO_L2_in_12__ap_done_global__q0;
  wire A_IO_L2_in_12__ap_start;
  wire A_IO_L2_in_12__ap_ready;
  wire A_IO_L2_in_12__ap_done;
  wire A_IO_L2_in_12__ap_idle;
  reg [1:0] A_IO_L2_in_12__state;
  wire A_IO_L2_in_13__ap_start_global__q0;
  wire A_IO_L2_in_13__is_done__q0;
  wire A_IO_L2_in_13__ap_done_global__q0;
  wire A_IO_L2_in_13__ap_start;
  wire A_IO_L2_in_13__ap_ready;
  wire A_IO_L2_in_13__ap_done;
  wire A_IO_L2_in_13__ap_idle;
  reg [1:0] A_IO_L2_in_13__state;
  wire A_IO_L2_in_14__ap_start_global__q0;
  wire A_IO_L2_in_14__is_done__q0;
  wire A_IO_L2_in_14__ap_done_global__q0;
  wire A_IO_L2_in_14__ap_start;
  wire A_IO_L2_in_14__ap_ready;
  wire A_IO_L2_in_14__ap_done;
  wire A_IO_L2_in_14__ap_idle;
  reg [1:0] A_IO_L2_in_14__state;
  wire A_IO_L2_in_15__ap_start_global__q0;
  wire A_IO_L2_in_15__is_done__q0;
  wire A_IO_L2_in_15__ap_done_global__q0;
  wire A_IO_L2_in_15__ap_start;
  wire A_IO_L2_in_15__ap_ready;
  wire A_IO_L2_in_15__ap_done;
  wire A_IO_L2_in_15__ap_idle;
  reg [1:0] A_IO_L2_in_15__state;
  wire A_IO_L2_in_16__ap_start_global__q0;
  wire A_IO_L2_in_16__is_done__q0;
  wire A_IO_L2_in_16__ap_done_global__q0;
  wire A_IO_L2_in_16__ap_start;
  wire A_IO_L2_in_16__ap_ready;
  wire A_IO_L2_in_16__ap_done;
  wire A_IO_L2_in_16__ap_idle;
  reg [1:0] A_IO_L2_in_16__state;
  wire A_IO_L2_in_boundary_0__ap_start_global__q0;
  wire A_IO_L2_in_boundary_0__is_done__q0;
  wire A_IO_L2_in_boundary_0__ap_done_global__q0;
  wire A_IO_L2_in_boundary_0__ap_start;
  wire A_IO_L2_in_boundary_0__ap_ready;
  wire A_IO_L2_in_boundary_0__ap_done;
  wire A_IO_L2_in_boundary_0__ap_idle;
  reg [1:0] A_IO_L2_in_boundary_0__state;
  wire A_IO_L3_in_0__ap_start_global__q0;
  wire A_IO_L3_in_0__is_done__q0;
  wire A_IO_L3_in_0__ap_done_global__q0;
  wire A_IO_L3_in_0__ap_start;
  wire A_IO_L3_in_0__ap_ready;
  wire A_IO_L3_in_0__ap_done;
  wire A_IO_L3_in_0__ap_idle;
  reg [1:0] A_IO_L3_in_0__state;
  wire [63:0] A_IO_L3_in_serialize_0___A__q0;
  wire A_IO_L3_in_serialize_0__ap_start_global__q0;
  wire A_IO_L3_in_serialize_0__is_done__q0;
  wire A_IO_L3_in_serialize_0__ap_done_global__q0;
  wire A_IO_L3_in_serialize_0__ap_start;
  wire A_IO_L3_in_serialize_0__ap_ready;
  wire A_IO_L3_in_serialize_0__ap_done;
  wire A_IO_L3_in_serialize_0__ap_idle;
  reg [1:0] A_IO_L3_in_serialize_0__state;
  wire A_PE_dummy_in_0__ap_start_global__q0;
  wire A_PE_dummy_in_0__is_done__q0;
  wire A_PE_dummy_in_0__ap_done_global__q0;
  wire A_PE_dummy_in_0__ap_start;
  wire A_PE_dummy_in_0__ap_ready;
  wire A_PE_dummy_in_0__ap_done;
  wire A_PE_dummy_in_0__ap_idle;
  reg [1:0] A_PE_dummy_in_0__state;
  wire A_PE_dummy_in_1__ap_start_global__q0;
  wire A_PE_dummy_in_1__is_done__q0;
  wire A_PE_dummy_in_1__ap_done_global__q0;
  wire A_PE_dummy_in_1__ap_start;
  wire A_PE_dummy_in_1__ap_ready;
  wire A_PE_dummy_in_1__ap_done;
  wire A_PE_dummy_in_1__ap_idle;
  reg [1:0] A_PE_dummy_in_1__state;
  wire A_PE_dummy_in_2__ap_start_global__q0;
  wire A_PE_dummy_in_2__is_done__q0;
  wire A_PE_dummy_in_2__ap_done_global__q0;
  wire A_PE_dummy_in_2__ap_start;
  wire A_PE_dummy_in_2__ap_ready;
  wire A_PE_dummy_in_2__ap_done;
  wire A_PE_dummy_in_2__ap_idle;
  reg [1:0] A_PE_dummy_in_2__state;
  wire A_PE_dummy_in_3__ap_start_global__q0;
  wire A_PE_dummy_in_3__is_done__q0;
  wire A_PE_dummy_in_3__ap_done_global__q0;
  wire A_PE_dummy_in_3__ap_start;
  wire A_PE_dummy_in_3__ap_ready;
  wire A_PE_dummy_in_3__ap_done;
  wire A_PE_dummy_in_3__ap_idle;
  reg [1:0] A_PE_dummy_in_3__state;
  wire A_PE_dummy_in_4__ap_start_global__q0;
  wire A_PE_dummy_in_4__is_done__q0;
  wire A_PE_dummy_in_4__ap_done_global__q0;
  wire A_PE_dummy_in_4__ap_start;
  wire A_PE_dummy_in_4__ap_ready;
  wire A_PE_dummy_in_4__ap_done;
  wire A_PE_dummy_in_4__ap_idle;
  reg [1:0] A_PE_dummy_in_4__state;
  wire A_PE_dummy_in_5__ap_start_global__q0;
  wire A_PE_dummy_in_5__is_done__q0;
  wire A_PE_dummy_in_5__ap_done_global__q0;
  wire A_PE_dummy_in_5__ap_start;
  wire A_PE_dummy_in_5__ap_ready;
  wire A_PE_dummy_in_5__ap_done;
  wire A_PE_dummy_in_5__ap_idle;
  reg [1:0] A_PE_dummy_in_5__state;
  wire A_PE_dummy_in_6__ap_start_global__q0;
  wire A_PE_dummy_in_6__is_done__q0;
  wire A_PE_dummy_in_6__ap_done_global__q0;
  wire A_PE_dummy_in_6__ap_start;
  wire A_PE_dummy_in_6__ap_ready;
  wire A_PE_dummy_in_6__ap_done;
  wire A_PE_dummy_in_6__ap_idle;
  reg [1:0] A_PE_dummy_in_6__state;
  wire A_PE_dummy_in_7__ap_start_global__q0;
  wire A_PE_dummy_in_7__is_done__q0;
  wire A_PE_dummy_in_7__ap_done_global__q0;
  wire A_PE_dummy_in_7__ap_start;
  wire A_PE_dummy_in_7__ap_ready;
  wire A_PE_dummy_in_7__ap_done;
  wire A_PE_dummy_in_7__ap_idle;
  reg [1:0] A_PE_dummy_in_7__state;
  wire A_PE_dummy_in_8__ap_start_global__q0;
  wire A_PE_dummy_in_8__is_done__q0;
  wire A_PE_dummy_in_8__ap_done_global__q0;
  wire A_PE_dummy_in_8__ap_start;
  wire A_PE_dummy_in_8__ap_ready;
  wire A_PE_dummy_in_8__ap_done;
  wire A_PE_dummy_in_8__ap_idle;
  reg [1:0] A_PE_dummy_in_8__state;
  wire A_PE_dummy_in_9__ap_start_global__q0;
  wire A_PE_dummy_in_9__is_done__q0;
  wire A_PE_dummy_in_9__ap_done_global__q0;
  wire A_PE_dummy_in_9__ap_start;
  wire A_PE_dummy_in_9__ap_ready;
  wire A_PE_dummy_in_9__ap_done;
  wire A_PE_dummy_in_9__ap_idle;
  reg [1:0] A_PE_dummy_in_9__state;
  wire A_PE_dummy_in_10__ap_start_global__q0;
  wire A_PE_dummy_in_10__is_done__q0;
  wire A_PE_dummy_in_10__ap_done_global__q0;
  wire A_PE_dummy_in_10__ap_start;
  wire A_PE_dummy_in_10__ap_ready;
  wire A_PE_dummy_in_10__ap_done;
  wire A_PE_dummy_in_10__ap_idle;
  reg [1:0] A_PE_dummy_in_10__state;
  wire A_PE_dummy_in_11__ap_start_global__q0;
  wire A_PE_dummy_in_11__is_done__q0;
  wire A_PE_dummy_in_11__ap_done_global__q0;
  wire A_PE_dummy_in_11__ap_start;
  wire A_PE_dummy_in_11__ap_ready;
  wire A_PE_dummy_in_11__ap_done;
  wire A_PE_dummy_in_11__ap_idle;
  reg [1:0] A_PE_dummy_in_11__state;
  wire A_PE_dummy_in_12__ap_start_global__q0;
  wire A_PE_dummy_in_12__is_done__q0;
  wire A_PE_dummy_in_12__ap_done_global__q0;
  wire A_PE_dummy_in_12__ap_start;
  wire A_PE_dummy_in_12__ap_ready;
  wire A_PE_dummy_in_12__ap_done;
  wire A_PE_dummy_in_12__ap_idle;
  reg [1:0] A_PE_dummy_in_12__state;
  wire A_PE_dummy_in_13__ap_start_global__q0;
  wire A_PE_dummy_in_13__is_done__q0;
  wire A_PE_dummy_in_13__ap_done_global__q0;
  wire A_PE_dummy_in_13__ap_start;
  wire A_PE_dummy_in_13__ap_ready;
  wire A_PE_dummy_in_13__ap_done;
  wire A_PE_dummy_in_13__ap_idle;
  reg [1:0] A_PE_dummy_in_13__state;
  wire A_PE_dummy_in_14__ap_start_global__q0;
  wire A_PE_dummy_in_14__is_done__q0;
  wire A_PE_dummy_in_14__ap_done_global__q0;
  wire A_PE_dummy_in_14__ap_start;
  wire A_PE_dummy_in_14__ap_ready;
  wire A_PE_dummy_in_14__ap_done;
  wire A_PE_dummy_in_14__ap_idle;
  reg [1:0] A_PE_dummy_in_14__state;
  wire A_PE_dummy_in_15__ap_start_global__q0;
  wire A_PE_dummy_in_15__is_done__q0;
  wire A_PE_dummy_in_15__ap_done_global__q0;
  wire A_PE_dummy_in_15__ap_start;
  wire A_PE_dummy_in_15__ap_ready;
  wire A_PE_dummy_in_15__ap_done;
  wire A_PE_dummy_in_15__ap_idle;
  reg [1:0] A_PE_dummy_in_15__state;
  wire A_PE_dummy_in_16__ap_start_global__q0;
  wire A_PE_dummy_in_16__is_done__q0;
  wire A_PE_dummy_in_16__ap_done_global__q0;
  wire A_PE_dummy_in_16__ap_start;
  wire A_PE_dummy_in_16__ap_ready;
  wire A_PE_dummy_in_16__ap_done;
  wire A_PE_dummy_in_16__ap_idle;
  reg [1:0] A_PE_dummy_in_16__state;
  wire A_PE_dummy_in_17__ap_start_global__q0;
  wire A_PE_dummy_in_17__is_done__q0;
  wire A_PE_dummy_in_17__ap_done_global__q0;
  wire A_PE_dummy_in_17__ap_start;
  wire A_PE_dummy_in_17__ap_ready;
  wire A_PE_dummy_in_17__ap_done;
  wire A_PE_dummy_in_17__ap_idle;
  reg [1:0] A_PE_dummy_in_17__state;
  wire B_IO_L2_in_0__ap_start_global__q0;
  wire B_IO_L2_in_0__is_done__q0;
  wire B_IO_L2_in_0__ap_done_global__q0;
  wire B_IO_L2_in_0__ap_start;
  wire B_IO_L2_in_0__ap_ready;
  wire B_IO_L2_in_0__ap_done;
  wire B_IO_L2_in_0__ap_idle;
  reg [1:0] B_IO_L2_in_0__state;
  wire B_IO_L2_in_1__ap_start_global__q0;
  wire B_IO_L2_in_1__is_done__q0;
  wire B_IO_L2_in_1__ap_done_global__q0;
  wire B_IO_L2_in_1__ap_start;
  wire B_IO_L2_in_1__ap_ready;
  wire B_IO_L2_in_1__ap_done;
  wire B_IO_L2_in_1__ap_idle;
  reg [1:0] B_IO_L2_in_1__state;
  wire B_IO_L2_in_2__ap_start_global__q0;
  wire B_IO_L2_in_2__is_done__q0;
  wire B_IO_L2_in_2__ap_done_global__q0;
  wire B_IO_L2_in_2__ap_start;
  wire B_IO_L2_in_2__ap_ready;
  wire B_IO_L2_in_2__ap_done;
  wire B_IO_L2_in_2__ap_idle;
  reg [1:0] B_IO_L2_in_2__state;
  wire B_IO_L2_in_3__ap_start_global__q0;
  wire B_IO_L2_in_3__is_done__q0;
  wire B_IO_L2_in_3__ap_done_global__q0;
  wire B_IO_L2_in_3__ap_start;
  wire B_IO_L2_in_3__ap_ready;
  wire B_IO_L2_in_3__ap_done;
  wire B_IO_L2_in_3__ap_idle;
  reg [1:0] B_IO_L2_in_3__state;
  wire B_IO_L2_in_4__ap_start_global__q0;
  wire B_IO_L2_in_4__is_done__q0;
  wire B_IO_L2_in_4__ap_done_global__q0;
  wire B_IO_L2_in_4__ap_start;
  wire B_IO_L2_in_4__ap_ready;
  wire B_IO_L2_in_4__ap_done;
  wire B_IO_L2_in_4__ap_idle;
  reg [1:0] B_IO_L2_in_4__state;
  wire B_IO_L2_in_5__ap_start_global__q0;
  wire B_IO_L2_in_5__is_done__q0;
  wire B_IO_L2_in_5__ap_done_global__q0;
  wire B_IO_L2_in_5__ap_start;
  wire B_IO_L2_in_5__ap_ready;
  wire B_IO_L2_in_5__ap_done;
  wire B_IO_L2_in_5__ap_idle;
  reg [1:0] B_IO_L2_in_5__state;
  wire B_IO_L2_in_6__ap_start_global__q0;
  wire B_IO_L2_in_6__is_done__q0;
  wire B_IO_L2_in_6__ap_done_global__q0;
  wire B_IO_L2_in_6__ap_start;
  wire B_IO_L2_in_6__ap_ready;
  wire B_IO_L2_in_6__ap_done;
  wire B_IO_L2_in_6__ap_idle;
  reg [1:0] B_IO_L2_in_6__state;
  wire B_IO_L2_in_7__ap_start_global__q0;
  wire B_IO_L2_in_7__is_done__q0;
  wire B_IO_L2_in_7__ap_done_global__q0;
  wire B_IO_L2_in_7__ap_start;
  wire B_IO_L2_in_7__ap_ready;
  wire B_IO_L2_in_7__ap_done;
  wire B_IO_L2_in_7__ap_idle;
  reg [1:0] B_IO_L2_in_7__state;
  wire B_IO_L2_in_8__ap_start_global__q0;
  wire B_IO_L2_in_8__is_done__q0;
  wire B_IO_L2_in_8__ap_done_global__q0;
  wire B_IO_L2_in_8__ap_start;
  wire B_IO_L2_in_8__ap_ready;
  wire B_IO_L2_in_8__ap_done;
  wire B_IO_L2_in_8__ap_idle;
  reg [1:0] B_IO_L2_in_8__state;
  wire B_IO_L2_in_9__ap_start_global__q0;
  wire B_IO_L2_in_9__is_done__q0;
  wire B_IO_L2_in_9__ap_done_global__q0;
  wire B_IO_L2_in_9__ap_start;
  wire B_IO_L2_in_9__ap_ready;
  wire B_IO_L2_in_9__ap_done;
  wire B_IO_L2_in_9__ap_idle;
  reg [1:0] B_IO_L2_in_9__state;
  wire B_IO_L2_in_10__ap_start_global__q0;
  wire B_IO_L2_in_10__is_done__q0;
  wire B_IO_L2_in_10__ap_done_global__q0;
  wire B_IO_L2_in_10__ap_start;
  wire B_IO_L2_in_10__ap_ready;
  wire B_IO_L2_in_10__ap_done;
  wire B_IO_L2_in_10__ap_idle;
  reg [1:0] B_IO_L2_in_10__state;
  wire B_IO_L2_in_11__ap_start_global__q0;
  wire B_IO_L2_in_11__is_done__q0;
  wire B_IO_L2_in_11__ap_done_global__q0;
  wire B_IO_L2_in_11__ap_start;
  wire B_IO_L2_in_11__ap_ready;
  wire B_IO_L2_in_11__ap_done;
  wire B_IO_L2_in_11__ap_idle;
  reg [1:0] B_IO_L2_in_11__state;
  wire B_IO_L2_in_12__ap_start_global__q0;
  wire B_IO_L2_in_12__is_done__q0;
  wire B_IO_L2_in_12__ap_done_global__q0;
  wire B_IO_L2_in_12__ap_start;
  wire B_IO_L2_in_12__ap_ready;
  wire B_IO_L2_in_12__ap_done;
  wire B_IO_L2_in_12__ap_idle;
  reg [1:0] B_IO_L2_in_12__state;
  wire B_IO_L2_in_13__ap_start_global__q0;
  wire B_IO_L2_in_13__is_done__q0;
  wire B_IO_L2_in_13__ap_done_global__q0;
  wire B_IO_L2_in_13__ap_start;
  wire B_IO_L2_in_13__ap_ready;
  wire B_IO_L2_in_13__ap_done;
  wire B_IO_L2_in_13__ap_idle;
  reg [1:0] B_IO_L2_in_13__state;
  wire B_IO_L2_in_14__ap_start_global__q0;
  wire B_IO_L2_in_14__is_done__q0;
  wire B_IO_L2_in_14__ap_done_global__q0;
  wire B_IO_L2_in_14__ap_start;
  wire B_IO_L2_in_14__ap_ready;
  wire B_IO_L2_in_14__ap_done;
  wire B_IO_L2_in_14__ap_idle;
  reg [1:0] B_IO_L2_in_14__state;
  wire B_IO_L2_in_15__ap_start_global__q0;
  wire B_IO_L2_in_15__is_done__q0;
  wire B_IO_L2_in_15__ap_done_global__q0;
  wire B_IO_L2_in_15__ap_start;
  wire B_IO_L2_in_15__ap_ready;
  wire B_IO_L2_in_15__ap_done;
  wire B_IO_L2_in_15__ap_idle;
  reg [1:0] B_IO_L2_in_15__state;
  wire B_IO_L2_in_boundary_0__ap_start_global__q0;
  wire B_IO_L2_in_boundary_0__is_done__q0;
  wire B_IO_L2_in_boundary_0__ap_done_global__q0;
  wire B_IO_L2_in_boundary_0__ap_start;
  wire B_IO_L2_in_boundary_0__ap_ready;
  wire B_IO_L2_in_boundary_0__ap_done;
  wire B_IO_L2_in_boundary_0__ap_idle;
  reg [1:0] B_IO_L2_in_boundary_0__state;
  wire B_IO_L3_in_0__ap_start_global__q0;
  wire B_IO_L3_in_0__is_done__q0;
  wire B_IO_L3_in_0__ap_done_global__q0;
  wire B_IO_L3_in_0__ap_start;
  wire B_IO_L3_in_0__ap_ready;
  wire B_IO_L3_in_0__ap_done;
  wire B_IO_L3_in_0__ap_idle;
  reg [1:0] B_IO_L3_in_0__state;
  wire [63:0] B_IO_L3_in_serialize_0___B__q0;
  wire B_IO_L3_in_serialize_0__ap_start_global__q0;
  wire B_IO_L3_in_serialize_0__is_done__q0;
  wire B_IO_L3_in_serialize_0__ap_done_global__q0;
  wire B_IO_L3_in_serialize_0__ap_start;
  wire B_IO_L3_in_serialize_0__ap_ready;
  wire B_IO_L3_in_serialize_0__ap_done;
  wire B_IO_L3_in_serialize_0__ap_idle;
  reg [1:0] B_IO_L3_in_serialize_0__state;
  wire B_PE_dummy_in_0__ap_start_global__q0;
  wire B_PE_dummy_in_0__is_done__q0;
  wire B_PE_dummy_in_0__ap_done_global__q0;
  wire B_PE_dummy_in_0__ap_start;
  wire B_PE_dummy_in_0__ap_ready;
  wire B_PE_dummy_in_0__ap_done;
  wire B_PE_dummy_in_0__ap_idle;
  reg [1:0] B_PE_dummy_in_0__state;
  wire B_PE_dummy_in_1__ap_start_global__q0;
  wire B_PE_dummy_in_1__is_done__q0;
  wire B_PE_dummy_in_1__ap_done_global__q0;
  wire B_PE_dummy_in_1__ap_start;
  wire B_PE_dummy_in_1__ap_ready;
  wire B_PE_dummy_in_1__ap_done;
  wire B_PE_dummy_in_1__ap_idle;
  reg [1:0] B_PE_dummy_in_1__state;
  wire B_PE_dummy_in_2__ap_start_global__q0;
  wire B_PE_dummy_in_2__is_done__q0;
  wire B_PE_dummy_in_2__ap_done_global__q0;
  wire B_PE_dummy_in_2__ap_start;
  wire B_PE_dummy_in_2__ap_ready;
  wire B_PE_dummy_in_2__ap_done;
  wire B_PE_dummy_in_2__ap_idle;
  reg [1:0] B_PE_dummy_in_2__state;
  wire B_PE_dummy_in_3__ap_start_global__q0;
  wire B_PE_dummy_in_3__is_done__q0;
  wire B_PE_dummy_in_3__ap_done_global__q0;
  wire B_PE_dummy_in_3__ap_start;
  wire B_PE_dummy_in_3__ap_ready;
  wire B_PE_dummy_in_3__ap_done;
  wire B_PE_dummy_in_3__ap_idle;
  reg [1:0] B_PE_dummy_in_3__state;
  wire B_PE_dummy_in_4__ap_start_global__q0;
  wire B_PE_dummy_in_4__is_done__q0;
  wire B_PE_dummy_in_4__ap_done_global__q0;
  wire B_PE_dummy_in_4__ap_start;
  wire B_PE_dummy_in_4__ap_ready;
  wire B_PE_dummy_in_4__ap_done;
  wire B_PE_dummy_in_4__ap_idle;
  reg [1:0] B_PE_dummy_in_4__state;
  wire B_PE_dummy_in_5__ap_start_global__q0;
  wire B_PE_dummy_in_5__is_done__q0;
  wire B_PE_dummy_in_5__ap_done_global__q0;
  wire B_PE_dummy_in_5__ap_start;
  wire B_PE_dummy_in_5__ap_ready;
  wire B_PE_dummy_in_5__ap_done;
  wire B_PE_dummy_in_5__ap_idle;
  reg [1:0] B_PE_dummy_in_5__state;
  wire B_PE_dummy_in_6__ap_start_global__q0;
  wire B_PE_dummy_in_6__is_done__q0;
  wire B_PE_dummy_in_6__ap_done_global__q0;
  wire B_PE_dummy_in_6__ap_start;
  wire B_PE_dummy_in_6__ap_ready;
  wire B_PE_dummy_in_6__ap_done;
  wire B_PE_dummy_in_6__ap_idle;
  reg [1:0] B_PE_dummy_in_6__state;
  wire B_PE_dummy_in_7__ap_start_global__q0;
  wire B_PE_dummy_in_7__is_done__q0;
  wire B_PE_dummy_in_7__ap_done_global__q0;
  wire B_PE_dummy_in_7__ap_start;
  wire B_PE_dummy_in_7__ap_ready;
  wire B_PE_dummy_in_7__ap_done;
  wire B_PE_dummy_in_7__ap_idle;
  reg [1:0] B_PE_dummy_in_7__state;
  wire B_PE_dummy_in_8__ap_start_global__q0;
  wire B_PE_dummy_in_8__is_done__q0;
  wire B_PE_dummy_in_8__ap_done_global__q0;
  wire B_PE_dummy_in_8__ap_start;
  wire B_PE_dummy_in_8__ap_ready;
  wire B_PE_dummy_in_8__ap_done;
  wire B_PE_dummy_in_8__ap_idle;
  reg [1:0] B_PE_dummy_in_8__state;
  wire B_PE_dummy_in_9__ap_start_global__q0;
  wire B_PE_dummy_in_9__is_done__q0;
  wire B_PE_dummy_in_9__ap_done_global__q0;
  wire B_PE_dummy_in_9__ap_start;
  wire B_PE_dummy_in_9__ap_ready;
  wire B_PE_dummy_in_9__ap_done;
  wire B_PE_dummy_in_9__ap_idle;
  reg [1:0] B_PE_dummy_in_9__state;
  wire B_PE_dummy_in_10__ap_start_global__q0;
  wire B_PE_dummy_in_10__is_done__q0;
  wire B_PE_dummy_in_10__ap_done_global__q0;
  wire B_PE_dummy_in_10__ap_start;
  wire B_PE_dummy_in_10__ap_ready;
  wire B_PE_dummy_in_10__ap_done;
  wire B_PE_dummy_in_10__ap_idle;
  reg [1:0] B_PE_dummy_in_10__state;
  wire B_PE_dummy_in_11__ap_start_global__q0;
  wire B_PE_dummy_in_11__is_done__q0;
  wire B_PE_dummy_in_11__ap_done_global__q0;
  wire B_PE_dummy_in_11__ap_start;
  wire B_PE_dummy_in_11__ap_ready;
  wire B_PE_dummy_in_11__ap_done;
  wire B_PE_dummy_in_11__ap_idle;
  reg [1:0] B_PE_dummy_in_11__state;
  wire B_PE_dummy_in_12__ap_start_global__q0;
  wire B_PE_dummy_in_12__is_done__q0;
  wire B_PE_dummy_in_12__ap_done_global__q0;
  wire B_PE_dummy_in_12__ap_start;
  wire B_PE_dummy_in_12__ap_ready;
  wire B_PE_dummy_in_12__ap_done;
  wire B_PE_dummy_in_12__ap_idle;
  reg [1:0] B_PE_dummy_in_12__state;
  wire B_PE_dummy_in_13__ap_start_global__q0;
  wire B_PE_dummy_in_13__is_done__q0;
  wire B_PE_dummy_in_13__ap_done_global__q0;
  wire B_PE_dummy_in_13__ap_start;
  wire B_PE_dummy_in_13__ap_ready;
  wire B_PE_dummy_in_13__ap_done;
  wire B_PE_dummy_in_13__ap_idle;
  reg [1:0] B_PE_dummy_in_13__state;
  wire B_PE_dummy_in_14__ap_start_global__q0;
  wire B_PE_dummy_in_14__is_done__q0;
  wire B_PE_dummy_in_14__ap_done_global__q0;
  wire B_PE_dummy_in_14__ap_start;
  wire B_PE_dummy_in_14__ap_ready;
  wire B_PE_dummy_in_14__ap_done;
  wire B_PE_dummy_in_14__ap_idle;
  reg [1:0] B_PE_dummy_in_14__state;
  wire B_PE_dummy_in_15__ap_start_global__q0;
  wire B_PE_dummy_in_15__is_done__q0;
  wire B_PE_dummy_in_15__ap_done_global__q0;
  wire B_PE_dummy_in_15__ap_start;
  wire B_PE_dummy_in_15__ap_ready;
  wire B_PE_dummy_in_15__ap_done;
  wire B_PE_dummy_in_15__ap_idle;
  reg [1:0] B_PE_dummy_in_15__state;
  wire B_PE_dummy_in_16__ap_start_global__q0;
  wire B_PE_dummy_in_16__is_done__q0;
  wire B_PE_dummy_in_16__ap_done_global__q0;
  wire B_PE_dummy_in_16__ap_start;
  wire B_PE_dummy_in_16__ap_ready;
  wire B_PE_dummy_in_16__ap_done;
  wire B_PE_dummy_in_16__ap_idle;
  reg [1:0] B_PE_dummy_in_16__state;
  wire C_drain_IO_L1_out_boundary_wrapper_0__ap_start_global__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_0__is_done__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_0__ap_done_global__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_0__ap_start;
  wire C_drain_IO_L1_out_boundary_wrapper_0__ap_ready;
  wire C_drain_IO_L1_out_boundary_wrapper_0__ap_done;
  wire C_drain_IO_L1_out_boundary_wrapper_0__ap_idle;
  reg [1:0] C_drain_IO_L1_out_boundary_wrapper_0__state;
  wire C_drain_IO_L1_out_boundary_wrapper_1__ap_start_global__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_1__is_done__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_1__ap_done_global__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_1__ap_start;
  wire C_drain_IO_L1_out_boundary_wrapper_1__ap_ready;
  wire C_drain_IO_L1_out_boundary_wrapper_1__ap_done;
  wire C_drain_IO_L1_out_boundary_wrapper_1__ap_idle;
  reg [1:0] C_drain_IO_L1_out_boundary_wrapper_1__state;
  wire C_drain_IO_L1_out_boundary_wrapper_2__ap_start_global__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_2__is_done__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_2__ap_done_global__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_2__ap_start;
  wire C_drain_IO_L1_out_boundary_wrapper_2__ap_ready;
  wire C_drain_IO_L1_out_boundary_wrapper_2__ap_done;
  wire C_drain_IO_L1_out_boundary_wrapper_2__ap_idle;
  reg [1:0] C_drain_IO_L1_out_boundary_wrapper_2__state;
  wire C_drain_IO_L1_out_boundary_wrapper_3__ap_start_global__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_3__is_done__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_3__ap_done_global__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_3__ap_start;
  wire C_drain_IO_L1_out_boundary_wrapper_3__ap_ready;
  wire C_drain_IO_L1_out_boundary_wrapper_3__ap_done;
  wire C_drain_IO_L1_out_boundary_wrapper_3__ap_idle;
  reg [1:0] C_drain_IO_L1_out_boundary_wrapper_3__state;
  wire C_drain_IO_L1_out_boundary_wrapper_4__ap_start_global__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_4__is_done__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_4__ap_done_global__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_4__ap_start;
  wire C_drain_IO_L1_out_boundary_wrapper_4__ap_ready;
  wire C_drain_IO_L1_out_boundary_wrapper_4__ap_done;
  wire C_drain_IO_L1_out_boundary_wrapper_4__ap_idle;
  reg [1:0] C_drain_IO_L1_out_boundary_wrapper_4__state;
  wire C_drain_IO_L1_out_boundary_wrapper_5__ap_start_global__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_5__is_done__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_5__ap_done_global__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_5__ap_start;
  wire C_drain_IO_L1_out_boundary_wrapper_5__ap_ready;
  wire C_drain_IO_L1_out_boundary_wrapper_5__ap_done;
  wire C_drain_IO_L1_out_boundary_wrapper_5__ap_idle;
  reg [1:0] C_drain_IO_L1_out_boundary_wrapper_5__state;
  wire C_drain_IO_L1_out_boundary_wrapper_6__ap_start_global__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_6__is_done__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_6__ap_done_global__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_6__ap_start;
  wire C_drain_IO_L1_out_boundary_wrapper_6__ap_ready;
  wire C_drain_IO_L1_out_boundary_wrapper_6__ap_done;
  wire C_drain_IO_L1_out_boundary_wrapper_6__ap_idle;
  reg [1:0] C_drain_IO_L1_out_boundary_wrapper_6__state;
  wire C_drain_IO_L1_out_boundary_wrapper_7__ap_start_global__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_7__is_done__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_7__ap_done_global__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_7__ap_start;
  wire C_drain_IO_L1_out_boundary_wrapper_7__ap_ready;
  wire C_drain_IO_L1_out_boundary_wrapper_7__ap_done;
  wire C_drain_IO_L1_out_boundary_wrapper_7__ap_idle;
  reg [1:0] C_drain_IO_L1_out_boundary_wrapper_7__state;
  wire C_drain_IO_L1_out_boundary_wrapper_8__ap_start_global__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_8__is_done__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_8__ap_done_global__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_8__ap_start;
  wire C_drain_IO_L1_out_boundary_wrapper_8__ap_ready;
  wire C_drain_IO_L1_out_boundary_wrapper_8__ap_done;
  wire C_drain_IO_L1_out_boundary_wrapper_8__ap_idle;
  reg [1:0] C_drain_IO_L1_out_boundary_wrapper_8__state;
  wire C_drain_IO_L1_out_boundary_wrapper_9__ap_start_global__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_9__is_done__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_9__ap_done_global__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_9__ap_start;
  wire C_drain_IO_L1_out_boundary_wrapper_9__ap_ready;
  wire C_drain_IO_L1_out_boundary_wrapper_9__ap_done;
  wire C_drain_IO_L1_out_boundary_wrapper_9__ap_idle;
  reg [1:0] C_drain_IO_L1_out_boundary_wrapper_9__state;
  wire C_drain_IO_L1_out_boundary_wrapper_10__ap_start_global__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_10__is_done__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_10__ap_done_global__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_10__ap_start;
  wire C_drain_IO_L1_out_boundary_wrapper_10__ap_ready;
  wire C_drain_IO_L1_out_boundary_wrapper_10__ap_done;
  wire C_drain_IO_L1_out_boundary_wrapper_10__ap_idle;
  reg [1:0] C_drain_IO_L1_out_boundary_wrapper_10__state;
  wire C_drain_IO_L1_out_boundary_wrapper_11__ap_start_global__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_11__is_done__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_11__ap_done_global__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_11__ap_start;
  wire C_drain_IO_L1_out_boundary_wrapper_11__ap_ready;
  wire C_drain_IO_L1_out_boundary_wrapper_11__ap_done;
  wire C_drain_IO_L1_out_boundary_wrapper_11__ap_idle;
  reg [1:0] C_drain_IO_L1_out_boundary_wrapper_11__state;
  wire C_drain_IO_L1_out_boundary_wrapper_12__ap_start_global__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_12__is_done__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_12__ap_done_global__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_12__ap_start;
  wire C_drain_IO_L1_out_boundary_wrapper_12__ap_ready;
  wire C_drain_IO_L1_out_boundary_wrapper_12__ap_done;
  wire C_drain_IO_L1_out_boundary_wrapper_12__ap_idle;
  reg [1:0] C_drain_IO_L1_out_boundary_wrapper_12__state;
  wire C_drain_IO_L1_out_boundary_wrapper_13__ap_start_global__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_13__is_done__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_13__ap_done_global__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_13__ap_start;
  wire C_drain_IO_L1_out_boundary_wrapper_13__ap_ready;
  wire C_drain_IO_L1_out_boundary_wrapper_13__ap_done;
  wire C_drain_IO_L1_out_boundary_wrapper_13__ap_idle;
  reg [1:0] C_drain_IO_L1_out_boundary_wrapper_13__state;
  wire C_drain_IO_L1_out_boundary_wrapper_14__ap_start_global__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_14__is_done__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_14__ap_done_global__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_14__ap_start;
  wire C_drain_IO_L1_out_boundary_wrapper_14__ap_ready;
  wire C_drain_IO_L1_out_boundary_wrapper_14__ap_done;
  wire C_drain_IO_L1_out_boundary_wrapper_14__ap_idle;
  reg [1:0] C_drain_IO_L1_out_boundary_wrapper_14__state;
  wire C_drain_IO_L1_out_boundary_wrapper_15__ap_start_global__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_15__is_done__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_15__ap_done_global__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_15__ap_start;
  wire C_drain_IO_L1_out_boundary_wrapper_15__ap_ready;
  wire C_drain_IO_L1_out_boundary_wrapper_15__ap_done;
  wire C_drain_IO_L1_out_boundary_wrapper_15__ap_idle;
  reg [1:0] C_drain_IO_L1_out_boundary_wrapper_15__state;
  wire C_drain_IO_L1_out_boundary_wrapper_16__ap_start_global__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_16__is_done__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_16__ap_done_global__q0;
  wire C_drain_IO_L1_out_boundary_wrapper_16__ap_start;
  wire C_drain_IO_L1_out_boundary_wrapper_16__ap_ready;
  wire C_drain_IO_L1_out_boundary_wrapper_16__ap_done;
  wire C_drain_IO_L1_out_boundary_wrapper_16__ap_idle;
  reg [1:0] C_drain_IO_L1_out_boundary_wrapper_16__state;
  wire C_drain_IO_L1_out_wrapper_0__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_0__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_0__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_0__ap_start;
  wire C_drain_IO_L1_out_wrapper_0__ap_ready;
  wire C_drain_IO_L1_out_wrapper_0__ap_done;
  wire C_drain_IO_L1_out_wrapper_0__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_0__state;
  wire C_drain_IO_L1_out_wrapper_1__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_1__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_1__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_1__ap_start;
  wire C_drain_IO_L1_out_wrapper_1__ap_ready;
  wire C_drain_IO_L1_out_wrapper_1__ap_done;
  wire C_drain_IO_L1_out_wrapper_1__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_1__state;
  wire C_drain_IO_L1_out_wrapper_2__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_2__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_2__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_2__ap_start;
  wire C_drain_IO_L1_out_wrapper_2__ap_ready;
  wire C_drain_IO_L1_out_wrapper_2__ap_done;
  wire C_drain_IO_L1_out_wrapper_2__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_2__state;
  wire C_drain_IO_L1_out_wrapper_3__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_3__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_3__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_3__ap_start;
  wire C_drain_IO_L1_out_wrapper_3__ap_ready;
  wire C_drain_IO_L1_out_wrapper_3__ap_done;
  wire C_drain_IO_L1_out_wrapper_3__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_3__state;
  wire C_drain_IO_L1_out_wrapper_4__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_4__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_4__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_4__ap_start;
  wire C_drain_IO_L1_out_wrapper_4__ap_ready;
  wire C_drain_IO_L1_out_wrapper_4__ap_done;
  wire C_drain_IO_L1_out_wrapper_4__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_4__state;
  wire C_drain_IO_L1_out_wrapper_5__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_5__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_5__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_5__ap_start;
  wire C_drain_IO_L1_out_wrapper_5__ap_ready;
  wire C_drain_IO_L1_out_wrapper_5__ap_done;
  wire C_drain_IO_L1_out_wrapper_5__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_5__state;
  wire C_drain_IO_L1_out_wrapper_6__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_6__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_6__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_6__ap_start;
  wire C_drain_IO_L1_out_wrapper_6__ap_ready;
  wire C_drain_IO_L1_out_wrapper_6__ap_done;
  wire C_drain_IO_L1_out_wrapper_6__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_6__state;
  wire C_drain_IO_L1_out_wrapper_7__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_7__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_7__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_7__ap_start;
  wire C_drain_IO_L1_out_wrapper_7__ap_ready;
  wire C_drain_IO_L1_out_wrapper_7__ap_done;
  wire C_drain_IO_L1_out_wrapper_7__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_7__state;
  wire C_drain_IO_L1_out_wrapper_8__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_8__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_8__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_8__ap_start;
  wire C_drain_IO_L1_out_wrapper_8__ap_ready;
  wire C_drain_IO_L1_out_wrapper_8__ap_done;
  wire C_drain_IO_L1_out_wrapper_8__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_8__state;
  wire C_drain_IO_L1_out_wrapper_9__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_9__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_9__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_9__ap_start;
  wire C_drain_IO_L1_out_wrapper_9__ap_ready;
  wire C_drain_IO_L1_out_wrapper_9__ap_done;
  wire C_drain_IO_L1_out_wrapper_9__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_9__state;
  wire C_drain_IO_L1_out_wrapper_10__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_10__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_10__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_10__ap_start;
  wire C_drain_IO_L1_out_wrapper_10__ap_ready;
  wire C_drain_IO_L1_out_wrapper_10__ap_done;
  wire C_drain_IO_L1_out_wrapper_10__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_10__state;
  wire C_drain_IO_L1_out_wrapper_11__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_11__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_11__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_11__ap_start;
  wire C_drain_IO_L1_out_wrapper_11__ap_ready;
  wire C_drain_IO_L1_out_wrapper_11__ap_done;
  wire C_drain_IO_L1_out_wrapper_11__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_11__state;
  wire C_drain_IO_L1_out_wrapper_12__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_12__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_12__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_12__ap_start;
  wire C_drain_IO_L1_out_wrapper_12__ap_ready;
  wire C_drain_IO_L1_out_wrapper_12__ap_done;
  wire C_drain_IO_L1_out_wrapper_12__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_12__state;
  wire C_drain_IO_L1_out_wrapper_13__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_13__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_13__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_13__ap_start;
  wire C_drain_IO_L1_out_wrapper_13__ap_ready;
  wire C_drain_IO_L1_out_wrapper_13__ap_done;
  wire C_drain_IO_L1_out_wrapper_13__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_13__state;
  wire C_drain_IO_L1_out_wrapper_14__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_14__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_14__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_14__ap_start;
  wire C_drain_IO_L1_out_wrapper_14__ap_ready;
  wire C_drain_IO_L1_out_wrapper_14__ap_done;
  wire C_drain_IO_L1_out_wrapper_14__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_14__state;
  wire C_drain_IO_L1_out_wrapper_15__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_15__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_15__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_15__ap_start;
  wire C_drain_IO_L1_out_wrapper_15__ap_ready;
  wire C_drain_IO_L1_out_wrapper_15__ap_done;
  wire C_drain_IO_L1_out_wrapper_15__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_15__state;
  wire C_drain_IO_L1_out_wrapper_16__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_16__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_16__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_16__ap_start;
  wire C_drain_IO_L1_out_wrapper_16__ap_ready;
  wire C_drain_IO_L1_out_wrapper_16__ap_done;
  wire C_drain_IO_L1_out_wrapper_16__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_16__state;
  wire C_drain_IO_L1_out_wrapper_17__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_17__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_17__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_17__ap_start;
  wire C_drain_IO_L1_out_wrapper_17__ap_ready;
  wire C_drain_IO_L1_out_wrapper_17__ap_done;
  wire C_drain_IO_L1_out_wrapper_17__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_17__state;
  wire C_drain_IO_L1_out_wrapper_18__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_18__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_18__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_18__ap_start;
  wire C_drain_IO_L1_out_wrapper_18__ap_ready;
  wire C_drain_IO_L1_out_wrapper_18__ap_done;
  wire C_drain_IO_L1_out_wrapper_18__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_18__state;
  wire C_drain_IO_L1_out_wrapper_19__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_19__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_19__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_19__ap_start;
  wire C_drain_IO_L1_out_wrapper_19__ap_ready;
  wire C_drain_IO_L1_out_wrapper_19__ap_done;
  wire C_drain_IO_L1_out_wrapper_19__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_19__state;
  wire C_drain_IO_L1_out_wrapper_20__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_20__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_20__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_20__ap_start;
  wire C_drain_IO_L1_out_wrapper_20__ap_ready;
  wire C_drain_IO_L1_out_wrapper_20__ap_done;
  wire C_drain_IO_L1_out_wrapper_20__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_20__state;
  wire C_drain_IO_L1_out_wrapper_21__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_21__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_21__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_21__ap_start;
  wire C_drain_IO_L1_out_wrapper_21__ap_ready;
  wire C_drain_IO_L1_out_wrapper_21__ap_done;
  wire C_drain_IO_L1_out_wrapper_21__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_21__state;
  wire C_drain_IO_L1_out_wrapper_22__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_22__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_22__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_22__ap_start;
  wire C_drain_IO_L1_out_wrapper_22__ap_ready;
  wire C_drain_IO_L1_out_wrapper_22__ap_done;
  wire C_drain_IO_L1_out_wrapper_22__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_22__state;
  wire C_drain_IO_L1_out_wrapper_23__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_23__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_23__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_23__ap_start;
  wire C_drain_IO_L1_out_wrapper_23__ap_ready;
  wire C_drain_IO_L1_out_wrapper_23__ap_done;
  wire C_drain_IO_L1_out_wrapper_23__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_23__state;
  wire C_drain_IO_L1_out_wrapper_24__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_24__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_24__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_24__ap_start;
  wire C_drain_IO_L1_out_wrapper_24__ap_ready;
  wire C_drain_IO_L1_out_wrapper_24__ap_done;
  wire C_drain_IO_L1_out_wrapper_24__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_24__state;
  wire C_drain_IO_L1_out_wrapper_25__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_25__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_25__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_25__ap_start;
  wire C_drain_IO_L1_out_wrapper_25__ap_ready;
  wire C_drain_IO_L1_out_wrapper_25__ap_done;
  wire C_drain_IO_L1_out_wrapper_25__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_25__state;
  wire C_drain_IO_L1_out_wrapper_26__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_26__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_26__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_26__ap_start;
  wire C_drain_IO_L1_out_wrapper_26__ap_ready;
  wire C_drain_IO_L1_out_wrapper_26__ap_done;
  wire C_drain_IO_L1_out_wrapper_26__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_26__state;
  wire C_drain_IO_L1_out_wrapper_27__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_27__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_27__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_27__ap_start;
  wire C_drain_IO_L1_out_wrapper_27__ap_ready;
  wire C_drain_IO_L1_out_wrapper_27__ap_done;
  wire C_drain_IO_L1_out_wrapper_27__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_27__state;
  wire C_drain_IO_L1_out_wrapper_28__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_28__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_28__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_28__ap_start;
  wire C_drain_IO_L1_out_wrapper_28__ap_ready;
  wire C_drain_IO_L1_out_wrapper_28__ap_done;
  wire C_drain_IO_L1_out_wrapper_28__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_28__state;
  wire C_drain_IO_L1_out_wrapper_29__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_29__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_29__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_29__ap_start;
  wire C_drain_IO_L1_out_wrapper_29__ap_ready;
  wire C_drain_IO_L1_out_wrapper_29__ap_done;
  wire C_drain_IO_L1_out_wrapper_29__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_29__state;
  wire C_drain_IO_L1_out_wrapper_30__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_30__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_30__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_30__ap_start;
  wire C_drain_IO_L1_out_wrapper_30__ap_ready;
  wire C_drain_IO_L1_out_wrapper_30__ap_done;
  wire C_drain_IO_L1_out_wrapper_30__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_30__state;
  wire C_drain_IO_L1_out_wrapper_31__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_31__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_31__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_31__ap_start;
  wire C_drain_IO_L1_out_wrapper_31__ap_ready;
  wire C_drain_IO_L1_out_wrapper_31__ap_done;
  wire C_drain_IO_L1_out_wrapper_31__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_31__state;
  wire C_drain_IO_L1_out_wrapper_32__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_32__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_32__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_32__ap_start;
  wire C_drain_IO_L1_out_wrapper_32__ap_ready;
  wire C_drain_IO_L1_out_wrapper_32__ap_done;
  wire C_drain_IO_L1_out_wrapper_32__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_32__state;
  wire C_drain_IO_L1_out_wrapper_33__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_33__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_33__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_33__ap_start;
  wire C_drain_IO_L1_out_wrapper_33__ap_ready;
  wire C_drain_IO_L1_out_wrapper_33__ap_done;
  wire C_drain_IO_L1_out_wrapper_33__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_33__state;
  wire C_drain_IO_L1_out_wrapper_34__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_34__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_34__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_34__ap_start;
  wire C_drain_IO_L1_out_wrapper_34__ap_ready;
  wire C_drain_IO_L1_out_wrapper_34__ap_done;
  wire C_drain_IO_L1_out_wrapper_34__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_34__state;
  wire C_drain_IO_L1_out_wrapper_35__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_35__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_35__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_35__ap_start;
  wire C_drain_IO_L1_out_wrapper_35__ap_ready;
  wire C_drain_IO_L1_out_wrapper_35__ap_done;
  wire C_drain_IO_L1_out_wrapper_35__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_35__state;
  wire C_drain_IO_L1_out_wrapper_36__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_36__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_36__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_36__ap_start;
  wire C_drain_IO_L1_out_wrapper_36__ap_ready;
  wire C_drain_IO_L1_out_wrapper_36__ap_done;
  wire C_drain_IO_L1_out_wrapper_36__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_36__state;
  wire C_drain_IO_L1_out_wrapper_37__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_37__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_37__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_37__ap_start;
  wire C_drain_IO_L1_out_wrapper_37__ap_ready;
  wire C_drain_IO_L1_out_wrapper_37__ap_done;
  wire C_drain_IO_L1_out_wrapper_37__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_37__state;
  wire C_drain_IO_L1_out_wrapper_38__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_38__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_38__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_38__ap_start;
  wire C_drain_IO_L1_out_wrapper_38__ap_ready;
  wire C_drain_IO_L1_out_wrapper_38__ap_done;
  wire C_drain_IO_L1_out_wrapper_38__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_38__state;
  wire C_drain_IO_L1_out_wrapper_39__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_39__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_39__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_39__ap_start;
  wire C_drain_IO_L1_out_wrapper_39__ap_ready;
  wire C_drain_IO_L1_out_wrapper_39__ap_done;
  wire C_drain_IO_L1_out_wrapper_39__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_39__state;
  wire C_drain_IO_L1_out_wrapper_40__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_40__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_40__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_40__ap_start;
  wire C_drain_IO_L1_out_wrapper_40__ap_ready;
  wire C_drain_IO_L1_out_wrapper_40__ap_done;
  wire C_drain_IO_L1_out_wrapper_40__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_40__state;
  wire C_drain_IO_L1_out_wrapper_41__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_41__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_41__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_41__ap_start;
  wire C_drain_IO_L1_out_wrapper_41__ap_ready;
  wire C_drain_IO_L1_out_wrapper_41__ap_done;
  wire C_drain_IO_L1_out_wrapper_41__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_41__state;
  wire C_drain_IO_L1_out_wrapper_42__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_42__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_42__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_42__ap_start;
  wire C_drain_IO_L1_out_wrapper_42__ap_ready;
  wire C_drain_IO_L1_out_wrapper_42__ap_done;
  wire C_drain_IO_L1_out_wrapper_42__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_42__state;
  wire C_drain_IO_L1_out_wrapper_43__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_43__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_43__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_43__ap_start;
  wire C_drain_IO_L1_out_wrapper_43__ap_ready;
  wire C_drain_IO_L1_out_wrapper_43__ap_done;
  wire C_drain_IO_L1_out_wrapper_43__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_43__state;
  wire C_drain_IO_L1_out_wrapper_44__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_44__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_44__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_44__ap_start;
  wire C_drain_IO_L1_out_wrapper_44__ap_ready;
  wire C_drain_IO_L1_out_wrapper_44__ap_done;
  wire C_drain_IO_L1_out_wrapper_44__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_44__state;
  wire C_drain_IO_L1_out_wrapper_45__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_45__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_45__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_45__ap_start;
  wire C_drain_IO_L1_out_wrapper_45__ap_ready;
  wire C_drain_IO_L1_out_wrapper_45__ap_done;
  wire C_drain_IO_L1_out_wrapper_45__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_45__state;
  wire C_drain_IO_L1_out_wrapper_46__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_46__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_46__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_46__ap_start;
  wire C_drain_IO_L1_out_wrapper_46__ap_ready;
  wire C_drain_IO_L1_out_wrapper_46__ap_done;
  wire C_drain_IO_L1_out_wrapper_46__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_46__state;
  wire C_drain_IO_L1_out_wrapper_47__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_47__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_47__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_47__ap_start;
  wire C_drain_IO_L1_out_wrapper_47__ap_ready;
  wire C_drain_IO_L1_out_wrapper_47__ap_done;
  wire C_drain_IO_L1_out_wrapper_47__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_47__state;
  wire C_drain_IO_L1_out_wrapper_48__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_48__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_48__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_48__ap_start;
  wire C_drain_IO_L1_out_wrapper_48__ap_ready;
  wire C_drain_IO_L1_out_wrapper_48__ap_done;
  wire C_drain_IO_L1_out_wrapper_48__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_48__state;
  wire C_drain_IO_L1_out_wrapper_49__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_49__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_49__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_49__ap_start;
  wire C_drain_IO_L1_out_wrapper_49__ap_ready;
  wire C_drain_IO_L1_out_wrapper_49__ap_done;
  wire C_drain_IO_L1_out_wrapper_49__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_49__state;
  wire C_drain_IO_L1_out_wrapper_50__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_50__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_50__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_50__ap_start;
  wire C_drain_IO_L1_out_wrapper_50__ap_ready;
  wire C_drain_IO_L1_out_wrapper_50__ap_done;
  wire C_drain_IO_L1_out_wrapper_50__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_50__state;
  wire C_drain_IO_L1_out_wrapper_51__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_51__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_51__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_51__ap_start;
  wire C_drain_IO_L1_out_wrapper_51__ap_ready;
  wire C_drain_IO_L1_out_wrapper_51__ap_done;
  wire C_drain_IO_L1_out_wrapper_51__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_51__state;
  wire C_drain_IO_L1_out_wrapper_52__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_52__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_52__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_52__ap_start;
  wire C_drain_IO_L1_out_wrapper_52__ap_ready;
  wire C_drain_IO_L1_out_wrapper_52__ap_done;
  wire C_drain_IO_L1_out_wrapper_52__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_52__state;
  wire C_drain_IO_L1_out_wrapper_53__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_53__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_53__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_53__ap_start;
  wire C_drain_IO_L1_out_wrapper_53__ap_ready;
  wire C_drain_IO_L1_out_wrapper_53__ap_done;
  wire C_drain_IO_L1_out_wrapper_53__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_53__state;
  wire C_drain_IO_L1_out_wrapper_54__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_54__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_54__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_54__ap_start;
  wire C_drain_IO_L1_out_wrapper_54__ap_ready;
  wire C_drain_IO_L1_out_wrapper_54__ap_done;
  wire C_drain_IO_L1_out_wrapper_54__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_54__state;
  wire C_drain_IO_L1_out_wrapper_55__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_55__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_55__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_55__ap_start;
  wire C_drain_IO_L1_out_wrapper_55__ap_ready;
  wire C_drain_IO_L1_out_wrapper_55__ap_done;
  wire C_drain_IO_L1_out_wrapper_55__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_55__state;
  wire C_drain_IO_L1_out_wrapper_56__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_56__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_56__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_56__ap_start;
  wire C_drain_IO_L1_out_wrapper_56__ap_ready;
  wire C_drain_IO_L1_out_wrapper_56__ap_done;
  wire C_drain_IO_L1_out_wrapper_56__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_56__state;
  wire C_drain_IO_L1_out_wrapper_57__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_57__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_57__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_57__ap_start;
  wire C_drain_IO_L1_out_wrapper_57__ap_ready;
  wire C_drain_IO_L1_out_wrapper_57__ap_done;
  wire C_drain_IO_L1_out_wrapper_57__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_57__state;
  wire C_drain_IO_L1_out_wrapper_58__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_58__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_58__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_58__ap_start;
  wire C_drain_IO_L1_out_wrapper_58__ap_ready;
  wire C_drain_IO_L1_out_wrapper_58__ap_done;
  wire C_drain_IO_L1_out_wrapper_58__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_58__state;
  wire C_drain_IO_L1_out_wrapper_59__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_59__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_59__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_59__ap_start;
  wire C_drain_IO_L1_out_wrapper_59__ap_ready;
  wire C_drain_IO_L1_out_wrapper_59__ap_done;
  wire C_drain_IO_L1_out_wrapper_59__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_59__state;
  wire C_drain_IO_L1_out_wrapper_60__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_60__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_60__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_60__ap_start;
  wire C_drain_IO_L1_out_wrapper_60__ap_ready;
  wire C_drain_IO_L1_out_wrapper_60__ap_done;
  wire C_drain_IO_L1_out_wrapper_60__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_60__state;
  wire C_drain_IO_L1_out_wrapper_61__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_61__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_61__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_61__ap_start;
  wire C_drain_IO_L1_out_wrapper_61__ap_ready;
  wire C_drain_IO_L1_out_wrapper_61__ap_done;
  wire C_drain_IO_L1_out_wrapper_61__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_61__state;
  wire C_drain_IO_L1_out_wrapper_62__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_62__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_62__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_62__ap_start;
  wire C_drain_IO_L1_out_wrapper_62__ap_ready;
  wire C_drain_IO_L1_out_wrapper_62__ap_done;
  wire C_drain_IO_L1_out_wrapper_62__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_62__state;
  wire C_drain_IO_L1_out_wrapper_63__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_63__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_63__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_63__ap_start;
  wire C_drain_IO_L1_out_wrapper_63__ap_ready;
  wire C_drain_IO_L1_out_wrapper_63__ap_done;
  wire C_drain_IO_L1_out_wrapper_63__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_63__state;
  wire C_drain_IO_L1_out_wrapper_64__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_64__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_64__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_64__ap_start;
  wire C_drain_IO_L1_out_wrapper_64__ap_ready;
  wire C_drain_IO_L1_out_wrapper_64__ap_done;
  wire C_drain_IO_L1_out_wrapper_64__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_64__state;
  wire C_drain_IO_L1_out_wrapper_65__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_65__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_65__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_65__ap_start;
  wire C_drain_IO_L1_out_wrapper_65__ap_ready;
  wire C_drain_IO_L1_out_wrapper_65__ap_done;
  wire C_drain_IO_L1_out_wrapper_65__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_65__state;
  wire C_drain_IO_L1_out_wrapper_66__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_66__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_66__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_66__ap_start;
  wire C_drain_IO_L1_out_wrapper_66__ap_ready;
  wire C_drain_IO_L1_out_wrapper_66__ap_done;
  wire C_drain_IO_L1_out_wrapper_66__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_66__state;
  wire C_drain_IO_L1_out_wrapper_67__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_67__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_67__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_67__ap_start;
  wire C_drain_IO_L1_out_wrapper_67__ap_ready;
  wire C_drain_IO_L1_out_wrapper_67__ap_done;
  wire C_drain_IO_L1_out_wrapper_67__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_67__state;
  wire C_drain_IO_L1_out_wrapper_68__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_68__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_68__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_68__ap_start;
  wire C_drain_IO_L1_out_wrapper_68__ap_ready;
  wire C_drain_IO_L1_out_wrapper_68__ap_done;
  wire C_drain_IO_L1_out_wrapper_68__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_68__state;
  wire C_drain_IO_L1_out_wrapper_69__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_69__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_69__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_69__ap_start;
  wire C_drain_IO_L1_out_wrapper_69__ap_ready;
  wire C_drain_IO_L1_out_wrapper_69__ap_done;
  wire C_drain_IO_L1_out_wrapper_69__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_69__state;
  wire C_drain_IO_L1_out_wrapper_70__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_70__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_70__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_70__ap_start;
  wire C_drain_IO_L1_out_wrapper_70__ap_ready;
  wire C_drain_IO_L1_out_wrapper_70__ap_done;
  wire C_drain_IO_L1_out_wrapper_70__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_70__state;
  wire C_drain_IO_L1_out_wrapper_71__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_71__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_71__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_71__ap_start;
  wire C_drain_IO_L1_out_wrapper_71__ap_ready;
  wire C_drain_IO_L1_out_wrapper_71__ap_done;
  wire C_drain_IO_L1_out_wrapper_71__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_71__state;
  wire C_drain_IO_L1_out_wrapper_72__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_72__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_72__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_72__ap_start;
  wire C_drain_IO_L1_out_wrapper_72__ap_ready;
  wire C_drain_IO_L1_out_wrapper_72__ap_done;
  wire C_drain_IO_L1_out_wrapper_72__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_72__state;
  wire C_drain_IO_L1_out_wrapper_73__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_73__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_73__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_73__ap_start;
  wire C_drain_IO_L1_out_wrapper_73__ap_ready;
  wire C_drain_IO_L1_out_wrapper_73__ap_done;
  wire C_drain_IO_L1_out_wrapper_73__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_73__state;
  wire C_drain_IO_L1_out_wrapper_74__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_74__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_74__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_74__ap_start;
  wire C_drain_IO_L1_out_wrapper_74__ap_ready;
  wire C_drain_IO_L1_out_wrapper_74__ap_done;
  wire C_drain_IO_L1_out_wrapper_74__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_74__state;
  wire C_drain_IO_L1_out_wrapper_75__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_75__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_75__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_75__ap_start;
  wire C_drain_IO_L1_out_wrapper_75__ap_ready;
  wire C_drain_IO_L1_out_wrapper_75__ap_done;
  wire C_drain_IO_L1_out_wrapper_75__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_75__state;
  wire C_drain_IO_L1_out_wrapper_76__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_76__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_76__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_76__ap_start;
  wire C_drain_IO_L1_out_wrapper_76__ap_ready;
  wire C_drain_IO_L1_out_wrapper_76__ap_done;
  wire C_drain_IO_L1_out_wrapper_76__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_76__state;
  wire C_drain_IO_L1_out_wrapper_77__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_77__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_77__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_77__ap_start;
  wire C_drain_IO_L1_out_wrapper_77__ap_ready;
  wire C_drain_IO_L1_out_wrapper_77__ap_done;
  wire C_drain_IO_L1_out_wrapper_77__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_77__state;
  wire C_drain_IO_L1_out_wrapper_78__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_78__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_78__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_78__ap_start;
  wire C_drain_IO_L1_out_wrapper_78__ap_ready;
  wire C_drain_IO_L1_out_wrapper_78__ap_done;
  wire C_drain_IO_L1_out_wrapper_78__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_78__state;
  wire C_drain_IO_L1_out_wrapper_79__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_79__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_79__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_79__ap_start;
  wire C_drain_IO_L1_out_wrapper_79__ap_ready;
  wire C_drain_IO_L1_out_wrapper_79__ap_done;
  wire C_drain_IO_L1_out_wrapper_79__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_79__state;
  wire C_drain_IO_L1_out_wrapper_80__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_80__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_80__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_80__ap_start;
  wire C_drain_IO_L1_out_wrapper_80__ap_ready;
  wire C_drain_IO_L1_out_wrapper_80__ap_done;
  wire C_drain_IO_L1_out_wrapper_80__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_80__state;
  wire C_drain_IO_L1_out_wrapper_81__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_81__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_81__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_81__ap_start;
  wire C_drain_IO_L1_out_wrapper_81__ap_ready;
  wire C_drain_IO_L1_out_wrapper_81__ap_done;
  wire C_drain_IO_L1_out_wrapper_81__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_81__state;
  wire C_drain_IO_L1_out_wrapper_82__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_82__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_82__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_82__ap_start;
  wire C_drain_IO_L1_out_wrapper_82__ap_ready;
  wire C_drain_IO_L1_out_wrapper_82__ap_done;
  wire C_drain_IO_L1_out_wrapper_82__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_82__state;
  wire C_drain_IO_L1_out_wrapper_83__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_83__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_83__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_83__ap_start;
  wire C_drain_IO_L1_out_wrapper_83__ap_ready;
  wire C_drain_IO_L1_out_wrapper_83__ap_done;
  wire C_drain_IO_L1_out_wrapper_83__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_83__state;
  wire C_drain_IO_L1_out_wrapper_84__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_84__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_84__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_84__ap_start;
  wire C_drain_IO_L1_out_wrapper_84__ap_ready;
  wire C_drain_IO_L1_out_wrapper_84__ap_done;
  wire C_drain_IO_L1_out_wrapper_84__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_84__state;
  wire C_drain_IO_L1_out_wrapper_85__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_85__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_85__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_85__ap_start;
  wire C_drain_IO_L1_out_wrapper_85__ap_ready;
  wire C_drain_IO_L1_out_wrapper_85__ap_done;
  wire C_drain_IO_L1_out_wrapper_85__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_85__state;
  wire C_drain_IO_L1_out_wrapper_86__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_86__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_86__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_86__ap_start;
  wire C_drain_IO_L1_out_wrapper_86__ap_ready;
  wire C_drain_IO_L1_out_wrapper_86__ap_done;
  wire C_drain_IO_L1_out_wrapper_86__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_86__state;
  wire C_drain_IO_L1_out_wrapper_87__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_87__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_87__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_87__ap_start;
  wire C_drain_IO_L1_out_wrapper_87__ap_ready;
  wire C_drain_IO_L1_out_wrapper_87__ap_done;
  wire C_drain_IO_L1_out_wrapper_87__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_87__state;
  wire C_drain_IO_L1_out_wrapper_88__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_88__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_88__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_88__ap_start;
  wire C_drain_IO_L1_out_wrapper_88__ap_ready;
  wire C_drain_IO_L1_out_wrapper_88__ap_done;
  wire C_drain_IO_L1_out_wrapper_88__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_88__state;
  wire C_drain_IO_L1_out_wrapper_89__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_89__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_89__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_89__ap_start;
  wire C_drain_IO_L1_out_wrapper_89__ap_ready;
  wire C_drain_IO_L1_out_wrapper_89__ap_done;
  wire C_drain_IO_L1_out_wrapper_89__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_89__state;
  wire C_drain_IO_L1_out_wrapper_90__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_90__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_90__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_90__ap_start;
  wire C_drain_IO_L1_out_wrapper_90__ap_ready;
  wire C_drain_IO_L1_out_wrapper_90__ap_done;
  wire C_drain_IO_L1_out_wrapper_90__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_90__state;
  wire C_drain_IO_L1_out_wrapper_91__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_91__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_91__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_91__ap_start;
  wire C_drain_IO_L1_out_wrapper_91__ap_ready;
  wire C_drain_IO_L1_out_wrapper_91__ap_done;
  wire C_drain_IO_L1_out_wrapper_91__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_91__state;
  wire C_drain_IO_L1_out_wrapper_92__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_92__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_92__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_92__ap_start;
  wire C_drain_IO_L1_out_wrapper_92__ap_ready;
  wire C_drain_IO_L1_out_wrapper_92__ap_done;
  wire C_drain_IO_L1_out_wrapper_92__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_92__state;
  wire C_drain_IO_L1_out_wrapper_93__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_93__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_93__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_93__ap_start;
  wire C_drain_IO_L1_out_wrapper_93__ap_ready;
  wire C_drain_IO_L1_out_wrapper_93__ap_done;
  wire C_drain_IO_L1_out_wrapper_93__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_93__state;
  wire C_drain_IO_L1_out_wrapper_94__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_94__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_94__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_94__ap_start;
  wire C_drain_IO_L1_out_wrapper_94__ap_ready;
  wire C_drain_IO_L1_out_wrapper_94__ap_done;
  wire C_drain_IO_L1_out_wrapper_94__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_94__state;
  wire C_drain_IO_L1_out_wrapper_95__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_95__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_95__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_95__ap_start;
  wire C_drain_IO_L1_out_wrapper_95__ap_ready;
  wire C_drain_IO_L1_out_wrapper_95__ap_done;
  wire C_drain_IO_L1_out_wrapper_95__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_95__state;
  wire C_drain_IO_L1_out_wrapper_96__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_96__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_96__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_96__ap_start;
  wire C_drain_IO_L1_out_wrapper_96__ap_ready;
  wire C_drain_IO_L1_out_wrapper_96__ap_done;
  wire C_drain_IO_L1_out_wrapper_96__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_96__state;
  wire C_drain_IO_L1_out_wrapper_97__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_97__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_97__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_97__ap_start;
  wire C_drain_IO_L1_out_wrapper_97__ap_ready;
  wire C_drain_IO_L1_out_wrapper_97__ap_done;
  wire C_drain_IO_L1_out_wrapper_97__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_97__state;
  wire C_drain_IO_L1_out_wrapper_98__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_98__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_98__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_98__ap_start;
  wire C_drain_IO_L1_out_wrapper_98__ap_ready;
  wire C_drain_IO_L1_out_wrapper_98__ap_done;
  wire C_drain_IO_L1_out_wrapper_98__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_98__state;
  wire C_drain_IO_L1_out_wrapper_99__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_99__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_99__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_99__ap_start;
  wire C_drain_IO_L1_out_wrapper_99__ap_ready;
  wire C_drain_IO_L1_out_wrapper_99__ap_done;
  wire C_drain_IO_L1_out_wrapper_99__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_99__state;
  wire C_drain_IO_L1_out_wrapper_100__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_100__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_100__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_100__ap_start;
  wire C_drain_IO_L1_out_wrapper_100__ap_ready;
  wire C_drain_IO_L1_out_wrapper_100__ap_done;
  wire C_drain_IO_L1_out_wrapper_100__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_100__state;
  wire C_drain_IO_L1_out_wrapper_101__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_101__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_101__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_101__ap_start;
  wire C_drain_IO_L1_out_wrapper_101__ap_ready;
  wire C_drain_IO_L1_out_wrapper_101__ap_done;
  wire C_drain_IO_L1_out_wrapper_101__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_101__state;
  wire C_drain_IO_L1_out_wrapper_102__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_102__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_102__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_102__ap_start;
  wire C_drain_IO_L1_out_wrapper_102__ap_ready;
  wire C_drain_IO_L1_out_wrapper_102__ap_done;
  wire C_drain_IO_L1_out_wrapper_102__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_102__state;
  wire C_drain_IO_L1_out_wrapper_103__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_103__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_103__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_103__ap_start;
  wire C_drain_IO_L1_out_wrapper_103__ap_ready;
  wire C_drain_IO_L1_out_wrapper_103__ap_done;
  wire C_drain_IO_L1_out_wrapper_103__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_103__state;
  wire C_drain_IO_L1_out_wrapper_104__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_104__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_104__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_104__ap_start;
  wire C_drain_IO_L1_out_wrapper_104__ap_ready;
  wire C_drain_IO_L1_out_wrapper_104__ap_done;
  wire C_drain_IO_L1_out_wrapper_104__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_104__state;
  wire C_drain_IO_L1_out_wrapper_105__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_105__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_105__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_105__ap_start;
  wire C_drain_IO_L1_out_wrapper_105__ap_ready;
  wire C_drain_IO_L1_out_wrapper_105__ap_done;
  wire C_drain_IO_L1_out_wrapper_105__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_105__state;
  wire C_drain_IO_L1_out_wrapper_106__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_106__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_106__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_106__ap_start;
  wire C_drain_IO_L1_out_wrapper_106__ap_ready;
  wire C_drain_IO_L1_out_wrapper_106__ap_done;
  wire C_drain_IO_L1_out_wrapper_106__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_106__state;
  wire C_drain_IO_L1_out_wrapper_107__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_107__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_107__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_107__ap_start;
  wire C_drain_IO_L1_out_wrapper_107__ap_ready;
  wire C_drain_IO_L1_out_wrapper_107__ap_done;
  wire C_drain_IO_L1_out_wrapper_107__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_107__state;
  wire C_drain_IO_L1_out_wrapper_108__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_108__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_108__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_108__ap_start;
  wire C_drain_IO_L1_out_wrapper_108__ap_ready;
  wire C_drain_IO_L1_out_wrapper_108__ap_done;
  wire C_drain_IO_L1_out_wrapper_108__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_108__state;
  wire C_drain_IO_L1_out_wrapper_109__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_109__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_109__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_109__ap_start;
  wire C_drain_IO_L1_out_wrapper_109__ap_ready;
  wire C_drain_IO_L1_out_wrapper_109__ap_done;
  wire C_drain_IO_L1_out_wrapper_109__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_109__state;
  wire C_drain_IO_L1_out_wrapper_110__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_110__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_110__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_110__ap_start;
  wire C_drain_IO_L1_out_wrapper_110__ap_ready;
  wire C_drain_IO_L1_out_wrapper_110__ap_done;
  wire C_drain_IO_L1_out_wrapper_110__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_110__state;
  wire C_drain_IO_L1_out_wrapper_111__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_111__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_111__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_111__ap_start;
  wire C_drain_IO_L1_out_wrapper_111__ap_ready;
  wire C_drain_IO_L1_out_wrapper_111__ap_done;
  wire C_drain_IO_L1_out_wrapper_111__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_111__state;
  wire C_drain_IO_L1_out_wrapper_112__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_112__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_112__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_112__ap_start;
  wire C_drain_IO_L1_out_wrapper_112__ap_ready;
  wire C_drain_IO_L1_out_wrapper_112__ap_done;
  wire C_drain_IO_L1_out_wrapper_112__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_112__state;
  wire C_drain_IO_L1_out_wrapper_113__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_113__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_113__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_113__ap_start;
  wire C_drain_IO_L1_out_wrapper_113__ap_ready;
  wire C_drain_IO_L1_out_wrapper_113__ap_done;
  wire C_drain_IO_L1_out_wrapper_113__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_113__state;
  wire C_drain_IO_L1_out_wrapper_114__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_114__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_114__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_114__ap_start;
  wire C_drain_IO_L1_out_wrapper_114__ap_ready;
  wire C_drain_IO_L1_out_wrapper_114__ap_done;
  wire C_drain_IO_L1_out_wrapper_114__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_114__state;
  wire C_drain_IO_L1_out_wrapper_115__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_115__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_115__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_115__ap_start;
  wire C_drain_IO_L1_out_wrapper_115__ap_ready;
  wire C_drain_IO_L1_out_wrapper_115__ap_done;
  wire C_drain_IO_L1_out_wrapper_115__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_115__state;
  wire C_drain_IO_L1_out_wrapper_116__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_116__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_116__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_116__ap_start;
  wire C_drain_IO_L1_out_wrapper_116__ap_ready;
  wire C_drain_IO_L1_out_wrapper_116__ap_done;
  wire C_drain_IO_L1_out_wrapper_116__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_116__state;
  wire C_drain_IO_L1_out_wrapper_117__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_117__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_117__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_117__ap_start;
  wire C_drain_IO_L1_out_wrapper_117__ap_ready;
  wire C_drain_IO_L1_out_wrapper_117__ap_done;
  wire C_drain_IO_L1_out_wrapper_117__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_117__state;
  wire C_drain_IO_L1_out_wrapper_118__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_118__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_118__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_118__ap_start;
  wire C_drain_IO_L1_out_wrapper_118__ap_ready;
  wire C_drain_IO_L1_out_wrapper_118__ap_done;
  wire C_drain_IO_L1_out_wrapper_118__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_118__state;
  wire C_drain_IO_L1_out_wrapper_119__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_119__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_119__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_119__ap_start;
  wire C_drain_IO_L1_out_wrapper_119__ap_ready;
  wire C_drain_IO_L1_out_wrapper_119__ap_done;
  wire C_drain_IO_L1_out_wrapper_119__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_119__state;
  wire C_drain_IO_L1_out_wrapper_120__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_120__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_120__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_120__ap_start;
  wire C_drain_IO_L1_out_wrapper_120__ap_ready;
  wire C_drain_IO_L1_out_wrapper_120__ap_done;
  wire C_drain_IO_L1_out_wrapper_120__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_120__state;
  wire C_drain_IO_L1_out_wrapper_121__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_121__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_121__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_121__ap_start;
  wire C_drain_IO_L1_out_wrapper_121__ap_ready;
  wire C_drain_IO_L1_out_wrapper_121__ap_done;
  wire C_drain_IO_L1_out_wrapper_121__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_121__state;
  wire C_drain_IO_L1_out_wrapper_122__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_122__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_122__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_122__ap_start;
  wire C_drain_IO_L1_out_wrapper_122__ap_ready;
  wire C_drain_IO_L1_out_wrapper_122__ap_done;
  wire C_drain_IO_L1_out_wrapper_122__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_122__state;
  wire C_drain_IO_L1_out_wrapper_123__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_123__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_123__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_123__ap_start;
  wire C_drain_IO_L1_out_wrapper_123__ap_ready;
  wire C_drain_IO_L1_out_wrapper_123__ap_done;
  wire C_drain_IO_L1_out_wrapper_123__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_123__state;
  wire C_drain_IO_L1_out_wrapper_124__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_124__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_124__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_124__ap_start;
  wire C_drain_IO_L1_out_wrapper_124__ap_ready;
  wire C_drain_IO_L1_out_wrapper_124__ap_done;
  wire C_drain_IO_L1_out_wrapper_124__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_124__state;
  wire C_drain_IO_L1_out_wrapper_125__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_125__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_125__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_125__ap_start;
  wire C_drain_IO_L1_out_wrapper_125__ap_ready;
  wire C_drain_IO_L1_out_wrapper_125__ap_done;
  wire C_drain_IO_L1_out_wrapper_125__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_125__state;
  wire C_drain_IO_L1_out_wrapper_126__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_126__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_126__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_126__ap_start;
  wire C_drain_IO_L1_out_wrapper_126__ap_ready;
  wire C_drain_IO_L1_out_wrapper_126__ap_done;
  wire C_drain_IO_L1_out_wrapper_126__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_126__state;
  wire C_drain_IO_L1_out_wrapper_127__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_127__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_127__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_127__ap_start;
  wire C_drain_IO_L1_out_wrapper_127__ap_ready;
  wire C_drain_IO_L1_out_wrapper_127__ap_done;
  wire C_drain_IO_L1_out_wrapper_127__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_127__state;
  wire C_drain_IO_L1_out_wrapper_128__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_128__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_128__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_128__ap_start;
  wire C_drain_IO_L1_out_wrapper_128__ap_ready;
  wire C_drain_IO_L1_out_wrapper_128__ap_done;
  wire C_drain_IO_L1_out_wrapper_128__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_128__state;
  wire C_drain_IO_L1_out_wrapper_129__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_129__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_129__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_129__ap_start;
  wire C_drain_IO_L1_out_wrapper_129__ap_ready;
  wire C_drain_IO_L1_out_wrapper_129__ap_done;
  wire C_drain_IO_L1_out_wrapper_129__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_129__state;
  wire C_drain_IO_L1_out_wrapper_130__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_130__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_130__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_130__ap_start;
  wire C_drain_IO_L1_out_wrapper_130__ap_ready;
  wire C_drain_IO_L1_out_wrapper_130__ap_done;
  wire C_drain_IO_L1_out_wrapper_130__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_130__state;
  wire C_drain_IO_L1_out_wrapper_131__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_131__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_131__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_131__ap_start;
  wire C_drain_IO_L1_out_wrapper_131__ap_ready;
  wire C_drain_IO_L1_out_wrapper_131__ap_done;
  wire C_drain_IO_L1_out_wrapper_131__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_131__state;
  wire C_drain_IO_L1_out_wrapper_132__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_132__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_132__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_132__ap_start;
  wire C_drain_IO_L1_out_wrapper_132__ap_ready;
  wire C_drain_IO_L1_out_wrapper_132__ap_done;
  wire C_drain_IO_L1_out_wrapper_132__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_132__state;
  wire C_drain_IO_L1_out_wrapper_133__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_133__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_133__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_133__ap_start;
  wire C_drain_IO_L1_out_wrapper_133__ap_ready;
  wire C_drain_IO_L1_out_wrapper_133__ap_done;
  wire C_drain_IO_L1_out_wrapper_133__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_133__state;
  wire C_drain_IO_L1_out_wrapper_134__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_134__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_134__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_134__ap_start;
  wire C_drain_IO_L1_out_wrapper_134__ap_ready;
  wire C_drain_IO_L1_out_wrapper_134__ap_done;
  wire C_drain_IO_L1_out_wrapper_134__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_134__state;
  wire C_drain_IO_L1_out_wrapper_135__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_135__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_135__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_135__ap_start;
  wire C_drain_IO_L1_out_wrapper_135__ap_ready;
  wire C_drain_IO_L1_out_wrapper_135__ap_done;
  wire C_drain_IO_L1_out_wrapper_135__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_135__state;
  wire C_drain_IO_L1_out_wrapper_136__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_136__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_136__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_136__ap_start;
  wire C_drain_IO_L1_out_wrapper_136__ap_ready;
  wire C_drain_IO_L1_out_wrapper_136__ap_done;
  wire C_drain_IO_L1_out_wrapper_136__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_136__state;
  wire C_drain_IO_L1_out_wrapper_137__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_137__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_137__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_137__ap_start;
  wire C_drain_IO_L1_out_wrapper_137__ap_ready;
  wire C_drain_IO_L1_out_wrapper_137__ap_done;
  wire C_drain_IO_L1_out_wrapper_137__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_137__state;
  wire C_drain_IO_L1_out_wrapper_138__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_138__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_138__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_138__ap_start;
  wire C_drain_IO_L1_out_wrapper_138__ap_ready;
  wire C_drain_IO_L1_out_wrapper_138__ap_done;
  wire C_drain_IO_L1_out_wrapper_138__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_138__state;
  wire C_drain_IO_L1_out_wrapper_139__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_139__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_139__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_139__ap_start;
  wire C_drain_IO_L1_out_wrapper_139__ap_ready;
  wire C_drain_IO_L1_out_wrapper_139__ap_done;
  wire C_drain_IO_L1_out_wrapper_139__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_139__state;
  wire C_drain_IO_L1_out_wrapper_140__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_140__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_140__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_140__ap_start;
  wire C_drain_IO_L1_out_wrapper_140__ap_ready;
  wire C_drain_IO_L1_out_wrapper_140__ap_done;
  wire C_drain_IO_L1_out_wrapper_140__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_140__state;
  wire C_drain_IO_L1_out_wrapper_141__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_141__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_141__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_141__ap_start;
  wire C_drain_IO_L1_out_wrapper_141__ap_ready;
  wire C_drain_IO_L1_out_wrapper_141__ap_done;
  wire C_drain_IO_L1_out_wrapper_141__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_141__state;
  wire C_drain_IO_L1_out_wrapper_142__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_142__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_142__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_142__ap_start;
  wire C_drain_IO_L1_out_wrapper_142__ap_ready;
  wire C_drain_IO_L1_out_wrapper_142__ap_done;
  wire C_drain_IO_L1_out_wrapper_142__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_142__state;
  wire C_drain_IO_L1_out_wrapper_143__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_143__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_143__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_143__ap_start;
  wire C_drain_IO_L1_out_wrapper_143__ap_ready;
  wire C_drain_IO_L1_out_wrapper_143__ap_done;
  wire C_drain_IO_L1_out_wrapper_143__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_143__state;
  wire C_drain_IO_L1_out_wrapper_144__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_144__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_144__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_144__ap_start;
  wire C_drain_IO_L1_out_wrapper_144__ap_ready;
  wire C_drain_IO_L1_out_wrapper_144__ap_done;
  wire C_drain_IO_L1_out_wrapper_144__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_144__state;
  wire C_drain_IO_L1_out_wrapper_145__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_145__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_145__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_145__ap_start;
  wire C_drain_IO_L1_out_wrapper_145__ap_ready;
  wire C_drain_IO_L1_out_wrapper_145__ap_done;
  wire C_drain_IO_L1_out_wrapper_145__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_145__state;
  wire C_drain_IO_L1_out_wrapper_146__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_146__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_146__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_146__ap_start;
  wire C_drain_IO_L1_out_wrapper_146__ap_ready;
  wire C_drain_IO_L1_out_wrapper_146__ap_done;
  wire C_drain_IO_L1_out_wrapper_146__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_146__state;
  wire C_drain_IO_L1_out_wrapper_147__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_147__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_147__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_147__ap_start;
  wire C_drain_IO_L1_out_wrapper_147__ap_ready;
  wire C_drain_IO_L1_out_wrapper_147__ap_done;
  wire C_drain_IO_L1_out_wrapper_147__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_147__state;
  wire C_drain_IO_L1_out_wrapper_148__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_148__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_148__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_148__ap_start;
  wire C_drain_IO_L1_out_wrapper_148__ap_ready;
  wire C_drain_IO_L1_out_wrapper_148__ap_done;
  wire C_drain_IO_L1_out_wrapper_148__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_148__state;
  wire C_drain_IO_L1_out_wrapper_149__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_149__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_149__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_149__ap_start;
  wire C_drain_IO_L1_out_wrapper_149__ap_ready;
  wire C_drain_IO_L1_out_wrapper_149__ap_done;
  wire C_drain_IO_L1_out_wrapper_149__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_149__state;
  wire C_drain_IO_L1_out_wrapper_150__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_150__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_150__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_150__ap_start;
  wire C_drain_IO_L1_out_wrapper_150__ap_ready;
  wire C_drain_IO_L1_out_wrapper_150__ap_done;
  wire C_drain_IO_L1_out_wrapper_150__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_150__state;
  wire C_drain_IO_L1_out_wrapper_151__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_151__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_151__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_151__ap_start;
  wire C_drain_IO_L1_out_wrapper_151__ap_ready;
  wire C_drain_IO_L1_out_wrapper_151__ap_done;
  wire C_drain_IO_L1_out_wrapper_151__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_151__state;
  wire C_drain_IO_L1_out_wrapper_152__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_152__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_152__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_152__ap_start;
  wire C_drain_IO_L1_out_wrapper_152__ap_ready;
  wire C_drain_IO_L1_out_wrapper_152__ap_done;
  wire C_drain_IO_L1_out_wrapper_152__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_152__state;
  wire C_drain_IO_L1_out_wrapper_153__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_153__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_153__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_153__ap_start;
  wire C_drain_IO_L1_out_wrapper_153__ap_ready;
  wire C_drain_IO_L1_out_wrapper_153__ap_done;
  wire C_drain_IO_L1_out_wrapper_153__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_153__state;
  wire C_drain_IO_L1_out_wrapper_154__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_154__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_154__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_154__ap_start;
  wire C_drain_IO_L1_out_wrapper_154__ap_ready;
  wire C_drain_IO_L1_out_wrapper_154__ap_done;
  wire C_drain_IO_L1_out_wrapper_154__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_154__state;
  wire C_drain_IO_L1_out_wrapper_155__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_155__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_155__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_155__ap_start;
  wire C_drain_IO_L1_out_wrapper_155__ap_ready;
  wire C_drain_IO_L1_out_wrapper_155__ap_done;
  wire C_drain_IO_L1_out_wrapper_155__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_155__state;
  wire C_drain_IO_L1_out_wrapper_156__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_156__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_156__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_156__ap_start;
  wire C_drain_IO_L1_out_wrapper_156__ap_ready;
  wire C_drain_IO_L1_out_wrapper_156__ap_done;
  wire C_drain_IO_L1_out_wrapper_156__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_156__state;
  wire C_drain_IO_L1_out_wrapper_157__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_157__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_157__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_157__ap_start;
  wire C_drain_IO_L1_out_wrapper_157__ap_ready;
  wire C_drain_IO_L1_out_wrapper_157__ap_done;
  wire C_drain_IO_L1_out_wrapper_157__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_157__state;
  wire C_drain_IO_L1_out_wrapper_158__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_158__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_158__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_158__ap_start;
  wire C_drain_IO_L1_out_wrapper_158__ap_ready;
  wire C_drain_IO_L1_out_wrapper_158__ap_done;
  wire C_drain_IO_L1_out_wrapper_158__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_158__state;
  wire C_drain_IO_L1_out_wrapper_159__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_159__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_159__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_159__ap_start;
  wire C_drain_IO_L1_out_wrapper_159__ap_ready;
  wire C_drain_IO_L1_out_wrapper_159__ap_done;
  wire C_drain_IO_L1_out_wrapper_159__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_159__state;
  wire C_drain_IO_L1_out_wrapper_160__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_160__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_160__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_160__ap_start;
  wire C_drain_IO_L1_out_wrapper_160__ap_ready;
  wire C_drain_IO_L1_out_wrapper_160__ap_done;
  wire C_drain_IO_L1_out_wrapper_160__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_160__state;
  wire C_drain_IO_L1_out_wrapper_161__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_161__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_161__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_161__ap_start;
  wire C_drain_IO_L1_out_wrapper_161__ap_ready;
  wire C_drain_IO_L1_out_wrapper_161__ap_done;
  wire C_drain_IO_L1_out_wrapper_161__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_161__state;
  wire C_drain_IO_L1_out_wrapper_162__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_162__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_162__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_162__ap_start;
  wire C_drain_IO_L1_out_wrapper_162__ap_ready;
  wire C_drain_IO_L1_out_wrapper_162__ap_done;
  wire C_drain_IO_L1_out_wrapper_162__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_162__state;
  wire C_drain_IO_L1_out_wrapper_163__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_163__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_163__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_163__ap_start;
  wire C_drain_IO_L1_out_wrapper_163__ap_ready;
  wire C_drain_IO_L1_out_wrapper_163__ap_done;
  wire C_drain_IO_L1_out_wrapper_163__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_163__state;
  wire C_drain_IO_L1_out_wrapper_164__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_164__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_164__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_164__ap_start;
  wire C_drain_IO_L1_out_wrapper_164__ap_ready;
  wire C_drain_IO_L1_out_wrapper_164__ap_done;
  wire C_drain_IO_L1_out_wrapper_164__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_164__state;
  wire C_drain_IO_L1_out_wrapper_165__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_165__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_165__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_165__ap_start;
  wire C_drain_IO_L1_out_wrapper_165__ap_ready;
  wire C_drain_IO_L1_out_wrapper_165__ap_done;
  wire C_drain_IO_L1_out_wrapper_165__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_165__state;
  wire C_drain_IO_L1_out_wrapper_166__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_166__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_166__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_166__ap_start;
  wire C_drain_IO_L1_out_wrapper_166__ap_ready;
  wire C_drain_IO_L1_out_wrapper_166__ap_done;
  wire C_drain_IO_L1_out_wrapper_166__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_166__state;
  wire C_drain_IO_L1_out_wrapper_167__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_167__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_167__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_167__ap_start;
  wire C_drain_IO_L1_out_wrapper_167__ap_ready;
  wire C_drain_IO_L1_out_wrapper_167__ap_done;
  wire C_drain_IO_L1_out_wrapper_167__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_167__state;
  wire C_drain_IO_L1_out_wrapper_168__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_168__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_168__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_168__ap_start;
  wire C_drain_IO_L1_out_wrapper_168__ap_ready;
  wire C_drain_IO_L1_out_wrapper_168__ap_done;
  wire C_drain_IO_L1_out_wrapper_168__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_168__state;
  wire C_drain_IO_L1_out_wrapper_169__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_169__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_169__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_169__ap_start;
  wire C_drain_IO_L1_out_wrapper_169__ap_ready;
  wire C_drain_IO_L1_out_wrapper_169__ap_done;
  wire C_drain_IO_L1_out_wrapper_169__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_169__state;
  wire C_drain_IO_L1_out_wrapper_170__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_170__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_170__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_170__ap_start;
  wire C_drain_IO_L1_out_wrapper_170__ap_ready;
  wire C_drain_IO_L1_out_wrapper_170__ap_done;
  wire C_drain_IO_L1_out_wrapper_170__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_170__state;
  wire C_drain_IO_L1_out_wrapper_171__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_171__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_171__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_171__ap_start;
  wire C_drain_IO_L1_out_wrapper_171__ap_ready;
  wire C_drain_IO_L1_out_wrapper_171__ap_done;
  wire C_drain_IO_L1_out_wrapper_171__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_171__state;
  wire C_drain_IO_L1_out_wrapper_172__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_172__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_172__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_172__ap_start;
  wire C_drain_IO_L1_out_wrapper_172__ap_ready;
  wire C_drain_IO_L1_out_wrapper_172__ap_done;
  wire C_drain_IO_L1_out_wrapper_172__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_172__state;
  wire C_drain_IO_L1_out_wrapper_173__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_173__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_173__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_173__ap_start;
  wire C_drain_IO_L1_out_wrapper_173__ap_ready;
  wire C_drain_IO_L1_out_wrapper_173__ap_done;
  wire C_drain_IO_L1_out_wrapper_173__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_173__state;
  wire C_drain_IO_L1_out_wrapper_174__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_174__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_174__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_174__ap_start;
  wire C_drain_IO_L1_out_wrapper_174__ap_ready;
  wire C_drain_IO_L1_out_wrapper_174__ap_done;
  wire C_drain_IO_L1_out_wrapper_174__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_174__state;
  wire C_drain_IO_L1_out_wrapper_175__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_175__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_175__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_175__ap_start;
  wire C_drain_IO_L1_out_wrapper_175__ap_ready;
  wire C_drain_IO_L1_out_wrapper_175__ap_done;
  wire C_drain_IO_L1_out_wrapper_175__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_175__state;
  wire C_drain_IO_L1_out_wrapper_176__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_176__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_176__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_176__ap_start;
  wire C_drain_IO_L1_out_wrapper_176__ap_ready;
  wire C_drain_IO_L1_out_wrapper_176__ap_done;
  wire C_drain_IO_L1_out_wrapper_176__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_176__state;
  wire C_drain_IO_L1_out_wrapper_177__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_177__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_177__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_177__ap_start;
  wire C_drain_IO_L1_out_wrapper_177__ap_ready;
  wire C_drain_IO_L1_out_wrapper_177__ap_done;
  wire C_drain_IO_L1_out_wrapper_177__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_177__state;
  wire C_drain_IO_L1_out_wrapper_178__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_178__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_178__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_178__ap_start;
  wire C_drain_IO_L1_out_wrapper_178__ap_ready;
  wire C_drain_IO_L1_out_wrapper_178__ap_done;
  wire C_drain_IO_L1_out_wrapper_178__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_178__state;
  wire C_drain_IO_L1_out_wrapper_179__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_179__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_179__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_179__ap_start;
  wire C_drain_IO_L1_out_wrapper_179__ap_ready;
  wire C_drain_IO_L1_out_wrapper_179__ap_done;
  wire C_drain_IO_L1_out_wrapper_179__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_179__state;
  wire C_drain_IO_L1_out_wrapper_180__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_180__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_180__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_180__ap_start;
  wire C_drain_IO_L1_out_wrapper_180__ap_ready;
  wire C_drain_IO_L1_out_wrapper_180__ap_done;
  wire C_drain_IO_L1_out_wrapper_180__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_180__state;
  wire C_drain_IO_L1_out_wrapper_181__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_181__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_181__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_181__ap_start;
  wire C_drain_IO_L1_out_wrapper_181__ap_ready;
  wire C_drain_IO_L1_out_wrapper_181__ap_done;
  wire C_drain_IO_L1_out_wrapper_181__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_181__state;
  wire C_drain_IO_L1_out_wrapper_182__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_182__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_182__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_182__ap_start;
  wire C_drain_IO_L1_out_wrapper_182__ap_ready;
  wire C_drain_IO_L1_out_wrapper_182__ap_done;
  wire C_drain_IO_L1_out_wrapper_182__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_182__state;
  wire C_drain_IO_L1_out_wrapper_183__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_183__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_183__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_183__ap_start;
  wire C_drain_IO_L1_out_wrapper_183__ap_ready;
  wire C_drain_IO_L1_out_wrapper_183__ap_done;
  wire C_drain_IO_L1_out_wrapper_183__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_183__state;
  wire C_drain_IO_L1_out_wrapper_184__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_184__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_184__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_184__ap_start;
  wire C_drain_IO_L1_out_wrapper_184__ap_ready;
  wire C_drain_IO_L1_out_wrapper_184__ap_done;
  wire C_drain_IO_L1_out_wrapper_184__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_184__state;
  wire C_drain_IO_L1_out_wrapper_185__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_185__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_185__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_185__ap_start;
  wire C_drain_IO_L1_out_wrapper_185__ap_ready;
  wire C_drain_IO_L1_out_wrapper_185__ap_done;
  wire C_drain_IO_L1_out_wrapper_185__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_185__state;
  wire C_drain_IO_L1_out_wrapper_186__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_186__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_186__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_186__ap_start;
  wire C_drain_IO_L1_out_wrapper_186__ap_ready;
  wire C_drain_IO_L1_out_wrapper_186__ap_done;
  wire C_drain_IO_L1_out_wrapper_186__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_186__state;
  wire C_drain_IO_L1_out_wrapper_187__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_187__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_187__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_187__ap_start;
  wire C_drain_IO_L1_out_wrapper_187__ap_ready;
  wire C_drain_IO_L1_out_wrapper_187__ap_done;
  wire C_drain_IO_L1_out_wrapper_187__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_187__state;
  wire C_drain_IO_L1_out_wrapper_188__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_188__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_188__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_188__ap_start;
  wire C_drain_IO_L1_out_wrapper_188__ap_ready;
  wire C_drain_IO_L1_out_wrapper_188__ap_done;
  wire C_drain_IO_L1_out_wrapper_188__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_188__state;
  wire C_drain_IO_L1_out_wrapper_189__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_189__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_189__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_189__ap_start;
  wire C_drain_IO_L1_out_wrapper_189__ap_ready;
  wire C_drain_IO_L1_out_wrapper_189__ap_done;
  wire C_drain_IO_L1_out_wrapper_189__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_189__state;
  wire C_drain_IO_L1_out_wrapper_190__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_190__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_190__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_190__ap_start;
  wire C_drain_IO_L1_out_wrapper_190__ap_ready;
  wire C_drain_IO_L1_out_wrapper_190__ap_done;
  wire C_drain_IO_L1_out_wrapper_190__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_190__state;
  wire C_drain_IO_L1_out_wrapper_191__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_191__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_191__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_191__ap_start;
  wire C_drain_IO_L1_out_wrapper_191__ap_ready;
  wire C_drain_IO_L1_out_wrapper_191__ap_done;
  wire C_drain_IO_L1_out_wrapper_191__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_191__state;
  wire C_drain_IO_L1_out_wrapper_192__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_192__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_192__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_192__ap_start;
  wire C_drain_IO_L1_out_wrapper_192__ap_ready;
  wire C_drain_IO_L1_out_wrapper_192__ap_done;
  wire C_drain_IO_L1_out_wrapper_192__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_192__state;
  wire C_drain_IO_L1_out_wrapper_193__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_193__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_193__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_193__ap_start;
  wire C_drain_IO_L1_out_wrapper_193__ap_ready;
  wire C_drain_IO_L1_out_wrapper_193__ap_done;
  wire C_drain_IO_L1_out_wrapper_193__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_193__state;
  wire C_drain_IO_L1_out_wrapper_194__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_194__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_194__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_194__ap_start;
  wire C_drain_IO_L1_out_wrapper_194__ap_ready;
  wire C_drain_IO_L1_out_wrapper_194__ap_done;
  wire C_drain_IO_L1_out_wrapper_194__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_194__state;
  wire C_drain_IO_L1_out_wrapper_195__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_195__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_195__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_195__ap_start;
  wire C_drain_IO_L1_out_wrapper_195__ap_ready;
  wire C_drain_IO_L1_out_wrapper_195__ap_done;
  wire C_drain_IO_L1_out_wrapper_195__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_195__state;
  wire C_drain_IO_L1_out_wrapper_196__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_196__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_196__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_196__ap_start;
  wire C_drain_IO_L1_out_wrapper_196__ap_ready;
  wire C_drain_IO_L1_out_wrapper_196__ap_done;
  wire C_drain_IO_L1_out_wrapper_196__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_196__state;
  wire C_drain_IO_L1_out_wrapper_197__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_197__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_197__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_197__ap_start;
  wire C_drain_IO_L1_out_wrapper_197__ap_ready;
  wire C_drain_IO_L1_out_wrapper_197__ap_done;
  wire C_drain_IO_L1_out_wrapper_197__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_197__state;
  wire C_drain_IO_L1_out_wrapper_198__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_198__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_198__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_198__ap_start;
  wire C_drain_IO_L1_out_wrapper_198__ap_ready;
  wire C_drain_IO_L1_out_wrapper_198__ap_done;
  wire C_drain_IO_L1_out_wrapper_198__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_198__state;
  wire C_drain_IO_L1_out_wrapper_199__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_199__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_199__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_199__ap_start;
  wire C_drain_IO_L1_out_wrapper_199__ap_ready;
  wire C_drain_IO_L1_out_wrapper_199__ap_done;
  wire C_drain_IO_L1_out_wrapper_199__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_199__state;
  wire C_drain_IO_L1_out_wrapper_200__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_200__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_200__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_200__ap_start;
  wire C_drain_IO_L1_out_wrapper_200__ap_ready;
  wire C_drain_IO_L1_out_wrapper_200__ap_done;
  wire C_drain_IO_L1_out_wrapper_200__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_200__state;
  wire C_drain_IO_L1_out_wrapper_201__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_201__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_201__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_201__ap_start;
  wire C_drain_IO_L1_out_wrapper_201__ap_ready;
  wire C_drain_IO_L1_out_wrapper_201__ap_done;
  wire C_drain_IO_L1_out_wrapper_201__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_201__state;
  wire C_drain_IO_L1_out_wrapper_202__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_202__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_202__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_202__ap_start;
  wire C_drain_IO_L1_out_wrapper_202__ap_ready;
  wire C_drain_IO_L1_out_wrapper_202__ap_done;
  wire C_drain_IO_L1_out_wrapper_202__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_202__state;
  wire C_drain_IO_L1_out_wrapper_203__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_203__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_203__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_203__ap_start;
  wire C_drain_IO_L1_out_wrapper_203__ap_ready;
  wire C_drain_IO_L1_out_wrapper_203__ap_done;
  wire C_drain_IO_L1_out_wrapper_203__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_203__state;
  wire C_drain_IO_L1_out_wrapper_204__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_204__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_204__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_204__ap_start;
  wire C_drain_IO_L1_out_wrapper_204__ap_ready;
  wire C_drain_IO_L1_out_wrapper_204__ap_done;
  wire C_drain_IO_L1_out_wrapper_204__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_204__state;
  wire C_drain_IO_L1_out_wrapper_205__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_205__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_205__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_205__ap_start;
  wire C_drain_IO_L1_out_wrapper_205__ap_ready;
  wire C_drain_IO_L1_out_wrapper_205__ap_done;
  wire C_drain_IO_L1_out_wrapper_205__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_205__state;
  wire C_drain_IO_L1_out_wrapper_206__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_206__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_206__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_206__ap_start;
  wire C_drain_IO_L1_out_wrapper_206__ap_ready;
  wire C_drain_IO_L1_out_wrapper_206__ap_done;
  wire C_drain_IO_L1_out_wrapper_206__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_206__state;
  wire C_drain_IO_L1_out_wrapper_207__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_207__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_207__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_207__ap_start;
  wire C_drain_IO_L1_out_wrapper_207__ap_ready;
  wire C_drain_IO_L1_out_wrapper_207__ap_done;
  wire C_drain_IO_L1_out_wrapper_207__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_207__state;
  wire C_drain_IO_L1_out_wrapper_208__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_208__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_208__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_208__ap_start;
  wire C_drain_IO_L1_out_wrapper_208__ap_ready;
  wire C_drain_IO_L1_out_wrapper_208__ap_done;
  wire C_drain_IO_L1_out_wrapper_208__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_208__state;
  wire C_drain_IO_L1_out_wrapper_209__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_209__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_209__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_209__ap_start;
  wire C_drain_IO_L1_out_wrapper_209__ap_ready;
  wire C_drain_IO_L1_out_wrapper_209__ap_done;
  wire C_drain_IO_L1_out_wrapper_209__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_209__state;
  wire C_drain_IO_L1_out_wrapper_210__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_210__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_210__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_210__ap_start;
  wire C_drain_IO_L1_out_wrapper_210__ap_ready;
  wire C_drain_IO_L1_out_wrapper_210__ap_done;
  wire C_drain_IO_L1_out_wrapper_210__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_210__state;
  wire C_drain_IO_L1_out_wrapper_211__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_211__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_211__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_211__ap_start;
  wire C_drain_IO_L1_out_wrapper_211__ap_ready;
  wire C_drain_IO_L1_out_wrapper_211__ap_done;
  wire C_drain_IO_L1_out_wrapper_211__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_211__state;
  wire C_drain_IO_L1_out_wrapper_212__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_212__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_212__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_212__ap_start;
  wire C_drain_IO_L1_out_wrapper_212__ap_ready;
  wire C_drain_IO_L1_out_wrapper_212__ap_done;
  wire C_drain_IO_L1_out_wrapper_212__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_212__state;
  wire C_drain_IO_L1_out_wrapper_213__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_213__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_213__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_213__ap_start;
  wire C_drain_IO_L1_out_wrapper_213__ap_ready;
  wire C_drain_IO_L1_out_wrapper_213__ap_done;
  wire C_drain_IO_L1_out_wrapper_213__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_213__state;
  wire C_drain_IO_L1_out_wrapper_214__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_214__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_214__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_214__ap_start;
  wire C_drain_IO_L1_out_wrapper_214__ap_ready;
  wire C_drain_IO_L1_out_wrapper_214__ap_done;
  wire C_drain_IO_L1_out_wrapper_214__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_214__state;
  wire C_drain_IO_L1_out_wrapper_215__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_215__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_215__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_215__ap_start;
  wire C_drain_IO_L1_out_wrapper_215__ap_ready;
  wire C_drain_IO_L1_out_wrapper_215__ap_done;
  wire C_drain_IO_L1_out_wrapper_215__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_215__state;
  wire C_drain_IO_L1_out_wrapper_216__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_216__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_216__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_216__ap_start;
  wire C_drain_IO_L1_out_wrapper_216__ap_ready;
  wire C_drain_IO_L1_out_wrapper_216__ap_done;
  wire C_drain_IO_L1_out_wrapper_216__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_216__state;
  wire C_drain_IO_L1_out_wrapper_217__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_217__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_217__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_217__ap_start;
  wire C_drain_IO_L1_out_wrapper_217__ap_ready;
  wire C_drain_IO_L1_out_wrapper_217__ap_done;
  wire C_drain_IO_L1_out_wrapper_217__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_217__state;
  wire C_drain_IO_L1_out_wrapper_218__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_218__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_218__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_218__ap_start;
  wire C_drain_IO_L1_out_wrapper_218__ap_ready;
  wire C_drain_IO_L1_out_wrapper_218__ap_done;
  wire C_drain_IO_L1_out_wrapper_218__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_218__state;
  wire C_drain_IO_L1_out_wrapper_219__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_219__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_219__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_219__ap_start;
  wire C_drain_IO_L1_out_wrapper_219__ap_ready;
  wire C_drain_IO_L1_out_wrapper_219__ap_done;
  wire C_drain_IO_L1_out_wrapper_219__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_219__state;
  wire C_drain_IO_L1_out_wrapper_220__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_220__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_220__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_220__ap_start;
  wire C_drain_IO_L1_out_wrapper_220__ap_ready;
  wire C_drain_IO_L1_out_wrapper_220__ap_done;
  wire C_drain_IO_L1_out_wrapper_220__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_220__state;
  wire C_drain_IO_L1_out_wrapper_221__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_221__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_221__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_221__ap_start;
  wire C_drain_IO_L1_out_wrapper_221__ap_ready;
  wire C_drain_IO_L1_out_wrapper_221__ap_done;
  wire C_drain_IO_L1_out_wrapper_221__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_221__state;
  wire C_drain_IO_L1_out_wrapper_222__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_222__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_222__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_222__ap_start;
  wire C_drain_IO_L1_out_wrapper_222__ap_ready;
  wire C_drain_IO_L1_out_wrapper_222__ap_done;
  wire C_drain_IO_L1_out_wrapper_222__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_222__state;
  wire C_drain_IO_L1_out_wrapper_223__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_223__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_223__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_223__ap_start;
  wire C_drain_IO_L1_out_wrapper_223__ap_ready;
  wire C_drain_IO_L1_out_wrapper_223__ap_done;
  wire C_drain_IO_L1_out_wrapper_223__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_223__state;
  wire C_drain_IO_L1_out_wrapper_224__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_224__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_224__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_224__ap_start;
  wire C_drain_IO_L1_out_wrapper_224__ap_ready;
  wire C_drain_IO_L1_out_wrapper_224__ap_done;
  wire C_drain_IO_L1_out_wrapper_224__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_224__state;
  wire C_drain_IO_L1_out_wrapper_225__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_225__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_225__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_225__ap_start;
  wire C_drain_IO_L1_out_wrapper_225__ap_ready;
  wire C_drain_IO_L1_out_wrapper_225__ap_done;
  wire C_drain_IO_L1_out_wrapper_225__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_225__state;
  wire C_drain_IO_L1_out_wrapper_226__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_226__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_226__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_226__ap_start;
  wire C_drain_IO_L1_out_wrapper_226__ap_ready;
  wire C_drain_IO_L1_out_wrapper_226__ap_done;
  wire C_drain_IO_L1_out_wrapper_226__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_226__state;
  wire C_drain_IO_L1_out_wrapper_227__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_227__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_227__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_227__ap_start;
  wire C_drain_IO_L1_out_wrapper_227__ap_ready;
  wire C_drain_IO_L1_out_wrapper_227__ap_done;
  wire C_drain_IO_L1_out_wrapper_227__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_227__state;
  wire C_drain_IO_L1_out_wrapper_228__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_228__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_228__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_228__ap_start;
  wire C_drain_IO_L1_out_wrapper_228__ap_ready;
  wire C_drain_IO_L1_out_wrapper_228__ap_done;
  wire C_drain_IO_L1_out_wrapper_228__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_228__state;
  wire C_drain_IO_L1_out_wrapper_229__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_229__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_229__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_229__ap_start;
  wire C_drain_IO_L1_out_wrapper_229__ap_ready;
  wire C_drain_IO_L1_out_wrapper_229__ap_done;
  wire C_drain_IO_L1_out_wrapper_229__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_229__state;
  wire C_drain_IO_L1_out_wrapper_230__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_230__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_230__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_230__ap_start;
  wire C_drain_IO_L1_out_wrapper_230__ap_ready;
  wire C_drain_IO_L1_out_wrapper_230__ap_done;
  wire C_drain_IO_L1_out_wrapper_230__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_230__state;
  wire C_drain_IO_L1_out_wrapper_231__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_231__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_231__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_231__ap_start;
  wire C_drain_IO_L1_out_wrapper_231__ap_ready;
  wire C_drain_IO_L1_out_wrapper_231__ap_done;
  wire C_drain_IO_L1_out_wrapper_231__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_231__state;
  wire C_drain_IO_L1_out_wrapper_232__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_232__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_232__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_232__ap_start;
  wire C_drain_IO_L1_out_wrapper_232__ap_ready;
  wire C_drain_IO_L1_out_wrapper_232__ap_done;
  wire C_drain_IO_L1_out_wrapper_232__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_232__state;
  wire C_drain_IO_L1_out_wrapper_233__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_233__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_233__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_233__ap_start;
  wire C_drain_IO_L1_out_wrapper_233__ap_ready;
  wire C_drain_IO_L1_out_wrapper_233__ap_done;
  wire C_drain_IO_L1_out_wrapper_233__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_233__state;
  wire C_drain_IO_L1_out_wrapper_234__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_234__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_234__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_234__ap_start;
  wire C_drain_IO_L1_out_wrapper_234__ap_ready;
  wire C_drain_IO_L1_out_wrapper_234__ap_done;
  wire C_drain_IO_L1_out_wrapper_234__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_234__state;
  wire C_drain_IO_L1_out_wrapper_235__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_235__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_235__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_235__ap_start;
  wire C_drain_IO_L1_out_wrapper_235__ap_ready;
  wire C_drain_IO_L1_out_wrapper_235__ap_done;
  wire C_drain_IO_L1_out_wrapper_235__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_235__state;
  wire C_drain_IO_L1_out_wrapper_236__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_236__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_236__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_236__ap_start;
  wire C_drain_IO_L1_out_wrapper_236__ap_ready;
  wire C_drain_IO_L1_out_wrapper_236__ap_done;
  wire C_drain_IO_L1_out_wrapper_236__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_236__state;
  wire C_drain_IO_L1_out_wrapper_237__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_237__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_237__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_237__ap_start;
  wire C_drain_IO_L1_out_wrapper_237__ap_ready;
  wire C_drain_IO_L1_out_wrapper_237__ap_done;
  wire C_drain_IO_L1_out_wrapper_237__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_237__state;
  wire C_drain_IO_L1_out_wrapper_238__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_238__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_238__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_238__ap_start;
  wire C_drain_IO_L1_out_wrapper_238__ap_ready;
  wire C_drain_IO_L1_out_wrapper_238__ap_done;
  wire C_drain_IO_L1_out_wrapper_238__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_238__state;
  wire C_drain_IO_L1_out_wrapper_239__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_239__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_239__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_239__ap_start;
  wire C_drain_IO_L1_out_wrapper_239__ap_ready;
  wire C_drain_IO_L1_out_wrapper_239__ap_done;
  wire C_drain_IO_L1_out_wrapper_239__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_239__state;
  wire C_drain_IO_L1_out_wrapper_240__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_240__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_240__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_240__ap_start;
  wire C_drain_IO_L1_out_wrapper_240__ap_ready;
  wire C_drain_IO_L1_out_wrapper_240__ap_done;
  wire C_drain_IO_L1_out_wrapper_240__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_240__state;
  wire C_drain_IO_L1_out_wrapper_241__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_241__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_241__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_241__ap_start;
  wire C_drain_IO_L1_out_wrapper_241__ap_ready;
  wire C_drain_IO_L1_out_wrapper_241__ap_done;
  wire C_drain_IO_L1_out_wrapper_241__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_241__state;
  wire C_drain_IO_L1_out_wrapper_242__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_242__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_242__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_242__ap_start;
  wire C_drain_IO_L1_out_wrapper_242__ap_ready;
  wire C_drain_IO_L1_out_wrapper_242__ap_done;
  wire C_drain_IO_L1_out_wrapper_242__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_242__state;
  wire C_drain_IO_L1_out_wrapper_243__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_243__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_243__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_243__ap_start;
  wire C_drain_IO_L1_out_wrapper_243__ap_ready;
  wire C_drain_IO_L1_out_wrapper_243__ap_done;
  wire C_drain_IO_L1_out_wrapper_243__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_243__state;
  wire C_drain_IO_L1_out_wrapper_244__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_244__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_244__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_244__ap_start;
  wire C_drain_IO_L1_out_wrapper_244__ap_ready;
  wire C_drain_IO_L1_out_wrapper_244__ap_done;
  wire C_drain_IO_L1_out_wrapper_244__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_244__state;
  wire C_drain_IO_L1_out_wrapper_245__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_245__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_245__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_245__ap_start;
  wire C_drain_IO_L1_out_wrapper_245__ap_ready;
  wire C_drain_IO_L1_out_wrapper_245__ap_done;
  wire C_drain_IO_L1_out_wrapper_245__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_245__state;
  wire C_drain_IO_L1_out_wrapper_246__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_246__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_246__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_246__ap_start;
  wire C_drain_IO_L1_out_wrapper_246__ap_ready;
  wire C_drain_IO_L1_out_wrapper_246__ap_done;
  wire C_drain_IO_L1_out_wrapper_246__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_246__state;
  wire C_drain_IO_L1_out_wrapper_247__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_247__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_247__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_247__ap_start;
  wire C_drain_IO_L1_out_wrapper_247__ap_ready;
  wire C_drain_IO_L1_out_wrapper_247__ap_done;
  wire C_drain_IO_L1_out_wrapper_247__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_247__state;
  wire C_drain_IO_L1_out_wrapper_248__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_248__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_248__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_248__ap_start;
  wire C_drain_IO_L1_out_wrapper_248__ap_ready;
  wire C_drain_IO_L1_out_wrapper_248__ap_done;
  wire C_drain_IO_L1_out_wrapper_248__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_248__state;
  wire C_drain_IO_L1_out_wrapper_249__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_249__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_249__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_249__ap_start;
  wire C_drain_IO_L1_out_wrapper_249__ap_ready;
  wire C_drain_IO_L1_out_wrapper_249__ap_done;
  wire C_drain_IO_L1_out_wrapper_249__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_249__state;
  wire C_drain_IO_L1_out_wrapper_250__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_250__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_250__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_250__ap_start;
  wire C_drain_IO_L1_out_wrapper_250__ap_ready;
  wire C_drain_IO_L1_out_wrapper_250__ap_done;
  wire C_drain_IO_L1_out_wrapper_250__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_250__state;
  wire C_drain_IO_L1_out_wrapper_251__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_251__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_251__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_251__ap_start;
  wire C_drain_IO_L1_out_wrapper_251__ap_ready;
  wire C_drain_IO_L1_out_wrapper_251__ap_done;
  wire C_drain_IO_L1_out_wrapper_251__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_251__state;
  wire C_drain_IO_L1_out_wrapper_252__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_252__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_252__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_252__ap_start;
  wire C_drain_IO_L1_out_wrapper_252__ap_ready;
  wire C_drain_IO_L1_out_wrapper_252__ap_done;
  wire C_drain_IO_L1_out_wrapper_252__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_252__state;
  wire C_drain_IO_L1_out_wrapper_253__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_253__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_253__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_253__ap_start;
  wire C_drain_IO_L1_out_wrapper_253__ap_ready;
  wire C_drain_IO_L1_out_wrapper_253__ap_done;
  wire C_drain_IO_L1_out_wrapper_253__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_253__state;
  wire C_drain_IO_L1_out_wrapper_254__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_254__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_254__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_254__ap_start;
  wire C_drain_IO_L1_out_wrapper_254__ap_ready;
  wire C_drain_IO_L1_out_wrapper_254__ap_done;
  wire C_drain_IO_L1_out_wrapper_254__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_254__state;
  wire C_drain_IO_L1_out_wrapper_255__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_255__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_255__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_255__ap_start;
  wire C_drain_IO_L1_out_wrapper_255__ap_ready;
  wire C_drain_IO_L1_out_wrapper_255__ap_done;
  wire C_drain_IO_L1_out_wrapper_255__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_255__state;
  wire C_drain_IO_L1_out_wrapper_256__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_256__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_256__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_256__ap_start;
  wire C_drain_IO_L1_out_wrapper_256__ap_ready;
  wire C_drain_IO_L1_out_wrapper_256__ap_done;
  wire C_drain_IO_L1_out_wrapper_256__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_256__state;
  wire C_drain_IO_L1_out_wrapper_257__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_257__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_257__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_257__ap_start;
  wire C_drain_IO_L1_out_wrapper_257__ap_ready;
  wire C_drain_IO_L1_out_wrapper_257__ap_done;
  wire C_drain_IO_L1_out_wrapper_257__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_257__state;
  wire C_drain_IO_L1_out_wrapper_258__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_258__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_258__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_258__ap_start;
  wire C_drain_IO_L1_out_wrapper_258__ap_ready;
  wire C_drain_IO_L1_out_wrapper_258__ap_done;
  wire C_drain_IO_L1_out_wrapper_258__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_258__state;
  wire C_drain_IO_L1_out_wrapper_259__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_259__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_259__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_259__ap_start;
  wire C_drain_IO_L1_out_wrapper_259__ap_ready;
  wire C_drain_IO_L1_out_wrapper_259__ap_done;
  wire C_drain_IO_L1_out_wrapper_259__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_259__state;
  wire C_drain_IO_L1_out_wrapper_260__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_260__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_260__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_260__ap_start;
  wire C_drain_IO_L1_out_wrapper_260__ap_ready;
  wire C_drain_IO_L1_out_wrapper_260__ap_done;
  wire C_drain_IO_L1_out_wrapper_260__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_260__state;
  wire C_drain_IO_L1_out_wrapper_261__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_261__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_261__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_261__ap_start;
  wire C_drain_IO_L1_out_wrapper_261__ap_ready;
  wire C_drain_IO_L1_out_wrapper_261__ap_done;
  wire C_drain_IO_L1_out_wrapper_261__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_261__state;
  wire C_drain_IO_L1_out_wrapper_262__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_262__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_262__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_262__ap_start;
  wire C_drain_IO_L1_out_wrapper_262__ap_ready;
  wire C_drain_IO_L1_out_wrapper_262__ap_done;
  wire C_drain_IO_L1_out_wrapper_262__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_262__state;
  wire C_drain_IO_L1_out_wrapper_263__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_263__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_263__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_263__ap_start;
  wire C_drain_IO_L1_out_wrapper_263__ap_ready;
  wire C_drain_IO_L1_out_wrapper_263__ap_done;
  wire C_drain_IO_L1_out_wrapper_263__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_263__state;
  wire C_drain_IO_L1_out_wrapper_264__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_264__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_264__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_264__ap_start;
  wire C_drain_IO_L1_out_wrapper_264__ap_ready;
  wire C_drain_IO_L1_out_wrapper_264__ap_done;
  wire C_drain_IO_L1_out_wrapper_264__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_264__state;
  wire C_drain_IO_L1_out_wrapper_265__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_265__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_265__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_265__ap_start;
  wire C_drain_IO_L1_out_wrapper_265__ap_ready;
  wire C_drain_IO_L1_out_wrapper_265__ap_done;
  wire C_drain_IO_L1_out_wrapper_265__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_265__state;
  wire C_drain_IO_L1_out_wrapper_266__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_266__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_266__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_266__ap_start;
  wire C_drain_IO_L1_out_wrapper_266__ap_ready;
  wire C_drain_IO_L1_out_wrapper_266__ap_done;
  wire C_drain_IO_L1_out_wrapper_266__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_266__state;
  wire C_drain_IO_L1_out_wrapper_267__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_267__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_267__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_267__ap_start;
  wire C_drain_IO_L1_out_wrapper_267__ap_ready;
  wire C_drain_IO_L1_out_wrapper_267__ap_done;
  wire C_drain_IO_L1_out_wrapper_267__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_267__state;
  wire C_drain_IO_L1_out_wrapper_268__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_268__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_268__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_268__ap_start;
  wire C_drain_IO_L1_out_wrapper_268__ap_ready;
  wire C_drain_IO_L1_out_wrapper_268__ap_done;
  wire C_drain_IO_L1_out_wrapper_268__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_268__state;
  wire C_drain_IO_L1_out_wrapper_269__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_269__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_269__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_269__ap_start;
  wire C_drain_IO_L1_out_wrapper_269__ap_ready;
  wire C_drain_IO_L1_out_wrapper_269__ap_done;
  wire C_drain_IO_L1_out_wrapper_269__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_269__state;
  wire C_drain_IO_L1_out_wrapper_270__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_270__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_270__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_270__ap_start;
  wire C_drain_IO_L1_out_wrapper_270__ap_ready;
  wire C_drain_IO_L1_out_wrapper_270__ap_done;
  wire C_drain_IO_L1_out_wrapper_270__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_270__state;
  wire C_drain_IO_L1_out_wrapper_271__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_271__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_271__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_271__ap_start;
  wire C_drain_IO_L1_out_wrapper_271__ap_ready;
  wire C_drain_IO_L1_out_wrapper_271__ap_done;
  wire C_drain_IO_L1_out_wrapper_271__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_271__state;
  wire C_drain_IO_L1_out_wrapper_272__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_272__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_272__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_272__ap_start;
  wire C_drain_IO_L1_out_wrapper_272__ap_ready;
  wire C_drain_IO_L1_out_wrapper_272__ap_done;
  wire C_drain_IO_L1_out_wrapper_272__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_272__state;
  wire C_drain_IO_L1_out_wrapper_273__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_273__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_273__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_273__ap_start;
  wire C_drain_IO_L1_out_wrapper_273__ap_ready;
  wire C_drain_IO_L1_out_wrapper_273__ap_done;
  wire C_drain_IO_L1_out_wrapper_273__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_273__state;
  wire C_drain_IO_L1_out_wrapper_274__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_274__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_274__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_274__ap_start;
  wire C_drain_IO_L1_out_wrapper_274__ap_ready;
  wire C_drain_IO_L1_out_wrapper_274__ap_done;
  wire C_drain_IO_L1_out_wrapper_274__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_274__state;
  wire C_drain_IO_L1_out_wrapper_275__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_275__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_275__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_275__ap_start;
  wire C_drain_IO_L1_out_wrapper_275__ap_ready;
  wire C_drain_IO_L1_out_wrapper_275__ap_done;
  wire C_drain_IO_L1_out_wrapper_275__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_275__state;
  wire C_drain_IO_L1_out_wrapper_276__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_276__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_276__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_276__ap_start;
  wire C_drain_IO_L1_out_wrapper_276__ap_ready;
  wire C_drain_IO_L1_out_wrapper_276__ap_done;
  wire C_drain_IO_L1_out_wrapper_276__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_276__state;
  wire C_drain_IO_L1_out_wrapper_277__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_277__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_277__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_277__ap_start;
  wire C_drain_IO_L1_out_wrapper_277__ap_ready;
  wire C_drain_IO_L1_out_wrapper_277__ap_done;
  wire C_drain_IO_L1_out_wrapper_277__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_277__state;
  wire C_drain_IO_L1_out_wrapper_278__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_278__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_278__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_278__ap_start;
  wire C_drain_IO_L1_out_wrapper_278__ap_ready;
  wire C_drain_IO_L1_out_wrapper_278__ap_done;
  wire C_drain_IO_L1_out_wrapper_278__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_278__state;
  wire C_drain_IO_L1_out_wrapper_279__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_279__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_279__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_279__ap_start;
  wire C_drain_IO_L1_out_wrapper_279__ap_ready;
  wire C_drain_IO_L1_out_wrapper_279__ap_done;
  wire C_drain_IO_L1_out_wrapper_279__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_279__state;
  wire C_drain_IO_L1_out_wrapper_280__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_280__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_280__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_280__ap_start;
  wire C_drain_IO_L1_out_wrapper_280__ap_ready;
  wire C_drain_IO_L1_out_wrapper_280__ap_done;
  wire C_drain_IO_L1_out_wrapper_280__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_280__state;
  wire C_drain_IO_L1_out_wrapper_281__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_281__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_281__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_281__ap_start;
  wire C_drain_IO_L1_out_wrapper_281__ap_ready;
  wire C_drain_IO_L1_out_wrapper_281__ap_done;
  wire C_drain_IO_L1_out_wrapper_281__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_281__state;
  wire C_drain_IO_L1_out_wrapper_282__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_282__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_282__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_282__ap_start;
  wire C_drain_IO_L1_out_wrapper_282__ap_ready;
  wire C_drain_IO_L1_out_wrapper_282__ap_done;
  wire C_drain_IO_L1_out_wrapper_282__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_282__state;
  wire C_drain_IO_L1_out_wrapper_283__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_283__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_283__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_283__ap_start;
  wire C_drain_IO_L1_out_wrapper_283__ap_ready;
  wire C_drain_IO_L1_out_wrapper_283__ap_done;
  wire C_drain_IO_L1_out_wrapper_283__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_283__state;
  wire C_drain_IO_L1_out_wrapper_284__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_284__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_284__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_284__ap_start;
  wire C_drain_IO_L1_out_wrapper_284__ap_ready;
  wire C_drain_IO_L1_out_wrapper_284__ap_done;
  wire C_drain_IO_L1_out_wrapper_284__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_284__state;
  wire C_drain_IO_L1_out_wrapper_285__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_285__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_285__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_285__ap_start;
  wire C_drain_IO_L1_out_wrapper_285__ap_ready;
  wire C_drain_IO_L1_out_wrapper_285__ap_done;
  wire C_drain_IO_L1_out_wrapper_285__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_285__state;
  wire C_drain_IO_L1_out_wrapper_286__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_286__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_286__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_286__ap_start;
  wire C_drain_IO_L1_out_wrapper_286__ap_ready;
  wire C_drain_IO_L1_out_wrapper_286__ap_done;
  wire C_drain_IO_L1_out_wrapper_286__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_286__state;
  wire C_drain_IO_L1_out_wrapper_287__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_287__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_287__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_287__ap_start;
  wire C_drain_IO_L1_out_wrapper_287__ap_ready;
  wire C_drain_IO_L1_out_wrapper_287__ap_done;
  wire C_drain_IO_L1_out_wrapper_287__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_287__state;
  wire C_drain_IO_L1_out_wrapper_288__ap_start_global__q0;
  wire C_drain_IO_L1_out_wrapper_288__is_done__q0;
  wire C_drain_IO_L1_out_wrapper_288__ap_done_global__q0;
  wire C_drain_IO_L1_out_wrapper_288__ap_start;
  wire C_drain_IO_L1_out_wrapper_288__ap_ready;
  wire C_drain_IO_L1_out_wrapper_288__ap_done;
  wire C_drain_IO_L1_out_wrapper_288__ap_idle;
  reg [1:0] C_drain_IO_L1_out_wrapper_288__state;
  wire C_drain_IO_L2_out_0__ap_start_global__q0;
  wire C_drain_IO_L2_out_0__is_done__q0;
  wire C_drain_IO_L2_out_0__ap_done_global__q0;
  wire C_drain_IO_L2_out_0__ap_start;
  wire C_drain_IO_L2_out_0__ap_ready;
  wire C_drain_IO_L2_out_0__ap_done;
  wire C_drain_IO_L2_out_0__ap_idle;
  reg [1:0] C_drain_IO_L2_out_0__state;
  wire C_drain_IO_L2_out_1__ap_start_global__q0;
  wire C_drain_IO_L2_out_1__is_done__q0;
  wire C_drain_IO_L2_out_1__ap_done_global__q0;
  wire C_drain_IO_L2_out_1__ap_start;
  wire C_drain_IO_L2_out_1__ap_ready;
  wire C_drain_IO_L2_out_1__ap_done;
  wire C_drain_IO_L2_out_1__ap_idle;
  reg [1:0] C_drain_IO_L2_out_1__state;
  wire C_drain_IO_L2_out_2__ap_start_global__q0;
  wire C_drain_IO_L2_out_2__is_done__q0;
  wire C_drain_IO_L2_out_2__ap_done_global__q0;
  wire C_drain_IO_L2_out_2__ap_start;
  wire C_drain_IO_L2_out_2__ap_ready;
  wire C_drain_IO_L2_out_2__ap_done;
  wire C_drain_IO_L2_out_2__ap_idle;
  reg [1:0] C_drain_IO_L2_out_2__state;
  wire C_drain_IO_L2_out_3__ap_start_global__q0;
  wire C_drain_IO_L2_out_3__is_done__q0;
  wire C_drain_IO_L2_out_3__ap_done_global__q0;
  wire C_drain_IO_L2_out_3__ap_start;
  wire C_drain_IO_L2_out_3__ap_ready;
  wire C_drain_IO_L2_out_3__ap_done;
  wire C_drain_IO_L2_out_3__ap_idle;
  reg [1:0] C_drain_IO_L2_out_3__state;
  wire C_drain_IO_L2_out_4__ap_start_global__q0;
  wire C_drain_IO_L2_out_4__is_done__q0;
  wire C_drain_IO_L2_out_4__ap_done_global__q0;
  wire C_drain_IO_L2_out_4__ap_start;
  wire C_drain_IO_L2_out_4__ap_ready;
  wire C_drain_IO_L2_out_4__ap_done;
  wire C_drain_IO_L2_out_4__ap_idle;
  reg [1:0] C_drain_IO_L2_out_4__state;
  wire C_drain_IO_L2_out_5__ap_start_global__q0;
  wire C_drain_IO_L2_out_5__is_done__q0;
  wire C_drain_IO_L2_out_5__ap_done_global__q0;
  wire C_drain_IO_L2_out_5__ap_start;
  wire C_drain_IO_L2_out_5__ap_ready;
  wire C_drain_IO_L2_out_5__ap_done;
  wire C_drain_IO_L2_out_5__ap_idle;
  reg [1:0] C_drain_IO_L2_out_5__state;
  wire C_drain_IO_L2_out_6__ap_start_global__q0;
  wire C_drain_IO_L2_out_6__is_done__q0;
  wire C_drain_IO_L2_out_6__ap_done_global__q0;
  wire C_drain_IO_L2_out_6__ap_start;
  wire C_drain_IO_L2_out_6__ap_ready;
  wire C_drain_IO_L2_out_6__ap_done;
  wire C_drain_IO_L2_out_6__ap_idle;
  reg [1:0] C_drain_IO_L2_out_6__state;
  wire C_drain_IO_L2_out_7__ap_start_global__q0;
  wire C_drain_IO_L2_out_7__is_done__q0;
  wire C_drain_IO_L2_out_7__ap_done_global__q0;
  wire C_drain_IO_L2_out_7__ap_start;
  wire C_drain_IO_L2_out_7__ap_ready;
  wire C_drain_IO_L2_out_7__ap_done;
  wire C_drain_IO_L2_out_7__ap_idle;
  reg [1:0] C_drain_IO_L2_out_7__state;
  wire C_drain_IO_L2_out_8__ap_start_global__q0;
  wire C_drain_IO_L2_out_8__is_done__q0;
  wire C_drain_IO_L2_out_8__ap_done_global__q0;
  wire C_drain_IO_L2_out_8__ap_start;
  wire C_drain_IO_L2_out_8__ap_ready;
  wire C_drain_IO_L2_out_8__ap_done;
  wire C_drain_IO_L2_out_8__ap_idle;
  reg [1:0] C_drain_IO_L2_out_8__state;
  wire C_drain_IO_L2_out_9__ap_start_global__q0;
  wire C_drain_IO_L2_out_9__is_done__q0;
  wire C_drain_IO_L2_out_9__ap_done_global__q0;
  wire C_drain_IO_L2_out_9__ap_start;
  wire C_drain_IO_L2_out_9__ap_ready;
  wire C_drain_IO_L2_out_9__ap_done;
  wire C_drain_IO_L2_out_9__ap_idle;
  reg [1:0] C_drain_IO_L2_out_9__state;
  wire C_drain_IO_L2_out_10__ap_start_global__q0;
  wire C_drain_IO_L2_out_10__is_done__q0;
  wire C_drain_IO_L2_out_10__ap_done_global__q0;
  wire C_drain_IO_L2_out_10__ap_start;
  wire C_drain_IO_L2_out_10__ap_ready;
  wire C_drain_IO_L2_out_10__ap_done;
  wire C_drain_IO_L2_out_10__ap_idle;
  reg [1:0] C_drain_IO_L2_out_10__state;
  wire C_drain_IO_L2_out_11__ap_start_global__q0;
  wire C_drain_IO_L2_out_11__is_done__q0;
  wire C_drain_IO_L2_out_11__ap_done_global__q0;
  wire C_drain_IO_L2_out_11__ap_start;
  wire C_drain_IO_L2_out_11__ap_ready;
  wire C_drain_IO_L2_out_11__ap_done;
  wire C_drain_IO_L2_out_11__ap_idle;
  reg [1:0] C_drain_IO_L2_out_11__state;
  wire C_drain_IO_L2_out_12__ap_start_global__q0;
  wire C_drain_IO_L2_out_12__is_done__q0;
  wire C_drain_IO_L2_out_12__ap_done_global__q0;
  wire C_drain_IO_L2_out_12__ap_start;
  wire C_drain_IO_L2_out_12__ap_ready;
  wire C_drain_IO_L2_out_12__ap_done;
  wire C_drain_IO_L2_out_12__ap_idle;
  reg [1:0] C_drain_IO_L2_out_12__state;
  wire C_drain_IO_L2_out_13__ap_start_global__q0;
  wire C_drain_IO_L2_out_13__is_done__q0;
  wire C_drain_IO_L2_out_13__ap_done_global__q0;
  wire C_drain_IO_L2_out_13__ap_start;
  wire C_drain_IO_L2_out_13__ap_ready;
  wire C_drain_IO_L2_out_13__ap_done;
  wire C_drain_IO_L2_out_13__ap_idle;
  reg [1:0] C_drain_IO_L2_out_13__state;
  wire C_drain_IO_L2_out_14__ap_start_global__q0;
  wire C_drain_IO_L2_out_14__is_done__q0;
  wire C_drain_IO_L2_out_14__ap_done_global__q0;
  wire C_drain_IO_L2_out_14__ap_start;
  wire C_drain_IO_L2_out_14__ap_ready;
  wire C_drain_IO_L2_out_14__ap_done;
  wire C_drain_IO_L2_out_14__ap_idle;
  reg [1:0] C_drain_IO_L2_out_14__state;
  wire C_drain_IO_L2_out_15__ap_start_global__q0;
  wire C_drain_IO_L2_out_15__is_done__q0;
  wire C_drain_IO_L2_out_15__ap_done_global__q0;
  wire C_drain_IO_L2_out_15__ap_start;
  wire C_drain_IO_L2_out_15__ap_ready;
  wire C_drain_IO_L2_out_15__ap_done;
  wire C_drain_IO_L2_out_15__ap_idle;
  reg [1:0] C_drain_IO_L2_out_15__state;
  wire C_drain_IO_L2_out_boundary_0__ap_start_global__q0;
  wire C_drain_IO_L2_out_boundary_0__is_done__q0;
  wire C_drain_IO_L2_out_boundary_0__ap_done_global__q0;
  wire C_drain_IO_L2_out_boundary_0__ap_start;
  wire C_drain_IO_L2_out_boundary_0__ap_ready;
  wire C_drain_IO_L2_out_boundary_0__ap_done;
  wire C_drain_IO_L2_out_boundary_0__ap_idle;
  reg [1:0] C_drain_IO_L2_out_boundary_0__state;
  wire C_drain_IO_L3_out_0__ap_start_global__q0;
  wire C_drain_IO_L3_out_0__is_done__q0;
  wire C_drain_IO_L3_out_0__ap_done_global__q0;
  wire C_drain_IO_L3_out_0__ap_start;
  wire C_drain_IO_L3_out_0__ap_ready;
  wire C_drain_IO_L3_out_0__ap_done;
  wire C_drain_IO_L3_out_0__ap_idle;
  reg [1:0] C_drain_IO_L3_out_0__state;
  wire [63:0] C_drain_IO_L3_out_serialize_0___C__q0;
  wire C_drain_IO_L3_out_serialize_0__ap_start_global__q0;
  wire C_drain_IO_L3_out_serialize_0__is_done__q0;
  wire C_drain_IO_L3_out_serialize_0__ap_done_global__q0;
  wire C_drain_IO_L3_out_serialize_0__ap_start;
  wire C_drain_IO_L3_out_serialize_0__ap_ready;
  wire C_drain_IO_L3_out_serialize_0__ap_done;
  wire C_drain_IO_L3_out_serialize_0__ap_idle;
  reg [1:0] C_drain_IO_L3_out_serialize_0__state;
  wire PE_wrapper_0__ap_start_global__q0;
  wire PE_wrapper_0__is_done__q0;
  wire PE_wrapper_0__ap_done_global__q0;
  wire PE_wrapper_0__ap_start;
  wire PE_wrapper_0__ap_ready;
  wire PE_wrapper_0__ap_done;
  wire PE_wrapper_0__ap_idle;
  reg [1:0] PE_wrapper_0__state;
  wire PE_wrapper_1__ap_start_global__q0;
  wire PE_wrapper_1__is_done__q0;
  wire PE_wrapper_1__ap_done_global__q0;
  wire PE_wrapper_1__ap_start;
  wire PE_wrapper_1__ap_ready;
  wire PE_wrapper_1__ap_done;
  wire PE_wrapper_1__ap_idle;
  reg [1:0] PE_wrapper_1__state;
  wire PE_wrapper_2__ap_start_global__q0;
  wire PE_wrapper_2__is_done__q0;
  wire PE_wrapper_2__ap_done_global__q0;
  wire PE_wrapper_2__ap_start;
  wire PE_wrapper_2__ap_ready;
  wire PE_wrapper_2__ap_done;
  wire PE_wrapper_2__ap_idle;
  reg [1:0] PE_wrapper_2__state;
  wire PE_wrapper_3__ap_start_global__q0;
  wire PE_wrapper_3__is_done__q0;
  wire PE_wrapper_3__ap_done_global__q0;
  wire PE_wrapper_3__ap_start;
  wire PE_wrapper_3__ap_ready;
  wire PE_wrapper_3__ap_done;
  wire PE_wrapper_3__ap_idle;
  reg [1:0] PE_wrapper_3__state;
  wire PE_wrapper_4__ap_start_global__q0;
  wire PE_wrapper_4__is_done__q0;
  wire PE_wrapper_4__ap_done_global__q0;
  wire PE_wrapper_4__ap_start;
  wire PE_wrapper_4__ap_ready;
  wire PE_wrapper_4__ap_done;
  wire PE_wrapper_4__ap_idle;
  reg [1:0] PE_wrapper_4__state;
  wire PE_wrapper_5__ap_start_global__q0;
  wire PE_wrapper_5__is_done__q0;
  wire PE_wrapper_5__ap_done_global__q0;
  wire PE_wrapper_5__ap_start;
  wire PE_wrapper_5__ap_ready;
  wire PE_wrapper_5__ap_done;
  wire PE_wrapper_5__ap_idle;
  reg [1:0] PE_wrapper_5__state;
  wire PE_wrapper_6__ap_start_global__q0;
  wire PE_wrapper_6__is_done__q0;
  wire PE_wrapper_6__ap_done_global__q0;
  wire PE_wrapper_6__ap_start;
  wire PE_wrapper_6__ap_ready;
  wire PE_wrapper_6__ap_done;
  wire PE_wrapper_6__ap_idle;
  reg [1:0] PE_wrapper_6__state;
  wire PE_wrapper_7__ap_start_global__q0;
  wire PE_wrapper_7__is_done__q0;
  wire PE_wrapper_7__ap_done_global__q0;
  wire PE_wrapper_7__ap_start;
  wire PE_wrapper_7__ap_ready;
  wire PE_wrapper_7__ap_done;
  wire PE_wrapper_7__ap_idle;
  reg [1:0] PE_wrapper_7__state;
  wire PE_wrapper_8__ap_start_global__q0;
  wire PE_wrapper_8__is_done__q0;
  wire PE_wrapper_8__ap_done_global__q0;
  wire PE_wrapper_8__ap_start;
  wire PE_wrapper_8__ap_ready;
  wire PE_wrapper_8__ap_done;
  wire PE_wrapper_8__ap_idle;
  reg [1:0] PE_wrapper_8__state;
  wire PE_wrapper_9__ap_start_global__q0;
  wire PE_wrapper_9__is_done__q0;
  wire PE_wrapper_9__ap_done_global__q0;
  wire PE_wrapper_9__ap_start;
  wire PE_wrapper_9__ap_ready;
  wire PE_wrapper_9__ap_done;
  wire PE_wrapper_9__ap_idle;
  reg [1:0] PE_wrapper_9__state;
  wire PE_wrapper_10__ap_start_global__q0;
  wire PE_wrapper_10__is_done__q0;
  wire PE_wrapper_10__ap_done_global__q0;
  wire PE_wrapper_10__ap_start;
  wire PE_wrapper_10__ap_ready;
  wire PE_wrapper_10__ap_done;
  wire PE_wrapper_10__ap_idle;
  reg [1:0] PE_wrapper_10__state;
  wire PE_wrapper_11__ap_start_global__q0;
  wire PE_wrapper_11__is_done__q0;
  wire PE_wrapper_11__ap_done_global__q0;
  wire PE_wrapper_11__ap_start;
  wire PE_wrapper_11__ap_ready;
  wire PE_wrapper_11__ap_done;
  wire PE_wrapper_11__ap_idle;
  reg [1:0] PE_wrapper_11__state;
  wire PE_wrapper_12__ap_start_global__q0;
  wire PE_wrapper_12__is_done__q0;
  wire PE_wrapper_12__ap_done_global__q0;
  wire PE_wrapper_12__ap_start;
  wire PE_wrapper_12__ap_ready;
  wire PE_wrapper_12__ap_done;
  wire PE_wrapper_12__ap_idle;
  reg [1:0] PE_wrapper_12__state;
  wire PE_wrapper_13__ap_start_global__q0;
  wire PE_wrapper_13__is_done__q0;
  wire PE_wrapper_13__ap_done_global__q0;
  wire PE_wrapper_13__ap_start;
  wire PE_wrapper_13__ap_ready;
  wire PE_wrapper_13__ap_done;
  wire PE_wrapper_13__ap_idle;
  reg [1:0] PE_wrapper_13__state;
  wire PE_wrapper_14__ap_start_global__q0;
  wire PE_wrapper_14__is_done__q0;
  wire PE_wrapper_14__ap_done_global__q0;
  wire PE_wrapper_14__ap_start;
  wire PE_wrapper_14__ap_ready;
  wire PE_wrapper_14__ap_done;
  wire PE_wrapper_14__ap_idle;
  reg [1:0] PE_wrapper_14__state;
  wire PE_wrapper_15__ap_start_global__q0;
  wire PE_wrapper_15__is_done__q0;
  wire PE_wrapper_15__ap_done_global__q0;
  wire PE_wrapper_15__ap_start;
  wire PE_wrapper_15__ap_ready;
  wire PE_wrapper_15__ap_done;
  wire PE_wrapper_15__ap_idle;
  reg [1:0] PE_wrapper_15__state;
  wire PE_wrapper_16__ap_start_global__q0;
  wire PE_wrapper_16__is_done__q0;
  wire PE_wrapper_16__ap_done_global__q0;
  wire PE_wrapper_16__ap_start;
  wire PE_wrapper_16__ap_ready;
  wire PE_wrapper_16__ap_done;
  wire PE_wrapper_16__ap_idle;
  reg [1:0] PE_wrapper_16__state;
  wire PE_wrapper_17__ap_start_global__q0;
  wire PE_wrapper_17__is_done__q0;
  wire PE_wrapper_17__ap_done_global__q0;
  wire PE_wrapper_17__ap_start;
  wire PE_wrapper_17__ap_ready;
  wire PE_wrapper_17__ap_done;
  wire PE_wrapper_17__ap_idle;
  reg [1:0] PE_wrapper_17__state;
  wire PE_wrapper_18__ap_start_global__q0;
  wire PE_wrapper_18__is_done__q0;
  wire PE_wrapper_18__ap_done_global__q0;
  wire PE_wrapper_18__ap_start;
  wire PE_wrapper_18__ap_ready;
  wire PE_wrapper_18__ap_done;
  wire PE_wrapper_18__ap_idle;
  reg [1:0] PE_wrapper_18__state;
  wire PE_wrapper_19__ap_start_global__q0;
  wire PE_wrapper_19__is_done__q0;
  wire PE_wrapper_19__ap_done_global__q0;
  wire PE_wrapper_19__ap_start;
  wire PE_wrapper_19__ap_ready;
  wire PE_wrapper_19__ap_done;
  wire PE_wrapper_19__ap_idle;
  reg [1:0] PE_wrapper_19__state;
  wire PE_wrapper_20__ap_start_global__q0;
  wire PE_wrapper_20__is_done__q0;
  wire PE_wrapper_20__ap_done_global__q0;
  wire PE_wrapper_20__ap_start;
  wire PE_wrapper_20__ap_ready;
  wire PE_wrapper_20__ap_done;
  wire PE_wrapper_20__ap_idle;
  reg [1:0] PE_wrapper_20__state;
  wire PE_wrapper_21__ap_start_global__q0;
  wire PE_wrapper_21__is_done__q0;
  wire PE_wrapper_21__ap_done_global__q0;
  wire PE_wrapper_21__ap_start;
  wire PE_wrapper_21__ap_ready;
  wire PE_wrapper_21__ap_done;
  wire PE_wrapper_21__ap_idle;
  reg [1:0] PE_wrapper_21__state;
  wire PE_wrapper_22__ap_start_global__q0;
  wire PE_wrapper_22__is_done__q0;
  wire PE_wrapper_22__ap_done_global__q0;
  wire PE_wrapper_22__ap_start;
  wire PE_wrapper_22__ap_ready;
  wire PE_wrapper_22__ap_done;
  wire PE_wrapper_22__ap_idle;
  reg [1:0] PE_wrapper_22__state;
  wire PE_wrapper_23__ap_start_global__q0;
  wire PE_wrapper_23__is_done__q0;
  wire PE_wrapper_23__ap_done_global__q0;
  wire PE_wrapper_23__ap_start;
  wire PE_wrapper_23__ap_ready;
  wire PE_wrapper_23__ap_done;
  wire PE_wrapper_23__ap_idle;
  reg [1:0] PE_wrapper_23__state;
  wire PE_wrapper_24__ap_start_global__q0;
  wire PE_wrapper_24__is_done__q0;
  wire PE_wrapper_24__ap_done_global__q0;
  wire PE_wrapper_24__ap_start;
  wire PE_wrapper_24__ap_ready;
  wire PE_wrapper_24__ap_done;
  wire PE_wrapper_24__ap_idle;
  reg [1:0] PE_wrapper_24__state;
  wire PE_wrapper_25__ap_start_global__q0;
  wire PE_wrapper_25__is_done__q0;
  wire PE_wrapper_25__ap_done_global__q0;
  wire PE_wrapper_25__ap_start;
  wire PE_wrapper_25__ap_ready;
  wire PE_wrapper_25__ap_done;
  wire PE_wrapper_25__ap_idle;
  reg [1:0] PE_wrapper_25__state;
  wire PE_wrapper_26__ap_start_global__q0;
  wire PE_wrapper_26__is_done__q0;
  wire PE_wrapper_26__ap_done_global__q0;
  wire PE_wrapper_26__ap_start;
  wire PE_wrapper_26__ap_ready;
  wire PE_wrapper_26__ap_done;
  wire PE_wrapper_26__ap_idle;
  reg [1:0] PE_wrapper_26__state;
  wire PE_wrapper_27__ap_start_global__q0;
  wire PE_wrapper_27__is_done__q0;
  wire PE_wrapper_27__ap_done_global__q0;
  wire PE_wrapper_27__ap_start;
  wire PE_wrapper_27__ap_ready;
  wire PE_wrapper_27__ap_done;
  wire PE_wrapper_27__ap_idle;
  reg [1:0] PE_wrapper_27__state;
  wire PE_wrapper_28__ap_start_global__q0;
  wire PE_wrapper_28__is_done__q0;
  wire PE_wrapper_28__ap_done_global__q0;
  wire PE_wrapper_28__ap_start;
  wire PE_wrapper_28__ap_ready;
  wire PE_wrapper_28__ap_done;
  wire PE_wrapper_28__ap_idle;
  reg [1:0] PE_wrapper_28__state;
  wire PE_wrapper_29__ap_start_global__q0;
  wire PE_wrapper_29__is_done__q0;
  wire PE_wrapper_29__ap_done_global__q0;
  wire PE_wrapper_29__ap_start;
  wire PE_wrapper_29__ap_ready;
  wire PE_wrapper_29__ap_done;
  wire PE_wrapper_29__ap_idle;
  reg [1:0] PE_wrapper_29__state;
  wire PE_wrapper_30__ap_start_global__q0;
  wire PE_wrapper_30__is_done__q0;
  wire PE_wrapper_30__ap_done_global__q0;
  wire PE_wrapper_30__ap_start;
  wire PE_wrapper_30__ap_ready;
  wire PE_wrapper_30__ap_done;
  wire PE_wrapper_30__ap_idle;
  reg [1:0] PE_wrapper_30__state;
  wire PE_wrapper_31__ap_start_global__q0;
  wire PE_wrapper_31__is_done__q0;
  wire PE_wrapper_31__ap_done_global__q0;
  wire PE_wrapper_31__ap_start;
  wire PE_wrapper_31__ap_ready;
  wire PE_wrapper_31__ap_done;
  wire PE_wrapper_31__ap_idle;
  reg [1:0] PE_wrapper_31__state;
  wire PE_wrapper_32__ap_start_global__q0;
  wire PE_wrapper_32__is_done__q0;
  wire PE_wrapper_32__ap_done_global__q0;
  wire PE_wrapper_32__ap_start;
  wire PE_wrapper_32__ap_ready;
  wire PE_wrapper_32__ap_done;
  wire PE_wrapper_32__ap_idle;
  reg [1:0] PE_wrapper_32__state;
  wire PE_wrapper_33__ap_start_global__q0;
  wire PE_wrapper_33__is_done__q0;
  wire PE_wrapper_33__ap_done_global__q0;
  wire PE_wrapper_33__ap_start;
  wire PE_wrapper_33__ap_ready;
  wire PE_wrapper_33__ap_done;
  wire PE_wrapper_33__ap_idle;
  reg [1:0] PE_wrapper_33__state;
  wire PE_wrapper_34__ap_start_global__q0;
  wire PE_wrapper_34__is_done__q0;
  wire PE_wrapper_34__ap_done_global__q0;
  wire PE_wrapper_34__ap_start;
  wire PE_wrapper_34__ap_ready;
  wire PE_wrapper_34__ap_done;
  wire PE_wrapper_34__ap_idle;
  reg [1:0] PE_wrapper_34__state;
  wire PE_wrapper_35__ap_start_global__q0;
  wire PE_wrapper_35__is_done__q0;
  wire PE_wrapper_35__ap_done_global__q0;
  wire PE_wrapper_35__ap_start;
  wire PE_wrapper_35__ap_ready;
  wire PE_wrapper_35__ap_done;
  wire PE_wrapper_35__ap_idle;
  reg [1:0] PE_wrapper_35__state;
  wire PE_wrapper_36__ap_start_global__q0;
  wire PE_wrapper_36__is_done__q0;
  wire PE_wrapper_36__ap_done_global__q0;
  wire PE_wrapper_36__ap_start;
  wire PE_wrapper_36__ap_ready;
  wire PE_wrapper_36__ap_done;
  wire PE_wrapper_36__ap_idle;
  reg [1:0] PE_wrapper_36__state;
  wire PE_wrapper_37__ap_start_global__q0;
  wire PE_wrapper_37__is_done__q0;
  wire PE_wrapper_37__ap_done_global__q0;
  wire PE_wrapper_37__ap_start;
  wire PE_wrapper_37__ap_ready;
  wire PE_wrapper_37__ap_done;
  wire PE_wrapper_37__ap_idle;
  reg [1:0] PE_wrapper_37__state;
  wire PE_wrapper_38__ap_start_global__q0;
  wire PE_wrapper_38__is_done__q0;
  wire PE_wrapper_38__ap_done_global__q0;
  wire PE_wrapper_38__ap_start;
  wire PE_wrapper_38__ap_ready;
  wire PE_wrapper_38__ap_done;
  wire PE_wrapper_38__ap_idle;
  reg [1:0] PE_wrapper_38__state;
  wire PE_wrapper_39__ap_start_global__q0;
  wire PE_wrapper_39__is_done__q0;
  wire PE_wrapper_39__ap_done_global__q0;
  wire PE_wrapper_39__ap_start;
  wire PE_wrapper_39__ap_ready;
  wire PE_wrapper_39__ap_done;
  wire PE_wrapper_39__ap_idle;
  reg [1:0] PE_wrapper_39__state;
  wire PE_wrapper_40__ap_start_global__q0;
  wire PE_wrapper_40__is_done__q0;
  wire PE_wrapper_40__ap_done_global__q0;
  wire PE_wrapper_40__ap_start;
  wire PE_wrapper_40__ap_ready;
  wire PE_wrapper_40__ap_done;
  wire PE_wrapper_40__ap_idle;
  reg [1:0] PE_wrapper_40__state;
  wire PE_wrapper_41__ap_start_global__q0;
  wire PE_wrapper_41__is_done__q0;
  wire PE_wrapper_41__ap_done_global__q0;
  wire PE_wrapper_41__ap_start;
  wire PE_wrapper_41__ap_ready;
  wire PE_wrapper_41__ap_done;
  wire PE_wrapper_41__ap_idle;
  reg [1:0] PE_wrapper_41__state;
  wire PE_wrapper_42__ap_start_global__q0;
  wire PE_wrapper_42__is_done__q0;
  wire PE_wrapper_42__ap_done_global__q0;
  wire PE_wrapper_42__ap_start;
  wire PE_wrapper_42__ap_ready;
  wire PE_wrapper_42__ap_done;
  wire PE_wrapper_42__ap_idle;
  reg [1:0] PE_wrapper_42__state;
  wire PE_wrapper_43__ap_start_global__q0;
  wire PE_wrapper_43__is_done__q0;
  wire PE_wrapper_43__ap_done_global__q0;
  wire PE_wrapper_43__ap_start;
  wire PE_wrapper_43__ap_ready;
  wire PE_wrapper_43__ap_done;
  wire PE_wrapper_43__ap_idle;
  reg [1:0] PE_wrapper_43__state;
  wire PE_wrapper_44__ap_start_global__q0;
  wire PE_wrapper_44__is_done__q0;
  wire PE_wrapper_44__ap_done_global__q0;
  wire PE_wrapper_44__ap_start;
  wire PE_wrapper_44__ap_ready;
  wire PE_wrapper_44__ap_done;
  wire PE_wrapper_44__ap_idle;
  reg [1:0] PE_wrapper_44__state;
  wire PE_wrapper_45__ap_start_global__q0;
  wire PE_wrapper_45__is_done__q0;
  wire PE_wrapper_45__ap_done_global__q0;
  wire PE_wrapper_45__ap_start;
  wire PE_wrapper_45__ap_ready;
  wire PE_wrapper_45__ap_done;
  wire PE_wrapper_45__ap_idle;
  reg [1:0] PE_wrapper_45__state;
  wire PE_wrapper_46__ap_start_global__q0;
  wire PE_wrapper_46__is_done__q0;
  wire PE_wrapper_46__ap_done_global__q0;
  wire PE_wrapper_46__ap_start;
  wire PE_wrapper_46__ap_ready;
  wire PE_wrapper_46__ap_done;
  wire PE_wrapper_46__ap_idle;
  reg [1:0] PE_wrapper_46__state;
  wire PE_wrapper_47__ap_start_global__q0;
  wire PE_wrapper_47__is_done__q0;
  wire PE_wrapper_47__ap_done_global__q0;
  wire PE_wrapper_47__ap_start;
  wire PE_wrapper_47__ap_ready;
  wire PE_wrapper_47__ap_done;
  wire PE_wrapper_47__ap_idle;
  reg [1:0] PE_wrapper_47__state;
  wire PE_wrapper_48__ap_start_global__q0;
  wire PE_wrapper_48__is_done__q0;
  wire PE_wrapper_48__ap_done_global__q0;
  wire PE_wrapper_48__ap_start;
  wire PE_wrapper_48__ap_ready;
  wire PE_wrapper_48__ap_done;
  wire PE_wrapper_48__ap_idle;
  reg [1:0] PE_wrapper_48__state;
  wire PE_wrapper_49__ap_start_global__q0;
  wire PE_wrapper_49__is_done__q0;
  wire PE_wrapper_49__ap_done_global__q0;
  wire PE_wrapper_49__ap_start;
  wire PE_wrapper_49__ap_ready;
  wire PE_wrapper_49__ap_done;
  wire PE_wrapper_49__ap_idle;
  reg [1:0] PE_wrapper_49__state;
  wire PE_wrapper_50__ap_start_global__q0;
  wire PE_wrapper_50__is_done__q0;
  wire PE_wrapper_50__ap_done_global__q0;
  wire PE_wrapper_50__ap_start;
  wire PE_wrapper_50__ap_ready;
  wire PE_wrapper_50__ap_done;
  wire PE_wrapper_50__ap_idle;
  reg [1:0] PE_wrapper_50__state;
  wire PE_wrapper_51__ap_start_global__q0;
  wire PE_wrapper_51__is_done__q0;
  wire PE_wrapper_51__ap_done_global__q0;
  wire PE_wrapper_51__ap_start;
  wire PE_wrapper_51__ap_ready;
  wire PE_wrapper_51__ap_done;
  wire PE_wrapper_51__ap_idle;
  reg [1:0] PE_wrapper_51__state;
  wire PE_wrapper_52__ap_start_global__q0;
  wire PE_wrapper_52__is_done__q0;
  wire PE_wrapper_52__ap_done_global__q0;
  wire PE_wrapper_52__ap_start;
  wire PE_wrapper_52__ap_ready;
  wire PE_wrapper_52__ap_done;
  wire PE_wrapper_52__ap_idle;
  reg [1:0] PE_wrapper_52__state;
  wire PE_wrapper_53__ap_start_global__q0;
  wire PE_wrapper_53__is_done__q0;
  wire PE_wrapper_53__ap_done_global__q0;
  wire PE_wrapper_53__ap_start;
  wire PE_wrapper_53__ap_ready;
  wire PE_wrapper_53__ap_done;
  wire PE_wrapper_53__ap_idle;
  reg [1:0] PE_wrapper_53__state;
  wire PE_wrapper_54__ap_start_global__q0;
  wire PE_wrapper_54__is_done__q0;
  wire PE_wrapper_54__ap_done_global__q0;
  wire PE_wrapper_54__ap_start;
  wire PE_wrapper_54__ap_ready;
  wire PE_wrapper_54__ap_done;
  wire PE_wrapper_54__ap_idle;
  reg [1:0] PE_wrapper_54__state;
  wire PE_wrapper_55__ap_start_global__q0;
  wire PE_wrapper_55__is_done__q0;
  wire PE_wrapper_55__ap_done_global__q0;
  wire PE_wrapper_55__ap_start;
  wire PE_wrapper_55__ap_ready;
  wire PE_wrapper_55__ap_done;
  wire PE_wrapper_55__ap_idle;
  reg [1:0] PE_wrapper_55__state;
  wire PE_wrapper_56__ap_start_global__q0;
  wire PE_wrapper_56__is_done__q0;
  wire PE_wrapper_56__ap_done_global__q0;
  wire PE_wrapper_56__ap_start;
  wire PE_wrapper_56__ap_ready;
  wire PE_wrapper_56__ap_done;
  wire PE_wrapper_56__ap_idle;
  reg [1:0] PE_wrapper_56__state;
  wire PE_wrapper_57__ap_start_global__q0;
  wire PE_wrapper_57__is_done__q0;
  wire PE_wrapper_57__ap_done_global__q0;
  wire PE_wrapper_57__ap_start;
  wire PE_wrapper_57__ap_ready;
  wire PE_wrapper_57__ap_done;
  wire PE_wrapper_57__ap_idle;
  reg [1:0] PE_wrapper_57__state;
  wire PE_wrapper_58__ap_start_global__q0;
  wire PE_wrapper_58__is_done__q0;
  wire PE_wrapper_58__ap_done_global__q0;
  wire PE_wrapper_58__ap_start;
  wire PE_wrapper_58__ap_ready;
  wire PE_wrapper_58__ap_done;
  wire PE_wrapper_58__ap_idle;
  reg [1:0] PE_wrapper_58__state;
  wire PE_wrapper_59__ap_start_global__q0;
  wire PE_wrapper_59__is_done__q0;
  wire PE_wrapper_59__ap_done_global__q0;
  wire PE_wrapper_59__ap_start;
  wire PE_wrapper_59__ap_ready;
  wire PE_wrapper_59__ap_done;
  wire PE_wrapper_59__ap_idle;
  reg [1:0] PE_wrapper_59__state;
  wire PE_wrapper_60__ap_start_global__q0;
  wire PE_wrapper_60__is_done__q0;
  wire PE_wrapper_60__ap_done_global__q0;
  wire PE_wrapper_60__ap_start;
  wire PE_wrapper_60__ap_ready;
  wire PE_wrapper_60__ap_done;
  wire PE_wrapper_60__ap_idle;
  reg [1:0] PE_wrapper_60__state;
  wire PE_wrapper_61__ap_start_global__q0;
  wire PE_wrapper_61__is_done__q0;
  wire PE_wrapper_61__ap_done_global__q0;
  wire PE_wrapper_61__ap_start;
  wire PE_wrapper_61__ap_ready;
  wire PE_wrapper_61__ap_done;
  wire PE_wrapper_61__ap_idle;
  reg [1:0] PE_wrapper_61__state;
  wire PE_wrapper_62__ap_start_global__q0;
  wire PE_wrapper_62__is_done__q0;
  wire PE_wrapper_62__ap_done_global__q0;
  wire PE_wrapper_62__ap_start;
  wire PE_wrapper_62__ap_ready;
  wire PE_wrapper_62__ap_done;
  wire PE_wrapper_62__ap_idle;
  reg [1:0] PE_wrapper_62__state;
  wire PE_wrapper_63__ap_start_global__q0;
  wire PE_wrapper_63__is_done__q0;
  wire PE_wrapper_63__ap_done_global__q0;
  wire PE_wrapper_63__ap_start;
  wire PE_wrapper_63__ap_ready;
  wire PE_wrapper_63__ap_done;
  wire PE_wrapper_63__ap_idle;
  reg [1:0] PE_wrapper_63__state;
  wire PE_wrapper_64__ap_start_global__q0;
  wire PE_wrapper_64__is_done__q0;
  wire PE_wrapper_64__ap_done_global__q0;
  wire PE_wrapper_64__ap_start;
  wire PE_wrapper_64__ap_ready;
  wire PE_wrapper_64__ap_done;
  wire PE_wrapper_64__ap_idle;
  reg [1:0] PE_wrapper_64__state;
  wire PE_wrapper_65__ap_start_global__q0;
  wire PE_wrapper_65__is_done__q0;
  wire PE_wrapper_65__ap_done_global__q0;
  wire PE_wrapper_65__ap_start;
  wire PE_wrapper_65__ap_ready;
  wire PE_wrapper_65__ap_done;
  wire PE_wrapper_65__ap_idle;
  reg [1:0] PE_wrapper_65__state;
  wire PE_wrapper_66__ap_start_global__q0;
  wire PE_wrapper_66__is_done__q0;
  wire PE_wrapper_66__ap_done_global__q0;
  wire PE_wrapper_66__ap_start;
  wire PE_wrapper_66__ap_ready;
  wire PE_wrapper_66__ap_done;
  wire PE_wrapper_66__ap_idle;
  reg [1:0] PE_wrapper_66__state;
  wire PE_wrapper_67__ap_start_global__q0;
  wire PE_wrapper_67__is_done__q0;
  wire PE_wrapper_67__ap_done_global__q0;
  wire PE_wrapper_67__ap_start;
  wire PE_wrapper_67__ap_ready;
  wire PE_wrapper_67__ap_done;
  wire PE_wrapper_67__ap_idle;
  reg [1:0] PE_wrapper_67__state;
  wire PE_wrapper_68__ap_start_global__q0;
  wire PE_wrapper_68__is_done__q0;
  wire PE_wrapper_68__ap_done_global__q0;
  wire PE_wrapper_68__ap_start;
  wire PE_wrapper_68__ap_ready;
  wire PE_wrapper_68__ap_done;
  wire PE_wrapper_68__ap_idle;
  reg [1:0] PE_wrapper_68__state;
  wire PE_wrapper_69__ap_start_global__q0;
  wire PE_wrapper_69__is_done__q0;
  wire PE_wrapper_69__ap_done_global__q0;
  wire PE_wrapper_69__ap_start;
  wire PE_wrapper_69__ap_ready;
  wire PE_wrapper_69__ap_done;
  wire PE_wrapper_69__ap_idle;
  reg [1:0] PE_wrapper_69__state;
  wire PE_wrapper_70__ap_start_global__q0;
  wire PE_wrapper_70__is_done__q0;
  wire PE_wrapper_70__ap_done_global__q0;
  wire PE_wrapper_70__ap_start;
  wire PE_wrapper_70__ap_ready;
  wire PE_wrapper_70__ap_done;
  wire PE_wrapper_70__ap_idle;
  reg [1:0] PE_wrapper_70__state;
  wire PE_wrapper_71__ap_start_global__q0;
  wire PE_wrapper_71__is_done__q0;
  wire PE_wrapper_71__ap_done_global__q0;
  wire PE_wrapper_71__ap_start;
  wire PE_wrapper_71__ap_ready;
  wire PE_wrapper_71__ap_done;
  wire PE_wrapper_71__ap_idle;
  reg [1:0] PE_wrapper_71__state;
  wire PE_wrapper_72__ap_start_global__q0;
  wire PE_wrapper_72__is_done__q0;
  wire PE_wrapper_72__ap_done_global__q0;
  wire PE_wrapper_72__ap_start;
  wire PE_wrapper_72__ap_ready;
  wire PE_wrapper_72__ap_done;
  wire PE_wrapper_72__ap_idle;
  reg [1:0] PE_wrapper_72__state;
  wire PE_wrapper_73__ap_start_global__q0;
  wire PE_wrapper_73__is_done__q0;
  wire PE_wrapper_73__ap_done_global__q0;
  wire PE_wrapper_73__ap_start;
  wire PE_wrapper_73__ap_ready;
  wire PE_wrapper_73__ap_done;
  wire PE_wrapper_73__ap_idle;
  reg [1:0] PE_wrapper_73__state;
  wire PE_wrapper_74__ap_start_global__q0;
  wire PE_wrapper_74__is_done__q0;
  wire PE_wrapper_74__ap_done_global__q0;
  wire PE_wrapper_74__ap_start;
  wire PE_wrapper_74__ap_ready;
  wire PE_wrapper_74__ap_done;
  wire PE_wrapper_74__ap_idle;
  reg [1:0] PE_wrapper_74__state;
  wire PE_wrapper_75__ap_start_global__q0;
  wire PE_wrapper_75__is_done__q0;
  wire PE_wrapper_75__ap_done_global__q0;
  wire PE_wrapper_75__ap_start;
  wire PE_wrapper_75__ap_ready;
  wire PE_wrapper_75__ap_done;
  wire PE_wrapper_75__ap_idle;
  reg [1:0] PE_wrapper_75__state;
  wire PE_wrapper_76__ap_start_global__q0;
  wire PE_wrapper_76__is_done__q0;
  wire PE_wrapper_76__ap_done_global__q0;
  wire PE_wrapper_76__ap_start;
  wire PE_wrapper_76__ap_ready;
  wire PE_wrapper_76__ap_done;
  wire PE_wrapper_76__ap_idle;
  reg [1:0] PE_wrapper_76__state;
  wire PE_wrapper_77__ap_start_global__q0;
  wire PE_wrapper_77__is_done__q0;
  wire PE_wrapper_77__ap_done_global__q0;
  wire PE_wrapper_77__ap_start;
  wire PE_wrapper_77__ap_ready;
  wire PE_wrapper_77__ap_done;
  wire PE_wrapper_77__ap_idle;
  reg [1:0] PE_wrapper_77__state;
  wire PE_wrapper_78__ap_start_global__q0;
  wire PE_wrapper_78__is_done__q0;
  wire PE_wrapper_78__ap_done_global__q0;
  wire PE_wrapper_78__ap_start;
  wire PE_wrapper_78__ap_ready;
  wire PE_wrapper_78__ap_done;
  wire PE_wrapper_78__ap_idle;
  reg [1:0] PE_wrapper_78__state;
  wire PE_wrapper_79__ap_start_global__q0;
  wire PE_wrapper_79__is_done__q0;
  wire PE_wrapper_79__ap_done_global__q0;
  wire PE_wrapper_79__ap_start;
  wire PE_wrapper_79__ap_ready;
  wire PE_wrapper_79__ap_done;
  wire PE_wrapper_79__ap_idle;
  reg [1:0] PE_wrapper_79__state;
  wire PE_wrapper_80__ap_start_global__q0;
  wire PE_wrapper_80__is_done__q0;
  wire PE_wrapper_80__ap_done_global__q0;
  wire PE_wrapper_80__ap_start;
  wire PE_wrapper_80__ap_ready;
  wire PE_wrapper_80__ap_done;
  wire PE_wrapper_80__ap_idle;
  reg [1:0] PE_wrapper_80__state;
  wire PE_wrapper_81__ap_start_global__q0;
  wire PE_wrapper_81__is_done__q0;
  wire PE_wrapper_81__ap_done_global__q0;
  wire PE_wrapper_81__ap_start;
  wire PE_wrapper_81__ap_ready;
  wire PE_wrapper_81__ap_done;
  wire PE_wrapper_81__ap_idle;
  reg [1:0] PE_wrapper_81__state;
  wire PE_wrapper_82__ap_start_global__q0;
  wire PE_wrapper_82__is_done__q0;
  wire PE_wrapper_82__ap_done_global__q0;
  wire PE_wrapper_82__ap_start;
  wire PE_wrapper_82__ap_ready;
  wire PE_wrapper_82__ap_done;
  wire PE_wrapper_82__ap_idle;
  reg [1:0] PE_wrapper_82__state;
  wire PE_wrapper_83__ap_start_global__q0;
  wire PE_wrapper_83__is_done__q0;
  wire PE_wrapper_83__ap_done_global__q0;
  wire PE_wrapper_83__ap_start;
  wire PE_wrapper_83__ap_ready;
  wire PE_wrapper_83__ap_done;
  wire PE_wrapper_83__ap_idle;
  reg [1:0] PE_wrapper_83__state;
  wire PE_wrapper_84__ap_start_global__q0;
  wire PE_wrapper_84__is_done__q0;
  wire PE_wrapper_84__ap_done_global__q0;
  wire PE_wrapper_84__ap_start;
  wire PE_wrapper_84__ap_ready;
  wire PE_wrapper_84__ap_done;
  wire PE_wrapper_84__ap_idle;
  reg [1:0] PE_wrapper_84__state;
  wire PE_wrapper_85__ap_start_global__q0;
  wire PE_wrapper_85__is_done__q0;
  wire PE_wrapper_85__ap_done_global__q0;
  wire PE_wrapper_85__ap_start;
  wire PE_wrapper_85__ap_ready;
  wire PE_wrapper_85__ap_done;
  wire PE_wrapper_85__ap_idle;
  reg [1:0] PE_wrapper_85__state;
  wire PE_wrapper_86__ap_start_global__q0;
  wire PE_wrapper_86__is_done__q0;
  wire PE_wrapper_86__ap_done_global__q0;
  wire PE_wrapper_86__ap_start;
  wire PE_wrapper_86__ap_ready;
  wire PE_wrapper_86__ap_done;
  wire PE_wrapper_86__ap_idle;
  reg [1:0] PE_wrapper_86__state;
  wire PE_wrapper_87__ap_start_global__q0;
  wire PE_wrapper_87__is_done__q0;
  wire PE_wrapper_87__ap_done_global__q0;
  wire PE_wrapper_87__ap_start;
  wire PE_wrapper_87__ap_ready;
  wire PE_wrapper_87__ap_done;
  wire PE_wrapper_87__ap_idle;
  reg [1:0] PE_wrapper_87__state;
  wire PE_wrapper_88__ap_start_global__q0;
  wire PE_wrapper_88__is_done__q0;
  wire PE_wrapper_88__ap_done_global__q0;
  wire PE_wrapper_88__ap_start;
  wire PE_wrapper_88__ap_ready;
  wire PE_wrapper_88__ap_done;
  wire PE_wrapper_88__ap_idle;
  reg [1:0] PE_wrapper_88__state;
  wire PE_wrapper_89__ap_start_global__q0;
  wire PE_wrapper_89__is_done__q0;
  wire PE_wrapper_89__ap_done_global__q0;
  wire PE_wrapper_89__ap_start;
  wire PE_wrapper_89__ap_ready;
  wire PE_wrapper_89__ap_done;
  wire PE_wrapper_89__ap_idle;
  reg [1:0] PE_wrapper_89__state;
  wire PE_wrapper_90__ap_start_global__q0;
  wire PE_wrapper_90__is_done__q0;
  wire PE_wrapper_90__ap_done_global__q0;
  wire PE_wrapper_90__ap_start;
  wire PE_wrapper_90__ap_ready;
  wire PE_wrapper_90__ap_done;
  wire PE_wrapper_90__ap_idle;
  reg [1:0] PE_wrapper_90__state;
  wire PE_wrapper_91__ap_start_global__q0;
  wire PE_wrapper_91__is_done__q0;
  wire PE_wrapper_91__ap_done_global__q0;
  wire PE_wrapper_91__ap_start;
  wire PE_wrapper_91__ap_ready;
  wire PE_wrapper_91__ap_done;
  wire PE_wrapper_91__ap_idle;
  reg [1:0] PE_wrapper_91__state;
  wire PE_wrapper_92__ap_start_global__q0;
  wire PE_wrapper_92__is_done__q0;
  wire PE_wrapper_92__ap_done_global__q0;
  wire PE_wrapper_92__ap_start;
  wire PE_wrapper_92__ap_ready;
  wire PE_wrapper_92__ap_done;
  wire PE_wrapper_92__ap_idle;
  reg [1:0] PE_wrapper_92__state;
  wire PE_wrapper_93__ap_start_global__q0;
  wire PE_wrapper_93__is_done__q0;
  wire PE_wrapper_93__ap_done_global__q0;
  wire PE_wrapper_93__ap_start;
  wire PE_wrapper_93__ap_ready;
  wire PE_wrapper_93__ap_done;
  wire PE_wrapper_93__ap_idle;
  reg [1:0] PE_wrapper_93__state;
  wire PE_wrapper_94__ap_start_global__q0;
  wire PE_wrapper_94__is_done__q0;
  wire PE_wrapper_94__ap_done_global__q0;
  wire PE_wrapper_94__ap_start;
  wire PE_wrapper_94__ap_ready;
  wire PE_wrapper_94__ap_done;
  wire PE_wrapper_94__ap_idle;
  reg [1:0] PE_wrapper_94__state;
  wire PE_wrapper_95__ap_start_global__q0;
  wire PE_wrapper_95__is_done__q0;
  wire PE_wrapper_95__ap_done_global__q0;
  wire PE_wrapper_95__ap_start;
  wire PE_wrapper_95__ap_ready;
  wire PE_wrapper_95__ap_done;
  wire PE_wrapper_95__ap_idle;
  reg [1:0] PE_wrapper_95__state;
  wire PE_wrapper_96__ap_start_global__q0;
  wire PE_wrapper_96__is_done__q0;
  wire PE_wrapper_96__ap_done_global__q0;
  wire PE_wrapper_96__ap_start;
  wire PE_wrapper_96__ap_ready;
  wire PE_wrapper_96__ap_done;
  wire PE_wrapper_96__ap_idle;
  reg [1:0] PE_wrapper_96__state;
  wire PE_wrapper_97__ap_start_global__q0;
  wire PE_wrapper_97__is_done__q0;
  wire PE_wrapper_97__ap_done_global__q0;
  wire PE_wrapper_97__ap_start;
  wire PE_wrapper_97__ap_ready;
  wire PE_wrapper_97__ap_done;
  wire PE_wrapper_97__ap_idle;
  reg [1:0] PE_wrapper_97__state;
  wire PE_wrapper_98__ap_start_global__q0;
  wire PE_wrapper_98__is_done__q0;
  wire PE_wrapper_98__ap_done_global__q0;
  wire PE_wrapper_98__ap_start;
  wire PE_wrapper_98__ap_ready;
  wire PE_wrapper_98__ap_done;
  wire PE_wrapper_98__ap_idle;
  reg [1:0] PE_wrapper_98__state;
  wire PE_wrapper_99__ap_start_global__q0;
  wire PE_wrapper_99__is_done__q0;
  wire PE_wrapper_99__ap_done_global__q0;
  wire PE_wrapper_99__ap_start;
  wire PE_wrapper_99__ap_ready;
  wire PE_wrapper_99__ap_done;
  wire PE_wrapper_99__ap_idle;
  reg [1:0] PE_wrapper_99__state;
  wire PE_wrapper_100__ap_start_global__q0;
  wire PE_wrapper_100__is_done__q0;
  wire PE_wrapper_100__ap_done_global__q0;
  wire PE_wrapper_100__ap_start;
  wire PE_wrapper_100__ap_ready;
  wire PE_wrapper_100__ap_done;
  wire PE_wrapper_100__ap_idle;
  reg [1:0] PE_wrapper_100__state;
  wire PE_wrapper_101__ap_start_global__q0;
  wire PE_wrapper_101__is_done__q0;
  wire PE_wrapper_101__ap_done_global__q0;
  wire PE_wrapper_101__ap_start;
  wire PE_wrapper_101__ap_ready;
  wire PE_wrapper_101__ap_done;
  wire PE_wrapper_101__ap_idle;
  reg [1:0] PE_wrapper_101__state;
  wire PE_wrapper_102__ap_start_global__q0;
  wire PE_wrapper_102__is_done__q0;
  wire PE_wrapper_102__ap_done_global__q0;
  wire PE_wrapper_102__ap_start;
  wire PE_wrapper_102__ap_ready;
  wire PE_wrapper_102__ap_done;
  wire PE_wrapper_102__ap_idle;
  reg [1:0] PE_wrapper_102__state;
  wire PE_wrapper_103__ap_start_global__q0;
  wire PE_wrapper_103__is_done__q0;
  wire PE_wrapper_103__ap_done_global__q0;
  wire PE_wrapper_103__ap_start;
  wire PE_wrapper_103__ap_ready;
  wire PE_wrapper_103__ap_done;
  wire PE_wrapper_103__ap_idle;
  reg [1:0] PE_wrapper_103__state;
  wire PE_wrapper_104__ap_start_global__q0;
  wire PE_wrapper_104__is_done__q0;
  wire PE_wrapper_104__ap_done_global__q0;
  wire PE_wrapper_104__ap_start;
  wire PE_wrapper_104__ap_ready;
  wire PE_wrapper_104__ap_done;
  wire PE_wrapper_104__ap_idle;
  reg [1:0] PE_wrapper_104__state;
  wire PE_wrapper_105__ap_start_global__q0;
  wire PE_wrapper_105__is_done__q0;
  wire PE_wrapper_105__ap_done_global__q0;
  wire PE_wrapper_105__ap_start;
  wire PE_wrapper_105__ap_ready;
  wire PE_wrapper_105__ap_done;
  wire PE_wrapper_105__ap_idle;
  reg [1:0] PE_wrapper_105__state;
  wire PE_wrapper_106__ap_start_global__q0;
  wire PE_wrapper_106__is_done__q0;
  wire PE_wrapper_106__ap_done_global__q0;
  wire PE_wrapper_106__ap_start;
  wire PE_wrapper_106__ap_ready;
  wire PE_wrapper_106__ap_done;
  wire PE_wrapper_106__ap_idle;
  reg [1:0] PE_wrapper_106__state;
  wire PE_wrapper_107__ap_start_global__q0;
  wire PE_wrapper_107__is_done__q0;
  wire PE_wrapper_107__ap_done_global__q0;
  wire PE_wrapper_107__ap_start;
  wire PE_wrapper_107__ap_ready;
  wire PE_wrapper_107__ap_done;
  wire PE_wrapper_107__ap_idle;
  reg [1:0] PE_wrapper_107__state;
  wire PE_wrapper_108__ap_start_global__q0;
  wire PE_wrapper_108__is_done__q0;
  wire PE_wrapper_108__ap_done_global__q0;
  wire PE_wrapper_108__ap_start;
  wire PE_wrapper_108__ap_ready;
  wire PE_wrapper_108__ap_done;
  wire PE_wrapper_108__ap_idle;
  reg [1:0] PE_wrapper_108__state;
  wire PE_wrapper_109__ap_start_global__q0;
  wire PE_wrapper_109__is_done__q0;
  wire PE_wrapper_109__ap_done_global__q0;
  wire PE_wrapper_109__ap_start;
  wire PE_wrapper_109__ap_ready;
  wire PE_wrapper_109__ap_done;
  wire PE_wrapper_109__ap_idle;
  reg [1:0] PE_wrapper_109__state;
  wire PE_wrapper_110__ap_start_global__q0;
  wire PE_wrapper_110__is_done__q0;
  wire PE_wrapper_110__ap_done_global__q0;
  wire PE_wrapper_110__ap_start;
  wire PE_wrapper_110__ap_ready;
  wire PE_wrapper_110__ap_done;
  wire PE_wrapper_110__ap_idle;
  reg [1:0] PE_wrapper_110__state;
  wire PE_wrapper_111__ap_start_global__q0;
  wire PE_wrapper_111__is_done__q0;
  wire PE_wrapper_111__ap_done_global__q0;
  wire PE_wrapper_111__ap_start;
  wire PE_wrapper_111__ap_ready;
  wire PE_wrapper_111__ap_done;
  wire PE_wrapper_111__ap_idle;
  reg [1:0] PE_wrapper_111__state;
  wire PE_wrapper_112__ap_start_global__q0;
  wire PE_wrapper_112__is_done__q0;
  wire PE_wrapper_112__ap_done_global__q0;
  wire PE_wrapper_112__ap_start;
  wire PE_wrapper_112__ap_ready;
  wire PE_wrapper_112__ap_done;
  wire PE_wrapper_112__ap_idle;
  reg [1:0] PE_wrapper_112__state;
  wire PE_wrapper_113__ap_start_global__q0;
  wire PE_wrapper_113__is_done__q0;
  wire PE_wrapper_113__ap_done_global__q0;
  wire PE_wrapper_113__ap_start;
  wire PE_wrapper_113__ap_ready;
  wire PE_wrapper_113__ap_done;
  wire PE_wrapper_113__ap_idle;
  reg [1:0] PE_wrapper_113__state;
  wire PE_wrapper_114__ap_start_global__q0;
  wire PE_wrapper_114__is_done__q0;
  wire PE_wrapper_114__ap_done_global__q0;
  wire PE_wrapper_114__ap_start;
  wire PE_wrapper_114__ap_ready;
  wire PE_wrapper_114__ap_done;
  wire PE_wrapper_114__ap_idle;
  reg [1:0] PE_wrapper_114__state;
  wire PE_wrapper_115__ap_start_global__q0;
  wire PE_wrapper_115__is_done__q0;
  wire PE_wrapper_115__ap_done_global__q0;
  wire PE_wrapper_115__ap_start;
  wire PE_wrapper_115__ap_ready;
  wire PE_wrapper_115__ap_done;
  wire PE_wrapper_115__ap_idle;
  reg [1:0] PE_wrapper_115__state;
  wire PE_wrapper_116__ap_start_global__q0;
  wire PE_wrapper_116__is_done__q0;
  wire PE_wrapper_116__ap_done_global__q0;
  wire PE_wrapper_116__ap_start;
  wire PE_wrapper_116__ap_ready;
  wire PE_wrapper_116__ap_done;
  wire PE_wrapper_116__ap_idle;
  reg [1:0] PE_wrapper_116__state;
  wire PE_wrapper_117__ap_start_global__q0;
  wire PE_wrapper_117__is_done__q0;
  wire PE_wrapper_117__ap_done_global__q0;
  wire PE_wrapper_117__ap_start;
  wire PE_wrapper_117__ap_ready;
  wire PE_wrapper_117__ap_done;
  wire PE_wrapper_117__ap_idle;
  reg [1:0] PE_wrapper_117__state;
  wire PE_wrapper_118__ap_start_global__q0;
  wire PE_wrapper_118__is_done__q0;
  wire PE_wrapper_118__ap_done_global__q0;
  wire PE_wrapper_118__ap_start;
  wire PE_wrapper_118__ap_ready;
  wire PE_wrapper_118__ap_done;
  wire PE_wrapper_118__ap_idle;
  reg [1:0] PE_wrapper_118__state;
  wire PE_wrapper_119__ap_start_global__q0;
  wire PE_wrapper_119__is_done__q0;
  wire PE_wrapper_119__ap_done_global__q0;
  wire PE_wrapper_119__ap_start;
  wire PE_wrapper_119__ap_ready;
  wire PE_wrapper_119__ap_done;
  wire PE_wrapper_119__ap_idle;
  reg [1:0] PE_wrapper_119__state;
  wire PE_wrapper_120__ap_start_global__q0;
  wire PE_wrapper_120__is_done__q0;
  wire PE_wrapper_120__ap_done_global__q0;
  wire PE_wrapper_120__ap_start;
  wire PE_wrapper_120__ap_ready;
  wire PE_wrapper_120__ap_done;
  wire PE_wrapper_120__ap_idle;
  reg [1:0] PE_wrapper_120__state;
  wire PE_wrapper_121__ap_start_global__q0;
  wire PE_wrapper_121__is_done__q0;
  wire PE_wrapper_121__ap_done_global__q0;
  wire PE_wrapper_121__ap_start;
  wire PE_wrapper_121__ap_ready;
  wire PE_wrapper_121__ap_done;
  wire PE_wrapper_121__ap_idle;
  reg [1:0] PE_wrapper_121__state;
  wire PE_wrapper_122__ap_start_global__q0;
  wire PE_wrapper_122__is_done__q0;
  wire PE_wrapper_122__ap_done_global__q0;
  wire PE_wrapper_122__ap_start;
  wire PE_wrapper_122__ap_ready;
  wire PE_wrapper_122__ap_done;
  wire PE_wrapper_122__ap_idle;
  reg [1:0] PE_wrapper_122__state;
  wire PE_wrapper_123__ap_start_global__q0;
  wire PE_wrapper_123__is_done__q0;
  wire PE_wrapper_123__ap_done_global__q0;
  wire PE_wrapper_123__ap_start;
  wire PE_wrapper_123__ap_ready;
  wire PE_wrapper_123__ap_done;
  wire PE_wrapper_123__ap_idle;
  reg [1:0] PE_wrapper_123__state;
  wire PE_wrapper_124__ap_start_global__q0;
  wire PE_wrapper_124__is_done__q0;
  wire PE_wrapper_124__ap_done_global__q0;
  wire PE_wrapper_124__ap_start;
  wire PE_wrapper_124__ap_ready;
  wire PE_wrapper_124__ap_done;
  wire PE_wrapper_124__ap_idle;
  reg [1:0] PE_wrapper_124__state;
  wire PE_wrapper_125__ap_start_global__q0;
  wire PE_wrapper_125__is_done__q0;
  wire PE_wrapper_125__ap_done_global__q0;
  wire PE_wrapper_125__ap_start;
  wire PE_wrapper_125__ap_ready;
  wire PE_wrapper_125__ap_done;
  wire PE_wrapper_125__ap_idle;
  reg [1:0] PE_wrapper_125__state;
  wire PE_wrapper_126__ap_start_global__q0;
  wire PE_wrapper_126__is_done__q0;
  wire PE_wrapper_126__ap_done_global__q0;
  wire PE_wrapper_126__ap_start;
  wire PE_wrapper_126__ap_ready;
  wire PE_wrapper_126__ap_done;
  wire PE_wrapper_126__ap_idle;
  reg [1:0] PE_wrapper_126__state;
  wire PE_wrapper_127__ap_start_global__q0;
  wire PE_wrapper_127__is_done__q0;
  wire PE_wrapper_127__ap_done_global__q0;
  wire PE_wrapper_127__ap_start;
  wire PE_wrapper_127__ap_ready;
  wire PE_wrapper_127__ap_done;
  wire PE_wrapper_127__ap_idle;
  reg [1:0] PE_wrapper_127__state;
  wire PE_wrapper_128__ap_start_global__q0;
  wire PE_wrapper_128__is_done__q0;
  wire PE_wrapper_128__ap_done_global__q0;
  wire PE_wrapper_128__ap_start;
  wire PE_wrapper_128__ap_ready;
  wire PE_wrapper_128__ap_done;
  wire PE_wrapper_128__ap_idle;
  reg [1:0] PE_wrapper_128__state;
  wire PE_wrapper_129__ap_start_global__q0;
  wire PE_wrapper_129__is_done__q0;
  wire PE_wrapper_129__ap_done_global__q0;
  wire PE_wrapper_129__ap_start;
  wire PE_wrapper_129__ap_ready;
  wire PE_wrapper_129__ap_done;
  wire PE_wrapper_129__ap_idle;
  reg [1:0] PE_wrapper_129__state;
  wire PE_wrapper_130__ap_start_global__q0;
  wire PE_wrapper_130__is_done__q0;
  wire PE_wrapper_130__ap_done_global__q0;
  wire PE_wrapper_130__ap_start;
  wire PE_wrapper_130__ap_ready;
  wire PE_wrapper_130__ap_done;
  wire PE_wrapper_130__ap_idle;
  reg [1:0] PE_wrapper_130__state;
  wire PE_wrapper_131__ap_start_global__q0;
  wire PE_wrapper_131__is_done__q0;
  wire PE_wrapper_131__ap_done_global__q0;
  wire PE_wrapper_131__ap_start;
  wire PE_wrapper_131__ap_ready;
  wire PE_wrapper_131__ap_done;
  wire PE_wrapper_131__ap_idle;
  reg [1:0] PE_wrapper_131__state;
  wire PE_wrapper_132__ap_start_global__q0;
  wire PE_wrapper_132__is_done__q0;
  wire PE_wrapper_132__ap_done_global__q0;
  wire PE_wrapper_132__ap_start;
  wire PE_wrapper_132__ap_ready;
  wire PE_wrapper_132__ap_done;
  wire PE_wrapper_132__ap_idle;
  reg [1:0] PE_wrapper_132__state;
  wire PE_wrapper_133__ap_start_global__q0;
  wire PE_wrapper_133__is_done__q0;
  wire PE_wrapper_133__ap_done_global__q0;
  wire PE_wrapper_133__ap_start;
  wire PE_wrapper_133__ap_ready;
  wire PE_wrapper_133__ap_done;
  wire PE_wrapper_133__ap_idle;
  reg [1:0] PE_wrapper_133__state;
  wire PE_wrapper_134__ap_start_global__q0;
  wire PE_wrapper_134__is_done__q0;
  wire PE_wrapper_134__ap_done_global__q0;
  wire PE_wrapper_134__ap_start;
  wire PE_wrapper_134__ap_ready;
  wire PE_wrapper_134__ap_done;
  wire PE_wrapper_134__ap_idle;
  reg [1:0] PE_wrapper_134__state;
  wire PE_wrapper_135__ap_start_global__q0;
  wire PE_wrapper_135__is_done__q0;
  wire PE_wrapper_135__ap_done_global__q0;
  wire PE_wrapper_135__ap_start;
  wire PE_wrapper_135__ap_ready;
  wire PE_wrapper_135__ap_done;
  wire PE_wrapper_135__ap_idle;
  reg [1:0] PE_wrapper_135__state;
  wire PE_wrapper_136__ap_start_global__q0;
  wire PE_wrapper_136__is_done__q0;
  wire PE_wrapper_136__ap_done_global__q0;
  wire PE_wrapper_136__ap_start;
  wire PE_wrapper_136__ap_ready;
  wire PE_wrapper_136__ap_done;
  wire PE_wrapper_136__ap_idle;
  reg [1:0] PE_wrapper_136__state;
  wire PE_wrapper_137__ap_start_global__q0;
  wire PE_wrapper_137__is_done__q0;
  wire PE_wrapper_137__ap_done_global__q0;
  wire PE_wrapper_137__ap_start;
  wire PE_wrapper_137__ap_ready;
  wire PE_wrapper_137__ap_done;
  wire PE_wrapper_137__ap_idle;
  reg [1:0] PE_wrapper_137__state;
  wire PE_wrapper_138__ap_start_global__q0;
  wire PE_wrapper_138__is_done__q0;
  wire PE_wrapper_138__ap_done_global__q0;
  wire PE_wrapper_138__ap_start;
  wire PE_wrapper_138__ap_ready;
  wire PE_wrapper_138__ap_done;
  wire PE_wrapper_138__ap_idle;
  reg [1:0] PE_wrapper_138__state;
  wire PE_wrapper_139__ap_start_global__q0;
  wire PE_wrapper_139__is_done__q0;
  wire PE_wrapper_139__ap_done_global__q0;
  wire PE_wrapper_139__ap_start;
  wire PE_wrapper_139__ap_ready;
  wire PE_wrapper_139__ap_done;
  wire PE_wrapper_139__ap_idle;
  reg [1:0] PE_wrapper_139__state;
  wire PE_wrapper_140__ap_start_global__q0;
  wire PE_wrapper_140__is_done__q0;
  wire PE_wrapper_140__ap_done_global__q0;
  wire PE_wrapper_140__ap_start;
  wire PE_wrapper_140__ap_ready;
  wire PE_wrapper_140__ap_done;
  wire PE_wrapper_140__ap_idle;
  reg [1:0] PE_wrapper_140__state;
  wire PE_wrapper_141__ap_start_global__q0;
  wire PE_wrapper_141__is_done__q0;
  wire PE_wrapper_141__ap_done_global__q0;
  wire PE_wrapper_141__ap_start;
  wire PE_wrapper_141__ap_ready;
  wire PE_wrapper_141__ap_done;
  wire PE_wrapper_141__ap_idle;
  reg [1:0] PE_wrapper_141__state;
  wire PE_wrapper_142__ap_start_global__q0;
  wire PE_wrapper_142__is_done__q0;
  wire PE_wrapper_142__ap_done_global__q0;
  wire PE_wrapper_142__ap_start;
  wire PE_wrapper_142__ap_ready;
  wire PE_wrapper_142__ap_done;
  wire PE_wrapper_142__ap_idle;
  reg [1:0] PE_wrapper_142__state;
  wire PE_wrapper_143__ap_start_global__q0;
  wire PE_wrapper_143__is_done__q0;
  wire PE_wrapper_143__ap_done_global__q0;
  wire PE_wrapper_143__ap_start;
  wire PE_wrapper_143__ap_ready;
  wire PE_wrapper_143__ap_done;
  wire PE_wrapper_143__ap_idle;
  reg [1:0] PE_wrapper_143__state;
  wire PE_wrapper_144__ap_start_global__q0;
  wire PE_wrapper_144__is_done__q0;
  wire PE_wrapper_144__ap_done_global__q0;
  wire PE_wrapper_144__ap_start;
  wire PE_wrapper_144__ap_ready;
  wire PE_wrapper_144__ap_done;
  wire PE_wrapper_144__ap_idle;
  reg [1:0] PE_wrapper_144__state;
  wire PE_wrapper_145__ap_start_global__q0;
  wire PE_wrapper_145__is_done__q0;
  wire PE_wrapper_145__ap_done_global__q0;
  wire PE_wrapper_145__ap_start;
  wire PE_wrapper_145__ap_ready;
  wire PE_wrapper_145__ap_done;
  wire PE_wrapper_145__ap_idle;
  reg [1:0] PE_wrapper_145__state;
  wire PE_wrapper_146__ap_start_global__q0;
  wire PE_wrapper_146__is_done__q0;
  wire PE_wrapper_146__ap_done_global__q0;
  wire PE_wrapper_146__ap_start;
  wire PE_wrapper_146__ap_ready;
  wire PE_wrapper_146__ap_done;
  wire PE_wrapper_146__ap_idle;
  reg [1:0] PE_wrapper_146__state;
  wire PE_wrapper_147__ap_start_global__q0;
  wire PE_wrapper_147__is_done__q0;
  wire PE_wrapper_147__ap_done_global__q0;
  wire PE_wrapper_147__ap_start;
  wire PE_wrapper_147__ap_ready;
  wire PE_wrapper_147__ap_done;
  wire PE_wrapper_147__ap_idle;
  reg [1:0] PE_wrapper_147__state;
  wire PE_wrapper_148__ap_start_global__q0;
  wire PE_wrapper_148__is_done__q0;
  wire PE_wrapper_148__ap_done_global__q0;
  wire PE_wrapper_148__ap_start;
  wire PE_wrapper_148__ap_ready;
  wire PE_wrapper_148__ap_done;
  wire PE_wrapper_148__ap_idle;
  reg [1:0] PE_wrapper_148__state;
  wire PE_wrapper_149__ap_start_global__q0;
  wire PE_wrapper_149__is_done__q0;
  wire PE_wrapper_149__ap_done_global__q0;
  wire PE_wrapper_149__ap_start;
  wire PE_wrapper_149__ap_ready;
  wire PE_wrapper_149__ap_done;
  wire PE_wrapper_149__ap_idle;
  reg [1:0] PE_wrapper_149__state;
  wire PE_wrapper_150__ap_start_global__q0;
  wire PE_wrapper_150__is_done__q0;
  wire PE_wrapper_150__ap_done_global__q0;
  wire PE_wrapper_150__ap_start;
  wire PE_wrapper_150__ap_ready;
  wire PE_wrapper_150__ap_done;
  wire PE_wrapper_150__ap_idle;
  reg [1:0] PE_wrapper_150__state;
  wire PE_wrapper_151__ap_start_global__q0;
  wire PE_wrapper_151__is_done__q0;
  wire PE_wrapper_151__ap_done_global__q0;
  wire PE_wrapper_151__ap_start;
  wire PE_wrapper_151__ap_ready;
  wire PE_wrapper_151__ap_done;
  wire PE_wrapper_151__ap_idle;
  reg [1:0] PE_wrapper_151__state;
  wire PE_wrapper_152__ap_start_global__q0;
  wire PE_wrapper_152__is_done__q0;
  wire PE_wrapper_152__ap_done_global__q0;
  wire PE_wrapper_152__ap_start;
  wire PE_wrapper_152__ap_ready;
  wire PE_wrapper_152__ap_done;
  wire PE_wrapper_152__ap_idle;
  reg [1:0] PE_wrapper_152__state;
  wire PE_wrapper_153__ap_start_global__q0;
  wire PE_wrapper_153__is_done__q0;
  wire PE_wrapper_153__ap_done_global__q0;
  wire PE_wrapper_153__ap_start;
  wire PE_wrapper_153__ap_ready;
  wire PE_wrapper_153__ap_done;
  wire PE_wrapper_153__ap_idle;
  reg [1:0] PE_wrapper_153__state;
  wire PE_wrapper_154__ap_start_global__q0;
  wire PE_wrapper_154__is_done__q0;
  wire PE_wrapper_154__ap_done_global__q0;
  wire PE_wrapper_154__ap_start;
  wire PE_wrapper_154__ap_ready;
  wire PE_wrapper_154__ap_done;
  wire PE_wrapper_154__ap_idle;
  reg [1:0] PE_wrapper_154__state;
  wire PE_wrapper_155__ap_start_global__q0;
  wire PE_wrapper_155__is_done__q0;
  wire PE_wrapper_155__ap_done_global__q0;
  wire PE_wrapper_155__ap_start;
  wire PE_wrapper_155__ap_ready;
  wire PE_wrapper_155__ap_done;
  wire PE_wrapper_155__ap_idle;
  reg [1:0] PE_wrapper_155__state;
  wire PE_wrapper_156__ap_start_global__q0;
  wire PE_wrapper_156__is_done__q0;
  wire PE_wrapper_156__ap_done_global__q0;
  wire PE_wrapper_156__ap_start;
  wire PE_wrapper_156__ap_ready;
  wire PE_wrapper_156__ap_done;
  wire PE_wrapper_156__ap_idle;
  reg [1:0] PE_wrapper_156__state;
  wire PE_wrapper_157__ap_start_global__q0;
  wire PE_wrapper_157__is_done__q0;
  wire PE_wrapper_157__ap_done_global__q0;
  wire PE_wrapper_157__ap_start;
  wire PE_wrapper_157__ap_ready;
  wire PE_wrapper_157__ap_done;
  wire PE_wrapper_157__ap_idle;
  reg [1:0] PE_wrapper_157__state;
  wire PE_wrapper_158__ap_start_global__q0;
  wire PE_wrapper_158__is_done__q0;
  wire PE_wrapper_158__ap_done_global__q0;
  wire PE_wrapper_158__ap_start;
  wire PE_wrapper_158__ap_ready;
  wire PE_wrapper_158__ap_done;
  wire PE_wrapper_158__ap_idle;
  reg [1:0] PE_wrapper_158__state;
  wire PE_wrapper_159__ap_start_global__q0;
  wire PE_wrapper_159__is_done__q0;
  wire PE_wrapper_159__ap_done_global__q0;
  wire PE_wrapper_159__ap_start;
  wire PE_wrapper_159__ap_ready;
  wire PE_wrapper_159__ap_done;
  wire PE_wrapper_159__ap_idle;
  reg [1:0] PE_wrapper_159__state;
  wire PE_wrapper_160__ap_start_global__q0;
  wire PE_wrapper_160__is_done__q0;
  wire PE_wrapper_160__ap_done_global__q0;
  wire PE_wrapper_160__ap_start;
  wire PE_wrapper_160__ap_ready;
  wire PE_wrapper_160__ap_done;
  wire PE_wrapper_160__ap_idle;
  reg [1:0] PE_wrapper_160__state;
  wire PE_wrapper_161__ap_start_global__q0;
  wire PE_wrapper_161__is_done__q0;
  wire PE_wrapper_161__ap_done_global__q0;
  wire PE_wrapper_161__ap_start;
  wire PE_wrapper_161__ap_ready;
  wire PE_wrapper_161__ap_done;
  wire PE_wrapper_161__ap_idle;
  reg [1:0] PE_wrapper_161__state;
  wire PE_wrapper_162__ap_start_global__q0;
  wire PE_wrapper_162__is_done__q0;
  wire PE_wrapper_162__ap_done_global__q0;
  wire PE_wrapper_162__ap_start;
  wire PE_wrapper_162__ap_ready;
  wire PE_wrapper_162__ap_done;
  wire PE_wrapper_162__ap_idle;
  reg [1:0] PE_wrapper_162__state;
  wire PE_wrapper_163__ap_start_global__q0;
  wire PE_wrapper_163__is_done__q0;
  wire PE_wrapper_163__ap_done_global__q0;
  wire PE_wrapper_163__ap_start;
  wire PE_wrapper_163__ap_ready;
  wire PE_wrapper_163__ap_done;
  wire PE_wrapper_163__ap_idle;
  reg [1:0] PE_wrapper_163__state;
  wire PE_wrapper_164__ap_start_global__q0;
  wire PE_wrapper_164__is_done__q0;
  wire PE_wrapper_164__ap_done_global__q0;
  wire PE_wrapper_164__ap_start;
  wire PE_wrapper_164__ap_ready;
  wire PE_wrapper_164__ap_done;
  wire PE_wrapper_164__ap_idle;
  reg [1:0] PE_wrapper_164__state;
  wire PE_wrapper_165__ap_start_global__q0;
  wire PE_wrapper_165__is_done__q0;
  wire PE_wrapper_165__ap_done_global__q0;
  wire PE_wrapper_165__ap_start;
  wire PE_wrapper_165__ap_ready;
  wire PE_wrapper_165__ap_done;
  wire PE_wrapper_165__ap_idle;
  reg [1:0] PE_wrapper_165__state;
  wire PE_wrapper_166__ap_start_global__q0;
  wire PE_wrapper_166__is_done__q0;
  wire PE_wrapper_166__ap_done_global__q0;
  wire PE_wrapper_166__ap_start;
  wire PE_wrapper_166__ap_ready;
  wire PE_wrapper_166__ap_done;
  wire PE_wrapper_166__ap_idle;
  reg [1:0] PE_wrapper_166__state;
  wire PE_wrapper_167__ap_start_global__q0;
  wire PE_wrapper_167__is_done__q0;
  wire PE_wrapper_167__ap_done_global__q0;
  wire PE_wrapper_167__ap_start;
  wire PE_wrapper_167__ap_ready;
  wire PE_wrapper_167__ap_done;
  wire PE_wrapper_167__ap_idle;
  reg [1:0] PE_wrapper_167__state;
  wire PE_wrapper_168__ap_start_global__q0;
  wire PE_wrapper_168__is_done__q0;
  wire PE_wrapper_168__ap_done_global__q0;
  wire PE_wrapper_168__ap_start;
  wire PE_wrapper_168__ap_ready;
  wire PE_wrapper_168__ap_done;
  wire PE_wrapper_168__ap_idle;
  reg [1:0] PE_wrapper_168__state;
  wire PE_wrapper_169__ap_start_global__q0;
  wire PE_wrapper_169__is_done__q0;
  wire PE_wrapper_169__ap_done_global__q0;
  wire PE_wrapper_169__ap_start;
  wire PE_wrapper_169__ap_ready;
  wire PE_wrapper_169__ap_done;
  wire PE_wrapper_169__ap_idle;
  reg [1:0] PE_wrapper_169__state;
  wire PE_wrapper_170__ap_start_global__q0;
  wire PE_wrapper_170__is_done__q0;
  wire PE_wrapper_170__ap_done_global__q0;
  wire PE_wrapper_170__ap_start;
  wire PE_wrapper_170__ap_ready;
  wire PE_wrapper_170__ap_done;
  wire PE_wrapper_170__ap_idle;
  reg [1:0] PE_wrapper_170__state;
  wire PE_wrapper_171__ap_start_global__q0;
  wire PE_wrapper_171__is_done__q0;
  wire PE_wrapper_171__ap_done_global__q0;
  wire PE_wrapper_171__ap_start;
  wire PE_wrapper_171__ap_ready;
  wire PE_wrapper_171__ap_done;
  wire PE_wrapper_171__ap_idle;
  reg [1:0] PE_wrapper_171__state;
  wire PE_wrapper_172__ap_start_global__q0;
  wire PE_wrapper_172__is_done__q0;
  wire PE_wrapper_172__ap_done_global__q0;
  wire PE_wrapper_172__ap_start;
  wire PE_wrapper_172__ap_ready;
  wire PE_wrapper_172__ap_done;
  wire PE_wrapper_172__ap_idle;
  reg [1:0] PE_wrapper_172__state;
  wire PE_wrapper_173__ap_start_global__q0;
  wire PE_wrapper_173__is_done__q0;
  wire PE_wrapper_173__ap_done_global__q0;
  wire PE_wrapper_173__ap_start;
  wire PE_wrapper_173__ap_ready;
  wire PE_wrapper_173__ap_done;
  wire PE_wrapper_173__ap_idle;
  reg [1:0] PE_wrapper_173__state;
  wire PE_wrapper_174__ap_start_global__q0;
  wire PE_wrapper_174__is_done__q0;
  wire PE_wrapper_174__ap_done_global__q0;
  wire PE_wrapper_174__ap_start;
  wire PE_wrapper_174__ap_ready;
  wire PE_wrapper_174__ap_done;
  wire PE_wrapper_174__ap_idle;
  reg [1:0] PE_wrapper_174__state;
  wire PE_wrapper_175__ap_start_global__q0;
  wire PE_wrapper_175__is_done__q0;
  wire PE_wrapper_175__ap_done_global__q0;
  wire PE_wrapper_175__ap_start;
  wire PE_wrapper_175__ap_ready;
  wire PE_wrapper_175__ap_done;
  wire PE_wrapper_175__ap_idle;
  reg [1:0] PE_wrapper_175__state;
  wire PE_wrapper_176__ap_start_global__q0;
  wire PE_wrapper_176__is_done__q0;
  wire PE_wrapper_176__ap_done_global__q0;
  wire PE_wrapper_176__ap_start;
  wire PE_wrapper_176__ap_ready;
  wire PE_wrapper_176__ap_done;
  wire PE_wrapper_176__ap_idle;
  reg [1:0] PE_wrapper_176__state;
  wire PE_wrapper_177__ap_start_global__q0;
  wire PE_wrapper_177__is_done__q0;
  wire PE_wrapper_177__ap_done_global__q0;
  wire PE_wrapper_177__ap_start;
  wire PE_wrapper_177__ap_ready;
  wire PE_wrapper_177__ap_done;
  wire PE_wrapper_177__ap_idle;
  reg [1:0] PE_wrapper_177__state;
  wire PE_wrapper_178__ap_start_global__q0;
  wire PE_wrapper_178__is_done__q0;
  wire PE_wrapper_178__ap_done_global__q0;
  wire PE_wrapper_178__ap_start;
  wire PE_wrapper_178__ap_ready;
  wire PE_wrapper_178__ap_done;
  wire PE_wrapper_178__ap_idle;
  reg [1:0] PE_wrapper_178__state;
  wire PE_wrapper_179__ap_start_global__q0;
  wire PE_wrapper_179__is_done__q0;
  wire PE_wrapper_179__ap_done_global__q0;
  wire PE_wrapper_179__ap_start;
  wire PE_wrapper_179__ap_ready;
  wire PE_wrapper_179__ap_done;
  wire PE_wrapper_179__ap_idle;
  reg [1:0] PE_wrapper_179__state;
  wire PE_wrapper_180__ap_start_global__q0;
  wire PE_wrapper_180__is_done__q0;
  wire PE_wrapper_180__ap_done_global__q0;
  wire PE_wrapper_180__ap_start;
  wire PE_wrapper_180__ap_ready;
  wire PE_wrapper_180__ap_done;
  wire PE_wrapper_180__ap_idle;
  reg [1:0] PE_wrapper_180__state;
  wire PE_wrapper_181__ap_start_global__q0;
  wire PE_wrapper_181__is_done__q0;
  wire PE_wrapper_181__ap_done_global__q0;
  wire PE_wrapper_181__ap_start;
  wire PE_wrapper_181__ap_ready;
  wire PE_wrapper_181__ap_done;
  wire PE_wrapper_181__ap_idle;
  reg [1:0] PE_wrapper_181__state;
  wire PE_wrapper_182__ap_start_global__q0;
  wire PE_wrapper_182__is_done__q0;
  wire PE_wrapper_182__ap_done_global__q0;
  wire PE_wrapper_182__ap_start;
  wire PE_wrapper_182__ap_ready;
  wire PE_wrapper_182__ap_done;
  wire PE_wrapper_182__ap_idle;
  reg [1:0] PE_wrapper_182__state;
  wire PE_wrapper_183__ap_start_global__q0;
  wire PE_wrapper_183__is_done__q0;
  wire PE_wrapper_183__ap_done_global__q0;
  wire PE_wrapper_183__ap_start;
  wire PE_wrapper_183__ap_ready;
  wire PE_wrapper_183__ap_done;
  wire PE_wrapper_183__ap_idle;
  reg [1:0] PE_wrapper_183__state;
  wire PE_wrapper_184__ap_start_global__q0;
  wire PE_wrapper_184__is_done__q0;
  wire PE_wrapper_184__ap_done_global__q0;
  wire PE_wrapper_184__ap_start;
  wire PE_wrapper_184__ap_ready;
  wire PE_wrapper_184__ap_done;
  wire PE_wrapper_184__ap_idle;
  reg [1:0] PE_wrapper_184__state;
  wire PE_wrapper_185__ap_start_global__q0;
  wire PE_wrapper_185__is_done__q0;
  wire PE_wrapper_185__ap_done_global__q0;
  wire PE_wrapper_185__ap_start;
  wire PE_wrapper_185__ap_ready;
  wire PE_wrapper_185__ap_done;
  wire PE_wrapper_185__ap_idle;
  reg [1:0] PE_wrapper_185__state;
  wire PE_wrapper_186__ap_start_global__q0;
  wire PE_wrapper_186__is_done__q0;
  wire PE_wrapper_186__ap_done_global__q0;
  wire PE_wrapper_186__ap_start;
  wire PE_wrapper_186__ap_ready;
  wire PE_wrapper_186__ap_done;
  wire PE_wrapper_186__ap_idle;
  reg [1:0] PE_wrapper_186__state;
  wire PE_wrapper_187__ap_start_global__q0;
  wire PE_wrapper_187__is_done__q0;
  wire PE_wrapper_187__ap_done_global__q0;
  wire PE_wrapper_187__ap_start;
  wire PE_wrapper_187__ap_ready;
  wire PE_wrapper_187__ap_done;
  wire PE_wrapper_187__ap_idle;
  reg [1:0] PE_wrapper_187__state;
  wire PE_wrapper_188__ap_start_global__q0;
  wire PE_wrapper_188__is_done__q0;
  wire PE_wrapper_188__ap_done_global__q0;
  wire PE_wrapper_188__ap_start;
  wire PE_wrapper_188__ap_ready;
  wire PE_wrapper_188__ap_done;
  wire PE_wrapper_188__ap_idle;
  reg [1:0] PE_wrapper_188__state;
  wire PE_wrapper_189__ap_start_global__q0;
  wire PE_wrapper_189__is_done__q0;
  wire PE_wrapper_189__ap_done_global__q0;
  wire PE_wrapper_189__ap_start;
  wire PE_wrapper_189__ap_ready;
  wire PE_wrapper_189__ap_done;
  wire PE_wrapper_189__ap_idle;
  reg [1:0] PE_wrapper_189__state;
  wire PE_wrapper_190__ap_start_global__q0;
  wire PE_wrapper_190__is_done__q0;
  wire PE_wrapper_190__ap_done_global__q0;
  wire PE_wrapper_190__ap_start;
  wire PE_wrapper_190__ap_ready;
  wire PE_wrapper_190__ap_done;
  wire PE_wrapper_190__ap_idle;
  reg [1:0] PE_wrapper_190__state;
  wire PE_wrapper_191__ap_start_global__q0;
  wire PE_wrapper_191__is_done__q0;
  wire PE_wrapper_191__ap_done_global__q0;
  wire PE_wrapper_191__ap_start;
  wire PE_wrapper_191__ap_ready;
  wire PE_wrapper_191__ap_done;
  wire PE_wrapper_191__ap_idle;
  reg [1:0] PE_wrapper_191__state;
  wire PE_wrapper_192__ap_start_global__q0;
  wire PE_wrapper_192__is_done__q0;
  wire PE_wrapper_192__ap_done_global__q0;
  wire PE_wrapper_192__ap_start;
  wire PE_wrapper_192__ap_ready;
  wire PE_wrapper_192__ap_done;
  wire PE_wrapper_192__ap_idle;
  reg [1:0] PE_wrapper_192__state;
  wire PE_wrapper_193__ap_start_global__q0;
  wire PE_wrapper_193__is_done__q0;
  wire PE_wrapper_193__ap_done_global__q0;
  wire PE_wrapper_193__ap_start;
  wire PE_wrapper_193__ap_ready;
  wire PE_wrapper_193__ap_done;
  wire PE_wrapper_193__ap_idle;
  reg [1:0] PE_wrapper_193__state;
  wire PE_wrapper_194__ap_start_global__q0;
  wire PE_wrapper_194__is_done__q0;
  wire PE_wrapper_194__ap_done_global__q0;
  wire PE_wrapper_194__ap_start;
  wire PE_wrapper_194__ap_ready;
  wire PE_wrapper_194__ap_done;
  wire PE_wrapper_194__ap_idle;
  reg [1:0] PE_wrapper_194__state;
  wire PE_wrapper_195__ap_start_global__q0;
  wire PE_wrapper_195__is_done__q0;
  wire PE_wrapper_195__ap_done_global__q0;
  wire PE_wrapper_195__ap_start;
  wire PE_wrapper_195__ap_ready;
  wire PE_wrapper_195__ap_done;
  wire PE_wrapper_195__ap_idle;
  reg [1:0] PE_wrapper_195__state;
  wire PE_wrapper_196__ap_start_global__q0;
  wire PE_wrapper_196__is_done__q0;
  wire PE_wrapper_196__ap_done_global__q0;
  wire PE_wrapper_196__ap_start;
  wire PE_wrapper_196__ap_ready;
  wire PE_wrapper_196__ap_done;
  wire PE_wrapper_196__ap_idle;
  reg [1:0] PE_wrapper_196__state;
  wire PE_wrapper_197__ap_start_global__q0;
  wire PE_wrapper_197__is_done__q0;
  wire PE_wrapper_197__ap_done_global__q0;
  wire PE_wrapper_197__ap_start;
  wire PE_wrapper_197__ap_ready;
  wire PE_wrapper_197__ap_done;
  wire PE_wrapper_197__ap_idle;
  reg [1:0] PE_wrapper_197__state;
  wire PE_wrapper_198__ap_start_global__q0;
  wire PE_wrapper_198__is_done__q0;
  wire PE_wrapper_198__ap_done_global__q0;
  wire PE_wrapper_198__ap_start;
  wire PE_wrapper_198__ap_ready;
  wire PE_wrapper_198__ap_done;
  wire PE_wrapper_198__ap_idle;
  reg [1:0] PE_wrapper_198__state;
  wire PE_wrapper_199__ap_start_global__q0;
  wire PE_wrapper_199__is_done__q0;
  wire PE_wrapper_199__ap_done_global__q0;
  wire PE_wrapper_199__ap_start;
  wire PE_wrapper_199__ap_ready;
  wire PE_wrapper_199__ap_done;
  wire PE_wrapper_199__ap_idle;
  reg [1:0] PE_wrapper_199__state;
  wire PE_wrapper_200__ap_start_global__q0;
  wire PE_wrapper_200__is_done__q0;
  wire PE_wrapper_200__ap_done_global__q0;
  wire PE_wrapper_200__ap_start;
  wire PE_wrapper_200__ap_ready;
  wire PE_wrapper_200__ap_done;
  wire PE_wrapper_200__ap_idle;
  reg [1:0] PE_wrapper_200__state;
  wire PE_wrapper_201__ap_start_global__q0;
  wire PE_wrapper_201__is_done__q0;
  wire PE_wrapper_201__ap_done_global__q0;
  wire PE_wrapper_201__ap_start;
  wire PE_wrapper_201__ap_ready;
  wire PE_wrapper_201__ap_done;
  wire PE_wrapper_201__ap_idle;
  reg [1:0] PE_wrapper_201__state;
  wire PE_wrapper_202__ap_start_global__q0;
  wire PE_wrapper_202__is_done__q0;
  wire PE_wrapper_202__ap_done_global__q0;
  wire PE_wrapper_202__ap_start;
  wire PE_wrapper_202__ap_ready;
  wire PE_wrapper_202__ap_done;
  wire PE_wrapper_202__ap_idle;
  reg [1:0] PE_wrapper_202__state;
  wire PE_wrapper_203__ap_start_global__q0;
  wire PE_wrapper_203__is_done__q0;
  wire PE_wrapper_203__ap_done_global__q0;
  wire PE_wrapper_203__ap_start;
  wire PE_wrapper_203__ap_ready;
  wire PE_wrapper_203__ap_done;
  wire PE_wrapper_203__ap_idle;
  reg [1:0] PE_wrapper_203__state;
  wire PE_wrapper_204__ap_start_global__q0;
  wire PE_wrapper_204__is_done__q0;
  wire PE_wrapper_204__ap_done_global__q0;
  wire PE_wrapper_204__ap_start;
  wire PE_wrapper_204__ap_ready;
  wire PE_wrapper_204__ap_done;
  wire PE_wrapper_204__ap_idle;
  reg [1:0] PE_wrapper_204__state;
  wire PE_wrapper_205__ap_start_global__q0;
  wire PE_wrapper_205__is_done__q0;
  wire PE_wrapper_205__ap_done_global__q0;
  wire PE_wrapper_205__ap_start;
  wire PE_wrapper_205__ap_ready;
  wire PE_wrapper_205__ap_done;
  wire PE_wrapper_205__ap_idle;
  reg [1:0] PE_wrapper_205__state;
  wire PE_wrapper_206__ap_start_global__q0;
  wire PE_wrapper_206__is_done__q0;
  wire PE_wrapper_206__ap_done_global__q0;
  wire PE_wrapper_206__ap_start;
  wire PE_wrapper_206__ap_ready;
  wire PE_wrapper_206__ap_done;
  wire PE_wrapper_206__ap_idle;
  reg [1:0] PE_wrapper_206__state;
  wire PE_wrapper_207__ap_start_global__q0;
  wire PE_wrapper_207__is_done__q0;
  wire PE_wrapper_207__ap_done_global__q0;
  wire PE_wrapper_207__ap_start;
  wire PE_wrapper_207__ap_ready;
  wire PE_wrapper_207__ap_done;
  wire PE_wrapper_207__ap_idle;
  reg [1:0] PE_wrapper_207__state;
  wire PE_wrapper_208__ap_start_global__q0;
  wire PE_wrapper_208__is_done__q0;
  wire PE_wrapper_208__ap_done_global__q0;
  wire PE_wrapper_208__ap_start;
  wire PE_wrapper_208__ap_ready;
  wire PE_wrapper_208__ap_done;
  wire PE_wrapper_208__ap_idle;
  reg [1:0] PE_wrapper_208__state;
  wire PE_wrapper_209__ap_start_global__q0;
  wire PE_wrapper_209__is_done__q0;
  wire PE_wrapper_209__ap_done_global__q0;
  wire PE_wrapper_209__ap_start;
  wire PE_wrapper_209__ap_ready;
  wire PE_wrapper_209__ap_done;
  wire PE_wrapper_209__ap_idle;
  reg [1:0] PE_wrapper_209__state;
  wire PE_wrapper_210__ap_start_global__q0;
  wire PE_wrapper_210__is_done__q0;
  wire PE_wrapper_210__ap_done_global__q0;
  wire PE_wrapper_210__ap_start;
  wire PE_wrapper_210__ap_ready;
  wire PE_wrapper_210__ap_done;
  wire PE_wrapper_210__ap_idle;
  reg [1:0] PE_wrapper_210__state;
  wire PE_wrapper_211__ap_start_global__q0;
  wire PE_wrapper_211__is_done__q0;
  wire PE_wrapper_211__ap_done_global__q0;
  wire PE_wrapper_211__ap_start;
  wire PE_wrapper_211__ap_ready;
  wire PE_wrapper_211__ap_done;
  wire PE_wrapper_211__ap_idle;
  reg [1:0] PE_wrapper_211__state;
  wire PE_wrapper_212__ap_start_global__q0;
  wire PE_wrapper_212__is_done__q0;
  wire PE_wrapper_212__ap_done_global__q0;
  wire PE_wrapper_212__ap_start;
  wire PE_wrapper_212__ap_ready;
  wire PE_wrapper_212__ap_done;
  wire PE_wrapper_212__ap_idle;
  reg [1:0] PE_wrapper_212__state;
  wire PE_wrapper_213__ap_start_global__q0;
  wire PE_wrapper_213__is_done__q0;
  wire PE_wrapper_213__ap_done_global__q0;
  wire PE_wrapper_213__ap_start;
  wire PE_wrapper_213__ap_ready;
  wire PE_wrapper_213__ap_done;
  wire PE_wrapper_213__ap_idle;
  reg [1:0] PE_wrapper_213__state;
  wire PE_wrapper_214__ap_start_global__q0;
  wire PE_wrapper_214__is_done__q0;
  wire PE_wrapper_214__ap_done_global__q0;
  wire PE_wrapper_214__ap_start;
  wire PE_wrapper_214__ap_ready;
  wire PE_wrapper_214__ap_done;
  wire PE_wrapper_214__ap_idle;
  reg [1:0] PE_wrapper_214__state;
  wire PE_wrapper_215__ap_start_global__q0;
  wire PE_wrapper_215__is_done__q0;
  wire PE_wrapper_215__ap_done_global__q0;
  wire PE_wrapper_215__ap_start;
  wire PE_wrapper_215__ap_ready;
  wire PE_wrapper_215__ap_done;
  wire PE_wrapper_215__ap_idle;
  reg [1:0] PE_wrapper_215__state;
  wire PE_wrapper_216__ap_start_global__q0;
  wire PE_wrapper_216__is_done__q0;
  wire PE_wrapper_216__ap_done_global__q0;
  wire PE_wrapper_216__ap_start;
  wire PE_wrapper_216__ap_ready;
  wire PE_wrapper_216__ap_done;
  wire PE_wrapper_216__ap_idle;
  reg [1:0] PE_wrapper_216__state;
  wire PE_wrapper_217__ap_start_global__q0;
  wire PE_wrapper_217__is_done__q0;
  wire PE_wrapper_217__ap_done_global__q0;
  wire PE_wrapper_217__ap_start;
  wire PE_wrapper_217__ap_ready;
  wire PE_wrapper_217__ap_done;
  wire PE_wrapper_217__ap_idle;
  reg [1:0] PE_wrapper_217__state;
  wire PE_wrapper_218__ap_start_global__q0;
  wire PE_wrapper_218__is_done__q0;
  wire PE_wrapper_218__ap_done_global__q0;
  wire PE_wrapper_218__ap_start;
  wire PE_wrapper_218__ap_ready;
  wire PE_wrapper_218__ap_done;
  wire PE_wrapper_218__ap_idle;
  reg [1:0] PE_wrapper_218__state;
  wire PE_wrapper_219__ap_start_global__q0;
  wire PE_wrapper_219__is_done__q0;
  wire PE_wrapper_219__ap_done_global__q0;
  wire PE_wrapper_219__ap_start;
  wire PE_wrapper_219__ap_ready;
  wire PE_wrapper_219__ap_done;
  wire PE_wrapper_219__ap_idle;
  reg [1:0] PE_wrapper_219__state;
  wire PE_wrapper_220__ap_start_global__q0;
  wire PE_wrapper_220__is_done__q0;
  wire PE_wrapper_220__ap_done_global__q0;
  wire PE_wrapper_220__ap_start;
  wire PE_wrapper_220__ap_ready;
  wire PE_wrapper_220__ap_done;
  wire PE_wrapper_220__ap_idle;
  reg [1:0] PE_wrapper_220__state;
  wire PE_wrapper_221__ap_start_global__q0;
  wire PE_wrapper_221__is_done__q0;
  wire PE_wrapper_221__ap_done_global__q0;
  wire PE_wrapper_221__ap_start;
  wire PE_wrapper_221__ap_ready;
  wire PE_wrapper_221__ap_done;
  wire PE_wrapper_221__ap_idle;
  reg [1:0] PE_wrapper_221__state;
  wire PE_wrapper_222__ap_start_global__q0;
  wire PE_wrapper_222__is_done__q0;
  wire PE_wrapper_222__ap_done_global__q0;
  wire PE_wrapper_222__ap_start;
  wire PE_wrapper_222__ap_ready;
  wire PE_wrapper_222__ap_done;
  wire PE_wrapper_222__ap_idle;
  reg [1:0] PE_wrapper_222__state;
  wire PE_wrapper_223__ap_start_global__q0;
  wire PE_wrapper_223__is_done__q0;
  wire PE_wrapper_223__ap_done_global__q0;
  wire PE_wrapper_223__ap_start;
  wire PE_wrapper_223__ap_ready;
  wire PE_wrapper_223__ap_done;
  wire PE_wrapper_223__ap_idle;
  reg [1:0] PE_wrapper_223__state;
  wire PE_wrapper_224__ap_start_global__q0;
  wire PE_wrapper_224__is_done__q0;
  wire PE_wrapper_224__ap_done_global__q0;
  wire PE_wrapper_224__ap_start;
  wire PE_wrapper_224__ap_ready;
  wire PE_wrapper_224__ap_done;
  wire PE_wrapper_224__ap_idle;
  reg [1:0] PE_wrapper_224__state;
  wire PE_wrapper_225__ap_start_global__q0;
  wire PE_wrapper_225__is_done__q0;
  wire PE_wrapper_225__ap_done_global__q0;
  wire PE_wrapper_225__ap_start;
  wire PE_wrapper_225__ap_ready;
  wire PE_wrapper_225__ap_done;
  wire PE_wrapper_225__ap_idle;
  reg [1:0] PE_wrapper_225__state;
  wire PE_wrapper_226__ap_start_global__q0;
  wire PE_wrapper_226__is_done__q0;
  wire PE_wrapper_226__ap_done_global__q0;
  wire PE_wrapper_226__ap_start;
  wire PE_wrapper_226__ap_ready;
  wire PE_wrapper_226__ap_done;
  wire PE_wrapper_226__ap_idle;
  reg [1:0] PE_wrapper_226__state;
  wire PE_wrapper_227__ap_start_global__q0;
  wire PE_wrapper_227__is_done__q0;
  wire PE_wrapper_227__ap_done_global__q0;
  wire PE_wrapper_227__ap_start;
  wire PE_wrapper_227__ap_ready;
  wire PE_wrapper_227__ap_done;
  wire PE_wrapper_227__ap_idle;
  reg [1:0] PE_wrapper_227__state;
  wire PE_wrapper_228__ap_start_global__q0;
  wire PE_wrapper_228__is_done__q0;
  wire PE_wrapper_228__ap_done_global__q0;
  wire PE_wrapper_228__ap_start;
  wire PE_wrapper_228__ap_ready;
  wire PE_wrapper_228__ap_done;
  wire PE_wrapper_228__ap_idle;
  reg [1:0] PE_wrapper_228__state;
  wire PE_wrapper_229__ap_start_global__q0;
  wire PE_wrapper_229__is_done__q0;
  wire PE_wrapper_229__ap_done_global__q0;
  wire PE_wrapper_229__ap_start;
  wire PE_wrapper_229__ap_ready;
  wire PE_wrapper_229__ap_done;
  wire PE_wrapper_229__ap_idle;
  reg [1:0] PE_wrapper_229__state;
  wire PE_wrapper_230__ap_start_global__q0;
  wire PE_wrapper_230__is_done__q0;
  wire PE_wrapper_230__ap_done_global__q0;
  wire PE_wrapper_230__ap_start;
  wire PE_wrapper_230__ap_ready;
  wire PE_wrapper_230__ap_done;
  wire PE_wrapper_230__ap_idle;
  reg [1:0] PE_wrapper_230__state;
  wire PE_wrapper_231__ap_start_global__q0;
  wire PE_wrapper_231__is_done__q0;
  wire PE_wrapper_231__ap_done_global__q0;
  wire PE_wrapper_231__ap_start;
  wire PE_wrapper_231__ap_ready;
  wire PE_wrapper_231__ap_done;
  wire PE_wrapper_231__ap_idle;
  reg [1:0] PE_wrapper_231__state;
  wire PE_wrapper_232__ap_start_global__q0;
  wire PE_wrapper_232__is_done__q0;
  wire PE_wrapper_232__ap_done_global__q0;
  wire PE_wrapper_232__ap_start;
  wire PE_wrapper_232__ap_ready;
  wire PE_wrapper_232__ap_done;
  wire PE_wrapper_232__ap_idle;
  reg [1:0] PE_wrapper_232__state;
  wire PE_wrapper_233__ap_start_global__q0;
  wire PE_wrapper_233__is_done__q0;
  wire PE_wrapper_233__ap_done_global__q0;
  wire PE_wrapper_233__ap_start;
  wire PE_wrapper_233__ap_ready;
  wire PE_wrapper_233__ap_done;
  wire PE_wrapper_233__ap_idle;
  reg [1:0] PE_wrapper_233__state;
  wire PE_wrapper_234__ap_start_global__q0;
  wire PE_wrapper_234__is_done__q0;
  wire PE_wrapper_234__ap_done_global__q0;
  wire PE_wrapper_234__ap_start;
  wire PE_wrapper_234__ap_ready;
  wire PE_wrapper_234__ap_done;
  wire PE_wrapper_234__ap_idle;
  reg [1:0] PE_wrapper_234__state;
  wire PE_wrapper_235__ap_start_global__q0;
  wire PE_wrapper_235__is_done__q0;
  wire PE_wrapper_235__ap_done_global__q0;
  wire PE_wrapper_235__ap_start;
  wire PE_wrapper_235__ap_ready;
  wire PE_wrapper_235__ap_done;
  wire PE_wrapper_235__ap_idle;
  reg [1:0] PE_wrapper_235__state;
  wire PE_wrapper_236__ap_start_global__q0;
  wire PE_wrapper_236__is_done__q0;
  wire PE_wrapper_236__ap_done_global__q0;
  wire PE_wrapper_236__ap_start;
  wire PE_wrapper_236__ap_ready;
  wire PE_wrapper_236__ap_done;
  wire PE_wrapper_236__ap_idle;
  reg [1:0] PE_wrapper_236__state;
  wire PE_wrapper_237__ap_start_global__q0;
  wire PE_wrapper_237__is_done__q0;
  wire PE_wrapper_237__ap_done_global__q0;
  wire PE_wrapper_237__ap_start;
  wire PE_wrapper_237__ap_ready;
  wire PE_wrapper_237__ap_done;
  wire PE_wrapper_237__ap_idle;
  reg [1:0] PE_wrapper_237__state;
  wire PE_wrapper_238__ap_start_global__q0;
  wire PE_wrapper_238__is_done__q0;
  wire PE_wrapper_238__ap_done_global__q0;
  wire PE_wrapper_238__ap_start;
  wire PE_wrapper_238__ap_ready;
  wire PE_wrapper_238__ap_done;
  wire PE_wrapper_238__ap_idle;
  reg [1:0] PE_wrapper_238__state;
  wire PE_wrapper_239__ap_start_global__q0;
  wire PE_wrapper_239__is_done__q0;
  wire PE_wrapper_239__ap_done_global__q0;
  wire PE_wrapper_239__ap_start;
  wire PE_wrapper_239__ap_ready;
  wire PE_wrapper_239__ap_done;
  wire PE_wrapper_239__ap_idle;
  reg [1:0] PE_wrapper_239__state;
  wire PE_wrapper_240__ap_start_global__q0;
  wire PE_wrapper_240__is_done__q0;
  wire PE_wrapper_240__ap_done_global__q0;
  wire PE_wrapper_240__ap_start;
  wire PE_wrapper_240__ap_ready;
  wire PE_wrapper_240__ap_done;
  wire PE_wrapper_240__ap_idle;
  reg [1:0] PE_wrapper_240__state;
  wire PE_wrapper_241__ap_start_global__q0;
  wire PE_wrapper_241__is_done__q0;
  wire PE_wrapper_241__ap_done_global__q0;
  wire PE_wrapper_241__ap_start;
  wire PE_wrapper_241__ap_ready;
  wire PE_wrapper_241__ap_done;
  wire PE_wrapper_241__ap_idle;
  reg [1:0] PE_wrapper_241__state;
  wire PE_wrapper_242__ap_start_global__q0;
  wire PE_wrapper_242__is_done__q0;
  wire PE_wrapper_242__ap_done_global__q0;
  wire PE_wrapper_242__ap_start;
  wire PE_wrapper_242__ap_ready;
  wire PE_wrapper_242__ap_done;
  wire PE_wrapper_242__ap_idle;
  reg [1:0] PE_wrapper_242__state;
  wire PE_wrapper_243__ap_start_global__q0;
  wire PE_wrapper_243__is_done__q0;
  wire PE_wrapper_243__ap_done_global__q0;
  wire PE_wrapper_243__ap_start;
  wire PE_wrapper_243__ap_ready;
  wire PE_wrapper_243__ap_done;
  wire PE_wrapper_243__ap_idle;
  reg [1:0] PE_wrapper_243__state;
  wire PE_wrapper_244__ap_start_global__q0;
  wire PE_wrapper_244__is_done__q0;
  wire PE_wrapper_244__ap_done_global__q0;
  wire PE_wrapper_244__ap_start;
  wire PE_wrapper_244__ap_ready;
  wire PE_wrapper_244__ap_done;
  wire PE_wrapper_244__ap_idle;
  reg [1:0] PE_wrapper_244__state;
  wire PE_wrapper_245__ap_start_global__q0;
  wire PE_wrapper_245__is_done__q0;
  wire PE_wrapper_245__ap_done_global__q0;
  wire PE_wrapper_245__ap_start;
  wire PE_wrapper_245__ap_ready;
  wire PE_wrapper_245__ap_done;
  wire PE_wrapper_245__ap_idle;
  reg [1:0] PE_wrapper_245__state;
  wire PE_wrapper_246__ap_start_global__q0;
  wire PE_wrapper_246__is_done__q0;
  wire PE_wrapper_246__ap_done_global__q0;
  wire PE_wrapper_246__ap_start;
  wire PE_wrapper_246__ap_ready;
  wire PE_wrapper_246__ap_done;
  wire PE_wrapper_246__ap_idle;
  reg [1:0] PE_wrapper_246__state;
  wire PE_wrapper_247__ap_start_global__q0;
  wire PE_wrapper_247__is_done__q0;
  wire PE_wrapper_247__ap_done_global__q0;
  wire PE_wrapper_247__ap_start;
  wire PE_wrapper_247__ap_ready;
  wire PE_wrapper_247__ap_done;
  wire PE_wrapper_247__ap_idle;
  reg [1:0] PE_wrapper_247__state;
  wire PE_wrapper_248__ap_start_global__q0;
  wire PE_wrapper_248__is_done__q0;
  wire PE_wrapper_248__ap_done_global__q0;
  wire PE_wrapper_248__ap_start;
  wire PE_wrapper_248__ap_ready;
  wire PE_wrapper_248__ap_done;
  wire PE_wrapper_248__ap_idle;
  reg [1:0] PE_wrapper_248__state;
  wire PE_wrapper_249__ap_start_global__q0;
  wire PE_wrapper_249__is_done__q0;
  wire PE_wrapper_249__ap_done_global__q0;
  wire PE_wrapper_249__ap_start;
  wire PE_wrapper_249__ap_ready;
  wire PE_wrapper_249__ap_done;
  wire PE_wrapper_249__ap_idle;
  reg [1:0] PE_wrapper_249__state;
  wire PE_wrapper_250__ap_start_global__q0;
  wire PE_wrapper_250__is_done__q0;
  wire PE_wrapper_250__ap_done_global__q0;
  wire PE_wrapper_250__ap_start;
  wire PE_wrapper_250__ap_ready;
  wire PE_wrapper_250__ap_done;
  wire PE_wrapper_250__ap_idle;
  reg [1:0] PE_wrapper_250__state;
  wire PE_wrapper_251__ap_start_global__q0;
  wire PE_wrapper_251__is_done__q0;
  wire PE_wrapper_251__ap_done_global__q0;
  wire PE_wrapper_251__ap_start;
  wire PE_wrapper_251__ap_ready;
  wire PE_wrapper_251__ap_done;
  wire PE_wrapper_251__ap_idle;
  reg [1:0] PE_wrapper_251__state;
  wire PE_wrapper_252__ap_start_global__q0;
  wire PE_wrapper_252__is_done__q0;
  wire PE_wrapper_252__ap_done_global__q0;
  wire PE_wrapper_252__ap_start;
  wire PE_wrapper_252__ap_ready;
  wire PE_wrapper_252__ap_done;
  wire PE_wrapper_252__ap_idle;
  reg [1:0] PE_wrapper_252__state;
  wire PE_wrapper_253__ap_start_global__q0;
  wire PE_wrapper_253__is_done__q0;
  wire PE_wrapper_253__ap_done_global__q0;
  wire PE_wrapper_253__ap_start;
  wire PE_wrapper_253__ap_ready;
  wire PE_wrapper_253__ap_done;
  wire PE_wrapper_253__ap_idle;
  reg [1:0] PE_wrapper_253__state;
  wire PE_wrapper_254__ap_start_global__q0;
  wire PE_wrapper_254__is_done__q0;
  wire PE_wrapper_254__ap_done_global__q0;
  wire PE_wrapper_254__ap_start;
  wire PE_wrapper_254__ap_ready;
  wire PE_wrapper_254__ap_done;
  wire PE_wrapper_254__ap_idle;
  reg [1:0] PE_wrapper_254__state;
  wire PE_wrapper_255__ap_start_global__q0;
  wire PE_wrapper_255__is_done__q0;
  wire PE_wrapper_255__ap_done_global__q0;
  wire PE_wrapper_255__ap_start;
  wire PE_wrapper_255__ap_ready;
  wire PE_wrapper_255__ap_done;
  wire PE_wrapper_255__ap_idle;
  reg [1:0] PE_wrapper_255__state;
  wire PE_wrapper_256__ap_start_global__q0;
  wire PE_wrapper_256__is_done__q0;
  wire PE_wrapper_256__ap_done_global__q0;
  wire PE_wrapper_256__ap_start;
  wire PE_wrapper_256__ap_ready;
  wire PE_wrapper_256__ap_done;
  wire PE_wrapper_256__ap_idle;
  reg [1:0] PE_wrapper_256__state;
  wire PE_wrapper_257__ap_start_global__q0;
  wire PE_wrapper_257__is_done__q0;
  wire PE_wrapper_257__ap_done_global__q0;
  wire PE_wrapper_257__ap_start;
  wire PE_wrapper_257__ap_ready;
  wire PE_wrapper_257__ap_done;
  wire PE_wrapper_257__ap_idle;
  reg [1:0] PE_wrapper_257__state;
  wire PE_wrapper_258__ap_start_global__q0;
  wire PE_wrapper_258__is_done__q0;
  wire PE_wrapper_258__ap_done_global__q0;
  wire PE_wrapper_258__ap_start;
  wire PE_wrapper_258__ap_ready;
  wire PE_wrapper_258__ap_done;
  wire PE_wrapper_258__ap_idle;
  reg [1:0] PE_wrapper_258__state;
  wire PE_wrapper_259__ap_start_global__q0;
  wire PE_wrapper_259__is_done__q0;
  wire PE_wrapper_259__ap_done_global__q0;
  wire PE_wrapper_259__ap_start;
  wire PE_wrapper_259__ap_ready;
  wire PE_wrapper_259__ap_done;
  wire PE_wrapper_259__ap_idle;
  reg [1:0] PE_wrapper_259__state;
  wire PE_wrapper_260__ap_start_global__q0;
  wire PE_wrapper_260__is_done__q0;
  wire PE_wrapper_260__ap_done_global__q0;
  wire PE_wrapper_260__ap_start;
  wire PE_wrapper_260__ap_ready;
  wire PE_wrapper_260__ap_done;
  wire PE_wrapper_260__ap_idle;
  reg [1:0] PE_wrapper_260__state;
  wire PE_wrapper_261__ap_start_global__q0;
  wire PE_wrapper_261__is_done__q0;
  wire PE_wrapper_261__ap_done_global__q0;
  wire PE_wrapper_261__ap_start;
  wire PE_wrapper_261__ap_ready;
  wire PE_wrapper_261__ap_done;
  wire PE_wrapper_261__ap_idle;
  reg [1:0] PE_wrapper_261__state;
  wire PE_wrapper_262__ap_start_global__q0;
  wire PE_wrapper_262__is_done__q0;
  wire PE_wrapper_262__ap_done_global__q0;
  wire PE_wrapper_262__ap_start;
  wire PE_wrapper_262__ap_ready;
  wire PE_wrapper_262__ap_done;
  wire PE_wrapper_262__ap_idle;
  reg [1:0] PE_wrapper_262__state;
  wire PE_wrapper_263__ap_start_global__q0;
  wire PE_wrapper_263__is_done__q0;
  wire PE_wrapper_263__ap_done_global__q0;
  wire PE_wrapper_263__ap_start;
  wire PE_wrapper_263__ap_ready;
  wire PE_wrapper_263__ap_done;
  wire PE_wrapper_263__ap_idle;
  reg [1:0] PE_wrapper_263__state;
  wire PE_wrapper_264__ap_start_global__q0;
  wire PE_wrapper_264__is_done__q0;
  wire PE_wrapper_264__ap_done_global__q0;
  wire PE_wrapper_264__ap_start;
  wire PE_wrapper_264__ap_ready;
  wire PE_wrapper_264__ap_done;
  wire PE_wrapper_264__ap_idle;
  reg [1:0] PE_wrapper_264__state;
  wire PE_wrapper_265__ap_start_global__q0;
  wire PE_wrapper_265__is_done__q0;
  wire PE_wrapper_265__ap_done_global__q0;
  wire PE_wrapper_265__ap_start;
  wire PE_wrapper_265__ap_ready;
  wire PE_wrapper_265__ap_done;
  wire PE_wrapper_265__ap_idle;
  reg [1:0] PE_wrapper_265__state;
  wire PE_wrapper_266__ap_start_global__q0;
  wire PE_wrapper_266__is_done__q0;
  wire PE_wrapper_266__ap_done_global__q0;
  wire PE_wrapper_266__ap_start;
  wire PE_wrapper_266__ap_ready;
  wire PE_wrapper_266__ap_done;
  wire PE_wrapper_266__ap_idle;
  reg [1:0] PE_wrapper_266__state;
  wire PE_wrapper_267__ap_start_global__q0;
  wire PE_wrapper_267__is_done__q0;
  wire PE_wrapper_267__ap_done_global__q0;
  wire PE_wrapper_267__ap_start;
  wire PE_wrapper_267__ap_ready;
  wire PE_wrapper_267__ap_done;
  wire PE_wrapper_267__ap_idle;
  reg [1:0] PE_wrapper_267__state;
  wire PE_wrapper_268__ap_start_global__q0;
  wire PE_wrapper_268__is_done__q0;
  wire PE_wrapper_268__ap_done_global__q0;
  wire PE_wrapper_268__ap_start;
  wire PE_wrapper_268__ap_ready;
  wire PE_wrapper_268__ap_done;
  wire PE_wrapper_268__ap_idle;
  reg [1:0] PE_wrapper_268__state;
  wire PE_wrapper_269__ap_start_global__q0;
  wire PE_wrapper_269__is_done__q0;
  wire PE_wrapper_269__ap_done_global__q0;
  wire PE_wrapper_269__ap_start;
  wire PE_wrapper_269__ap_ready;
  wire PE_wrapper_269__ap_done;
  wire PE_wrapper_269__ap_idle;
  reg [1:0] PE_wrapper_269__state;
  wire PE_wrapper_270__ap_start_global__q0;
  wire PE_wrapper_270__is_done__q0;
  wire PE_wrapper_270__ap_done_global__q0;
  wire PE_wrapper_270__ap_start;
  wire PE_wrapper_270__ap_ready;
  wire PE_wrapper_270__ap_done;
  wire PE_wrapper_270__ap_idle;
  reg [1:0] PE_wrapper_270__state;
  wire PE_wrapper_271__ap_start_global__q0;
  wire PE_wrapper_271__is_done__q0;
  wire PE_wrapper_271__ap_done_global__q0;
  wire PE_wrapper_271__ap_start;
  wire PE_wrapper_271__ap_ready;
  wire PE_wrapper_271__ap_done;
  wire PE_wrapper_271__ap_idle;
  reg [1:0] PE_wrapper_271__state;
  wire PE_wrapper_272__ap_start_global__q0;
  wire PE_wrapper_272__is_done__q0;
  wire PE_wrapper_272__ap_done_global__q0;
  wire PE_wrapper_272__ap_start;
  wire PE_wrapper_272__ap_ready;
  wire PE_wrapper_272__ap_done;
  wire PE_wrapper_272__ap_idle;
  reg [1:0] PE_wrapper_272__state;
  wire PE_wrapper_273__ap_start_global__q0;
  wire PE_wrapper_273__is_done__q0;
  wire PE_wrapper_273__ap_done_global__q0;
  wire PE_wrapper_273__ap_start;
  wire PE_wrapper_273__ap_ready;
  wire PE_wrapper_273__ap_done;
  wire PE_wrapper_273__ap_idle;
  reg [1:0] PE_wrapper_273__state;
  wire PE_wrapper_274__ap_start_global__q0;
  wire PE_wrapper_274__is_done__q0;
  wire PE_wrapper_274__ap_done_global__q0;
  wire PE_wrapper_274__ap_start;
  wire PE_wrapper_274__ap_ready;
  wire PE_wrapper_274__ap_done;
  wire PE_wrapper_274__ap_idle;
  reg [1:0] PE_wrapper_274__state;
  wire PE_wrapper_275__ap_start_global__q0;
  wire PE_wrapper_275__is_done__q0;
  wire PE_wrapper_275__ap_done_global__q0;
  wire PE_wrapper_275__ap_start;
  wire PE_wrapper_275__ap_ready;
  wire PE_wrapper_275__ap_done;
  wire PE_wrapper_275__ap_idle;
  reg [1:0] PE_wrapper_275__state;
  wire PE_wrapper_276__ap_start_global__q0;
  wire PE_wrapper_276__is_done__q0;
  wire PE_wrapper_276__ap_done_global__q0;
  wire PE_wrapper_276__ap_start;
  wire PE_wrapper_276__ap_ready;
  wire PE_wrapper_276__ap_done;
  wire PE_wrapper_276__ap_idle;
  reg [1:0] PE_wrapper_276__state;
  wire PE_wrapper_277__ap_start_global__q0;
  wire PE_wrapper_277__is_done__q0;
  wire PE_wrapper_277__ap_done_global__q0;
  wire PE_wrapper_277__ap_start;
  wire PE_wrapper_277__ap_ready;
  wire PE_wrapper_277__ap_done;
  wire PE_wrapper_277__ap_idle;
  reg [1:0] PE_wrapper_277__state;
  wire PE_wrapper_278__ap_start_global__q0;
  wire PE_wrapper_278__is_done__q0;
  wire PE_wrapper_278__ap_done_global__q0;
  wire PE_wrapper_278__ap_start;
  wire PE_wrapper_278__ap_ready;
  wire PE_wrapper_278__ap_done;
  wire PE_wrapper_278__ap_idle;
  reg [1:0] PE_wrapper_278__state;
  wire PE_wrapper_279__ap_start_global__q0;
  wire PE_wrapper_279__is_done__q0;
  wire PE_wrapper_279__ap_done_global__q0;
  wire PE_wrapper_279__ap_start;
  wire PE_wrapper_279__ap_ready;
  wire PE_wrapper_279__ap_done;
  wire PE_wrapper_279__ap_idle;
  reg [1:0] PE_wrapper_279__state;
  wire PE_wrapper_280__ap_start_global__q0;
  wire PE_wrapper_280__is_done__q0;
  wire PE_wrapper_280__ap_done_global__q0;
  wire PE_wrapper_280__ap_start;
  wire PE_wrapper_280__ap_ready;
  wire PE_wrapper_280__ap_done;
  wire PE_wrapper_280__ap_idle;
  reg [1:0] PE_wrapper_280__state;
  wire PE_wrapper_281__ap_start_global__q0;
  wire PE_wrapper_281__is_done__q0;
  wire PE_wrapper_281__ap_done_global__q0;
  wire PE_wrapper_281__ap_start;
  wire PE_wrapper_281__ap_ready;
  wire PE_wrapper_281__ap_done;
  wire PE_wrapper_281__ap_idle;
  reg [1:0] PE_wrapper_281__state;
  wire PE_wrapper_282__ap_start_global__q0;
  wire PE_wrapper_282__is_done__q0;
  wire PE_wrapper_282__ap_done_global__q0;
  wire PE_wrapper_282__ap_start;
  wire PE_wrapper_282__ap_ready;
  wire PE_wrapper_282__ap_done;
  wire PE_wrapper_282__ap_idle;
  reg [1:0] PE_wrapper_282__state;
  wire PE_wrapper_283__ap_start_global__q0;
  wire PE_wrapper_283__is_done__q0;
  wire PE_wrapper_283__ap_done_global__q0;
  wire PE_wrapper_283__ap_start;
  wire PE_wrapper_283__ap_ready;
  wire PE_wrapper_283__ap_done;
  wire PE_wrapper_283__ap_idle;
  reg [1:0] PE_wrapper_283__state;
  wire PE_wrapper_284__ap_start_global__q0;
  wire PE_wrapper_284__is_done__q0;
  wire PE_wrapper_284__ap_done_global__q0;
  wire PE_wrapper_284__ap_start;
  wire PE_wrapper_284__ap_ready;
  wire PE_wrapper_284__ap_done;
  wire PE_wrapper_284__ap_idle;
  reg [1:0] PE_wrapper_284__state;
  wire PE_wrapper_285__ap_start_global__q0;
  wire PE_wrapper_285__is_done__q0;
  wire PE_wrapper_285__ap_done_global__q0;
  wire PE_wrapper_285__ap_start;
  wire PE_wrapper_285__ap_ready;
  wire PE_wrapper_285__ap_done;
  wire PE_wrapper_285__ap_idle;
  reg [1:0] PE_wrapper_285__state;
  wire PE_wrapper_286__ap_start_global__q0;
  wire PE_wrapper_286__is_done__q0;
  wire PE_wrapper_286__ap_done_global__q0;
  wire PE_wrapper_286__ap_start;
  wire PE_wrapper_286__ap_ready;
  wire PE_wrapper_286__ap_done;
  wire PE_wrapper_286__ap_idle;
  reg [1:0] PE_wrapper_286__state;
  wire PE_wrapper_287__ap_start_global__q0;
  wire PE_wrapper_287__is_done__q0;
  wire PE_wrapper_287__ap_done_global__q0;
  wire PE_wrapper_287__ap_start;
  wire PE_wrapper_287__ap_ready;
  wire PE_wrapper_287__ap_done;
  wire PE_wrapper_287__ap_idle;
  reg [1:0] PE_wrapper_287__state;
  wire PE_wrapper_288__ap_start_global__q0;
  wire PE_wrapper_288__is_done__q0;
  wire PE_wrapper_288__ap_done_global__q0;
  wire PE_wrapper_288__ap_start;
  wire PE_wrapper_288__ap_ready;
  wire PE_wrapper_288__ap_done;
  wire PE_wrapper_288__ap_idle;
  reg [1:0] PE_wrapper_288__state;
  wire PE_wrapper_289__ap_start_global__q0;
  wire PE_wrapper_289__is_done__q0;
  wire PE_wrapper_289__ap_done_global__q0;
  wire PE_wrapper_289__ap_start;
  wire PE_wrapper_289__ap_ready;
  wire PE_wrapper_289__ap_done;
  wire PE_wrapper_289__ap_idle;
  reg [1:0] PE_wrapper_289__state;
  wire PE_wrapper_290__ap_start_global__q0;
  wire PE_wrapper_290__is_done__q0;
  wire PE_wrapper_290__ap_done_global__q0;
  wire PE_wrapper_290__ap_start;
  wire PE_wrapper_290__ap_ready;
  wire PE_wrapper_290__ap_done;
  wire PE_wrapper_290__ap_idle;
  reg [1:0] PE_wrapper_290__state;
  wire PE_wrapper_291__ap_start_global__q0;
  wire PE_wrapper_291__is_done__q0;
  wire PE_wrapper_291__ap_done_global__q0;
  wire PE_wrapper_291__ap_start;
  wire PE_wrapper_291__ap_ready;
  wire PE_wrapper_291__ap_done;
  wire PE_wrapper_291__ap_idle;
  reg [1:0] PE_wrapper_291__state;
  wire PE_wrapper_292__ap_start_global__q0;
  wire PE_wrapper_292__is_done__q0;
  wire PE_wrapper_292__ap_done_global__q0;
  wire PE_wrapper_292__ap_start;
  wire PE_wrapper_292__ap_ready;
  wire PE_wrapper_292__ap_done;
  wire PE_wrapper_292__ap_idle;
  reg [1:0] PE_wrapper_292__state;
  wire PE_wrapper_293__ap_start_global__q0;
  wire PE_wrapper_293__is_done__q0;
  wire PE_wrapper_293__ap_done_global__q0;
  wire PE_wrapper_293__ap_start;
  wire PE_wrapper_293__ap_ready;
  wire PE_wrapper_293__ap_done;
  wire PE_wrapper_293__ap_idle;
  reg [1:0] PE_wrapper_293__state;
  wire PE_wrapper_294__ap_start_global__q0;
  wire PE_wrapper_294__is_done__q0;
  wire PE_wrapper_294__ap_done_global__q0;
  wire PE_wrapper_294__ap_start;
  wire PE_wrapper_294__ap_ready;
  wire PE_wrapper_294__ap_done;
  wire PE_wrapper_294__ap_idle;
  reg [1:0] PE_wrapper_294__state;
  wire PE_wrapper_295__ap_start_global__q0;
  wire PE_wrapper_295__is_done__q0;
  wire PE_wrapper_295__ap_done_global__q0;
  wire PE_wrapper_295__ap_start;
  wire PE_wrapper_295__ap_ready;
  wire PE_wrapper_295__ap_done;
  wire PE_wrapper_295__ap_idle;
  reg [1:0] PE_wrapper_295__state;
  wire PE_wrapper_296__ap_start_global__q0;
  wire PE_wrapper_296__is_done__q0;
  wire PE_wrapper_296__ap_done_global__q0;
  wire PE_wrapper_296__ap_start;
  wire PE_wrapper_296__ap_ready;
  wire PE_wrapper_296__ap_done;
  wire PE_wrapper_296__ap_idle;
  reg [1:0] PE_wrapper_296__state;
  wire PE_wrapper_297__ap_start_global__q0;
  wire PE_wrapper_297__is_done__q0;
  wire PE_wrapper_297__ap_done_global__q0;
  wire PE_wrapper_297__ap_start;
  wire PE_wrapper_297__ap_ready;
  wire PE_wrapper_297__ap_done;
  wire PE_wrapper_297__ap_idle;
  reg [1:0] PE_wrapper_297__state;
  wire PE_wrapper_298__ap_start_global__q0;
  wire PE_wrapper_298__is_done__q0;
  wire PE_wrapper_298__ap_done_global__q0;
  wire PE_wrapper_298__ap_start;
  wire PE_wrapper_298__ap_ready;
  wire PE_wrapper_298__ap_done;
  wire PE_wrapper_298__ap_idle;
  reg [1:0] PE_wrapper_298__state;
  wire PE_wrapper_299__ap_start_global__q0;
  wire PE_wrapper_299__is_done__q0;
  wire PE_wrapper_299__ap_done_global__q0;
  wire PE_wrapper_299__ap_start;
  wire PE_wrapper_299__ap_ready;
  wire PE_wrapper_299__ap_done;
  wire PE_wrapper_299__ap_idle;
  reg [1:0] PE_wrapper_299__state;
  wire PE_wrapper_300__ap_start_global__q0;
  wire PE_wrapper_300__is_done__q0;
  wire PE_wrapper_300__ap_done_global__q0;
  wire PE_wrapper_300__ap_start;
  wire PE_wrapper_300__ap_ready;
  wire PE_wrapper_300__ap_done;
  wire PE_wrapper_300__ap_idle;
  reg [1:0] PE_wrapper_300__state;
  wire PE_wrapper_301__ap_start_global__q0;
  wire PE_wrapper_301__is_done__q0;
  wire PE_wrapper_301__ap_done_global__q0;
  wire PE_wrapper_301__ap_start;
  wire PE_wrapper_301__ap_ready;
  wire PE_wrapper_301__ap_done;
  wire PE_wrapper_301__ap_idle;
  reg [1:0] PE_wrapper_301__state;
  wire PE_wrapper_302__ap_start_global__q0;
  wire PE_wrapper_302__is_done__q0;
  wire PE_wrapper_302__ap_done_global__q0;
  wire PE_wrapper_302__ap_start;
  wire PE_wrapper_302__ap_ready;
  wire PE_wrapper_302__ap_done;
  wire PE_wrapper_302__ap_idle;
  reg [1:0] PE_wrapper_302__state;
  wire PE_wrapper_303__ap_start_global__q0;
  wire PE_wrapper_303__is_done__q0;
  wire PE_wrapper_303__ap_done_global__q0;
  wire PE_wrapper_303__ap_start;
  wire PE_wrapper_303__ap_ready;
  wire PE_wrapper_303__ap_done;
  wire PE_wrapper_303__ap_idle;
  reg [1:0] PE_wrapper_303__state;
  wire PE_wrapper_304__ap_start_global__q0;
  wire PE_wrapper_304__is_done__q0;
  wire PE_wrapper_304__ap_done_global__q0;
  wire PE_wrapper_304__ap_start;
  wire PE_wrapper_304__ap_ready;
  wire PE_wrapper_304__ap_done;
  wire PE_wrapper_304__ap_idle;
  reg [1:0] PE_wrapper_304__state;
  wire PE_wrapper_305__ap_start_global__q0;
  wire PE_wrapper_305__is_done__q0;
  wire PE_wrapper_305__ap_done_global__q0;
  wire PE_wrapper_305__ap_start;
  wire PE_wrapper_305__ap_ready;
  wire PE_wrapper_305__ap_done;
  wire PE_wrapper_305__ap_idle;
  reg [1:0] PE_wrapper_305__state;
  reg [1:0] tapa_state;
  reg [0:0] countdown;
  wire ap_start__q0;
  wire ap_done__q0;
  assign A_IO_L2_in_0__ap_start_global__q0 = ap_start__q0;
  assign A_IO_L2_in_0__is_done__q0 = (A_IO_L2_in_0__state == 2'b10);
  assign A_IO_L2_in_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      A_IO_L2_in_0__state <= 2'b00;
    end else begin
      if(A_IO_L2_in_0__state == 2'b00) begin
        if(A_IO_L2_in_0__ap_start_global__q0) begin
          A_IO_L2_in_0__state <= 2'b01;
        end 
      end 
      if(A_IO_L2_in_0__state == 2'b01) begin
        if(A_IO_L2_in_0__ap_ready) begin
          if(A_IO_L2_in_0__ap_done) begin
            A_IO_L2_in_0__state <= 2'b10;
          end else begin
            A_IO_L2_in_0__state <= 2'b11;
          end
        end 
      end 
      if(A_IO_L2_in_0__state == 2'b11) begin
        if(A_IO_L2_in_0__ap_done) begin
          A_IO_L2_in_0__state <= 2'b10;
        end 
      end 
      if(A_IO_L2_in_0__state == 2'b10) begin
        if(A_IO_L2_in_0__ap_done_global__q0) begin
          A_IO_L2_in_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign A_IO_L2_in_0__ap_start = (A_IO_L2_in_0__state == 2'b01);
  assign A_IO_L2_in_1__ap_start_global__q0 = ap_start__q0;
  assign A_IO_L2_in_1__is_done__q0 = (A_IO_L2_in_1__state == 2'b10);
  assign A_IO_L2_in_1__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      A_IO_L2_in_1__state <= 2'b00;
    end else begin
      if(A_IO_L2_in_1__state == 2'b00) begin
        if(A_IO_L2_in_1__ap_start_global__q0) begin
          A_IO_L2_in_1__state <= 2'b01;
        end 
      end 
      if(A_IO_L2_in_1__state == 2'b01) begin
        if(A_IO_L2_in_1__ap_ready) begin
          if(A_IO_L2_in_1__ap_done) begin
            A_IO_L2_in_1__state <= 2'b10;
          end else begin
            A_IO_L2_in_1__state <= 2'b11;
          end
        end 
      end 
      if(A_IO_L2_in_1__state == 2'b11) begin
        if(A_IO_L2_in_1__ap_done) begin
          A_IO_L2_in_1__state <= 2'b10;
        end 
      end 
      if(A_IO_L2_in_1__state == 2'b10) begin
        if(A_IO_L2_in_1__ap_done_global__q0) begin
          A_IO_L2_in_1__state <= 2'b00;
        end 
      end 
    end
  end

  assign A_IO_L2_in_1__ap_start = (A_IO_L2_in_1__state == 2'b01);
  assign A_IO_L2_in_2__ap_start_global__q0 = ap_start__q0;
  assign A_IO_L2_in_2__is_done__q0 = (A_IO_L2_in_2__state == 2'b10);
  assign A_IO_L2_in_2__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      A_IO_L2_in_2__state <= 2'b00;
    end else begin
      if(A_IO_L2_in_2__state == 2'b00) begin
        if(A_IO_L2_in_2__ap_start_global__q0) begin
          A_IO_L2_in_2__state <= 2'b01;
        end 
      end 
      if(A_IO_L2_in_2__state == 2'b01) begin
        if(A_IO_L2_in_2__ap_ready) begin
          if(A_IO_L2_in_2__ap_done) begin
            A_IO_L2_in_2__state <= 2'b10;
          end else begin
            A_IO_L2_in_2__state <= 2'b11;
          end
        end 
      end 
      if(A_IO_L2_in_2__state == 2'b11) begin
        if(A_IO_L2_in_2__ap_done) begin
          A_IO_L2_in_2__state <= 2'b10;
        end 
      end 
      if(A_IO_L2_in_2__state == 2'b10) begin
        if(A_IO_L2_in_2__ap_done_global__q0) begin
          A_IO_L2_in_2__state <= 2'b00;
        end 
      end 
    end
  end

  assign A_IO_L2_in_2__ap_start = (A_IO_L2_in_2__state == 2'b01);
  assign A_IO_L2_in_3__ap_start_global__q0 = ap_start__q0;
  assign A_IO_L2_in_3__is_done__q0 = (A_IO_L2_in_3__state == 2'b10);
  assign A_IO_L2_in_3__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      A_IO_L2_in_3__state <= 2'b00;
    end else begin
      if(A_IO_L2_in_3__state == 2'b00) begin
        if(A_IO_L2_in_3__ap_start_global__q0) begin
          A_IO_L2_in_3__state <= 2'b01;
        end 
      end 
      if(A_IO_L2_in_3__state == 2'b01) begin
        if(A_IO_L2_in_3__ap_ready) begin
          if(A_IO_L2_in_3__ap_done) begin
            A_IO_L2_in_3__state <= 2'b10;
          end else begin
            A_IO_L2_in_3__state <= 2'b11;
          end
        end 
      end 
      if(A_IO_L2_in_3__state == 2'b11) begin
        if(A_IO_L2_in_3__ap_done) begin
          A_IO_L2_in_3__state <= 2'b10;
        end 
      end 
      if(A_IO_L2_in_3__state == 2'b10) begin
        if(A_IO_L2_in_3__ap_done_global__q0) begin
          A_IO_L2_in_3__state <= 2'b00;
        end 
      end 
    end
  end

  assign A_IO_L2_in_3__ap_start = (A_IO_L2_in_3__state == 2'b01);
  assign A_IO_L2_in_4__ap_start_global__q0 = ap_start__q0;
  assign A_IO_L2_in_4__is_done__q0 = (A_IO_L2_in_4__state == 2'b10);
  assign A_IO_L2_in_4__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      A_IO_L2_in_4__state <= 2'b00;
    end else begin
      if(A_IO_L2_in_4__state == 2'b00) begin
        if(A_IO_L2_in_4__ap_start_global__q0) begin
          A_IO_L2_in_4__state <= 2'b01;
        end 
      end 
      if(A_IO_L2_in_4__state == 2'b01) begin
        if(A_IO_L2_in_4__ap_ready) begin
          if(A_IO_L2_in_4__ap_done) begin
            A_IO_L2_in_4__state <= 2'b10;
          end else begin
            A_IO_L2_in_4__state <= 2'b11;
          end
        end 
      end 
      if(A_IO_L2_in_4__state == 2'b11) begin
        if(A_IO_L2_in_4__ap_done) begin
          A_IO_L2_in_4__state <= 2'b10;
        end 
      end 
      if(A_IO_L2_in_4__state == 2'b10) begin
        if(A_IO_L2_in_4__ap_done_global__q0) begin
          A_IO_L2_in_4__state <= 2'b00;
        end 
      end 
    end
  end

  assign A_IO_L2_in_4__ap_start = (A_IO_L2_in_4__state == 2'b01);
  assign A_IO_L2_in_5__ap_start_global__q0 = ap_start__q0;
  assign A_IO_L2_in_5__is_done__q0 = (A_IO_L2_in_5__state == 2'b10);
  assign A_IO_L2_in_5__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      A_IO_L2_in_5__state <= 2'b00;
    end else begin
      if(A_IO_L2_in_5__state == 2'b00) begin
        if(A_IO_L2_in_5__ap_start_global__q0) begin
          A_IO_L2_in_5__state <= 2'b01;
        end 
      end 
      if(A_IO_L2_in_5__state == 2'b01) begin
        if(A_IO_L2_in_5__ap_ready) begin
          if(A_IO_L2_in_5__ap_done) begin
            A_IO_L2_in_5__state <= 2'b10;
          end else begin
            A_IO_L2_in_5__state <= 2'b11;
          end
        end 
      end 
      if(A_IO_L2_in_5__state == 2'b11) begin
        if(A_IO_L2_in_5__ap_done) begin
          A_IO_L2_in_5__state <= 2'b10;
        end 
      end 
      if(A_IO_L2_in_5__state == 2'b10) begin
        if(A_IO_L2_in_5__ap_done_global__q0) begin
          A_IO_L2_in_5__state <= 2'b00;
        end 
      end 
    end
  end

  assign A_IO_L2_in_5__ap_start = (A_IO_L2_in_5__state == 2'b01);
  assign A_IO_L2_in_6__ap_start_global__q0 = ap_start__q0;
  assign A_IO_L2_in_6__is_done__q0 = (A_IO_L2_in_6__state == 2'b10);
  assign A_IO_L2_in_6__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      A_IO_L2_in_6__state <= 2'b00;
    end else begin
      if(A_IO_L2_in_6__state == 2'b00) begin
        if(A_IO_L2_in_6__ap_start_global__q0) begin
          A_IO_L2_in_6__state <= 2'b01;
        end 
      end 
      if(A_IO_L2_in_6__state == 2'b01) begin
        if(A_IO_L2_in_6__ap_ready) begin
          if(A_IO_L2_in_6__ap_done) begin
            A_IO_L2_in_6__state <= 2'b10;
          end else begin
            A_IO_L2_in_6__state <= 2'b11;
          end
        end 
      end 
      if(A_IO_L2_in_6__state == 2'b11) begin
        if(A_IO_L2_in_6__ap_done) begin
          A_IO_L2_in_6__state <= 2'b10;
        end 
      end 
      if(A_IO_L2_in_6__state == 2'b10) begin
        if(A_IO_L2_in_6__ap_done_global__q0) begin
          A_IO_L2_in_6__state <= 2'b00;
        end 
      end 
    end
  end

  assign A_IO_L2_in_6__ap_start = (A_IO_L2_in_6__state == 2'b01);
  assign A_IO_L2_in_7__ap_start_global__q0 = ap_start__q0;
  assign A_IO_L2_in_7__is_done__q0 = (A_IO_L2_in_7__state == 2'b10);
  assign A_IO_L2_in_7__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      A_IO_L2_in_7__state <= 2'b00;
    end else begin
      if(A_IO_L2_in_7__state == 2'b00) begin
        if(A_IO_L2_in_7__ap_start_global__q0) begin
          A_IO_L2_in_7__state <= 2'b01;
        end 
      end 
      if(A_IO_L2_in_7__state == 2'b01) begin
        if(A_IO_L2_in_7__ap_ready) begin
          if(A_IO_L2_in_7__ap_done) begin
            A_IO_L2_in_7__state <= 2'b10;
          end else begin
            A_IO_L2_in_7__state <= 2'b11;
          end
        end 
      end 
      if(A_IO_L2_in_7__state == 2'b11) begin
        if(A_IO_L2_in_7__ap_done) begin
          A_IO_L2_in_7__state <= 2'b10;
        end 
      end 
      if(A_IO_L2_in_7__state == 2'b10) begin
        if(A_IO_L2_in_7__ap_done_global__q0) begin
          A_IO_L2_in_7__state <= 2'b00;
        end 
      end 
    end
  end

  assign A_IO_L2_in_7__ap_start = (A_IO_L2_in_7__state == 2'b01);
  assign A_IO_L2_in_8__ap_start_global__q0 = ap_start__q0;
  assign A_IO_L2_in_8__is_done__q0 = (A_IO_L2_in_8__state == 2'b10);
  assign A_IO_L2_in_8__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      A_IO_L2_in_8__state <= 2'b00;
    end else begin
      if(A_IO_L2_in_8__state == 2'b00) begin
        if(A_IO_L2_in_8__ap_start_global__q0) begin
          A_IO_L2_in_8__state <= 2'b01;
        end 
      end 
      if(A_IO_L2_in_8__state == 2'b01) begin
        if(A_IO_L2_in_8__ap_ready) begin
          if(A_IO_L2_in_8__ap_done) begin
            A_IO_L2_in_8__state <= 2'b10;
          end else begin
            A_IO_L2_in_8__state <= 2'b11;
          end
        end 
      end 
      if(A_IO_L2_in_8__state == 2'b11) begin
        if(A_IO_L2_in_8__ap_done) begin
          A_IO_L2_in_8__state <= 2'b10;
        end 
      end 
      if(A_IO_L2_in_8__state == 2'b10) begin
        if(A_IO_L2_in_8__ap_done_global__q0) begin
          A_IO_L2_in_8__state <= 2'b00;
        end 
      end 
    end
  end

  assign A_IO_L2_in_8__ap_start = (A_IO_L2_in_8__state == 2'b01);
  assign A_IO_L2_in_9__ap_start_global__q0 = ap_start__q0;
  assign A_IO_L2_in_9__is_done__q0 = (A_IO_L2_in_9__state == 2'b10);
  assign A_IO_L2_in_9__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      A_IO_L2_in_9__state <= 2'b00;
    end else begin
      if(A_IO_L2_in_9__state == 2'b00) begin
        if(A_IO_L2_in_9__ap_start_global__q0) begin
          A_IO_L2_in_9__state <= 2'b01;
        end 
      end 
      if(A_IO_L2_in_9__state == 2'b01) begin
        if(A_IO_L2_in_9__ap_ready) begin
          if(A_IO_L2_in_9__ap_done) begin
            A_IO_L2_in_9__state <= 2'b10;
          end else begin
            A_IO_L2_in_9__state <= 2'b11;
          end
        end 
      end 
      if(A_IO_L2_in_9__state == 2'b11) begin
        if(A_IO_L2_in_9__ap_done) begin
          A_IO_L2_in_9__state <= 2'b10;
        end 
      end 
      if(A_IO_L2_in_9__state == 2'b10) begin
        if(A_IO_L2_in_9__ap_done_global__q0) begin
          A_IO_L2_in_9__state <= 2'b00;
        end 
      end 
    end
  end

  assign A_IO_L2_in_9__ap_start = (A_IO_L2_in_9__state == 2'b01);
  assign A_IO_L2_in_10__ap_start_global__q0 = ap_start__q0;
  assign A_IO_L2_in_10__is_done__q0 = (A_IO_L2_in_10__state == 2'b10);
  assign A_IO_L2_in_10__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      A_IO_L2_in_10__state <= 2'b00;
    end else begin
      if(A_IO_L2_in_10__state == 2'b00) begin
        if(A_IO_L2_in_10__ap_start_global__q0) begin
          A_IO_L2_in_10__state <= 2'b01;
        end 
      end 
      if(A_IO_L2_in_10__state == 2'b01) begin
        if(A_IO_L2_in_10__ap_ready) begin
          if(A_IO_L2_in_10__ap_done) begin
            A_IO_L2_in_10__state <= 2'b10;
          end else begin
            A_IO_L2_in_10__state <= 2'b11;
          end
        end 
      end 
      if(A_IO_L2_in_10__state == 2'b11) begin
        if(A_IO_L2_in_10__ap_done) begin
          A_IO_L2_in_10__state <= 2'b10;
        end 
      end 
      if(A_IO_L2_in_10__state == 2'b10) begin
        if(A_IO_L2_in_10__ap_done_global__q0) begin
          A_IO_L2_in_10__state <= 2'b00;
        end 
      end 
    end
  end

  assign A_IO_L2_in_10__ap_start = (A_IO_L2_in_10__state == 2'b01);
  assign A_IO_L2_in_11__ap_start_global__q0 = ap_start__q0;
  assign A_IO_L2_in_11__is_done__q0 = (A_IO_L2_in_11__state == 2'b10);
  assign A_IO_L2_in_11__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      A_IO_L2_in_11__state <= 2'b00;
    end else begin
      if(A_IO_L2_in_11__state == 2'b00) begin
        if(A_IO_L2_in_11__ap_start_global__q0) begin
          A_IO_L2_in_11__state <= 2'b01;
        end 
      end 
      if(A_IO_L2_in_11__state == 2'b01) begin
        if(A_IO_L2_in_11__ap_ready) begin
          if(A_IO_L2_in_11__ap_done) begin
            A_IO_L2_in_11__state <= 2'b10;
          end else begin
            A_IO_L2_in_11__state <= 2'b11;
          end
        end 
      end 
      if(A_IO_L2_in_11__state == 2'b11) begin
        if(A_IO_L2_in_11__ap_done) begin
          A_IO_L2_in_11__state <= 2'b10;
        end 
      end 
      if(A_IO_L2_in_11__state == 2'b10) begin
        if(A_IO_L2_in_11__ap_done_global__q0) begin
          A_IO_L2_in_11__state <= 2'b00;
        end 
      end 
    end
  end

  assign A_IO_L2_in_11__ap_start = (A_IO_L2_in_11__state == 2'b01);
  assign A_IO_L2_in_12__ap_start_global__q0 = ap_start__q0;
  assign A_IO_L2_in_12__is_done__q0 = (A_IO_L2_in_12__state == 2'b10);
  assign A_IO_L2_in_12__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      A_IO_L2_in_12__state <= 2'b00;
    end else begin
      if(A_IO_L2_in_12__state == 2'b00) begin
        if(A_IO_L2_in_12__ap_start_global__q0) begin
          A_IO_L2_in_12__state <= 2'b01;
        end 
      end 
      if(A_IO_L2_in_12__state == 2'b01) begin
        if(A_IO_L2_in_12__ap_ready) begin
          if(A_IO_L2_in_12__ap_done) begin
            A_IO_L2_in_12__state <= 2'b10;
          end else begin
            A_IO_L2_in_12__state <= 2'b11;
          end
        end 
      end 
      if(A_IO_L2_in_12__state == 2'b11) begin
        if(A_IO_L2_in_12__ap_done) begin
          A_IO_L2_in_12__state <= 2'b10;
        end 
      end 
      if(A_IO_L2_in_12__state == 2'b10) begin
        if(A_IO_L2_in_12__ap_done_global__q0) begin
          A_IO_L2_in_12__state <= 2'b00;
        end 
      end 
    end
  end

  assign A_IO_L2_in_12__ap_start = (A_IO_L2_in_12__state == 2'b01);
  assign A_IO_L2_in_13__ap_start_global__q0 = ap_start__q0;
  assign A_IO_L2_in_13__is_done__q0 = (A_IO_L2_in_13__state == 2'b10);
  assign A_IO_L2_in_13__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      A_IO_L2_in_13__state <= 2'b00;
    end else begin
      if(A_IO_L2_in_13__state == 2'b00) begin
        if(A_IO_L2_in_13__ap_start_global__q0) begin
          A_IO_L2_in_13__state <= 2'b01;
        end 
      end 
      if(A_IO_L2_in_13__state == 2'b01) begin
        if(A_IO_L2_in_13__ap_ready) begin
          if(A_IO_L2_in_13__ap_done) begin
            A_IO_L2_in_13__state <= 2'b10;
          end else begin
            A_IO_L2_in_13__state <= 2'b11;
          end
        end 
      end 
      if(A_IO_L2_in_13__state == 2'b11) begin
        if(A_IO_L2_in_13__ap_done) begin
          A_IO_L2_in_13__state <= 2'b10;
        end 
      end 
      if(A_IO_L2_in_13__state == 2'b10) begin
        if(A_IO_L2_in_13__ap_done_global__q0) begin
          A_IO_L2_in_13__state <= 2'b00;
        end 
      end 
    end
  end

  assign A_IO_L2_in_13__ap_start = (A_IO_L2_in_13__state == 2'b01);
  assign A_IO_L2_in_14__ap_start_global__q0 = ap_start__q0;
  assign A_IO_L2_in_14__is_done__q0 = (A_IO_L2_in_14__state == 2'b10);
  assign A_IO_L2_in_14__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      A_IO_L2_in_14__state <= 2'b00;
    end else begin
      if(A_IO_L2_in_14__state == 2'b00) begin
        if(A_IO_L2_in_14__ap_start_global__q0) begin
          A_IO_L2_in_14__state <= 2'b01;
        end 
      end 
      if(A_IO_L2_in_14__state == 2'b01) begin
        if(A_IO_L2_in_14__ap_ready) begin
          if(A_IO_L2_in_14__ap_done) begin
            A_IO_L2_in_14__state <= 2'b10;
          end else begin
            A_IO_L2_in_14__state <= 2'b11;
          end
        end 
      end 
      if(A_IO_L2_in_14__state == 2'b11) begin
        if(A_IO_L2_in_14__ap_done) begin
          A_IO_L2_in_14__state <= 2'b10;
        end 
      end 
      if(A_IO_L2_in_14__state == 2'b10) begin
        if(A_IO_L2_in_14__ap_done_global__q0) begin
          A_IO_L2_in_14__state <= 2'b00;
        end 
      end 
    end
  end

  assign A_IO_L2_in_14__ap_start = (A_IO_L2_in_14__state == 2'b01);
  assign A_IO_L2_in_15__ap_start_global__q0 = ap_start__q0;
  assign A_IO_L2_in_15__is_done__q0 = (A_IO_L2_in_15__state == 2'b10);
  assign A_IO_L2_in_15__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      A_IO_L2_in_15__state <= 2'b00;
    end else begin
      if(A_IO_L2_in_15__state == 2'b00) begin
        if(A_IO_L2_in_15__ap_start_global__q0) begin
          A_IO_L2_in_15__state <= 2'b01;
        end 
      end 
      if(A_IO_L2_in_15__state == 2'b01) begin
        if(A_IO_L2_in_15__ap_ready) begin
          if(A_IO_L2_in_15__ap_done) begin
            A_IO_L2_in_15__state <= 2'b10;
          end else begin
            A_IO_L2_in_15__state <= 2'b11;
          end
        end 
      end 
      if(A_IO_L2_in_15__state == 2'b11) begin
        if(A_IO_L2_in_15__ap_done) begin
          A_IO_L2_in_15__state <= 2'b10;
        end 
      end 
      if(A_IO_L2_in_15__state == 2'b10) begin
        if(A_IO_L2_in_15__ap_done_global__q0) begin
          A_IO_L2_in_15__state <= 2'b00;
        end 
      end 
    end
  end

  assign A_IO_L2_in_15__ap_start = (A_IO_L2_in_15__state == 2'b01);
  assign A_IO_L2_in_16__ap_start_global__q0 = ap_start__q0;
  assign A_IO_L2_in_16__is_done__q0 = (A_IO_L2_in_16__state == 2'b10);
  assign A_IO_L2_in_16__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      A_IO_L2_in_16__state <= 2'b00;
    end else begin
      if(A_IO_L2_in_16__state == 2'b00) begin
        if(A_IO_L2_in_16__ap_start_global__q0) begin
          A_IO_L2_in_16__state <= 2'b01;
        end 
      end 
      if(A_IO_L2_in_16__state == 2'b01) begin
        if(A_IO_L2_in_16__ap_ready) begin
          if(A_IO_L2_in_16__ap_done) begin
            A_IO_L2_in_16__state <= 2'b10;
          end else begin
            A_IO_L2_in_16__state <= 2'b11;
          end
        end 
      end 
      if(A_IO_L2_in_16__state == 2'b11) begin
        if(A_IO_L2_in_16__ap_done) begin
          A_IO_L2_in_16__state <= 2'b10;
        end 
      end 
      if(A_IO_L2_in_16__state == 2'b10) begin
        if(A_IO_L2_in_16__ap_done_global__q0) begin
          A_IO_L2_in_16__state <= 2'b00;
        end 
      end 
    end
  end

  assign A_IO_L2_in_16__ap_start = (A_IO_L2_in_16__state == 2'b01);
  assign A_IO_L2_in_boundary_0__ap_start_global__q0 = ap_start__q0;
  assign A_IO_L2_in_boundary_0__is_done__q0 = (A_IO_L2_in_boundary_0__state == 2'b10);
  assign A_IO_L2_in_boundary_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      A_IO_L2_in_boundary_0__state <= 2'b00;
    end else begin
      if(A_IO_L2_in_boundary_0__state == 2'b00) begin
        if(A_IO_L2_in_boundary_0__ap_start_global__q0) begin
          A_IO_L2_in_boundary_0__state <= 2'b01;
        end 
      end 
      if(A_IO_L2_in_boundary_0__state == 2'b01) begin
        if(A_IO_L2_in_boundary_0__ap_ready) begin
          if(A_IO_L2_in_boundary_0__ap_done) begin
            A_IO_L2_in_boundary_0__state <= 2'b10;
          end else begin
            A_IO_L2_in_boundary_0__state <= 2'b11;
          end
        end 
      end 
      if(A_IO_L2_in_boundary_0__state == 2'b11) begin
        if(A_IO_L2_in_boundary_0__ap_done) begin
          A_IO_L2_in_boundary_0__state <= 2'b10;
        end 
      end 
      if(A_IO_L2_in_boundary_0__state == 2'b10) begin
        if(A_IO_L2_in_boundary_0__ap_done_global__q0) begin
          A_IO_L2_in_boundary_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign A_IO_L2_in_boundary_0__ap_start = (A_IO_L2_in_boundary_0__state == 2'b01);
  assign A_IO_L3_in_0__ap_start_global__q0 = ap_start__q0;
  assign A_IO_L3_in_0__is_done__q0 = (A_IO_L3_in_0__state == 2'b10);
  assign A_IO_L3_in_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      A_IO_L3_in_0__state <= 2'b00;
    end else begin
      if(A_IO_L3_in_0__state == 2'b00) begin
        if(A_IO_L3_in_0__ap_start_global__q0) begin
          A_IO_L3_in_0__state <= 2'b01;
        end 
      end 
      if(A_IO_L3_in_0__state == 2'b01) begin
        if(A_IO_L3_in_0__ap_ready) begin
          if(A_IO_L3_in_0__ap_done) begin
            A_IO_L3_in_0__state <= 2'b10;
          end else begin
            A_IO_L3_in_0__state <= 2'b11;
          end
        end 
      end 
      if(A_IO_L3_in_0__state == 2'b11) begin
        if(A_IO_L3_in_0__ap_done) begin
          A_IO_L3_in_0__state <= 2'b10;
        end 
      end 
      if(A_IO_L3_in_0__state == 2'b10) begin
        if(A_IO_L3_in_0__ap_done_global__q0) begin
          A_IO_L3_in_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign A_IO_L3_in_0__ap_start = (A_IO_L3_in_0__state == 2'b01);
  assign A_IO_L3_in_serialize_0___A__q0 = A;
  assign A_IO_L3_in_serialize_0__ap_start_global__q0 = ap_start__q0;
  assign A_IO_L3_in_serialize_0__is_done__q0 = (A_IO_L3_in_serialize_0__state == 2'b10);
  assign A_IO_L3_in_serialize_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      A_IO_L3_in_serialize_0__state <= 2'b00;
    end else begin
      if(A_IO_L3_in_serialize_0__state == 2'b00) begin
        if(A_IO_L3_in_serialize_0__ap_start_global__q0) begin
          A_IO_L3_in_serialize_0__state <= 2'b01;
        end 
      end 
      if(A_IO_L3_in_serialize_0__state == 2'b01) begin
        if(A_IO_L3_in_serialize_0__ap_ready) begin
          if(A_IO_L3_in_serialize_0__ap_done) begin
            A_IO_L3_in_serialize_0__state <= 2'b10;
          end else begin
            A_IO_L3_in_serialize_0__state <= 2'b11;
          end
        end 
      end 
      if(A_IO_L3_in_serialize_0__state == 2'b11) begin
        if(A_IO_L3_in_serialize_0__ap_done) begin
          A_IO_L3_in_serialize_0__state <= 2'b10;
        end 
      end 
      if(A_IO_L3_in_serialize_0__state == 2'b10) begin
        if(A_IO_L3_in_serialize_0__ap_done_global__q0) begin
          A_IO_L3_in_serialize_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign A_IO_L3_in_serialize_0__ap_start = (A_IO_L3_in_serialize_0__state == 2'b01);
  assign A_PE_dummy_in_0__ap_start_global__q0 = ap_start__q0;
  assign A_PE_dummy_in_0__is_done__q0 = (A_PE_dummy_in_0__state == 2'b10);
  assign A_PE_dummy_in_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      A_PE_dummy_in_0__state <= 2'b00;
    end else begin
      if(A_PE_dummy_in_0__state == 2'b00) begin
        if(A_PE_dummy_in_0__ap_start_global__q0) begin
          A_PE_dummy_in_0__state <= 2'b01;
        end 
      end 
      if(A_PE_dummy_in_0__state == 2'b01) begin
        if(A_PE_dummy_in_0__ap_ready) begin
          if(A_PE_dummy_in_0__ap_done) begin
            A_PE_dummy_in_0__state <= 2'b10;
          end else begin
            A_PE_dummy_in_0__state <= 2'b11;
          end
        end 
      end 
      if(A_PE_dummy_in_0__state == 2'b11) begin
        if(A_PE_dummy_in_0__ap_done) begin
          A_PE_dummy_in_0__state <= 2'b10;
        end 
      end 
      if(A_PE_dummy_in_0__state == 2'b10) begin
        if(A_PE_dummy_in_0__ap_done_global__q0) begin
          A_PE_dummy_in_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign A_PE_dummy_in_0__ap_start = (A_PE_dummy_in_0__state == 2'b01);
  assign A_PE_dummy_in_1__ap_start_global__q0 = ap_start__q0;
  assign A_PE_dummy_in_1__is_done__q0 = (A_PE_dummy_in_1__state == 2'b10);
  assign A_PE_dummy_in_1__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      A_PE_dummy_in_1__state <= 2'b00;
    end else begin
      if(A_PE_dummy_in_1__state == 2'b00) begin
        if(A_PE_dummy_in_1__ap_start_global__q0) begin
          A_PE_dummy_in_1__state <= 2'b01;
        end 
      end 
      if(A_PE_dummy_in_1__state == 2'b01) begin
        if(A_PE_dummy_in_1__ap_ready) begin
          if(A_PE_dummy_in_1__ap_done) begin
            A_PE_dummy_in_1__state <= 2'b10;
          end else begin
            A_PE_dummy_in_1__state <= 2'b11;
          end
        end 
      end 
      if(A_PE_dummy_in_1__state == 2'b11) begin
        if(A_PE_dummy_in_1__ap_done) begin
          A_PE_dummy_in_1__state <= 2'b10;
        end 
      end 
      if(A_PE_dummy_in_1__state == 2'b10) begin
        if(A_PE_dummy_in_1__ap_done_global__q0) begin
          A_PE_dummy_in_1__state <= 2'b00;
        end 
      end 
    end
  end

  assign A_PE_dummy_in_1__ap_start = (A_PE_dummy_in_1__state == 2'b01);
  assign A_PE_dummy_in_2__ap_start_global__q0 = ap_start__q0;
  assign A_PE_dummy_in_2__is_done__q0 = (A_PE_dummy_in_2__state == 2'b10);
  assign A_PE_dummy_in_2__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      A_PE_dummy_in_2__state <= 2'b00;
    end else begin
      if(A_PE_dummy_in_2__state == 2'b00) begin
        if(A_PE_dummy_in_2__ap_start_global__q0) begin
          A_PE_dummy_in_2__state <= 2'b01;
        end 
      end 
      if(A_PE_dummy_in_2__state == 2'b01) begin
        if(A_PE_dummy_in_2__ap_ready) begin
          if(A_PE_dummy_in_2__ap_done) begin
            A_PE_dummy_in_2__state <= 2'b10;
          end else begin
            A_PE_dummy_in_2__state <= 2'b11;
          end
        end 
      end 
      if(A_PE_dummy_in_2__state == 2'b11) begin
        if(A_PE_dummy_in_2__ap_done) begin
          A_PE_dummy_in_2__state <= 2'b10;
        end 
      end 
      if(A_PE_dummy_in_2__state == 2'b10) begin
        if(A_PE_dummy_in_2__ap_done_global__q0) begin
          A_PE_dummy_in_2__state <= 2'b00;
        end 
      end 
    end
  end

  assign A_PE_dummy_in_2__ap_start = (A_PE_dummy_in_2__state == 2'b01);
  assign A_PE_dummy_in_3__ap_start_global__q0 = ap_start__q0;
  assign A_PE_dummy_in_3__is_done__q0 = (A_PE_dummy_in_3__state == 2'b10);
  assign A_PE_dummy_in_3__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      A_PE_dummy_in_3__state <= 2'b00;
    end else begin
      if(A_PE_dummy_in_3__state == 2'b00) begin
        if(A_PE_dummy_in_3__ap_start_global__q0) begin
          A_PE_dummy_in_3__state <= 2'b01;
        end 
      end 
      if(A_PE_dummy_in_3__state == 2'b01) begin
        if(A_PE_dummy_in_3__ap_ready) begin
          if(A_PE_dummy_in_3__ap_done) begin
            A_PE_dummy_in_3__state <= 2'b10;
          end else begin
            A_PE_dummy_in_3__state <= 2'b11;
          end
        end 
      end 
      if(A_PE_dummy_in_3__state == 2'b11) begin
        if(A_PE_dummy_in_3__ap_done) begin
          A_PE_dummy_in_3__state <= 2'b10;
        end 
      end 
      if(A_PE_dummy_in_3__state == 2'b10) begin
        if(A_PE_dummy_in_3__ap_done_global__q0) begin
          A_PE_dummy_in_3__state <= 2'b00;
        end 
      end 
    end
  end

  assign A_PE_dummy_in_3__ap_start = (A_PE_dummy_in_3__state == 2'b01);
  assign A_PE_dummy_in_4__ap_start_global__q0 = ap_start__q0;
  assign A_PE_dummy_in_4__is_done__q0 = (A_PE_dummy_in_4__state == 2'b10);
  assign A_PE_dummy_in_4__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      A_PE_dummy_in_4__state <= 2'b00;
    end else begin
      if(A_PE_dummy_in_4__state == 2'b00) begin
        if(A_PE_dummy_in_4__ap_start_global__q0) begin
          A_PE_dummy_in_4__state <= 2'b01;
        end 
      end 
      if(A_PE_dummy_in_4__state == 2'b01) begin
        if(A_PE_dummy_in_4__ap_ready) begin
          if(A_PE_dummy_in_4__ap_done) begin
            A_PE_dummy_in_4__state <= 2'b10;
          end else begin
            A_PE_dummy_in_4__state <= 2'b11;
          end
        end 
      end 
      if(A_PE_dummy_in_4__state == 2'b11) begin
        if(A_PE_dummy_in_4__ap_done) begin
          A_PE_dummy_in_4__state <= 2'b10;
        end 
      end 
      if(A_PE_dummy_in_4__state == 2'b10) begin
        if(A_PE_dummy_in_4__ap_done_global__q0) begin
          A_PE_dummy_in_4__state <= 2'b00;
        end 
      end 
    end
  end

  assign A_PE_dummy_in_4__ap_start = (A_PE_dummy_in_4__state == 2'b01);
  assign A_PE_dummy_in_5__ap_start_global__q0 = ap_start__q0;
  assign A_PE_dummy_in_5__is_done__q0 = (A_PE_dummy_in_5__state == 2'b10);
  assign A_PE_dummy_in_5__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      A_PE_dummy_in_5__state <= 2'b00;
    end else begin
      if(A_PE_dummy_in_5__state == 2'b00) begin
        if(A_PE_dummy_in_5__ap_start_global__q0) begin
          A_PE_dummy_in_5__state <= 2'b01;
        end 
      end 
      if(A_PE_dummy_in_5__state == 2'b01) begin
        if(A_PE_dummy_in_5__ap_ready) begin
          if(A_PE_dummy_in_5__ap_done) begin
            A_PE_dummy_in_5__state <= 2'b10;
          end else begin
            A_PE_dummy_in_5__state <= 2'b11;
          end
        end 
      end 
      if(A_PE_dummy_in_5__state == 2'b11) begin
        if(A_PE_dummy_in_5__ap_done) begin
          A_PE_dummy_in_5__state <= 2'b10;
        end 
      end 
      if(A_PE_dummy_in_5__state == 2'b10) begin
        if(A_PE_dummy_in_5__ap_done_global__q0) begin
          A_PE_dummy_in_5__state <= 2'b00;
        end 
      end 
    end
  end

  assign A_PE_dummy_in_5__ap_start = (A_PE_dummy_in_5__state == 2'b01);
  assign A_PE_dummy_in_6__ap_start_global__q0 = ap_start__q0;
  assign A_PE_dummy_in_6__is_done__q0 = (A_PE_dummy_in_6__state == 2'b10);
  assign A_PE_dummy_in_6__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      A_PE_dummy_in_6__state <= 2'b00;
    end else begin
      if(A_PE_dummy_in_6__state == 2'b00) begin
        if(A_PE_dummy_in_6__ap_start_global__q0) begin
          A_PE_dummy_in_6__state <= 2'b01;
        end 
      end 
      if(A_PE_dummy_in_6__state == 2'b01) begin
        if(A_PE_dummy_in_6__ap_ready) begin
          if(A_PE_dummy_in_6__ap_done) begin
            A_PE_dummy_in_6__state <= 2'b10;
          end else begin
            A_PE_dummy_in_6__state <= 2'b11;
          end
        end 
      end 
      if(A_PE_dummy_in_6__state == 2'b11) begin
        if(A_PE_dummy_in_6__ap_done) begin
          A_PE_dummy_in_6__state <= 2'b10;
        end 
      end 
      if(A_PE_dummy_in_6__state == 2'b10) begin
        if(A_PE_dummy_in_6__ap_done_global__q0) begin
          A_PE_dummy_in_6__state <= 2'b00;
        end 
      end 
    end
  end

  assign A_PE_dummy_in_6__ap_start = (A_PE_dummy_in_6__state == 2'b01);
  assign A_PE_dummy_in_7__ap_start_global__q0 = ap_start__q0;
  assign A_PE_dummy_in_7__is_done__q0 = (A_PE_dummy_in_7__state == 2'b10);
  assign A_PE_dummy_in_7__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      A_PE_dummy_in_7__state <= 2'b00;
    end else begin
      if(A_PE_dummy_in_7__state == 2'b00) begin
        if(A_PE_dummy_in_7__ap_start_global__q0) begin
          A_PE_dummy_in_7__state <= 2'b01;
        end 
      end 
      if(A_PE_dummy_in_7__state == 2'b01) begin
        if(A_PE_dummy_in_7__ap_ready) begin
          if(A_PE_dummy_in_7__ap_done) begin
            A_PE_dummy_in_7__state <= 2'b10;
          end else begin
            A_PE_dummy_in_7__state <= 2'b11;
          end
        end 
      end 
      if(A_PE_dummy_in_7__state == 2'b11) begin
        if(A_PE_dummy_in_7__ap_done) begin
          A_PE_dummy_in_7__state <= 2'b10;
        end 
      end 
      if(A_PE_dummy_in_7__state == 2'b10) begin
        if(A_PE_dummy_in_7__ap_done_global__q0) begin
          A_PE_dummy_in_7__state <= 2'b00;
        end 
      end 
    end
  end

  assign A_PE_dummy_in_7__ap_start = (A_PE_dummy_in_7__state == 2'b01);
  assign A_PE_dummy_in_8__ap_start_global__q0 = ap_start__q0;
  assign A_PE_dummy_in_8__is_done__q0 = (A_PE_dummy_in_8__state == 2'b10);
  assign A_PE_dummy_in_8__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      A_PE_dummy_in_8__state <= 2'b00;
    end else begin
      if(A_PE_dummy_in_8__state == 2'b00) begin
        if(A_PE_dummy_in_8__ap_start_global__q0) begin
          A_PE_dummy_in_8__state <= 2'b01;
        end 
      end 
      if(A_PE_dummy_in_8__state == 2'b01) begin
        if(A_PE_dummy_in_8__ap_ready) begin
          if(A_PE_dummy_in_8__ap_done) begin
            A_PE_dummy_in_8__state <= 2'b10;
          end else begin
            A_PE_dummy_in_8__state <= 2'b11;
          end
        end 
      end 
      if(A_PE_dummy_in_8__state == 2'b11) begin
        if(A_PE_dummy_in_8__ap_done) begin
          A_PE_dummy_in_8__state <= 2'b10;
        end 
      end 
      if(A_PE_dummy_in_8__state == 2'b10) begin
        if(A_PE_dummy_in_8__ap_done_global__q0) begin
          A_PE_dummy_in_8__state <= 2'b00;
        end 
      end 
    end
  end

  assign A_PE_dummy_in_8__ap_start = (A_PE_dummy_in_8__state == 2'b01);
  assign A_PE_dummy_in_9__ap_start_global__q0 = ap_start__q0;
  assign A_PE_dummy_in_9__is_done__q0 = (A_PE_dummy_in_9__state == 2'b10);
  assign A_PE_dummy_in_9__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      A_PE_dummy_in_9__state <= 2'b00;
    end else begin
      if(A_PE_dummy_in_9__state == 2'b00) begin
        if(A_PE_dummy_in_9__ap_start_global__q0) begin
          A_PE_dummy_in_9__state <= 2'b01;
        end 
      end 
      if(A_PE_dummy_in_9__state == 2'b01) begin
        if(A_PE_dummy_in_9__ap_ready) begin
          if(A_PE_dummy_in_9__ap_done) begin
            A_PE_dummy_in_9__state <= 2'b10;
          end else begin
            A_PE_dummy_in_9__state <= 2'b11;
          end
        end 
      end 
      if(A_PE_dummy_in_9__state == 2'b11) begin
        if(A_PE_dummy_in_9__ap_done) begin
          A_PE_dummy_in_9__state <= 2'b10;
        end 
      end 
      if(A_PE_dummy_in_9__state == 2'b10) begin
        if(A_PE_dummy_in_9__ap_done_global__q0) begin
          A_PE_dummy_in_9__state <= 2'b00;
        end 
      end 
    end
  end

  assign A_PE_dummy_in_9__ap_start = (A_PE_dummy_in_9__state == 2'b01);
  assign A_PE_dummy_in_10__ap_start_global__q0 = ap_start__q0;
  assign A_PE_dummy_in_10__is_done__q0 = (A_PE_dummy_in_10__state == 2'b10);
  assign A_PE_dummy_in_10__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      A_PE_dummy_in_10__state <= 2'b00;
    end else begin
      if(A_PE_dummy_in_10__state == 2'b00) begin
        if(A_PE_dummy_in_10__ap_start_global__q0) begin
          A_PE_dummy_in_10__state <= 2'b01;
        end 
      end 
      if(A_PE_dummy_in_10__state == 2'b01) begin
        if(A_PE_dummy_in_10__ap_ready) begin
          if(A_PE_dummy_in_10__ap_done) begin
            A_PE_dummy_in_10__state <= 2'b10;
          end else begin
            A_PE_dummy_in_10__state <= 2'b11;
          end
        end 
      end 
      if(A_PE_dummy_in_10__state == 2'b11) begin
        if(A_PE_dummy_in_10__ap_done) begin
          A_PE_dummy_in_10__state <= 2'b10;
        end 
      end 
      if(A_PE_dummy_in_10__state == 2'b10) begin
        if(A_PE_dummy_in_10__ap_done_global__q0) begin
          A_PE_dummy_in_10__state <= 2'b00;
        end 
      end 
    end
  end

  assign A_PE_dummy_in_10__ap_start = (A_PE_dummy_in_10__state == 2'b01);
  assign A_PE_dummy_in_11__ap_start_global__q0 = ap_start__q0;
  assign A_PE_dummy_in_11__is_done__q0 = (A_PE_dummy_in_11__state == 2'b10);
  assign A_PE_dummy_in_11__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      A_PE_dummy_in_11__state <= 2'b00;
    end else begin
      if(A_PE_dummy_in_11__state == 2'b00) begin
        if(A_PE_dummy_in_11__ap_start_global__q0) begin
          A_PE_dummy_in_11__state <= 2'b01;
        end 
      end 
      if(A_PE_dummy_in_11__state == 2'b01) begin
        if(A_PE_dummy_in_11__ap_ready) begin
          if(A_PE_dummy_in_11__ap_done) begin
            A_PE_dummy_in_11__state <= 2'b10;
          end else begin
            A_PE_dummy_in_11__state <= 2'b11;
          end
        end 
      end 
      if(A_PE_dummy_in_11__state == 2'b11) begin
        if(A_PE_dummy_in_11__ap_done) begin
          A_PE_dummy_in_11__state <= 2'b10;
        end 
      end 
      if(A_PE_dummy_in_11__state == 2'b10) begin
        if(A_PE_dummy_in_11__ap_done_global__q0) begin
          A_PE_dummy_in_11__state <= 2'b00;
        end 
      end 
    end
  end

  assign A_PE_dummy_in_11__ap_start = (A_PE_dummy_in_11__state == 2'b01);
  assign A_PE_dummy_in_12__ap_start_global__q0 = ap_start__q0;
  assign A_PE_dummy_in_12__is_done__q0 = (A_PE_dummy_in_12__state == 2'b10);
  assign A_PE_dummy_in_12__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      A_PE_dummy_in_12__state <= 2'b00;
    end else begin
      if(A_PE_dummy_in_12__state == 2'b00) begin
        if(A_PE_dummy_in_12__ap_start_global__q0) begin
          A_PE_dummy_in_12__state <= 2'b01;
        end 
      end 
      if(A_PE_dummy_in_12__state == 2'b01) begin
        if(A_PE_dummy_in_12__ap_ready) begin
          if(A_PE_dummy_in_12__ap_done) begin
            A_PE_dummy_in_12__state <= 2'b10;
          end else begin
            A_PE_dummy_in_12__state <= 2'b11;
          end
        end 
      end 
      if(A_PE_dummy_in_12__state == 2'b11) begin
        if(A_PE_dummy_in_12__ap_done) begin
          A_PE_dummy_in_12__state <= 2'b10;
        end 
      end 
      if(A_PE_dummy_in_12__state == 2'b10) begin
        if(A_PE_dummy_in_12__ap_done_global__q0) begin
          A_PE_dummy_in_12__state <= 2'b00;
        end 
      end 
    end
  end

  assign A_PE_dummy_in_12__ap_start = (A_PE_dummy_in_12__state == 2'b01);
  assign A_PE_dummy_in_13__ap_start_global__q0 = ap_start__q0;
  assign A_PE_dummy_in_13__is_done__q0 = (A_PE_dummy_in_13__state == 2'b10);
  assign A_PE_dummy_in_13__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      A_PE_dummy_in_13__state <= 2'b00;
    end else begin
      if(A_PE_dummy_in_13__state == 2'b00) begin
        if(A_PE_dummy_in_13__ap_start_global__q0) begin
          A_PE_dummy_in_13__state <= 2'b01;
        end 
      end 
      if(A_PE_dummy_in_13__state == 2'b01) begin
        if(A_PE_dummy_in_13__ap_ready) begin
          if(A_PE_dummy_in_13__ap_done) begin
            A_PE_dummy_in_13__state <= 2'b10;
          end else begin
            A_PE_dummy_in_13__state <= 2'b11;
          end
        end 
      end 
      if(A_PE_dummy_in_13__state == 2'b11) begin
        if(A_PE_dummy_in_13__ap_done) begin
          A_PE_dummy_in_13__state <= 2'b10;
        end 
      end 
      if(A_PE_dummy_in_13__state == 2'b10) begin
        if(A_PE_dummy_in_13__ap_done_global__q0) begin
          A_PE_dummy_in_13__state <= 2'b00;
        end 
      end 
    end
  end

  assign A_PE_dummy_in_13__ap_start = (A_PE_dummy_in_13__state == 2'b01);
  assign A_PE_dummy_in_14__ap_start_global__q0 = ap_start__q0;
  assign A_PE_dummy_in_14__is_done__q0 = (A_PE_dummy_in_14__state == 2'b10);
  assign A_PE_dummy_in_14__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      A_PE_dummy_in_14__state <= 2'b00;
    end else begin
      if(A_PE_dummy_in_14__state == 2'b00) begin
        if(A_PE_dummy_in_14__ap_start_global__q0) begin
          A_PE_dummy_in_14__state <= 2'b01;
        end 
      end 
      if(A_PE_dummy_in_14__state == 2'b01) begin
        if(A_PE_dummy_in_14__ap_ready) begin
          if(A_PE_dummy_in_14__ap_done) begin
            A_PE_dummy_in_14__state <= 2'b10;
          end else begin
            A_PE_dummy_in_14__state <= 2'b11;
          end
        end 
      end 
      if(A_PE_dummy_in_14__state == 2'b11) begin
        if(A_PE_dummy_in_14__ap_done) begin
          A_PE_dummy_in_14__state <= 2'b10;
        end 
      end 
      if(A_PE_dummy_in_14__state == 2'b10) begin
        if(A_PE_dummy_in_14__ap_done_global__q0) begin
          A_PE_dummy_in_14__state <= 2'b00;
        end 
      end 
    end
  end

  assign A_PE_dummy_in_14__ap_start = (A_PE_dummy_in_14__state == 2'b01);
  assign A_PE_dummy_in_15__ap_start_global__q0 = ap_start__q0;
  assign A_PE_dummy_in_15__is_done__q0 = (A_PE_dummy_in_15__state == 2'b10);
  assign A_PE_dummy_in_15__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      A_PE_dummy_in_15__state <= 2'b00;
    end else begin
      if(A_PE_dummy_in_15__state == 2'b00) begin
        if(A_PE_dummy_in_15__ap_start_global__q0) begin
          A_PE_dummy_in_15__state <= 2'b01;
        end 
      end 
      if(A_PE_dummy_in_15__state == 2'b01) begin
        if(A_PE_dummy_in_15__ap_ready) begin
          if(A_PE_dummy_in_15__ap_done) begin
            A_PE_dummy_in_15__state <= 2'b10;
          end else begin
            A_PE_dummy_in_15__state <= 2'b11;
          end
        end 
      end 
      if(A_PE_dummy_in_15__state == 2'b11) begin
        if(A_PE_dummy_in_15__ap_done) begin
          A_PE_dummy_in_15__state <= 2'b10;
        end 
      end 
      if(A_PE_dummy_in_15__state == 2'b10) begin
        if(A_PE_dummy_in_15__ap_done_global__q0) begin
          A_PE_dummy_in_15__state <= 2'b00;
        end 
      end 
    end
  end

  assign A_PE_dummy_in_15__ap_start = (A_PE_dummy_in_15__state == 2'b01);
  assign A_PE_dummy_in_16__ap_start_global__q0 = ap_start__q0;
  assign A_PE_dummy_in_16__is_done__q0 = (A_PE_dummy_in_16__state == 2'b10);
  assign A_PE_dummy_in_16__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      A_PE_dummy_in_16__state <= 2'b00;
    end else begin
      if(A_PE_dummy_in_16__state == 2'b00) begin
        if(A_PE_dummy_in_16__ap_start_global__q0) begin
          A_PE_dummy_in_16__state <= 2'b01;
        end 
      end 
      if(A_PE_dummy_in_16__state == 2'b01) begin
        if(A_PE_dummy_in_16__ap_ready) begin
          if(A_PE_dummy_in_16__ap_done) begin
            A_PE_dummy_in_16__state <= 2'b10;
          end else begin
            A_PE_dummy_in_16__state <= 2'b11;
          end
        end 
      end 
      if(A_PE_dummy_in_16__state == 2'b11) begin
        if(A_PE_dummy_in_16__ap_done) begin
          A_PE_dummy_in_16__state <= 2'b10;
        end 
      end 
      if(A_PE_dummy_in_16__state == 2'b10) begin
        if(A_PE_dummy_in_16__ap_done_global__q0) begin
          A_PE_dummy_in_16__state <= 2'b00;
        end 
      end 
    end
  end

  assign A_PE_dummy_in_16__ap_start = (A_PE_dummy_in_16__state == 2'b01);
  assign A_PE_dummy_in_17__ap_start_global__q0 = ap_start__q0;
  assign A_PE_dummy_in_17__is_done__q0 = (A_PE_dummy_in_17__state == 2'b10);
  assign A_PE_dummy_in_17__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      A_PE_dummy_in_17__state <= 2'b00;
    end else begin
      if(A_PE_dummy_in_17__state == 2'b00) begin
        if(A_PE_dummy_in_17__ap_start_global__q0) begin
          A_PE_dummy_in_17__state <= 2'b01;
        end 
      end 
      if(A_PE_dummy_in_17__state == 2'b01) begin
        if(A_PE_dummy_in_17__ap_ready) begin
          if(A_PE_dummy_in_17__ap_done) begin
            A_PE_dummy_in_17__state <= 2'b10;
          end else begin
            A_PE_dummy_in_17__state <= 2'b11;
          end
        end 
      end 
      if(A_PE_dummy_in_17__state == 2'b11) begin
        if(A_PE_dummy_in_17__ap_done) begin
          A_PE_dummy_in_17__state <= 2'b10;
        end 
      end 
      if(A_PE_dummy_in_17__state == 2'b10) begin
        if(A_PE_dummy_in_17__ap_done_global__q0) begin
          A_PE_dummy_in_17__state <= 2'b00;
        end 
      end 
    end
  end

  assign A_PE_dummy_in_17__ap_start = (A_PE_dummy_in_17__state == 2'b01);
  assign B_IO_L2_in_0__ap_start_global__q0 = ap_start__q0;
  assign B_IO_L2_in_0__is_done__q0 = (B_IO_L2_in_0__state == 2'b10);
  assign B_IO_L2_in_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      B_IO_L2_in_0__state <= 2'b00;
    end else begin
      if(B_IO_L2_in_0__state == 2'b00) begin
        if(B_IO_L2_in_0__ap_start_global__q0) begin
          B_IO_L2_in_0__state <= 2'b01;
        end 
      end 
      if(B_IO_L2_in_0__state == 2'b01) begin
        if(B_IO_L2_in_0__ap_ready) begin
          if(B_IO_L2_in_0__ap_done) begin
            B_IO_L2_in_0__state <= 2'b10;
          end else begin
            B_IO_L2_in_0__state <= 2'b11;
          end
        end 
      end 
      if(B_IO_L2_in_0__state == 2'b11) begin
        if(B_IO_L2_in_0__ap_done) begin
          B_IO_L2_in_0__state <= 2'b10;
        end 
      end 
      if(B_IO_L2_in_0__state == 2'b10) begin
        if(B_IO_L2_in_0__ap_done_global__q0) begin
          B_IO_L2_in_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign B_IO_L2_in_0__ap_start = (B_IO_L2_in_0__state == 2'b01);
  assign B_IO_L2_in_1__ap_start_global__q0 = ap_start__q0;
  assign B_IO_L2_in_1__is_done__q0 = (B_IO_L2_in_1__state == 2'b10);
  assign B_IO_L2_in_1__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      B_IO_L2_in_1__state <= 2'b00;
    end else begin
      if(B_IO_L2_in_1__state == 2'b00) begin
        if(B_IO_L2_in_1__ap_start_global__q0) begin
          B_IO_L2_in_1__state <= 2'b01;
        end 
      end 
      if(B_IO_L2_in_1__state == 2'b01) begin
        if(B_IO_L2_in_1__ap_ready) begin
          if(B_IO_L2_in_1__ap_done) begin
            B_IO_L2_in_1__state <= 2'b10;
          end else begin
            B_IO_L2_in_1__state <= 2'b11;
          end
        end 
      end 
      if(B_IO_L2_in_1__state == 2'b11) begin
        if(B_IO_L2_in_1__ap_done) begin
          B_IO_L2_in_1__state <= 2'b10;
        end 
      end 
      if(B_IO_L2_in_1__state == 2'b10) begin
        if(B_IO_L2_in_1__ap_done_global__q0) begin
          B_IO_L2_in_1__state <= 2'b00;
        end 
      end 
    end
  end

  assign B_IO_L2_in_1__ap_start = (B_IO_L2_in_1__state == 2'b01);
  assign B_IO_L2_in_2__ap_start_global__q0 = ap_start__q0;
  assign B_IO_L2_in_2__is_done__q0 = (B_IO_L2_in_2__state == 2'b10);
  assign B_IO_L2_in_2__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      B_IO_L2_in_2__state <= 2'b00;
    end else begin
      if(B_IO_L2_in_2__state == 2'b00) begin
        if(B_IO_L2_in_2__ap_start_global__q0) begin
          B_IO_L2_in_2__state <= 2'b01;
        end 
      end 
      if(B_IO_L2_in_2__state == 2'b01) begin
        if(B_IO_L2_in_2__ap_ready) begin
          if(B_IO_L2_in_2__ap_done) begin
            B_IO_L2_in_2__state <= 2'b10;
          end else begin
            B_IO_L2_in_2__state <= 2'b11;
          end
        end 
      end 
      if(B_IO_L2_in_2__state == 2'b11) begin
        if(B_IO_L2_in_2__ap_done) begin
          B_IO_L2_in_2__state <= 2'b10;
        end 
      end 
      if(B_IO_L2_in_2__state == 2'b10) begin
        if(B_IO_L2_in_2__ap_done_global__q0) begin
          B_IO_L2_in_2__state <= 2'b00;
        end 
      end 
    end
  end

  assign B_IO_L2_in_2__ap_start = (B_IO_L2_in_2__state == 2'b01);
  assign B_IO_L2_in_3__ap_start_global__q0 = ap_start__q0;
  assign B_IO_L2_in_3__is_done__q0 = (B_IO_L2_in_3__state == 2'b10);
  assign B_IO_L2_in_3__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      B_IO_L2_in_3__state <= 2'b00;
    end else begin
      if(B_IO_L2_in_3__state == 2'b00) begin
        if(B_IO_L2_in_3__ap_start_global__q0) begin
          B_IO_L2_in_3__state <= 2'b01;
        end 
      end 
      if(B_IO_L2_in_3__state == 2'b01) begin
        if(B_IO_L2_in_3__ap_ready) begin
          if(B_IO_L2_in_3__ap_done) begin
            B_IO_L2_in_3__state <= 2'b10;
          end else begin
            B_IO_L2_in_3__state <= 2'b11;
          end
        end 
      end 
      if(B_IO_L2_in_3__state == 2'b11) begin
        if(B_IO_L2_in_3__ap_done) begin
          B_IO_L2_in_3__state <= 2'b10;
        end 
      end 
      if(B_IO_L2_in_3__state == 2'b10) begin
        if(B_IO_L2_in_3__ap_done_global__q0) begin
          B_IO_L2_in_3__state <= 2'b00;
        end 
      end 
    end
  end

  assign B_IO_L2_in_3__ap_start = (B_IO_L2_in_3__state == 2'b01);
  assign B_IO_L2_in_4__ap_start_global__q0 = ap_start__q0;
  assign B_IO_L2_in_4__is_done__q0 = (B_IO_L2_in_4__state == 2'b10);
  assign B_IO_L2_in_4__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      B_IO_L2_in_4__state <= 2'b00;
    end else begin
      if(B_IO_L2_in_4__state == 2'b00) begin
        if(B_IO_L2_in_4__ap_start_global__q0) begin
          B_IO_L2_in_4__state <= 2'b01;
        end 
      end 
      if(B_IO_L2_in_4__state == 2'b01) begin
        if(B_IO_L2_in_4__ap_ready) begin
          if(B_IO_L2_in_4__ap_done) begin
            B_IO_L2_in_4__state <= 2'b10;
          end else begin
            B_IO_L2_in_4__state <= 2'b11;
          end
        end 
      end 
      if(B_IO_L2_in_4__state == 2'b11) begin
        if(B_IO_L2_in_4__ap_done) begin
          B_IO_L2_in_4__state <= 2'b10;
        end 
      end 
      if(B_IO_L2_in_4__state == 2'b10) begin
        if(B_IO_L2_in_4__ap_done_global__q0) begin
          B_IO_L2_in_4__state <= 2'b00;
        end 
      end 
    end
  end

  assign B_IO_L2_in_4__ap_start = (B_IO_L2_in_4__state == 2'b01);
  assign B_IO_L2_in_5__ap_start_global__q0 = ap_start__q0;
  assign B_IO_L2_in_5__is_done__q0 = (B_IO_L2_in_5__state == 2'b10);
  assign B_IO_L2_in_5__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      B_IO_L2_in_5__state <= 2'b00;
    end else begin
      if(B_IO_L2_in_5__state == 2'b00) begin
        if(B_IO_L2_in_5__ap_start_global__q0) begin
          B_IO_L2_in_5__state <= 2'b01;
        end 
      end 
      if(B_IO_L2_in_5__state == 2'b01) begin
        if(B_IO_L2_in_5__ap_ready) begin
          if(B_IO_L2_in_5__ap_done) begin
            B_IO_L2_in_5__state <= 2'b10;
          end else begin
            B_IO_L2_in_5__state <= 2'b11;
          end
        end 
      end 
      if(B_IO_L2_in_5__state == 2'b11) begin
        if(B_IO_L2_in_5__ap_done) begin
          B_IO_L2_in_5__state <= 2'b10;
        end 
      end 
      if(B_IO_L2_in_5__state == 2'b10) begin
        if(B_IO_L2_in_5__ap_done_global__q0) begin
          B_IO_L2_in_5__state <= 2'b00;
        end 
      end 
    end
  end

  assign B_IO_L2_in_5__ap_start = (B_IO_L2_in_5__state == 2'b01);
  assign B_IO_L2_in_6__ap_start_global__q0 = ap_start__q0;
  assign B_IO_L2_in_6__is_done__q0 = (B_IO_L2_in_6__state == 2'b10);
  assign B_IO_L2_in_6__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      B_IO_L2_in_6__state <= 2'b00;
    end else begin
      if(B_IO_L2_in_6__state == 2'b00) begin
        if(B_IO_L2_in_6__ap_start_global__q0) begin
          B_IO_L2_in_6__state <= 2'b01;
        end 
      end 
      if(B_IO_L2_in_6__state == 2'b01) begin
        if(B_IO_L2_in_6__ap_ready) begin
          if(B_IO_L2_in_6__ap_done) begin
            B_IO_L2_in_6__state <= 2'b10;
          end else begin
            B_IO_L2_in_6__state <= 2'b11;
          end
        end 
      end 
      if(B_IO_L2_in_6__state == 2'b11) begin
        if(B_IO_L2_in_6__ap_done) begin
          B_IO_L2_in_6__state <= 2'b10;
        end 
      end 
      if(B_IO_L2_in_6__state == 2'b10) begin
        if(B_IO_L2_in_6__ap_done_global__q0) begin
          B_IO_L2_in_6__state <= 2'b00;
        end 
      end 
    end
  end

  assign B_IO_L2_in_6__ap_start = (B_IO_L2_in_6__state == 2'b01);
  assign B_IO_L2_in_7__ap_start_global__q0 = ap_start__q0;
  assign B_IO_L2_in_7__is_done__q0 = (B_IO_L2_in_7__state == 2'b10);
  assign B_IO_L2_in_7__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      B_IO_L2_in_7__state <= 2'b00;
    end else begin
      if(B_IO_L2_in_7__state == 2'b00) begin
        if(B_IO_L2_in_7__ap_start_global__q0) begin
          B_IO_L2_in_7__state <= 2'b01;
        end 
      end 
      if(B_IO_L2_in_7__state == 2'b01) begin
        if(B_IO_L2_in_7__ap_ready) begin
          if(B_IO_L2_in_7__ap_done) begin
            B_IO_L2_in_7__state <= 2'b10;
          end else begin
            B_IO_L2_in_7__state <= 2'b11;
          end
        end 
      end 
      if(B_IO_L2_in_7__state == 2'b11) begin
        if(B_IO_L2_in_7__ap_done) begin
          B_IO_L2_in_7__state <= 2'b10;
        end 
      end 
      if(B_IO_L2_in_7__state == 2'b10) begin
        if(B_IO_L2_in_7__ap_done_global__q0) begin
          B_IO_L2_in_7__state <= 2'b00;
        end 
      end 
    end
  end

  assign B_IO_L2_in_7__ap_start = (B_IO_L2_in_7__state == 2'b01);
  assign B_IO_L2_in_8__ap_start_global__q0 = ap_start__q0;
  assign B_IO_L2_in_8__is_done__q0 = (B_IO_L2_in_8__state == 2'b10);
  assign B_IO_L2_in_8__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      B_IO_L2_in_8__state <= 2'b00;
    end else begin
      if(B_IO_L2_in_8__state == 2'b00) begin
        if(B_IO_L2_in_8__ap_start_global__q0) begin
          B_IO_L2_in_8__state <= 2'b01;
        end 
      end 
      if(B_IO_L2_in_8__state == 2'b01) begin
        if(B_IO_L2_in_8__ap_ready) begin
          if(B_IO_L2_in_8__ap_done) begin
            B_IO_L2_in_8__state <= 2'b10;
          end else begin
            B_IO_L2_in_8__state <= 2'b11;
          end
        end 
      end 
      if(B_IO_L2_in_8__state == 2'b11) begin
        if(B_IO_L2_in_8__ap_done) begin
          B_IO_L2_in_8__state <= 2'b10;
        end 
      end 
      if(B_IO_L2_in_8__state == 2'b10) begin
        if(B_IO_L2_in_8__ap_done_global__q0) begin
          B_IO_L2_in_8__state <= 2'b00;
        end 
      end 
    end
  end

  assign B_IO_L2_in_8__ap_start = (B_IO_L2_in_8__state == 2'b01);
  assign B_IO_L2_in_9__ap_start_global__q0 = ap_start__q0;
  assign B_IO_L2_in_9__is_done__q0 = (B_IO_L2_in_9__state == 2'b10);
  assign B_IO_L2_in_9__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      B_IO_L2_in_9__state <= 2'b00;
    end else begin
      if(B_IO_L2_in_9__state == 2'b00) begin
        if(B_IO_L2_in_9__ap_start_global__q0) begin
          B_IO_L2_in_9__state <= 2'b01;
        end 
      end 
      if(B_IO_L2_in_9__state == 2'b01) begin
        if(B_IO_L2_in_9__ap_ready) begin
          if(B_IO_L2_in_9__ap_done) begin
            B_IO_L2_in_9__state <= 2'b10;
          end else begin
            B_IO_L2_in_9__state <= 2'b11;
          end
        end 
      end 
      if(B_IO_L2_in_9__state == 2'b11) begin
        if(B_IO_L2_in_9__ap_done) begin
          B_IO_L2_in_9__state <= 2'b10;
        end 
      end 
      if(B_IO_L2_in_9__state == 2'b10) begin
        if(B_IO_L2_in_9__ap_done_global__q0) begin
          B_IO_L2_in_9__state <= 2'b00;
        end 
      end 
    end
  end

  assign B_IO_L2_in_9__ap_start = (B_IO_L2_in_9__state == 2'b01);
  assign B_IO_L2_in_10__ap_start_global__q0 = ap_start__q0;
  assign B_IO_L2_in_10__is_done__q0 = (B_IO_L2_in_10__state == 2'b10);
  assign B_IO_L2_in_10__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      B_IO_L2_in_10__state <= 2'b00;
    end else begin
      if(B_IO_L2_in_10__state == 2'b00) begin
        if(B_IO_L2_in_10__ap_start_global__q0) begin
          B_IO_L2_in_10__state <= 2'b01;
        end 
      end 
      if(B_IO_L2_in_10__state == 2'b01) begin
        if(B_IO_L2_in_10__ap_ready) begin
          if(B_IO_L2_in_10__ap_done) begin
            B_IO_L2_in_10__state <= 2'b10;
          end else begin
            B_IO_L2_in_10__state <= 2'b11;
          end
        end 
      end 
      if(B_IO_L2_in_10__state == 2'b11) begin
        if(B_IO_L2_in_10__ap_done) begin
          B_IO_L2_in_10__state <= 2'b10;
        end 
      end 
      if(B_IO_L2_in_10__state == 2'b10) begin
        if(B_IO_L2_in_10__ap_done_global__q0) begin
          B_IO_L2_in_10__state <= 2'b00;
        end 
      end 
    end
  end

  assign B_IO_L2_in_10__ap_start = (B_IO_L2_in_10__state == 2'b01);
  assign B_IO_L2_in_11__ap_start_global__q0 = ap_start__q0;
  assign B_IO_L2_in_11__is_done__q0 = (B_IO_L2_in_11__state == 2'b10);
  assign B_IO_L2_in_11__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      B_IO_L2_in_11__state <= 2'b00;
    end else begin
      if(B_IO_L2_in_11__state == 2'b00) begin
        if(B_IO_L2_in_11__ap_start_global__q0) begin
          B_IO_L2_in_11__state <= 2'b01;
        end 
      end 
      if(B_IO_L2_in_11__state == 2'b01) begin
        if(B_IO_L2_in_11__ap_ready) begin
          if(B_IO_L2_in_11__ap_done) begin
            B_IO_L2_in_11__state <= 2'b10;
          end else begin
            B_IO_L2_in_11__state <= 2'b11;
          end
        end 
      end 
      if(B_IO_L2_in_11__state == 2'b11) begin
        if(B_IO_L2_in_11__ap_done) begin
          B_IO_L2_in_11__state <= 2'b10;
        end 
      end 
      if(B_IO_L2_in_11__state == 2'b10) begin
        if(B_IO_L2_in_11__ap_done_global__q0) begin
          B_IO_L2_in_11__state <= 2'b00;
        end 
      end 
    end
  end

  assign B_IO_L2_in_11__ap_start = (B_IO_L2_in_11__state == 2'b01);
  assign B_IO_L2_in_12__ap_start_global__q0 = ap_start__q0;
  assign B_IO_L2_in_12__is_done__q0 = (B_IO_L2_in_12__state == 2'b10);
  assign B_IO_L2_in_12__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      B_IO_L2_in_12__state <= 2'b00;
    end else begin
      if(B_IO_L2_in_12__state == 2'b00) begin
        if(B_IO_L2_in_12__ap_start_global__q0) begin
          B_IO_L2_in_12__state <= 2'b01;
        end 
      end 
      if(B_IO_L2_in_12__state == 2'b01) begin
        if(B_IO_L2_in_12__ap_ready) begin
          if(B_IO_L2_in_12__ap_done) begin
            B_IO_L2_in_12__state <= 2'b10;
          end else begin
            B_IO_L2_in_12__state <= 2'b11;
          end
        end 
      end 
      if(B_IO_L2_in_12__state == 2'b11) begin
        if(B_IO_L2_in_12__ap_done) begin
          B_IO_L2_in_12__state <= 2'b10;
        end 
      end 
      if(B_IO_L2_in_12__state == 2'b10) begin
        if(B_IO_L2_in_12__ap_done_global__q0) begin
          B_IO_L2_in_12__state <= 2'b00;
        end 
      end 
    end
  end

  assign B_IO_L2_in_12__ap_start = (B_IO_L2_in_12__state == 2'b01);
  assign B_IO_L2_in_13__ap_start_global__q0 = ap_start__q0;
  assign B_IO_L2_in_13__is_done__q0 = (B_IO_L2_in_13__state == 2'b10);
  assign B_IO_L2_in_13__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      B_IO_L2_in_13__state <= 2'b00;
    end else begin
      if(B_IO_L2_in_13__state == 2'b00) begin
        if(B_IO_L2_in_13__ap_start_global__q0) begin
          B_IO_L2_in_13__state <= 2'b01;
        end 
      end 
      if(B_IO_L2_in_13__state == 2'b01) begin
        if(B_IO_L2_in_13__ap_ready) begin
          if(B_IO_L2_in_13__ap_done) begin
            B_IO_L2_in_13__state <= 2'b10;
          end else begin
            B_IO_L2_in_13__state <= 2'b11;
          end
        end 
      end 
      if(B_IO_L2_in_13__state == 2'b11) begin
        if(B_IO_L2_in_13__ap_done) begin
          B_IO_L2_in_13__state <= 2'b10;
        end 
      end 
      if(B_IO_L2_in_13__state == 2'b10) begin
        if(B_IO_L2_in_13__ap_done_global__q0) begin
          B_IO_L2_in_13__state <= 2'b00;
        end 
      end 
    end
  end

  assign B_IO_L2_in_13__ap_start = (B_IO_L2_in_13__state == 2'b01);
  assign B_IO_L2_in_14__ap_start_global__q0 = ap_start__q0;
  assign B_IO_L2_in_14__is_done__q0 = (B_IO_L2_in_14__state == 2'b10);
  assign B_IO_L2_in_14__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      B_IO_L2_in_14__state <= 2'b00;
    end else begin
      if(B_IO_L2_in_14__state == 2'b00) begin
        if(B_IO_L2_in_14__ap_start_global__q0) begin
          B_IO_L2_in_14__state <= 2'b01;
        end 
      end 
      if(B_IO_L2_in_14__state == 2'b01) begin
        if(B_IO_L2_in_14__ap_ready) begin
          if(B_IO_L2_in_14__ap_done) begin
            B_IO_L2_in_14__state <= 2'b10;
          end else begin
            B_IO_L2_in_14__state <= 2'b11;
          end
        end 
      end 
      if(B_IO_L2_in_14__state == 2'b11) begin
        if(B_IO_L2_in_14__ap_done) begin
          B_IO_L2_in_14__state <= 2'b10;
        end 
      end 
      if(B_IO_L2_in_14__state == 2'b10) begin
        if(B_IO_L2_in_14__ap_done_global__q0) begin
          B_IO_L2_in_14__state <= 2'b00;
        end 
      end 
    end
  end

  assign B_IO_L2_in_14__ap_start = (B_IO_L2_in_14__state == 2'b01);
  assign B_IO_L2_in_15__ap_start_global__q0 = ap_start__q0;
  assign B_IO_L2_in_15__is_done__q0 = (B_IO_L2_in_15__state == 2'b10);
  assign B_IO_L2_in_15__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      B_IO_L2_in_15__state <= 2'b00;
    end else begin
      if(B_IO_L2_in_15__state == 2'b00) begin
        if(B_IO_L2_in_15__ap_start_global__q0) begin
          B_IO_L2_in_15__state <= 2'b01;
        end 
      end 
      if(B_IO_L2_in_15__state == 2'b01) begin
        if(B_IO_L2_in_15__ap_ready) begin
          if(B_IO_L2_in_15__ap_done) begin
            B_IO_L2_in_15__state <= 2'b10;
          end else begin
            B_IO_L2_in_15__state <= 2'b11;
          end
        end 
      end 
      if(B_IO_L2_in_15__state == 2'b11) begin
        if(B_IO_L2_in_15__ap_done) begin
          B_IO_L2_in_15__state <= 2'b10;
        end 
      end 
      if(B_IO_L2_in_15__state == 2'b10) begin
        if(B_IO_L2_in_15__ap_done_global__q0) begin
          B_IO_L2_in_15__state <= 2'b00;
        end 
      end 
    end
  end

  assign B_IO_L2_in_15__ap_start = (B_IO_L2_in_15__state == 2'b01);
  assign B_IO_L2_in_boundary_0__ap_start_global__q0 = ap_start__q0;
  assign B_IO_L2_in_boundary_0__is_done__q0 = (B_IO_L2_in_boundary_0__state == 2'b10);
  assign B_IO_L2_in_boundary_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      B_IO_L2_in_boundary_0__state <= 2'b00;
    end else begin
      if(B_IO_L2_in_boundary_0__state == 2'b00) begin
        if(B_IO_L2_in_boundary_0__ap_start_global__q0) begin
          B_IO_L2_in_boundary_0__state <= 2'b01;
        end 
      end 
      if(B_IO_L2_in_boundary_0__state == 2'b01) begin
        if(B_IO_L2_in_boundary_0__ap_ready) begin
          if(B_IO_L2_in_boundary_0__ap_done) begin
            B_IO_L2_in_boundary_0__state <= 2'b10;
          end else begin
            B_IO_L2_in_boundary_0__state <= 2'b11;
          end
        end 
      end 
      if(B_IO_L2_in_boundary_0__state == 2'b11) begin
        if(B_IO_L2_in_boundary_0__ap_done) begin
          B_IO_L2_in_boundary_0__state <= 2'b10;
        end 
      end 
      if(B_IO_L2_in_boundary_0__state == 2'b10) begin
        if(B_IO_L2_in_boundary_0__ap_done_global__q0) begin
          B_IO_L2_in_boundary_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign B_IO_L2_in_boundary_0__ap_start = (B_IO_L2_in_boundary_0__state == 2'b01);
  assign B_IO_L3_in_0__ap_start_global__q0 = ap_start__q0;
  assign B_IO_L3_in_0__is_done__q0 = (B_IO_L3_in_0__state == 2'b10);
  assign B_IO_L3_in_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      B_IO_L3_in_0__state <= 2'b00;
    end else begin
      if(B_IO_L3_in_0__state == 2'b00) begin
        if(B_IO_L3_in_0__ap_start_global__q0) begin
          B_IO_L3_in_0__state <= 2'b01;
        end 
      end 
      if(B_IO_L3_in_0__state == 2'b01) begin
        if(B_IO_L3_in_0__ap_ready) begin
          if(B_IO_L3_in_0__ap_done) begin
            B_IO_L3_in_0__state <= 2'b10;
          end else begin
            B_IO_L3_in_0__state <= 2'b11;
          end
        end 
      end 
      if(B_IO_L3_in_0__state == 2'b11) begin
        if(B_IO_L3_in_0__ap_done) begin
          B_IO_L3_in_0__state <= 2'b10;
        end 
      end 
      if(B_IO_L3_in_0__state == 2'b10) begin
        if(B_IO_L3_in_0__ap_done_global__q0) begin
          B_IO_L3_in_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign B_IO_L3_in_0__ap_start = (B_IO_L3_in_0__state == 2'b01);
  assign B_IO_L3_in_serialize_0___B__q0 = B;
  assign B_IO_L3_in_serialize_0__ap_start_global__q0 = ap_start__q0;
  assign B_IO_L3_in_serialize_0__is_done__q0 = (B_IO_L3_in_serialize_0__state == 2'b10);
  assign B_IO_L3_in_serialize_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      B_IO_L3_in_serialize_0__state <= 2'b00;
    end else begin
      if(B_IO_L3_in_serialize_0__state == 2'b00) begin
        if(B_IO_L3_in_serialize_0__ap_start_global__q0) begin
          B_IO_L3_in_serialize_0__state <= 2'b01;
        end 
      end 
      if(B_IO_L3_in_serialize_0__state == 2'b01) begin
        if(B_IO_L3_in_serialize_0__ap_ready) begin
          if(B_IO_L3_in_serialize_0__ap_done) begin
            B_IO_L3_in_serialize_0__state <= 2'b10;
          end else begin
            B_IO_L3_in_serialize_0__state <= 2'b11;
          end
        end 
      end 
      if(B_IO_L3_in_serialize_0__state == 2'b11) begin
        if(B_IO_L3_in_serialize_0__ap_done) begin
          B_IO_L3_in_serialize_0__state <= 2'b10;
        end 
      end 
      if(B_IO_L3_in_serialize_0__state == 2'b10) begin
        if(B_IO_L3_in_serialize_0__ap_done_global__q0) begin
          B_IO_L3_in_serialize_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign B_IO_L3_in_serialize_0__ap_start = (B_IO_L3_in_serialize_0__state == 2'b01);
  assign B_PE_dummy_in_0__ap_start_global__q0 = ap_start__q0;
  assign B_PE_dummy_in_0__is_done__q0 = (B_PE_dummy_in_0__state == 2'b10);
  assign B_PE_dummy_in_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      B_PE_dummy_in_0__state <= 2'b00;
    end else begin
      if(B_PE_dummy_in_0__state == 2'b00) begin
        if(B_PE_dummy_in_0__ap_start_global__q0) begin
          B_PE_dummy_in_0__state <= 2'b01;
        end 
      end 
      if(B_PE_dummy_in_0__state == 2'b01) begin
        if(B_PE_dummy_in_0__ap_ready) begin
          if(B_PE_dummy_in_0__ap_done) begin
            B_PE_dummy_in_0__state <= 2'b10;
          end else begin
            B_PE_dummy_in_0__state <= 2'b11;
          end
        end 
      end 
      if(B_PE_dummy_in_0__state == 2'b11) begin
        if(B_PE_dummy_in_0__ap_done) begin
          B_PE_dummy_in_0__state <= 2'b10;
        end 
      end 
      if(B_PE_dummy_in_0__state == 2'b10) begin
        if(B_PE_dummy_in_0__ap_done_global__q0) begin
          B_PE_dummy_in_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign B_PE_dummy_in_0__ap_start = (B_PE_dummy_in_0__state == 2'b01);
  assign B_PE_dummy_in_1__ap_start_global__q0 = ap_start__q0;
  assign B_PE_dummy_in_1__is_done__q0 = (B_PE_dummy_in_1__state == 2'b10);
  assign B_PE_dummy_in_1__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      B_PE_dummy_in_1__state <= 2'b00;
    end else begin
      if(B_PE_dummy_in_1__state == 2'b00) begin
        if(B_PE_dummy_in_1__ap_start_global__q0) begin
          B_PE_dummy_in_1__state <= 2'b01;
        end 
      end 
      if(B_PE_dummy_in_1__state == 2'b01) begin
        if(B_PE_dummy_in_1__ap_ready) begin
          if(B_PE_dummy_in_1__ap_done) begin
            B_PE_dummy_in_1__state <= 2'b10;
          end else begin
            B_PE_dummy_in_1__state <= 2'b11;
          end
        end 
      end 
      if(B_PE_dummy_in_1__state == 2'b11) begin
        if(B_PE_dummy_in_1__ap_done) begin
          B_PE_dummy_in_1__state <= 2'b10;
        end 
      end 
      if(B_PE_dummy_in_1__state == 2'b10) begin
        if(B_PE_dummy_in_1__ap_done_global__q0) begin
          B_PE_dummy_in_1__state <= 2'b00;
        end 
      end 
    end
  end

  assign B_PE_dummy_in_1__ap_start = (B_PE_dummy_in_1__state == 2'b01);
  assign B_PE_dummy_in_2__ap_start_global__q0 = ap_start__q0;
  assign B_PE_dummy_in_2__is_done__q0 = (B_PE_dummy_in_2__state == 2'b10);
  assign B_PE_dummy_in_2__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      B_PE_dummy_in_2__state <= 2'b00;
    end else begin
      if(B_PE_dummy_in_2__state == 2'b00) begin
        if(B_PE_dummy_in_2__ap_start_global__q0) begin
          B_PE_dummy_in_2__state <= 2'b01;
        end 
      end 
      if(B_PE_dummy_in_2__state == 2'b01) begin
        if(B_PE_dummy_in_2__ap_ready) begin
          if(B_PE_dummy_in_2__ap_done) begin
            B_PE_dummy_in_2__state <= 2'b10;
          end else begin
            B_PE_dummy_in_2__state <= 2'b11;
          end
        end 
      end 
      if(B_PE_dummy_in_2__state == 2'b11) begin
        if(B_PE_dummy_in_2__ap_done) begin
          B_PE_dummy_in_2__state <= 2'b10;
        end 
      end 
      if(B_PE_dummy_in_2__state == 2'b10) begin
        if(B_PE_dummy_in_2__ap_done_global__q0) begin
          B_PE_dummy_in_2__state <= 2'b00;
        end 
      end 
    end
  end

  assign B_PE_dummy_in_2__ap_start = (B_PE_dummy_in_2__state == 2'b01);
  assign B_PE_dummy_in_3__ap_start_global__q0 = ap_start__q0;
  assign B_PE_dummy_in_3__is_done__q0 = (B_PE_dummy_in_3__state == 2'b10);
  assign B_PE_dummy_in_3__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      B_PE_dummy_in_3__state <= 2'b00;
    end else begin
      if(B_PE_dummy_in_3__state == 2'b00) begin
        if(B_PE_dummy_in_3__ap_start_global__q0) begin
          B_PE_dummy_in_3__state <= 2'b01;
        end 
      end 
      if(B_PE_dummy_in_3__state == 2'b01) begin
        if(B_PE_dummy_in_3__ap_ready) begin
          if(B_PE_dummy_in_3__ap_done) begin
            B_PE_dummy_in_3__state <= 2'b10;
          end else begin
            B_PE_dummy_in_3__state <= 2'b11;
          end
        end 
      end 
      if(B_PE_dummy_in_3__state == 2'b11) begin
        if(B_PE_dummy_in_3__ap_done) begin
          B_PE_dummy_in_3__state <= 2'b10;
        end 
      end 
      if(B_PE_dummy_in_3__state == 2'b10) begin
        if(B_PE_dummy_in_3__ap_done_global__q0) begin
          B_PE_dummy_in_3__state <= 2'b00;
        end 
      end 
    end
  end

  assign B_PE_dummy_in_3__ap_start = (B_PE_dummy_in_3__state == 2'b01);
  assign B_PE_dummy_in_4__ap_start_global__q0 = ap_start__q0;
  assign B_PE_dummy_in_4__is_done__q0 = (B_PE_dummy_in_4__state == 2'b10);
  assign B_PE_dummy_in_4__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      B_PE_dummy_in_4__state <= 2'b00;
    end else begin
      if(B_PE_dummy_in_4__state == 2'b00) begin
        if(B_PE_dummy_in_4__ap_start_global__q0) begin
          B_PE_dummy_in_4__state <= 2'b01;
        end 
      end 
      if(B_PE_dummy_in_4__state == 2'b01) begin
        if(B_PE_dummy_in_4__ap_ready) begin
          if(B_PE_dummy_in_4__ap_done) begin
            B_PE_dummy_in_4__state <= 2'b10;
          end else begin
            B_PE_dummy_in_4__state <= 2'b11;
          end
        end 
      end 
      if(B_PE_dummy_in_4__state == 2'b11) begin
        if(B_PE_dummy_in_4__ap_done) begin
          B_PE_dummy_in_4__state <= 2'b10;
        end 
      end 
      if(B_PE_dummy_in_4__state == 2'b10) begin
        if(B_PE_dummy_in_4__ap_done_global__q0) begin
          B_PE_dummy_in_4__state <= 2'b00;
        end 
      end 
    end
  end

  assign B_PE_dummy_in_4__ap_start = (B_PE_dummy_in_4__state == 2'b01);
  assign B_PE_dummy_in_5__ap_start_global__q0 = ap_start__q0;
  assign B_PE_dummy_in_5__is_done__q0 = (B_PE_dummy_in_5__state == 2'b10);
  assign B_PE_dummy_in_5__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      B_PE_dummy_in_5__state <= 2'b00;
    end else begin
      if(B_PE_dummy_in_5__state == 2'b00) begin
        if(B_PE_dummy_in_5__ap_start_global__q0) begin
          B_PE_dummy_in_5__state <= 2'b01;
        end 
      end 
      if(B_PE_dummy_in_5__state == 2'b01) begin
        if(B_PE_dummy_in_5__ap_ready) begin
          if(B_PE_dummy_in_5__ap_done) begin
            B_PE_dummy_in_5__state <= 2'b10;
          end else begin
            B_PE_dummy_in_5__state <= 2'b11;
          end
        end 
      end 
      if(B_PE_dummy_in_5__state == 2'b11) begin
        if(B_PE_dummy_in_5__ap_done) begin
          B_PE_dummy_in_5__state <= 2'b10;
        end 
      end 
      if(B_PE_dummy_in_5__state == 2'b10) begin
        if(B_PE_dummy_in_5__ap_done_global__q0) begin
          B_PE_dummy_in_5__state <= 2'b00;
        end 
      end 
    end
  end

  assign B_PE_dummy_in_5__ap_start = (B_PE_dummy_in_5__state == 2'b01);
  assign B_PE_dummy_in_6__ap_start_global__q0 = ap_start__q0;
  assign B_PE_dummy_in_6__is_done__q0 = (B_PE_dummy_in_6__state == 2'b10);
  assign B_PE_dummy_in_6__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      B_PE_dummy_in_6__state <= 2'b00;
    end else begin
      if(B_PE_dummy_in_6__state == 2'b00) begin
        if(B_PE_dummy_in_6__ap_start_global__q0) begin
          B_PE_dummy_in_6__state <= 2'b01;
        end 
      end 
      if(B_PE_dummy_in_6__state == 2'b01) begin
        if(B_PE_dummy_in_6__ap_ready) begin
          if(B_PE_dummy_in_6__ap_done) begin
            B_PE_dummy_in_6__state <= 2'b10;
          end else begin
            B_PE_dummy_in_6__state <= 2'b11;
          end
        end 
      end 
      if(B_PE_dummy_in_6__state == 2'b11) begin
        if(B_PE_dummy_in_6__ap_done) begin
          B_PE_dummy_in_6__state <= 2'b10;
        end 
      end 
      if(B_PE_dummy_in_6__state == 2'b10) begin
        if(B_PE_dummy_in_6__ap_done_global__q0) begin
          B_PE_dummy_in_6__state <= 2'b00;
        end 
      end 
    end
  end

  assign B_PE_dummy_in_6__ap_start = (B_PE_dummy_in_6__state == 2'b01);
  assign B_PE_dummy_in_7__ap_start_global__q0 = ap_start__q0;
  assign B_PE_dummy_in_7__is_done__q0 = (B_PE_dummy_in_7__state == 2'b10);
  assign B_PE_dummy_in_7__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      B_PE_dummy_in_7__state <= 2'b00;
    end else begin
      if(B_PE_dummy_in_7__state == 2'b00) begin
        if(B_PE_dummy_in_7__ap_start_global__q0) begin
          B_PE_dummy_in_7__state <= 2'b01;
        end 
      end 
      if(B_PE_dummy_in_7__state == 2'b01) begin
        if(B_PE_dummy_in_7__ap_ready) begin
          if(B_PE_dummy_in_7__ap_done) begin
            B_PE_dummy_in_7__state <= 2'b10;
          end else begin
            B_PE_dummy_in_7__state <= 2'b11;
          end
        end 
      end 
      if(B_PE_dummy_in_7__state == 2'b11) begin
        if(B_PE_dummy_in_7__ap_done) begin
          B_PE_dummy_in_7__state <= 2'b10;
        end 
      end 
      if(B_PE_dummy_in_7__state == 2'b10) begin
        if(B_PE_dummy_in_7__ap_done_global__q0) begin
          B_PE_dummy_in_7__state <= 2'b00;
        end 
      end 
    end
  end

  assign B_PE_dummy_in_7__ap_start = (B_PE_dummy_in_7__state == 2'b01);
  assign B_PE_dummy_in_8__ap_start_global__q0 = ap_start__q0;
  assign B_PE_dummy_in_8__is_done__q0 = (B_PE_dummy_in_8__state == 2'b10);
  assign B_PE_dummy_in_8__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      B_PE_dummy_in_8__state <= 2'b00;
    end else begin
      if(B_PE_dummy_in_8__state == 2'b00) begin
        if(B_PE_dummy_in_8__ap_start_global__q0) begin
          B_PE_dummy_in_8__state <= 2'b01;
        end 
      end 
      if(B_PE_dummy_in_8__state == 2'b01) begin
        if(B_PE_dummy_in_8__ap_ready) begin
          if(B_PE_dummy_in_8__ap_done) begin
            B_PE_dummy_in_8__state <= 2'b10;
          end else begin
            B_PE_dummy_in_8__state <= 2'b11;
          end
        end 
      end 
      if(B_PE_dummy_in_8__state == 2'b11) begin
        if(B_PE_dummy_in_8__ap_done) begin
          B_PE_dummy_in_8__state <= 2'b10;
        end 
      end 
      if(B_PE_dummy_in_8__state == 2'b10) begin
        if(B_PE_dummy_in_8__ap_done_global__q0) begin
          B_PE_dummy_in_8__state <= 2'b00;
        end 
      end 
    end
  end

  assign B_PE_dummy_in_8__ap_start = (B_PE_dummy_in_8__state == 2'b01);
  assign B_PE_dummy_in_9__ap_start_global__q0 = ap_start__q0;
  assign B_PE_dummy_in_9__is_done__q0 = (B_PE_dummy_in_9__state == 2'b10);
  assign B_PE_dummy_in_9__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      B_PE_dummy_in_9__state <= 2'b00;
    end else begin
      if(B_PE_dummy_in_9__state == 2'b00) begin
        if(B_PE_dummy_in_9__ap_start_global__q0) begin
          B_PE_dummy_in_9__state <= 2'b01;
        end 
      end 
      if(B_PE_dummy_in_9__state == 2'b01) begin
        if(B_PE_dummy_in_9__ap_ready) begin
          if(B_PE_dummy_in_9__ap_done) begin
            B_PE_dummy_in_9__state <= 2'b10;
          end else begin
            B_PE_dummy_in_9__state <= 2'b11;
          end
        end 
      end 
      if(B_PE_dummy_in_9__state == 2'b11) begin
        if(B_PE_dummy_in_9__ap_done) begin
          B_PE_dummy_in_9__state <= 2'b10;
        end 
      end 
      if(B_PE_dummy_in_9__state == 2'b10) begin
        if(B_PE_dummy_in_9__ap_done_global__q0) begin
          B_PE_dummy_in_9__state <= 2'b00;
        end 
      end 
    end
  end

  assign B_PE_dummy_in_9__ap_start = (B_PE_dummy_in_9__state == 2'b01);
  assign B_PE_dummy_in_10__ap_start_global__q0 = ap_start__q0;
  assign B_PE_dummy_in_10__is_done__q0 = (B_PE_dummy_in_10__state == 2'b10);
  assign B_PE_dummy_in_10__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      B_PE_dummy_in_10__state <= 2'b00;
    end else begin
      if(B_PE_dummy_in_10__state == 2'b00) begin
        if(B_PE_dummy_in_10__ap_start_global__q0) begin
          B_PE_dummy_in_10__state <= 2'b01;
        end 
      end 
      if(B_PE_dummy_in_10__state == 2'b01) begin
        if(B_PE_dummy_in_10__ap_ready) begin
          if(B_PE_dummy_in_10__ap_done) begin
            B_PE_dummy_in_10__state <= 2'b10;
          end else begin
            B_PE_dummy_in_10__state <= 2'b11;
          end
        end 
      end 
      if(B_PE_dummy_in_10__state == 2'b11) begin
        if(B_PE_dummy_in_10__ap_done) begin
          B_PE_dummy_in_10__state <= 2'b10;
        end 
      end 
      if(B_PE_dummy_in_10__state == 2'b10) begin
        if(B_PE_dummy_in_10__ap_done_global__q0) begin
          B_PE_dummy_in_10__state <= 2'b00;
        end 
      end 
    end
  end

  assign B_PE_dummy_in_10__ap_start = (B_PE_dummy_in_10__state == 2'b01);
  assign B_PE_dummy_in_11__ap_start_global__q0 = ap_start__q0;
  assign B_PE_dummy_in_11__is_done__q0 = (B_PE_dummy_in_11__state == 2'b10);
  assign B_PE_dummy_in_11__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      B_PE_dummy_in_11__state <= 2'b00;
    end else begin
      if(B_PE_dummy_in_11__state == 2'b00) begin
        if(B_PE_dummy_in_11__ap_start_global__q0) begin
          B_PE_dummy_in_11__state <= 2'b01;
        end 
      end 
      if(B_PE_dummy_in_11__state == 2'b01) begin
        if(B_PE_dummy_in_11__ap_ready) begin
          if(B_PE_dummy_in_11__ap_done) begin
            B_PE_dummy_in_11__state <= 2'b10;
          end else begin
            B_PE_dummy_in_11__state <= 2'b11;
          end
        end 
      end 
      if(B_PE_dummy_in_11__state == 2'b11) begin
        if(B_PE_dummy_in_11__ap_done) begin
          B_PE_dummy_in_11__state <= 2'b10;
        end 
      end 
      if(B_PE_dummy_in_11__state == 2'b10) begin
        if(B_PE_dummy_in_11__ap_done_global__q0) begin
          B_PE_dummy_in_11__state <= 2'b00;
        end 
      end 
    end
  end

  assign B_PE_dummy_in_11__ap_start = (B_PE_dummy_in_11__state == 2'b01);
  assign B_PE_dummy_in_12__ap_start_global__q0 = ap_start__q0;
  assign B_PE_dummy_in_12__is_done__q0 = (B_PE_dummy_in_12__state == 2'b10);
  assign B_PE_dummy_in_12__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      B_PE_dummy_in_12__state <= 2'b00;
    end else begin
      if(B_PE_dummy_in_12__state == 2'b00) begin
        if(B_PE_dummy_in_12__ap_start_global__q0) begin
          B_PE_dummy_in_12__state <= 2'b01;
        end 
      end 
      if(B_PE_dummy_in_12__state == 2'b01) begin
        if(B_PE_dummy_in_12__ap_ready) begin
          if(B_PE_dummy_in_12__ap_done) begin
            B_PE_dummy_in_12__state <= 2'b10;
          end else begin
            B_PE_dummy_in_12__state <= 2'b11;
          end
        end 
      end 
      if(B_PE_dummy_in_12__state == 2'b11) begin
        if(B_PE_dummy_in_12__ap_done) begin
          B_PE_dummy_in_12__state <= 2'b10;
        end 
      end 
      if(B_PE_dummy_in_12__state == 2'b10) begin
        if(B_PE_dummy_in_12__ap_done_global__q0) begin
          B_PE_dummy_in_12__state <= 2'b00;
        end 
      end 
    end
  end

  assign B_PE_dummy_in_12__ap_start = (B_PE_dummy_in_12__state == 2'b01);
  assign B_PE_dummy_in_13__ap_start_global__q0 = ap_start__q0;
  assign B_PE_dummy_in_13__is_done__q0 = (B_PE_dummy_in_13__state == 2'b10);
  assign B_PE_dummy_in_13__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      B_PE_dummy_in_13__state <= 2'b00;
    end else begin
      if(B_PE_dummy_in_13__state == 2'b00) begin
        if(B_PE_dummy_in_13__ap_start_global__q0) begin
          B_PE_dummy_in_13__state <= 2'b01;
        end 
      end 
      if(B_PE_dummy_in_13__state == 2'b01) begin
        if(B_PE_dummy_in_13__ap_ready) begin
          if(B_PE_dummy_in_13__ap_done) begin
            B_PE_dummy_in_13__state <= 2'b10;
          end else begin
            B_PE_dummy_in_13__state <= 2'b11;
          end
        end 
      end 
      if(B_PE_dummy_in_13__state == 2'b11) begin
        if(B_PE_dummy_in_13__ap_done) begin
          B_PE_dummy_in_13__state <= 2'b10;
        end 
      end 
      if(B_PE_dummy_in_13__state == 2'b10) begin
        if(B_PE_dummy_in_13__ap_done_global__q0) begin
          B_PE_dummy_in_13__state <= 2'b00;
        end 
      end 
    end
  end

  assign B_PE_dummy_in_13__ap_start = (B_PE_dummy_in_13__state == 2'b01);
  assign B_PE_dummy_in_14__ap_start_global__q0 = ap_start__q0;
  assign B_PE_dummy_in_14__is_done__q0 = (B_PE_dummy_in_14__state == 2'b10);
  assign B_PE_dummy_in_14__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      B_PE_dummy_in_14__state <= 2'b00;
    end else begin
      if(B_PE_dummy_in_14__state == 2'b00) begin
        if(B_PE_dummy_in_14__ap_start_global__q0) begin
          B_PE_dummy_in_14__state <= 2'b01;
        end 
      end 
      if(B_PE_dummy_in_14__state == 2'b01) begin
        if(B_PE_dummy_in_14__ap_ready) begin
          if(B_PE_dummy_in_14__ap_done) begin
            B_PE_dummy_in_14__state <= 2'b10;
          end else begin
            B_PE_dummy_in_14__state <= 2'b11;
          end
        end 
      end 
      if(B_PE_dummy_in_14__state == 2'b11) begin
        if(B_PE_dummy_in_14__ap_done) begin
          B_PE_dummy_in_14__state <= 2'b10;
        end 
      end 
      if(B_PE_dummy_in_14__state == 2'b10) begin
        if(B_PE_dummy_in_14__ap_done_global__q0) begin
          B_PE_dummy_in_14__state <= 2'b00;
        end 
      end 
    end
  end

  assign B_PE_dummy_in_14__ap_start = (B_PE_dummy_in_14__state == 2'b01);
  assign B_PE_dummy_in_15__ap_start_global__q0 = ap_start__q0;
  assign B_PE_dummy_in_15__is_done__q0 = (B_PE_dummy_in_15__state == 2'b10);
  assign B_PE_dummy_in_15__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      B_PE_dummy_in_15__state <= 2'b00;
    end else begin
      if(B_PE_dummy_in_15__state == 2'b00) begin
        if(B_PE_dummy_in_15__ap_start_global__q0) begin
          B_PE_dummy_in_15__state <= 2'b01;
        end 
      end 
      if(B_PE_dummy_in_15__state == 2'b01) begin
        if(B_PE_dummy_in_15__ap_ready) begin
          if(B_PE_dummy_in_15__ap_done) begin
            B_PE_dummy_in_15__state <= 2'b10;
          end else begin
            B_PE_dummy_in_15__state <= 2'b11;
          end
        end 
      end 
      if(B_PE_dummy_in_15__state == 2'b11) begin
        if(B_PE_dummy_in_15__ap_done) begin
          B_PE_dummy_in_15__state <= 2'b10;
        end 
      end 
      if(B_PE_dummy_in_15__state == 2'b10) begin
        if(B_PE_dummy_in_15__ap_done_global__q0) begin
          B_PE_dummy_in_15__state <= 2'b00;
        end 
      end 
    end
  end

  assign B_PE_dummy_in_15__ap_start = (B_PE_dummy_in_15__state == 2'b01);
  assign B_PE_dummy_in_16__ap_start_global__q0 = ap_start__q0;
  assign B_PE_dummy_in_16__is_done__q0 = (B_PE_dummy_in_16__state == 2'b10);
  assign B_PE_dummy_in_16__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      B_PE_dummy_in_16__state <= 2'b00;
    end else begin
      if(B_PE_dummy_in_16__state == 2'b00) begin
        if(B_PE_dummy_in_16__ap_start_global__q0) begin
          B_PE_dummy_in_16__state <= 2'b01;
        end 
      end 
      if(B_PE_dummy_in_16__state == 2'b01) begin
        if(B_PE_dummy_in_16__ap_ready) begin
          if(B_PE_dummy_in_16__ap_done) begin
            B_PE_dummy_in_16__state <= 2'b10;
          end else begin
            B_PE_dummy_in_16__state <= 2'b11;
          end
        end 
      end 
      if(B_PE_dummy_in_16__state == 2'b11) begin
        if(B_PE_dummy_in_16__ap_done) begin
          B_PE_dummy_in_16__state <= 2'b10;
        end 
      end 
      if(B_PE_dummy_in_16__state == 2'b10) begin
        if(B_PE_dummy_in_16__ap_done_global__q0) begin
          B_PE_dummy_in_16__state <= 2'b00;
        end 
      end 
    end
  end

  assign B_PE_dummy_in_16__ap_start = (B_PE_dummy_in_16__state == 2'b01);
  assign C_drain_IO_L1_out_boundary_wrapper_0__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_boundary_wrapper_0__is_done__q0 = (C_drain_IO_L1_out_boundary_wrapper_0__state == 2'b10);
  assign C_drain_IO_L1_out_boundary_wrapper_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_boundary_wrapper_0__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_boundary_wrapper_0__state == 2'b00) begin
        if(C_drain_IO_L1_out_boundary_wrapper_0__ap_start_global__q0) begin
          C_drain_IO_L1_out_boundary_wrapper_0__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_0__state == 2'b01) begin
        if(C_drain_IO_L1_out_boundary_wrapper_0__ap_ready) begin
          if(C_drain_IO_L1_out_boundary_wrapper_0__ap_done) begin
            C_drain_IO_L1_out_boundary_wrapper_0__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_boundary_wrapper_0__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_0__state == 2'b11) begin
        if(C_drain_IO_L1_out_boundary_wrapper_0__ap_done) begin
          C_drain_IO_L1_out_boundary_wrapper_0__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_0__state == 2'b10) begin
        if(C_drain_IO_L1_out_boundary_wrapper_0__ap_done_global__q0) begin
          C_drain_IO_L1_out_boundary_wrapper_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_boundary_wrapper_0__ap_start = (C_drain_IO_L1_out_boundary_wrapper_0__state == 2'b01);
  assign C_drain_IO_L1_out_boundary_wrapper_1__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_boundary_wrapper_1__is_done__q0 = (C_drain_IO_L1_out_boundary_wrapper_1__state == 2'b10);
  assign C_drain_IO_L1_out_boundary_wrapper_1__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_boundary_wrapper_1__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_boundary_wrapper_1__state == 2'b00) begin
        if(C_drain_IO_L1_out_boundary_wrapper_1__ap_start_global__q0) begin
          C_drain_IO_L1_out_boundary_wrapper_1__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_1__state == 2'b01) begin
        if(C_drain_IO_L1_out_boundary_wrapper_1__ap_ready) begin
          if(C_drain_IO_L1_out_boundary_wrapper_1__ap_done) begin
            C_drain_IO_L1_out_boundary_wrapper_1__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_boundary_wrapper_1__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_1__state == 2'b11) begin
        if(C_drain_IO_L1_out_boundary_wrapper_1__ap_done) begin
          C_drain_IO_L1_out_boundary_wrapper_1__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_1__state == 2'b10) begin
        if(C_drain_IO_L1_out_boundary_wrapper_1__ap_done_global__q0) begin
          C_drain_IO_L1_out_boundary_wrapper_1__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_boundary_wrapper_1__ap_start = (C_drain_IO_L1_out_boundary_wrapper_1__state == 2'b01);
  assign C_drain_IO_L1_out_boundary_wrapper_2__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_boundary_wrapper_2__is_done__q0 = (C_drain_IO_L1_out_boundary_wrapper_2__state == 2'b10);
  assign C_drain_IO_L1_out_boundary_wrapper_2__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_boundary_wrapper_2__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_boundary_wrapper_2__state == 2'b00) begin
        if(C_drain_IO_L1_out_boundary_wrapper_2__ap_start_global__q0) begin
          C_drain_IO_L1_out_boundary_wrapper_2__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_2__state == 2'b01) begin
        if(C_drain_IO_L1_out_boundary_wrapper_2__ap_ready) begin
          if(C_drain_IO_L1_out_boundary_wrapper_2__ap_done) begin
            C_drain_IO_L1_out_boundary_wrapper_2__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_boundary_wrapper_2__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_2__state == 2'b11) begin
        if(C_drain_IO_L1_out_boundary_wrapper_2__ap_done) begin
          C_drain_IO_L1_out_boundary_wrapper_2__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_2__state == 2'b10) begin
        if(C_drain_IO_L1_out_boundary_wrapper_2__ap_done_global__q0) begin
          C_drain_IO_L1_out_boundary_wrapper_2__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_boundary_wrapper_2__ap_start = (C_drain_IO_L1_out_boundary_wrapper_2__state == 2'b01);
  assign C_drain_IO_L1_out_boundary_wrapper_3__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_boundary_wrapper_3__is_done__q0 = (C_drain_IO_L1_out_boundary_wrapper_3__state == 2'b10);
  assign C_drain_IO_L1_out_boundary_wrapper_3__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_boundary_wrapper_3__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_boundary_wrapper_3__state == 2'b00) begin
        if(C_drain_IO_L1_out_boundary_wrapper_3__ap_start_global__q0) begin
          C_drain_IO_L1_out_boundary_wrapper_3__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_3__state == 2'b01) begin
        if(C_drain_IO_L1_out_boundary_wrapper_3__ap_ready) begin
          if(C_drain_IO_L1_out_boundary_wrapper_3__ap_done) begin
            C_drain_IO_L1_out_boundary_wrapper_3__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_boundary_wrapper_3__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_3__state == 2'b11) begin
        if(C_drain_IO_L1_out_boundary_wrapper_3__ap_done) begin
          C_drain_IO_L1_out_boundary_wrapper_3__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_3__state == 2'b10) begin
        if(C_drain_IO_L1_out_boundary_wrapper_3__ap_done_global__q0) begin
          C_drain_IO_L1_out_boundary_wrapper_3__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_boundary_wrapper_3__ap_start = (C_drain_IO_L1_out_boundary_wrapper_3__state == 2'b01);
  assign C_drain_IO_L1_out_boundary_wrapper_4__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_boundary_wrapper_4__is_done__q0 = (C_drain_IO_L1_out_boundary_wrapper_4__state == 2'b10);
  assign C_drain_IO_L1_out_boundary_wrapper_4__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_boundary_wrapper_4__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_boundary_wrapper_4__state == 2'b00) begin
        if(C_drain_IO_L1_out_boundary_wrapper_4__ap_start_global__q0) begin
          C_drain_IO_L1_out_boundary_wrapper_4__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_4__state == 2'b01) begin
        if(C_drain_IO_L1_out_boundary_wrapper_4__ap_ready) begin
          if(C_drain_IO_L1_out_boundary_wrapper_4__ap_done) begin
            C_drain_IO_L1_out_boundary_wrapper_4__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_boundary_wrapper_4__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_4__state == 2'b11) begin
        if(C_drain_IO_L1_out_boundary_wrapper_4__ap_done) begin
          C_drain_IO_L1_out_boundary_wrapper_4__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_4__state == 2'b10) begin
        if(C_drain_IO_L1_out_boundary_wrapper_4__ap_done_global__q0) begin
          C_drain_IO_L1_out_boundary_wrapper_4__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_boundary_wrapper_4__ap_start = (C_drain_IO_L1_out_boundary_wrapper_4__state == 2'b01);
  assign C_drain_IO_L1_out_boundary_wrapper_5__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_boundary_wrapper_5__is_done__q0 = (C_drain_IO_L1_out_boundary_wrapper_5__state == 2'b10);
  assign C_drain_IO_L1_out_boundary_wrapper_5__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_boundary_wrapper_5__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_boundary_wrapper_5__state == 2'b00) begin
        if(C_drain_IO_L1_out_boundary_wrapper_5__ap_start_global__q0) begin
          C_drain_IO_L1_out_boundary_wrapper_5__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_5__state == 2'b01) begin
        if(C_drain_IO_L1_out_boundary_wrapper_5__ap_ready) begin
          if(C_drain_IO_L1_out_boundary_wrapper_5__ap_done) begin
            C_drain_IO_L1_out_boundary_wrapper_5__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_boundary_wrapper_5__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_5__state == 2'b11) begin
        if(C_drain_IO_L1_out_boundary_wrapper_5__ap_done) begin
          C_drain_IO_L1_out_boundary_wrapper_5__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_5__state == 2'b10) begin
        if(C_drain_IO_L1_out_boundary_wrapper_5__ap_done_global__q0) begin
          C_drain_IO_L1_out_boundary_wrapper_5__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_boundary_wrapper_5__ap_start = (C_drain_IO_L1_out_boundary_wrapper_5__state == 2'b01);
  assign C_drain_IO_L1_out_boundary_wrapper_6__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_boundary_wrapper_6__is_done__q0 = (C_drain_IO_L1_out_boundary_wrapper_6__state == 2'b10);
  assign C_drain_IO_L1_out_boundary_wrapper_6__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_boundary_wrapper_6__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_boundary_wrapper_6__state == 2'b00) begin
        if(C_drain_IO_L1_out_boundary_wrapper_6__ap_start_global__q0) begin
          C_drain_IO_L1_out_boundary_wrapper_6__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_6__state == 2'b01) begin
        if(C_drain_IO_L1_out_boundary_wrapper_6__ap_ready) begin
          if(C_drain_IO_L1_out_boundary_wrapper_6__ap_done) begin
            C_drain_IO_L1_out_boundary_wrapper_6__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_boundary_wrapper_6__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_6__state == 2'b11) begin
        if(C_drain_IO_L1_out_boundary_wrapper_6__ap_done) begin
          C_drain_IO_L1_out_boundary_wrapper_6__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_6__state == 2'b10) begin
        if(C_drain_IO_L1_out_boundary_wrapper_6__ap_done_global__q0) begin
          C_drain_IO_L1_out_boundary_wrapper_6__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_boundary_wrapper_6__ap_start = (C_drain_IO_L1_out_boundary_wrapper_6__state == 2'b01);
  assign C_drain_IO_L1_out_boundary_wrapper_7__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_boundary_wrapper_7__is_done__q0 = (C_drain_IO_L1_out_boundary_wrapper_7__state == 2'b10);
  assign C_drain_IO_L1_out_boundary_wrapper_7__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_boundary_wrapper_7__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_boundary_wrapper_7__state == 2'b00) begin
        if(C_drain_IO_L1_out_boundary_wrapper_7__ap_start_global__q0) begin
          C_drain_IO_L1_out_boundary_wrapper_7__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_7__state == 2'b01) begin
        if(C_drain_IO_L1_out_boundary_wrapper_7__ap_ready) begin
          if(C_drain_IO_L1_out_boundary_wrapper_7__ap_done) begin
            C_drain_IO_L1_out_boundary_wrapper_7__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_boundary_wrapper_7__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_7__state == 2'b11) begin
        if(C_drain_IO_L1_out_boundary_wrapper_7__ap_done) begin
          C_drain_IO_L1_out_boundary_wrapper_7__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_7__state == 2'b10) begin
        if(C_drain_IO_L1_out_boundary_wrapper_7__ap_done_global__q0) begin
          C_drain_IO_L1_out_boundary_wrapper_7__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_boundary_wrapper_7__ap_start = (C_drain_IO_L1_out_boundary_wrapper_7__state == 2'b01);
  assign C_drain_IO_L1_out_boundary_wrapper_8__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_boundary_wrapper_8__is_done__q0 = (C_drain_IO_L1_out_boundary_wrapper_8__state == 2'b10);
  assign C_drain_IO_L1_out_boundary_wrapper_8__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_boundary_wrapper_8__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_boundary_wrapper_8__state == 2'b00) begin
        if(C_drain_IO_L1_out_boundary_wrapper_8__ap_start_global__q0) begin
          C_drain_IO_L1_out_boundary_wrapper_8__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_8__state == 2'b01) begin
        if(C_drain_IO_L1_out_boundary_wrapper_8__ap_ready) begin
          if(C_drain_IO_L1_out_boundary_wrapper_8__ap_done) begin
            C_drain_IO_L1_out_boundary_wrapper_8__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_boundary_wrapper_8__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_8__state == 2'b11) begin
        if(C_drain_IO_L1_out_boundary_wrapper_8__ap_done) begin
          C_drain_IO_L1_out_boundary_wrapper_8__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_8__state == 2'b10) begin
        if(C_drain_IO_L1_out_boundary_wrapper_8__ap_done_global__q0) begin
          C_drain_IO_L1_out_boundary_wrapper_8__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_boundary_wrapper_8__ap_start = (C_drain_IO_L1_out_boundary_wrapper_8__state == 2'b01);
  assign C_drain_IO_L1_out_boundary_wrapper_9__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_boundary_wrapper_9__is_done__q0 = (C_drain_IO_L1_out_boundary_wrapper_9__state == 2'b10);
  assign C_drain_IO_L1_out_boundary_wrapper_9__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_boundary_wrapper_9__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_boundary_wrapper_9__state == 2'b00) begin
        if(C_drain_IO_L1_out_boundary_wrapper_9__ap_start_global__q0) begin
          C_drain_IO_L1_out_boundary_wrapper_9__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_9__state == 2'b01) begin
        if(C_drain_IO_L1_out_boundary_wrapper_9__ap_ready) begin
          if(C_drain_IO_L1_out_boundary_wrapper_9__ap_done) begin
            C_drain_IO_L1_out_boundary_wrapper_9__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_boundary_wrapper_9__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_9__state == 2'b11) begin
        if(C_drain_IO_L1_out_boundary_wrapper_9__ap_done) begin
          C_drain_IO_L1_out_boundary_wrapper_9__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_9__state == 2'b10) begin
        if(C_drain_IO_L1_out_boundary_wrapper_9__ap_done_global__q0) begin
          C_drain_IO_L1_out_boundary_wrapper_9__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_boundary_wrapper_9__ap_start = (C_drain_IO_L1_out_boundary_wrapper_9__state == 2'b01);
  assign C_drain_IO_L1_out_boundary_wrapper_10__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_boundary_wrapper_10__is_done__q0 = (C_drain_IO_L1_out_boundary_wrapper_10__state == 2'b10);
  assign C_drain_IO_L1_out_boundary_wrapper_10__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_boundary_wrapper_10__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_boundary_wrapper_10__state == 2'b00) begin
        if(C_drain_IO_L1_out_boundary_wrapper_10__ap_start_global__q0) begin
          C_drain_IO_L1_out_boundary_wrapper_10__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_10__state == 2'b01) begin
        if(C_drain_IO_L1_out_boundary_wrapper_10__ap_ready) begin
          if(C_drain_IO_L1_out_boundary_wrapper_10__ap_done) begin
            C_drain_IO_L1_out_boundary_wrapper_10__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_boundary_wrapper_10__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_10__state == 2'b11) begin
        if(C_drain_IO_L1_out_boundary_wrapper_10__ap_done) begin
          C_drain_IO_L1_out_boundary_wrapper_10__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_10__state == 2'b10) begin
        if(C_drain_IO_L1_out_boundary_wrapper_10__ap_done_global__q0) begin
          C_drain_IO_L1_out_boundary_wrapper_10__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_boundary_wrapper_10__ap_start = (C_drain_IO_L1_out_boundary_wrapper_10__state == 2'b01);
  assign C_drain_IO_L1_out_boundary_wrapper_11__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_boundary_wrapper_11__is_done__q0 = (C_drain_IO_L1_out_boundary_wrapper_11__state == 2'b10);
  assign C_drain_IO_L1_out_boundary_wrapper_11__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_boundary_wrapper_11__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_boundary_wrapper_11__state == 2'b00) begin
        if(C_drain_IO_L1_out_boundary_wrapper_11__ap_start_global__q0) begin
          C_drain_IO_L1_out_boundary_wrapper_11__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_11__state == 2'b01) begin
        if(C_drain_IO_L1_out_boundary_wrapper_11__ap_ready) begin
          if(C_drain_IO_L1_out_boundary_wrapper_11__ap_done) begin
            C_drain_IO_L1_out_boundary_wrapper_11__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_boundary_wrapper_11__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_11__state == 2'b11) begin
        if(C_drain_IO_L1_out_boundary_wrapper_11__ap_done) begin
          C_drain_IO_L1_out_boundary_wrapper_11__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_11__state == 2'b10) begin
        if(C_drain_IO_L1_out_boundary_wrapper_11__ap_done_global__q0) begin
          C_drain_IO_L1_out_boundary_wrapper_11__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_boundary_wrapper_11__ap_start = (C_drain_IO_L1_out_boundary_wrapper_11__state == 2'b01);
  assign C_drain_IO_L1_out_boundary_wrapper_12__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_boundary_wrapper_12__is_done__q0 = (C_drain_IO_L1_out_boundary_wrapper_12__state == 2'b10);
  assign C_drain_IO_L1_out_boundary_wrapper_12__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_boundary_wrapper_12__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_boundary_wrapper_12__state == 2'b00) begin
        if(C_drain_IO_L1_out_boundary_wrapper_12__ap_start_global__q0) begin
          C_drain_IO_L1_out_boundary_wrapper_12__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_12__state == 2'b01) begin
        if(C_drain_IO_L1_out_boundary_wrapper_12__ap_ready) begin
          if(C_drain_IO_L1_out_boundary_wrapper_12__ap_done) begin
            C_drain_IO_L1_out_boundary_wrapper_12__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_boundary_wrapper_12__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_12__state == 2'b11) begin
        if(C_drain_IO_L1_out_boundary_wrapper_12__ap_done) begin
          C_drain_IO_L1_out_boundary_wrapper_12__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_12__state == 2'b10) begin
        if(C_drain_IO_L1_out_boundary_wrapper_12__ap_done_global__q0) begin
          C_drain_IO_L1_out_boundary_wrapper_12__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_boundary_wrapper_12__ap_start = (C_drain_IO_L1_out_boundary_wrapper_12__state == 2'b01);
  assign C_drain_IO_L1_out_boundary_wrapper_13__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_boundary_wrapper_13__is_done__q0 = (C_drain_IO_L1_out_boundary_wrapper_13__state == 2'b10);
  assign C_drain_IO_L1_out_boundary_wrapper_13__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_boundary_wrapper_13__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_boundary_wrapper_13__state == 2'b00) begin
        if(C_drain_IO_L1_out_boundary_wrapper_13__ap_start_global__q0) begin
          C_drain_IO_L1_out_boundary_wrapper_13__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_13__state == 2'b01) begin
        if(C_drain_IO_L1_out_boundary_wrapper_13__ap_ready) begin
          if(C_drain_IO_L1_out_boundary_wrapper_13__ap_done) begin
            C_drain_IO_L1_out_boundary_wrapper_13__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_boundary_wrapper_13__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_13__state == 2'b11) begin
        if(C_drain_IO_L1_out_boundary_wrapper_13__ap_done) begin
          C_drain_IO_L1_out_boundary_wrapper_13__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_13__state == 2'b10) begin
        if(C_drain_IO_L1_out_boundary_wrapper_13__ap_done_global__q0) begin
          C_drain_IO_L1_out_boundary_wrapper_13__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_boundary_wrapper_13__ap_start = (C_drain_IO_L1_out_boundary_wrapper_13__state == 2'b01);
  assign C_drain_IO_L1_out_boundary_wrapper_14__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_boundary_wrapper_14__is_done__q0 = (C_drain_IO_L1_out_boundary_wrapper_14__state == 2'b10);
  assign C_drain_IO_L1_out_boundary_wrapper_14__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_boundary_wrapper_14__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_boundary_wrapper_14__state == 2'b00) begin
        if(C_drain_IO_L1_out_boundary_wrapper_14__ap_start_global__q0) begin
          C_drain_IO_L1_out_boundary_wrapper_14__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_14__state == 2'b01) begin
        if(C_drain_IO_L1_out_boundary_wrapper_14__ap_ready) begin
          if(C_drain_IO_L1_out_boundary_wrapper_14__ap_done) begin
            C_drain_IO_L1_out_boundary_wrapper_14__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_boundary_wrapper_14__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_14__state == 2'b11) begin
        if(C_drain_IO_L1_out_boundary_wrapper_14__ap_done) begin
          C_drain_IO_L1_out_boundary_wrapper_14__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_14__state == 2'b10) begin
        if(C_drain_IO_L1_out_boundary_wrapper_14__ap_done_global__q0) begin
          C_drain_IO_L1_out_boundary_wrapper_14__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_boundary_wrapper_14__ap_start = (C_drain_IO_L1_out_boundary_wrapper_14__state == 2'b01);
  assign C_drain_IO_L1_out_boundary_wrapper_15__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_boundary_wrapper_15__is_done__q0 = (C_drain_IO_L1_out_boundary_wrapper_15__state == 2'b10);
  assign C_drain_IO_L1_out_boundary_wrapper_15__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_boundary_wrapper_15__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_boundary_wrapper_15__state == 2'b00) begin
        if(C_drain_IO_L1_out_boundary_wrapper_15__ap_start_global__q0) begin
          C_drain_IO_L1_out_boundary_wrapper_15__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_15__state == 2'b01) begin
        if(C_drain_IO_L1_out_boundary_wrapper_15__ap_ready) begin
          if(C_drain_IO_L1_out_boundary_wrapper_15__ap_done) begin
            C_drain_IO_L1_out_boundary_wrapper_15__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_boundary_wrapper_15__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_15__state == 2'b11) begin
        if(C_drain_IO_L1_out_boundary_wrapper_15__ap_done) begin
          C_drain_IO_L1_out_boundary_wrapper_15__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_15__state == 2'b10) begin
        if(C_drain_IO_L1_out_boundary_wrapper_15__ap_done_global__q0) begin
          C_drain_IO_L1_out_boundary_wrapper_15__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_boundary_wrapper_15__ap_start = (C_drain_IO_L1_out_boundary_wrapper_15__state == 2'b01);
  assign C_drain_IO_L1_out_boundary_wrapper_16__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_boundary_wrapper_16__is_done__q0 = (C_drain_IO_L1_out_boundary_wrapper_16__state == 2'b10);
  assign C_drain_IO_L1_out_boundary_wrapper_16__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_boundary_wrapper_16__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_boundary_wrapper_16__state == 2'b00) begin
        if(C_drain_IO_L1_out_boundary_wrapper_16__ap_start_global__q0) begin
          C_drain_IO_L1_out_boundary_wrapper_16__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_16__state == 2'b01) begin
        if(C_drain_IO_L1_out_boundary_wrapper_16__ap_ready) begin
          if(C_drain_IO_L1_out_boundary_wrapper_16__ap_done) begin
            C_drain_IO_L1_out_boundary_wrapper_16__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_boundary_wrapper_16__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_16__state == 2'b11) begin
        if(C_drain_IO_L1_out_boundary_wrapper_16__ap_done) begin
          C_drain_IO_L1_out_boundary_wrapper_16__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_boundary_wrapper_16__state == 2'b10) begin
        if(C_drain_IO_L1_out_boundary_wrapper_16__ap_done_global__q0) begin
          C_drain_IO_L1_out_boundary_wrapper_16__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_boundary_wrapper_16__ap_start = (C_drain_IO_L1_out_boundary_wrapper_16__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_0__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_0__is_done__q0 = (C_drain_IO_L1_out_wrapper_0__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_0__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_0__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_0__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_0__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_0__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_0__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_0__ap_done) begin
            C_drain_IO_L1_out_wrapper_0__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_0__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_0__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_0__ap_done) begin
          C_drain_IO_L1_out_wrapper_0__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_0__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_0__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_0__ap_start = (C_drain_IO_L1_out_wrapper_0__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_1__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_1__is_done__q0 = (C_drain_IO_L1_out_wrapper_1__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_1__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_1__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_1__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_1__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_1__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_1__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_1__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_1__ap_done) begin
            C_drain_IO_L1_out_wrapper_1__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_1__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_1__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_1__ap_done) begin
          C_drain_IO_L1_out_wrapper_1__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_1__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_1__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_1__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_1__ap_start = (C_drain_IO_L1_out_wrapper_1__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_2__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_2__is_done__q0 = (C_drain_IO_L1_out_wrapper_2__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_2__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_2__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_2__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_2__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_2__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_2__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_2__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_2__ap_done) begin
            C_drain_IO_L1_out_wrapper_2__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_2__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_2__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_2__ap_done) begin
          C_drain_IO_L1_out_wrapper_2__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_2__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_2__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_2__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_2__ap_start = (C_drain_IO_L1_out_wrapper_2__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_3__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_3__is_done__q0 = (C_drain_IO_L1_out_wrapper_3__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_3__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_3__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_3__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_3__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_3__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_3__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_3__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_3__ap_done) begin
            C_drain_IO_L1_out_wrapper_3__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_3__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_3__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_3__ap_done) begin
          C_drain_IO_L1_out_wrapper_3__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_3__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_3__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_3__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_3__ap_start = (C_drain_IO_L1_out_wrapper_3__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_4__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_4__is_done__q0 = (C_drain_IO_L1_out_wrapper_4__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_4__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_4__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_4__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_4__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_4__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_4__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_4__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_4__ap_done) begin
            C_drain_IO_L1_out_wrapper_4__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_4__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_4__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_4__ap_done) begin
          C_drain_IO_L1_out_wrapper_4__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_4__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_4__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_4__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_4__ap_start = (C_drain_IO_L1_out_wrapper_4__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_5__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_5__is_done__q0 = (C_drain_IO_L1_out_wrapper_5__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_5__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_5__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_5__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_5__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_5__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_5__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_5__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_5__ap_done) begin
            C_drain_IO_L1_out_wrapper_5__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_5__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_5__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_5__ap_done) begin
          C_drain_IO_L1_out_wrapper_5__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_5__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_5__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_5__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_5__ap_start = (C_drain_IO_L1_out_wrapper_5__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_6__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_6__is_done__q0 = (C_drain_IO_L1_out_wrapper_6__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_6__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_6__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_6__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_6__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_6__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_6__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_6__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_6__ap_done) begin
            C_drain_IO_L1_out_wrapper_6__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_6__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_6__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_6__ap_done) begin
          C_drain_IO_L1_out_wrapper_6__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_6__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_6__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_6__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_6__ap_start = (C_drain_IO_L1_out_wrapper_6__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_7__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_7__is_done__q0 = (C_drain_IO_L1_out_wrapper_7__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_7__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_7__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_7__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_7__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_7__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_7__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_7__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_7__ap_done) begin
            C_drain_IO_L1_out_wrapper_7__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_7__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_7__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_7__ap_done) begin
          C_drain_IO_L1_out_wrapper_7__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_7__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_7__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_7__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_7__ap_start = (C_drain_IO_L1_out_wrapper_7__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_8__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_8__is_done__q0 = (C_drain_IO_L1_out_wrapper_8__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_8__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_8__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_8__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_8__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_8__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_8__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_8__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_8__ap_done) begin
            C_drain_IO_L1_out_wrapper_8__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_8__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_8__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_8__ap_done) begin
          C_drain_IO_L1_out_wrapper_8__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_8__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_8__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_8__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_8__ap_start = (C_drain_IO_L1_out_wrapper_8__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_9__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_9__is_done__q0 = (C_drain_IO_L1_out_wrapper_9__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_9__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_9__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_9__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_9__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_9__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_9__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_9__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_9__ap_done) begin
            C_drain_IO_L1_out_wrapper_9__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_9__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_9__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_9__ap_done) begin
          C_drain_IO_L1_out_wrapper_9__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_9__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_9__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_9__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_9__ap_start = (C_drain_IO_L1_out_wrapper_9__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_10__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_10__is_done__q0 = (C_drain_IO_L1_out_wrapper_10__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_10__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_10__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_10__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_10__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_10__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_10__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_10__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_10__ap_done) begin
            C_drain_IO_L1_out_wrapper_10__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_10__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_10__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_10__ap_done) begin
          C_drain_IO_L1_out_wrapper_10__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_10__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_10__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_10__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_10__ap_start = (C_drain_IO_L1_out_wrapper_10__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_11__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_11__is_done__q0 = (C_drain_IO_L1_out_wrapper_11__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_11__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_11__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_11__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_11__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_11__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_11__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_11__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_11__ap_done) begin
            C_drain_IO_L1_out_wrapper_11__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_11__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_11__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_11__ap_done) begin
          C_drain_IO_L1_out_wrapper_11__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_11__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_11__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_11__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_11__ap_start = (C_drain_IO_L1_out_wrapper_11__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_12__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_12__is_done__q0 = (C_drain_IO_L1_out_wrapper_12__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_12__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_12__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_12__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_12__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_12__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_12__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_12__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_12__ap_done) begin
            C_drain_IO_L1_out_wrapper_12__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_12__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_12__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_12__ap_done) begin
          C_drain_IO_L1_out_wrapper_12__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_12__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_12__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_12__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_12__ap_start = (C_drain_IO_L1_out_wrapper_12__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_13__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_13__is_done__q0 = (C_drain_IO_L1_out_wrapper_13__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_13__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_13__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_13__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_13__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_13__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_13__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_13__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_13__ap_done) begin
            C_drain_IO_L1_out_wrapper_13__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_13__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_13__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_13__ap_done) begin
          C_drain_IO_L1_out_wrapper_13__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_13__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_13__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_13__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_13__ap_start = (C_drain_IO_L1_out_wrapper_13__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_14__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_14__is_done__q0 = (C_drain_IO_L1_out_wrapper_14__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_14__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_14__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_14__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_14__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_14__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_14__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_14__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_14__ap_done) begin
            C_drain_IO_L1_out_wrapper_14__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_14__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_14__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_14__ap_done) begin
          C_drain_IO_L1_out_wrapper_14__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_14__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_14__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_14__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_14__ap_start = (C_drain_IO_L1_out_wrapper_14__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_15__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_15__is_done__q0 = (C_drain_IO_L1_out_wrapper_15__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_15__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_15__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_15__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_15__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_15__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_15__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_15__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_15__ap_done) begin
            C_drain_IO_L1_out_wrapper_15__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_15__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_15__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_15__ap_done) begin
          C_drain_IO_L1_out_wrapper_15__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_15__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_15__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_15__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_15__ap_start = (C_drain_IO_L1_out_wrapper_15__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_16__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_16__is_done__q0 = (C_drain_IO_L1_out_wrapper_16__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_16__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_16__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_16__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_16__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_16__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_16__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_16__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_16__ap_done) begin
            C_drain_IO_L1_out_wrapper_16__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_16__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_16__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_16__ap_done) begin
          C_drain_IO_L1_out_wrapper_16__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_16__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_16__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_16__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_16__ap_start = (C_drain_IO_L1_out_wrapper_16__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_17__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_17__is_done__q0 = (C_drain_IO_L1_out_wrapper_17__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_17__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_17__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_17__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_17__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_17__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_17__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_17__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_17__ap_done) begin
            C_drain_IO_L1_out_wrapper_17__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_17__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_17__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_17__ap_done) begin
          C_drain_IO_L1_out_wrapper_17__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_17__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_17__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_17__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_17__ap_start = (C_drain_IO_L1_out_wrapper_17__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_18__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_18__is_done__q0 = (C_drain_IO_L1_out_wrapper_18__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_18__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_18__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_18__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_18__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_18__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_18__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_18__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_18__ap_done) begin
            C_drain_IO_L1_out_wrapper_18__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_18__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_18__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_18__ap_done) begin
          C_drain_IO_L1_out_wrapper_18__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_18__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_18__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_18__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_18__ap_start = (C_drain_IO_L1_out_wrapper_18__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_19__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_19__is_done__q0 = (C_drain_IO_L1_out_wrapper_19__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_19__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_19__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_19__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_19__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_19__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_19__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_19__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_19__ap_done) begin
            C_drain_IO_L1_out_wrapper_19__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_19__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_19__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_19__ap_done) begin
          C_drain_IO_L1_out_wrapper_19__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_19__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_19__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_19__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_19__ap_start = (C_drain_IO_L1_out_wrapper_19__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_20__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_20__is_done__q0 = (C_drain_IO_L1_out_wrapper_20__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_20__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_20__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_20__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_20__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_20__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_20__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_20__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_20__ap_done) begin
            C_drain_IO_L1_out_wrapper_20__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_20__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_20__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_20__ap_done) begin
          C_drain_IO_L1_out_wrapper_20__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_20__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_20__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_20__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_20__ap_start = (C_drain_IO_L1_out_wrapper_20__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_21__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_21__is_done__q0 = (C_drain_IO_L1_out_wrapper_21__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_21__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_21__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_21__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_21__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_21__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_21__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_21__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_21__ap_done) begin
            C_drain_IO_L1_out_wrapper_21__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_21__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_21__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_21__ap_done) begin
          C_drain_IO_L1_out_wrapper_21__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_21__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_21__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_21__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_21__ap_start = (C_drain_IO_L1_out_wrapper_21__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_22__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_22__is_done__q0 = (C_drain_IO_L1_out_wrapper_22__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_22__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_22__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_22__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_22__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_22__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_22__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_22__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_22__ap_done) begin
            C_drain_IO_L1_out_wrapper_22__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_22__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_22__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_22__ap_done) begin
          C_drain_IO_L1_out_wrapper_22__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_22__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_22__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_22__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_22__ap_start = (C_drain_IO_L1_out_wrapper_22__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_23__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_23__is_done__q0 = (C_drain_IO_L1_out_wrapper_23__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_23__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_23__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_23__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_23__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_23__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_23__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_23__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_23__ap_done) begin
            C_drain_IO_L1_out_wrapper_23__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_23__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_23__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_23__ap_done) begin
          C_drain_IO_L1_out_wrapper_23__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_23__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_23__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_23__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_23__ap_start = (C_drain_IO_L1_out_wrapper_23__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_24__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_24__is_done__q0 = (C_drain_IO_L1_out_wrapper_24__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_24__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_24__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_24__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_24__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_24__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_24__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_24__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_24__ap_done) begin
            C_drain_IO_L1_out_wrapper_24__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_24__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_24__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_24__ap_done) begin
          C_drain_IO_L1_out_wrapper_24__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_24__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_24__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_24__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_24__ap_start = (C_drain_IO_L1_out_wrapper_24__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_25__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_25__is_done__q0 = (C_drain_IO_L1_out_wrapper_25__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_25__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_25__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_25__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_25__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_25__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_25__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_25__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_25__ap_done) begin
            C_drain_IO_L1_out_wrapper_25__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_25__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_25__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_25__ap_done) begin
          C_drain_IO_L1_out_wrapper_25__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_25__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_25__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_25__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_25__ap_start = (C_drain_IO_L1_out_wrapper_25__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_26__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_26__is_done__q0 = (C_drain_IO_L1_out_wrapper_26__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_26__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_26__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_26__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_26__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_26__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_26__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_26__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_26__ap_done) begin
            C_drain_IO_L1_out_wrapper_26__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_26__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_26__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_26__ap_done) begin
          C_drain_IO_L1_out_wrapper_26__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_26__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_26__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_26__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_26__ap_start = (C_drain_IO_L1_out_wrapper_26__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_27__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_27__is_done__q0 = (C_drain_IO_L1_out_wrapper_27__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_27__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_27__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_27__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_27__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_27__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_27__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_27__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_27__ap_done) begin
            C_drain_IO_L1_out_wrapper_27__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_27__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_27__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_27__ap_done) begin
          C_drain_IO_L1_out_wrapper_27__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_27__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_27__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_27__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_27__ap_start = (C_drain_IO_L1_out_wrapper_27__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_28__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_28__is_done__q0 = (C_drain_IO_L1_out_wrapper_28__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_28__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_28__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_28__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_28__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_28__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_28__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_28__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_28__ap_done) begin
            C_drain_IO_L1_out_wrapper_28__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_28__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_28__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_28__ap_done) begin
          C_drain_IO_L1_out_wrapper_28__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_28__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_28__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_28__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_28__ap_start = (C_drain_IO_L1_out_wrapper_28__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_29__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_29__is_done__q0 = (C_drain_IO_L1_out_wrapper_29__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_29__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_29__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_29__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_29__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_29__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_29__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_29__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_29__ap_done) begin
            C_drain_IO_L1_out_wrapper_29__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_29__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_29__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_29__ap_done) begin
          C_drain_IO_L1_out_wrapper_29__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_29__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_29__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_29__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_29__ap_start = (C_drain_IO_L1_out_wrapper_29__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_30__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_30__is_done__q0 = (C_drain_IO_L1_out_wrapper_30__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_30__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_30__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_30__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_30__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_30__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_30__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_30__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_30__ap_done) begin
            C_drain_IO_L1_out_wrapper_30__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_30__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_30__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_30__ap_done) begin
          C_drain_IO_L1_out_wrapper_30__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_30__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_30__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_30__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_30__ap_start = (C_drain_IO_L1_out_wrapper_30__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_31__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_31__is_done__q0 = (C_drain_IO_L1_out_wrapper_31__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_31__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_31__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_31__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_31__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_31__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_31__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_31__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_31__ap_done) begin
            C_drain_IO_L1_out_wrapper_31__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_31__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_31__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_31__ap_done) begin
          C_drain_IO_L1_out_wrapper_31__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_31__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_31__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_31__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_31__ap_start = (C_drain_IO_L1_out_wrapper_31__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_32__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_32__is_done__q0 = (C_drain_IO_L1_out_wrapper_32__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_32__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_32__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_32__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_32__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_32__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_32__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_32__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_32__ap_done) begin
            C_drain_IO_L1_out_wrapper_32__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_32__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_32__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_32__ap_done) begin
          C_drain_IO_L1_out_wrapper_32__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_32__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_32__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_32__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_32__ap_start = (C_drain_IO_L1_out_wrapper_32__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_33__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_33__is_done__q0 = (C_drain_IO_L1_out_wrapper_33__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_33__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_33__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_33__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_33__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_33__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_33__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_33__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_33__ap_done) begin
            C_drain_IO_L1_out_wrapper_33__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_33__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_33__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_33__ap_done) begin
          C_drain_IO_L1_out_wrapper_33__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_33__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_33__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_33__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_33__ap_start = (C_drain_IO_L1_out_wrapper_33__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_34__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_34__is_done__q0 = (C_drain_IO_L1_out_wrapper_34__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_34__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_34__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_34__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_34__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_34__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_34__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_34__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_34__ap_done) begin
            C_drain_IO_L1_out_wrapper_34__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_34__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_34__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_34__ap_done) begin
          C_drain_IO_L1_out_wrapper_34__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_34__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_34__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_34__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_34__ap_start = (C_drain_IO_L1_out_wrapper_34__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_35__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_35__is_done__q0 = (C_drain_IO_L1_out_wrapper_35__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_35__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_35__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_35__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_35__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_35__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_35__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_35__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_35__ap_done) begin
            C_drain_IO_L1_out_wrapper_35__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_35__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_35__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_35__ap_done) begin
          C_drain_IO_L1_out_wrapper_35__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_35__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_35__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_35__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_35__ap_start = (C_drain_IO_L1_out_wrapper_35__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_36__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_36__is_done__q0 = (C_drain_IO_L1_out_wrapper_36__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_36__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_36__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_36__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_36__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_36__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_36__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_36__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_36__ap_done) begin
            C_drain_IO_L1_out_wrapper_36__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_36__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_36__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_36__ap_done) begin
          C_drain_IO_L1_out_wrapper_36__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_36__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_36__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_36__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_36__ap_start = (C_drain_IO_L1_out_wrapper_36__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_37__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_37__is_done__q0 = (C_drain_IO_L1_out_wrapper_37__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_37__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_37__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_37__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_37__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_37__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_37__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_37__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_37__ap_done) begin
            C_drain_IO_L1_out_wrapper_37__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_37__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_37__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_37__ap_done) begin
          C_drain_IO_L1_out_wrapper_37__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_37__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_37__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_37__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_37__ap_start = (C_drain_IO_L1_out_wrapper_37__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_38__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_38__is_done__q0 = (C_drain_IO_L1_out_wrapper_38__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_38__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_38__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_38__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_38__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_38__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_38__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_38__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_38__ap_done) begin
            C_drain_IO_L1_out_wrapper_38__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_38__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_38__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_38__ap_done) begin
          C_drain_IO_L1_out_wrapper_38__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_38__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_38__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_38__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_38__ap_start = (C_drain_IO_L1_out_wrapper_38__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_39__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_39__is_done__q0 = (C_drain_IO_L1_out_wrapper_39__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_39__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_39__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_39__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_39__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_39__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_39__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_39__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_39__ap_done) begin
            C_drain_IO_L1_out_wrapper_39__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_39__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_39__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_39__ap_done) begin
          C_drain_IO_L1_out_wrapper_39__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_39__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_39__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_39__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_39__ap_start = (C_drain_IO_L1_out_wrapper_39__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_40__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_40__is_done__q0 = (C_drain_IO_L1_out_wrapper_40__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_40__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_40__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_40__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_40__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_40__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_40__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_40__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_40__ap_done) begin
            C_drain_IO_L1_out_wrapper_40__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_40__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_40__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_40__ap_done) begin
          C_drain_IO_L1_out_wrapper_40__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_40__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_40__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_40__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_40__ap_start = (C_drain_IO_L1_out_wrapper_40__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_41__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_41__is_done__q0 = (C_drain_IO_L1_out_wrapper_41__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_41__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_41__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_41__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_41__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_41__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_41__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_41__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_41__ap_done) begin
            C_drain_IO_L1_out_wrapper_41__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_41__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_41__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_41__ap_done) begin
          C_drain_IO_L1_out_wrapper_41__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_41__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_41__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_41__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_41__ap_start = (C_drain_IO_L1_out_wrapper_41__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_42__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_42__is_done__q0 = (C_drain_IO_L1_out_wrapper_42__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_42__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_42__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_42__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_42__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_42__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_42__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_42__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_42__ap_done) begin
            C_drain_IO_L1_out_wrapper_42__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_42__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_42__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_42__ap_done) begin
          C_drain_IO_L1_out_wrapper_42__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_42__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_42__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_42__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_42__ap_start = (C_drain_IO_L1_out_wrapper_42__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_43__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_43__is_done__q0 = (C_drain_IO_L1_out_wrapper_43__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_43__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_43__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_43__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_43__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_43__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_43__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_43__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_43__ap_done) begin
            C_drain_IO_L1_out_wrapper_43__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_43__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_43__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_43__ap_done) begin
          C_drain_IO_L1_out_wrapper_43__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_43__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_43__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_43__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_43__ap_start = (C_drain_IO_L1_out_wrapper_43__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_44__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_44__is_done__q0 = (C_drain_IO_L1_out_wrapper_44__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_44__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_44__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_44__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_44__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_44__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_44__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_44__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_44__ap_done) begin
            C_drain_IO_L1_out_wrapper_44__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_44__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_44__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_44__ap_done) begin
          C_drain_IO_L1_out_wrapper_44__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_44__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_44__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_44__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_44__ap_start = (C_drain_IO_L1_out_wrapper_44__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_45__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_45__is_done__q0 = (C_drain_IO_L1_out_wrapper_45__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_45__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_45__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_45__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_45__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_45__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_45__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_45__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_45__ap_done) begin
            C_drain_IO_L1_out_wrapper_45__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_45__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_45__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_45__ap_done) begin
          C_drain_IO_L1_out_wrapper_45__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_45__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_45__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_45__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_45__ap_start = (C_drain_IO_L1_out_wrapper_45__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_46__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_46__is_done__q0 = (C_drain_IO_L1_out_wrapper_46__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_46__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_46__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_46__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_46__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_46__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_46__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_46__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_46__ap_done) begin
            C_drain_IO_L1_out_wrapper_46__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_46__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_46__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_46__ap_done) begin
          C_drain_IO_L1_out_wrapper_46__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_46__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_46__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_46__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_46__ap_start = (C_drain_IO_L1_out_wrapper_46__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_47__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_47__is_done__q0 = (C_drain_IO_L1_out_wrapper_47__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_47__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_47__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_47__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_47__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_47__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_47__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_47__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_47__ap_done) begin
            C_drain_IO_L1_out_wrapper_47__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_47__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_47__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_47__ap_done) begin
          C_drain_IO_L1_out_wrapper_47__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_47__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_47__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_47__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_47__ap_start = (C_drain_IO_L1_out_wrapper_47__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_48__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_48__is_done__q0 = (C_drain_IO_L1_out_wrapper_48__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_48__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_48__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_48__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_48__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_48__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_48__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_48__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_48__ap_done) begin
            C_drain_IO_L1_out_wrapper_48__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_48__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_48__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_48__ap_done) begin
          C_drain_IO_L1_out_wrapper_48__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_48__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_48__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_48__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_48__ap_start = (C_drain_IO_L1_out_wrapper_48__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_49__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_49__is_done__q0 = (C_drain_IO_L1_out_wrapper_49__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_49__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_49__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_49__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_49__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_49__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_49__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_49__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_49__ap_done) begin
            C_drain_IO_L1_out_wrapper_49__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_49__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_49__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_49__ap_done) begin
          C_drain_IO_L1_out_wrapper_49__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_49__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_49__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_49__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_49__ap_start = (C_drain_IO_L1_out_wrapper_49__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_50__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_50__is_done__q0 = (C_drain_IO_L1_out_wrapper_50__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_50__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_50__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_50__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_50__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_50__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_50__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_50__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_50__ap_done) begin
            C_drain_IO_L1_out_wrapper_50__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_50__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_50__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_50__ap_done) begin
          C_drain_IO_L1_out_wrapper_50__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_50__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_50__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_50__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_50__ap_start = (C_drain_IO_L1_out_wrapper_50__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_51__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_51__is_done__q0 = (C_drain_IO_L1_out_wrapper_51__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_51__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_51__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_51__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_51__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_51__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_51__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_51__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_51__ap_done) begin
            C_drain_IO_L1_out_wrapper_51__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_51__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_51__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_51__ap_done) begin
          C_drain_IO_L1_out_wrapper_51__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_51__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_51__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_51__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_51__ap_start = (C_drain_IO_L1_out_wrapper_51__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_52__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_52__is_done__q0 = (C_drain_IO_L1_out_wrapper_52__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_52__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_52__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_52__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_52__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_52__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_52__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_52__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_52__ap_done) begin
            C_drain_IO_L1_out_wrapper_52__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_52__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_52__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_52__ap_done) begin
          C_drain_IO_L1_out_wrapper_52__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_52__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_52__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_52__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_52__ap_start = (C_drain_IO_L1_out_wrapper_52__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_53__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_53__is_done__q0 = (C_drain_IO_L1_out_wrapper_53__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_53__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_53__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_53__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_53__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_53__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_53__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_53__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_53__ap_done) begin
            C_drain_IO_L1_out_wrapper_53__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_53__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_53__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_53__ap_done) begin
          C_drain_IO_L1_out_wrapper_53__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_53__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_53__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_53__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_53__ap_start = (C_drain_IO_L1_out_wrapper_53__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_54__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_54__is_done__q0 = (C_drain_IO_L1_out_wrapper_54__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_54__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_54__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_54__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_54__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_54__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_54__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_54__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_54__ap_done) begin
            C_drain_IO_L1_out_wrapper_54__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_54__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_54__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_54__ap_done) begin
          C_drain_IO_L1_out_wrapper_54__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_54__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_54__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_54__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_54__ap_start = (C_drain_IO_L1_out_wrapper_54__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_55__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_55__is_done__q0 = (C_drain_IO_L1_out_wrapper_55__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_55__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_55__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_55__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_55__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_55__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_55__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_55__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_55__ap_done) begin
            C_drain_IO_L1_out_wrapper_55__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_55__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_55__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_55__ap_done) begin
          C_drain_IO_L1_out_wrapper_55__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_55__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_55__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_55__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_55__ap_start = (C_drain_IO_L1_out_wrapper_55__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_56__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_56__is_done__q0 = (C_drain_IO_L1_out_wrapper_56__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_56__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_56__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_56__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_56__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_56__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_56__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_56__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_56__ap_done) begin
            C_drain_IO_L1_out_wrapper_56__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_56__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_56__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_56__ap_done) begin
          C_drain_IO_L1_out_wrapper_56__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_56__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_56__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_56__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_56__ap_start = (C_drain_IO_L1_out_wrapper_56__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_57__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_57__is_done__q0 = (C_drain_IO_L1_out_wrapper_57__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_57__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_57__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_57__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_57__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_57__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_57__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_57__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_57__ap_done) begin
            C_drain_IO_L1_out_wrapper_57__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_57__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_57__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_57__ap_done) begin
          C_drain_IO_L1_out_wrapper_57__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_57__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_57__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_57__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_57__ap_start = (C_drain_IO_L1_out_wrapper_57__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_58__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_58__is_done__q0 = (C_drain_IO_L1_out_wrapper_58__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_58__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_58__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_58__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_58__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_58__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_58__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_58__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_58__ap_done) begin
            C_drain_IO_L1_out_wrapper_58__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_58__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_58__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_58__ap_done) begin
          C_drain_IO_L1_out_wrapper_58__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_58__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_58__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_58__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_58__ap_start = (C_drain_IO_L1_out_wrapper_58__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_59__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_59__is_done__q0 = (C_drain_IO_L1_out_wrapper_59__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_59__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_59__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_59__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_59__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_59__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_59__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_59__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_59__ap_done) begin
            C_drain_IO_L1_out_wrapper_59__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_59__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_59__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_59__ap_done) begin
          C_drain_IO_L1_out_wrapper_59__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_59__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_59__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_59__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_59__ap_start = (C_drain_IO_L1_out_wrapper_59__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_60__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_60__is_done__q0 = (C_drain_IO_L1_out_wrapper_60__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_60__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_60__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_60__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_60__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_60__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_60__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_60__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_60__ap_done) begin
            C_drain_IO_L1_out_wrapper_60__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_60__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_60__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_60__ap_done) begin
          C_drain_IO_L1_out_wrapper_60__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_60__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_60__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_60__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_60__ap_start = (C_drain_IO_L1_out_wrapper_60__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_61__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_61__is_done__q0 = (C_drain_IO_L1_out_wrapper_61__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_61__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_61__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_61__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_61__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_61__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_61__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_61__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_61__ap_done) begin
            C_drain_IO_L1_out_wrapper_61__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_61__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_61__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_61__ap_done) begin
          C_drain_IO_L1_out_wrapper_61__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_61__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_61__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_61__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_61__ap_start = (C_drain_IO_L1_out_wrapper_61__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_62__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_62__is_done__q0 = (C_drain_IO_L1_out_wrapper_62__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_62__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_62__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_62__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_62__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_62__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_62__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_62__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_62__ap_done) begin
            C_drain_IO_L1_out_wrapper_62__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_62__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_62__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_62__ap_done) begin
          C_drain_IO_L1_out_wrapper_62__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_62__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_62__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_62__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_62__ap_start = (C_drain_IO_L1_out_wrapper_62__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_63__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_63__is_done__q0 = (C_drain_IO_L1_out_wrapper_63__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_63__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_63__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_63__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_63__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_63__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_63__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_63__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_63__ap_done) begin
            C_drain_IO_L1_out_wrapper_63__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_63__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_63__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_63__ap_done) begin
          C_drain_IO_L1_out_wrapper_63__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_63__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_63__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_63__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_63__ap_start = (C_drain_IO_L1_out_wrapper_63__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_64__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_64__is_done__q0 = (C_drain_IO_L1_out_wrapper_64__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_64__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_64__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_64__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_64__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_64__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_64__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_64__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_64__ap_done) begin
            C_drain_IO_L1_out_wrapper_64__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_64__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_64__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_64__ap_done) begin
          C_drain_IO_L1_out_wrapper_64__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_64__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_64__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_64__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_64__ap_start = (C_drain_IO_L1_out_wrapper_64__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_65__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_65__is_done__q0 = (C_drain_IO_L1_out_wrapper_65__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_65__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_65__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_65__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_65__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_65__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_65__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_65__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_65__ap_done) begin
            C_drain_IO_L1_out_wrapper_65__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_65__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_65__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_65__ap_done) begin
          C_drain_IO_L1_out_wrapper_65__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_65__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_65__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_65__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_65__ap_start = (C_drain_IO_L1_out_wrapper_65__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_66__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_66__is_done__q0 = (C_drain_IO_L1_out_wrapper_66__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_66__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_66__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_66__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_66__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_66__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_66__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_66__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_66__ap_done) begin
            C_drain_IO_L1_out_wrapper_66__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_66__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_66__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_66__ap_done) begin
          C_drain_IO_L1_out_wrapper_66__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_66__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_66__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_66__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_66__ap_start = (C_drain_IO_L1_out_wrapper_66__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_67__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_67__is_done__q0 = (C_drain_IO_L1_out_wrapper_67__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_67__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_67__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_67__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_67__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_67__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_67__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_67__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_67__ap_done) begin
            C_drain_IO_L1_out_wrapper_67__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_67__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_67__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_67__ap_done) begin
          C_drain_IO_L1_out_wrapper_67__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_67__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_67__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_67__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_67__ap_start = (C_drain_IO_L1_out_wrapper_67__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_68__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_68__is_done__q0 = (C_drain_IO_L1_out_wrapper_68__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_68__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_68__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_68__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_68__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_68__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_68__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_68__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_68__ap_done) begin
            C_drain_IO_L1_out_wrapper_68__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_68__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_68__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_68__ap_done) begin
          C_drain_IO_L1_out_wrapper_68__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_68__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_68__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_68__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_68__ap_start = (C_drain_IO_L1_out_wrapper_68__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_69__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_69__is_done__q0 = (C_drain_IO_L1_out_wrapper_69__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_69__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_69__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_69__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_69__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_69__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_69__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_69__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_69__ap_done) begin
            C_drain_IO_L1_out_wrapper_69__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_69__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_69__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_69__ap_done) begin
          C_drain_IO_L1_out_wrapper_69__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_69__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_69__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_69__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_69__ap_start = (C_drain_IO_L1_out_wrapper_69__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_70__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_70__is_done__q0 = (C_drain_IO_L1_out_wrapper_70__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_70__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_70__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_70__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_70__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_70__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_70__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_70__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_70__ap_done) begin
            C_drain_IO_L1_out_wrapper_70__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_70__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_70__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_70__ap_done) begin
          C_drain_IO_L1_out_wrapper_70__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_70__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_70__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_70__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_70__ap_start = (C_drain_IO_L1_out_wrapper_70__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_71__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_71__is_done__q0 = (C_drain_IO_L1_out_wrapper_71__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_71__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_71__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_71__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_71__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_71__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_71__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_71__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_71__ap_done) begin
            C_drain_IO_L1_out_wrapper_71__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_71__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_71__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_71__ap_done) begin
          C_drain_IO_L1_out_wrapper_71__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_71__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_71__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_71__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_71__ap_start = (C_drain_IO_L1_out_wrapper_71__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_72__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_72__is_done__q0 = (C_drain_IO_L1_out_wrapper_72__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_72__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_72__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_72__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_72__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_72__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_72__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_72__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_72__ap_done) begin
            C_drain_IO_L1_out_wrapper_72__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_72__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_72__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_72__ap_done) begin
          C_drain_IO_L1_out_wrapper_72__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_72__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_72__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_72__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_72__ap_start = (C_drain_IO_L1_out_wrapper_72__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_73__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_73__is_done__q0 = (C_drain_IO_L1_out_wrapper_73__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_73__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_73__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_73__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_73__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_73__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_73__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_73__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_73__ap_done) begin
            C_drain_IO_L1_out_wrapper_73__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_73__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_73__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_73__ap_done) begin
          C_drain_IO_L1_out_wrapper_73__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_73__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_73__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_73__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_73__ap_start = (C_drain_IO_L1_out_wrapper_73__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_74__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_74__is_done__q0 = (C_drain_IO_L1_out_wrapper_74__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_74__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_74__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_74__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_74__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_74__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_74__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_74__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_74__ap_done) begin
            C_drain_IO_L1_out_wrapper_74__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_74__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_74__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_74__ap_done) begin
          C_drain_IO_L1_out_wrapper_74__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_74__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_74__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_74__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_74__ap_start = (C_drain_IO_L1_out_wrapper_74__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_75__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_75__is_done__q0 = (C_drain_IO_L1_out_wrapper_75__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_75__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_75__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_75__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_75__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_75__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_75__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_75__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_75__ap_done) begin
            C_drain_IO_L1_out_wrapper_75__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_75__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_75__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_75__ap_done) begin
          C_drain_IO_L1_out_wrapper_75__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_75__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_75__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_75__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_75__ap_start = (C_drain_IO_L1_out_wrapper_75__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_76__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_76__is_done__q0 = (C_drain_IO_L1_out_wrapper_76__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_76__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_76__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_76__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_76__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_76__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_76__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_76__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_76__ap_done) begin
            C_drain_IO_L1_out_wrapper_76__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_76__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_76__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_76__ap_done) begin
          C_drain_IO_L1_out_wrapper_76__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_76__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_76__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_76__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_76__ap_start = (C_drain_IO_L1_out_wrapper_76__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_77__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_77__is_done__q0 = (C_drain_IO_L1_out_wrapper_77__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_77__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_77__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_77__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_77__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_77__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_77__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_77__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_77__ap_done) begin
            C_drain_IO_L1_out_wrapper_77__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_77__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_77__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_77__ap_done) begin
          C_drain_IO_L1_out_wrapper_77__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_77__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_77__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_77__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_77__ap_start = (C_drain_IO_L1_out_wrapper_77__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_78__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_78__is_done__q0 = (C_drain_IO_L1_out_wrapper_78__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_78__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_78__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_78__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_78__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_78__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_78__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_78__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_78__ap_done) begin
            C_drain_IO_L1_out_wrapper_78__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_78__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_78__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_78__ap_done) begin
          C_drain_IO_L1_out_wrapper_78__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_78__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_78__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_78__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_78__ap_start = (C_drain_IO_L1_out_wrapper_78__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_79__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_79__is_done__q0 = (C_drain_IO_L1_out_wrapper_79__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_79__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_79__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_79__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_79__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_79__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_79__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_79__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_79__ap_done) begin
            C_drain_IO_L1_out_wrapper_79__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_79__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_79__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_79__ap_done) begin
          C_drain_IO_L1_out_wrapper_79__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_79__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_79__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_79__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_79__ap_start = (C_drain_IO_L1_out_wrapper_79__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_80__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_80__is_done__q0 = (C_drain_IO_L1_out_wrapper_80__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_80__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_80__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_80__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_80__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_80__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_80__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_80__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_80__ap_done) begin
            C_drain_IO_L1_out_wrapper_80__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_80__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_80__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_80__ap_done) begin
          C_drain_IO_L1_out_wrapper_80__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_80__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_80__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_80__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_80__ap_start = (C_drain_IO_L1_out_wrapper_80__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_81__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_81__is_done__q0 = (C_drain_IO_L1_out_wrapper_81__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_81__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_81__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_81__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_81__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_81__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_81__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_81__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_81__ap_done) begin
            C_drain_IO_L1_out_wrapper_81__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_81__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_81__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_81__ap_done) begin
          C_drain_IO_L1_out_wrapper_81__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_81__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_81__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_81__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_81__ap_start = (C_drain_IO_L1_out_wrapper_81__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_82__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_82__is_done__q0 = (C_drain_IO_L1_out_wrapper_82__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_82__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_82__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_82__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_82__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_82__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_82__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_82__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_82__ap_done) begin
            C_drain_IO_L1_out_wrapper_82__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_82__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_82__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_82__ap_done) begin
          C_drain_IO_L1_out_wrapper_82__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_82__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_82__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_82__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_82__ap_start = (C_drain_IO_L1_out_wrapper_82__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_83__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_83__is_done__q0 = (C_drain_IO_L1_out_wrapper_83__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_83__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_83__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_83__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_83__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_83__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_83__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_83__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_83__ap_done) begin
            C_drain_IO_L1_out_wrapper_83__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_83__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_83__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_83__ap_done) begin
          C_drain_IO_L1_out_wrapper_83__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_83__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_83__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_83__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_83__ap_start = (C_drain_IO_L1_out_wrapper_83__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_84__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_84__is_done__q0 = (C_drain_IO_L1_out_wrapper_84__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_84__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_84__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_84__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_84__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_84__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_84__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_84__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_84__ap_done) begin
            C_drain_IO_L1_out_wrapper_84__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_84__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_84__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_84__ap_done) begin
          C_drain_IO_L1_out_wrapper_84__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_84__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_84__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_84__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_84__ap_start = (C_drain_IO_L1_out_wrapper_84__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_85__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_85__is_done__q0 = (C_drain_IO_L1_out_wrapper_85__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_85__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_85__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_85__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_85__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_85__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_85__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_85__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_85__ap_done) begin
            C_drain_IO_L1_out_wrapper_85__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_85__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_85__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_85__ap_done) begin
          C_drain_IO_L1_out_wrapper_85__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_85__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_85__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_85__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_85__ap_start = (C_drain_IO_L1_out_wrapper_85__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_86__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_86__is_done__q0 = (C_drain_IO_L1_out_wrapper_86__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_86__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_86__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_86__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_86__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_86__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_86__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_86__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_86__ap_done) begin
            C_drain_IO_L1_out_wrapper_86__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_86__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_86__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_86__ap_done) begin
          C_drain_IO_L1_out_wrapper_86__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_86__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_86__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_86__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_86__ap_start = (C_drain_IO_L1_out_wrapper_86__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_87__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_87__is_done__q0 = (C_drain_IO_L1_out_wrapper_87__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_87__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_87__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_87__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_87__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_87__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_87__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_87__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_87__ap_done) begin
            C_drain_IO_L1_out_wrapper_87__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_87__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_87__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_87__ap_done) begin
          C_drain_IO_L1_out_wrapper_87__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_87__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_87__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_87__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_87__ap_start = (C_drain_IO_L1_out_wrapper_87__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_88__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_88__is_done__q0 = (C_drain_IO_L1_out_wrapper_88__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_88__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_88__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_88__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_88__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_88__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_88__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_88__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_88__ap_done) begin
            C_drain_IO_L1_out_wrapper_88__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_88__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_88__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_88__ap_done) begin
          C_drain_IO_L1_out_wrapper_88__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_88__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_88__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_88__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_88__ap_start = (C_drain_IO_L1_out_wrapper_88__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_89__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_89__is_done__q0 = (C_drain_IO_L1_out_wrapper_89__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_89__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_89__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_89__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_89__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_89__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_89__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_89__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_89__ap_done) begin
            C_drain_IO_L1_out_wrapper_89__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_89__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_89__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_89__ap_done) begin
          C_drain_IO_L1_out_wrapper_89__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_89__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_89__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_89__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_89__ap_start = (C_drain_IO_L1_out_wrapper_89__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_90__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_90__is_done__q0 = (C_drain_IO_L1_out_wrapper_90__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_90__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_90__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_90__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_90__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_90__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_90__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_90__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_90__ap_done) begin
            C_drain_IO_L1_out_wrapper_90__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_90__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_90__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_90__ap_done) begin
          C_drain_IO_L1_out_wrapper_90__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_90__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_90__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_90__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_90__ap_start = (C_drain_IO_L1_out_wrapper_90__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_91__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_91__is_done__q0 = (C_drain_IO_L1_out_wrapper_91__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_91__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_91__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_91__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_91__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_91__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_91__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_91__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_91__ap_done) begin
            C_drain_IO_L1_out_wrapper_91__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_91__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_91__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_91__ap_done) begin
          C_drain_IO_L1_out_wrapper_91__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_91__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_91__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_91__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_91__ap_start = (C_drain_IO_L1_out_wrapper_91__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_92__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_92__is_done__q0 = (C_drain_IO_L1_out_wrapper_92__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_92__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_92__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_92__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_92__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_92__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_92__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_92__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_92__ap_done) begin
            C_drain_IO_L1_out_wrapper_92__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_92__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_92__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_92__ap_done) begin
          C_drain_IO_L1_out_wrapper_92__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_92__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_92__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_92__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_92__ap_start = (C_drain_IO_L1_out_wrapper_92__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_93__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_93__is_done__q0 = (C_drain_IO_L1_out_wrapper_93__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_93__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_93__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_93__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_93__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_93__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_93__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_93__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_93__ap_done) begin
            C_drain_IO_L1_out_wrapper_93__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_93__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_93__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_93__ap_done) begin
          C_drain_IO_L1_out_wrapper_93__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_93__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_93__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_93__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_93__ap_start = (C_drain_IO_L1_out_wrapper_93__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_94__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_94__is_done__q0 = (C_drain_IO_L1_out_wrapper_94__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_94__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_94__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_94__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_94__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_94__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_94__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_94__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_94__ap_done) begin
            C_drain_IO_L1_out_wrapper_94__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_94__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_94__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_94__ap_done) begin
          C_drain_IO_L1_out_wrapper_94__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_94__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_94__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_94__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_94__ap_start = (C_drain_IO_L1_out_wrapper_94__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_95__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_95__is_done__q0 = (C_drain_IO_L1_out_wrapper_95__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_95__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_95__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_95__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_95__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_95__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_95__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_95__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_95__ap_done) begin
            C_drain_IO_L1_out_wrapper_95__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_95__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_95__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_95__ap_done) begin
          C_drain_IO_L1_out_wrapper_95__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_95__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_95__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_95__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_95__ap_start = (C_drain_IO_L1_out_wrapper_95__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_96__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_96__is_done__q0 = (C_drain_IO_L1_out_wrapper_96__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_96__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_96__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_96__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_96__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_96__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_96__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_96__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_96__ap_done) begin
            C_drain_IO_L1_out_wrapper_96__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_96__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_96__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_96__ap_done) begin
          C_drain_IO_L1_out_wrapper_96__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_96__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_96__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_96__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_96__ap_start = (C_drain_IO_L1_out_wrapper_96__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_97__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_97__is_done__q0 = (C_drain_IO_L1_out_wrapper_97__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_97__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_97__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_97__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_97__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_97__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_97__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_97__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_97__ap_done) begin
            C_drain_IO_L1_out_wrapper_97__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_97__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_97__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_97__ap_done) begin
          C_drain_IO_L1_out_wrapper_97__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_97__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_97__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_97__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_97__ap_start = (C_drain_IO_L1_out_wrapper_97__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_98__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_98__is_done__q0 = (C_drain_IO_L1_out_wrapper_98__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_98__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_98__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_98__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_98__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_98__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_98__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_98__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_98__ap_done) begin
            C_drain_IO_L1_out_wrapper_98__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_98__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_98__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_98__ap_done) begin
          C_drain_IO_L1_out_wrapper_98__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_98__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_98__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_98__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_98__ap_start = (C_drain_IO_L1_out_wrapper_98__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_99__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_99__is_done__q0 = (C_drain_IO_L1_out_wrapper_99__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_99__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_99__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_99__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_99__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_99__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_99__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_99__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_99__ap_done) begin
            C_drain_IO_L1_out_wrapper_99__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_99__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_99__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_99__ap_done) begin
          C_drain_IO_L1_out_wrapper_99__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_99__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_99__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_99__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_99__ap_start = (C_drain_IO_L1_out_wrapper_99__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_100__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_100__is_done__q0 = (C_drain_IO_L1_out_wrapper_100__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_100__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_100__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_100__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_100__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_100__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_100__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_100__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_100__ap_done) begin
            C_drain_IO_L1_out_wrapper_100__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_100__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_100__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_100__ap_done) begin
          C_drain_IO_L1_out_wrapper_100__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_100__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_100__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_100__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_100__ap_start = (C_drain_IO_L1_out_wrapper_100__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_101__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_101__is_done__q0 = (C_drain_IO_L1_out_wrapper_101__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_101__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_101__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_101__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_101__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_101__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_101__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_101__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_101__ap_done) begin
            C_drain_IO_L1_out_wrapper_101__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_101__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_101__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_101__ap_done) begin
          C_drain_IO_L1_out_wrapper_101__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_101__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_101__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_101__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_101__ap_start = (C_drain_IO_L1_out_wrapper_101__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_102__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_102__is_done__q0 = (C_drain_IO_L1_out_wrapper_102__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_102__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_102__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_102__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_102__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_102__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_102__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_102__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_102__ap_done) begin
            C_drain_IO_L1_out_wrapper_102__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_102__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_102__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_102__ap_done) begin
          C_drain_IO_L1_out_wrapper_102__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_102__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_102__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_102__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_102__ap_start = (C_drain_IO_L1_out_wrapper_102__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_103__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_103__is_done__q0 = (C_drain_IO_L1_out_wrapper_103__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_103__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_103__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_103__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_103__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_103__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_103__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_103__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_103__ap_done) begin
            C_drain_IO_L1_out_wrapper_103__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_103__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_103__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_103__ap_done) begin
          C_drain_IO_L1_out_wrapper_103__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_103__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_103__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_103__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_103__ap_start = (C_drain_IO_L1_out_wrapper_103__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_104__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_104__is_done__q0 = (C_drain_IO_L1_out_wrapper_104__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_104__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_104__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_104__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_104__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_104__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_104__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_104__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_104__ap_done) begin
            C_drain_IO_L1_out_wrapper_104__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_104__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_104__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_104__ap_done) begin
          C_drain_IO_L1_out_wrapper_104__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_104__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_104__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_104__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_104__ap_start = (C_drain_IO_L1_out_wrapper_104__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_105__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_105__is_done__q0 = (C_drain_IO_L1_out_wrapper_105__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_105__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_105__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_105__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_105__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_105__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_105__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_105__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_105__ap_done) begin
            C_drain_IO_L1_out_wrapper_105__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_105__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_105__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_105__ap_done) begin
          C_drain_IO_L1_out_wrapper_105__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_105__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_105__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_105__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_105__ap_start = (C_drain_IO_L1_out_wrapper_105__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_106__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_106__is_done__q0 = (C_drain_IO_L1_out_wrapper_106__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_106__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_106__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_106__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_106__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_106__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_106__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_106__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_106__ap_done) begin
            C_drain_IO_L1_out_wrapper_106__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_106__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_106__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_106__ap_done) begin
          C_drain_IO_L1_out_wrapper_106__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_106__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_106__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_106__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_106__ap_start = (C_drain_IO_L1_out_wrapper_106__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_107__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_107__is_done__q0 = (C_drain_IO_L1_out_wrapper_107__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_107__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_107__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_107__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_107__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_107__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_107__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_107__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_107__ap_done) begin
            C_drain_IO_L1_out_wrapper_107__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_107__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_107__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_107__ap_done) begin
          C_drain_IO_L1_out_wrapper_107__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_107__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_107__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_107__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_107__ap_start = (C_drain_IO_L1_out_wrapper_107__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_108__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_108__is_done__q0 = (C_drain_IO_L1_out_wrapper_108__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_108__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_108__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_108__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_108__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_108__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_108__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_108__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_108__ap_done) begin
            C_drain_IO_L1_out_wrapper_108__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_108__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_108__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_108__ap_done) begin
          C_drain_IO_L1_out_wrapper_108__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_108__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_108__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_108__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_108__ap_start = (C_drain_IO_L1_out_wrapper_108__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_109__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_109__is_done__q0 = (C_drain_IO_L1_out_wrapper_109__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_109__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_109__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_109__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_109__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_109__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_109__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_109__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_109__ap_done) begin
            C_drain_IO_L1_out_wrapper_109__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_109__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_109__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_109__ap_done) begin
          C_drain_IO_L1_out_wrapper_109__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_109__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_109__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_109__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_109__ap_start = (C_drain_IO_L1_out_wrapper_109__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_110__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_110__is_done__q0 = (C_drain_IO_L1_out_wrapper_110__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_110__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_110__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_110__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_110__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_110__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_110__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_110__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_110__ap_done) begin
            C_drain_IO_L1_out_wrapper_110__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_110__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_110__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_110__ap_done) begin
          C_drain_IO_L1_out_wrapper_110__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_110__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_110__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_110__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_110__ap_start = (C_drain_IO_L1_out_wrapper_110__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_111__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_111__is_done__q0 = (C_drain_IO_L1_out_wrapper_111__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_111__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_111__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_111__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_111__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_111__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_111__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_111__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_111__ap_done) begin
            C_drain_IO_L1_out_wrapper_111__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_111__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_111__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_111__ap_done) begin
          C_drain_IO_L1_out_wrapper_111__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_111__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_111__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_111__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_111__ap_start = (C_drain_IO_L1_out_wrapper_111__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_112__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_112__is_done__q0 = (C_drain_IO_L1_out_wrapper_112__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_112__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_112__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_112__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_112__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_112__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_112__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_112__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_112__ap_done) begin
            C_drain_IO_L1_out_wrapper_112__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_112__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_112__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_112__ap_done) begin
          C_drain_IO_L1_out_wrapper_112__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_112__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_112__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_112__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_112__ap_start = (C_drain_IO_L1_out_wrapper_112__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_113__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_113__is_done__q0 = (C_drain_IO_L1_out_wrapper_113__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_113__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_113__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_113__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_113__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_113__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_113__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_113__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_113__ap_done) begin
            C_drain_IO_L1_out_wrapper_113__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_113__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_113__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_113__ap_done) begin
          C_drain_IO_L1_out_wrapper_113__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_113__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_113__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_113__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_113__ap_start = (C_drain_IO_L1_out_wrapper_113__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_114__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_114__is_done__q0 = (C_drain_IO_L1_out_wrapper_114__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_114__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_114__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_114__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_114__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_114__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_114__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_114__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_114__ap_done) begin
            C_drain_IO_L1_out_wrapper_114__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_114__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_114__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_114__ap_done) begin
          C_drain_IO_L1_out_wrapper_114__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_114__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_114__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_114__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_114__ap_start = (C_drain_IO_L1_out_wrapper_114__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_115__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_115__is_done__q0 = (C_drain_IO_L1_out_wrapper_115__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_115__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_115__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_115__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_115__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_115__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_115__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_115__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_115__ap_done) begin
            C_drain_IO_L1_out_wrapper_115__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_115__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_115__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_115__ap_done) begin
          C_drain_IO_L1_out_wrapper_115__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_115__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_115__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_115__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_115__ap_start = (C_drain_IO_L1_out_wrapper_115__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_116__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_116__is_done__q0 = (C_drain_IO_L1_out_wrapper_116__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_116__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_116__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_116__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_116__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_116__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_116__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_116__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_116__ap_done) begin
            C_drain_IO_L1_out_wrapper_116__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_116__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_116__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_116__ap_done) begin
          C_drain_IO_L1_out_wrapper_116__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_116__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_116__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_116__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_116__ap_start = (C_drain_IO_L1_out_wrapper_116__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_117__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_117__is_done__q0 = (C_drain_IO_L1_out_wrapper_117__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_117__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_117__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_117__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_117__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_117__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_117__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_117__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_117__ap_done) begin
            C_drain_IO_L1_out_wrapper_117__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_117__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_117__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_117__ap_done) begin
          C_drain_IO_L1_out_wrapper_117__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_117__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_117__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_117__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_117__ap_start = (C_drain_IO_L1_out_wrapper_117__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_118__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_118__is_done__q0 = (C_drain_IO_L1_out_wrapper_118__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_118__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_118__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_118__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_118__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_118__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_118__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_118__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_118__ap_done) begin
            C_drain_IO_L1_out_wrapper_118__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_118__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_118__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_118__ap_done) begin
          C_drain_IO_L1_out_wrapper_118__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_118__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_118__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_118__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_118__ap_start = (C_drain_IO_L1_out_wrapper_118__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_119__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_119__is_done__q0 = (C_drain_IO_L1_out_wrapper_119__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_119__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_119__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_119__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_119__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_119__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_119__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_119__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_119__ap_done) begin
            C_drain_IO_L1_out_wrapper_119__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_119__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_119__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_119__ap_done) begin
          C_drain_IO_L1_out_wrapper_119__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_119__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_119__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_119__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_119__ap_start = (C_drain_IO_L1_out_wrapper_119__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_120__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_120__is_done__q0 = (C_drain_IO_L1_out_wrapper_120__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_120__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_120__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_120__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_120__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_120__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_120__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_120__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_120__ap_done) begin
            C_drain_IO_L1_out_wrapper_120__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_120__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_120__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_120__ap_done) begin
          C_drain_IO_L1_out_wrapper_120__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_120__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_120__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_120__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_120__ap_start = (C_drain_IO_L1_out_wrapper_120__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_121__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_121__is_done__q0 = (C_drain_IO_L1_out_wrapper_121__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_121__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_121__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_121__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_121__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_121__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_121__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_121__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_121__ap_done) begin
            C_drain_IO_L1_out_wrapper_121__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_121__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_121__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_121__ap_done) begin
          C_drain_IO_L1_out_wrapper_121__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_121__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_121__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_121__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_121__ap_start = (C_drain_IO_L1_out_wrapper_121__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_122__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_122__is_done__q0 = (C_drain_IO_L1_out_wrapper_122__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_122__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_122__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_122__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_122__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_122__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_122__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_122__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_122__ap_done) begin
            C_drain_IO_L1_out_wrapper_122__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_122__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_122__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_122__ap_done) begin
          C_drain_IO_L1_out_wrapper_122__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_122__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_122__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_122__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_122__ap_start = (C_drain_IO_L1_out_wrapper_122__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_123__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_123__is_done__q0 = (C_drain_IO_L1_out_wrapper_123__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_123__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_123__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_123__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_123__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_123__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_123__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_123__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_123__ap_done) begin
            C_drain_IO_L1_out_wrapper_123__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_123__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_123__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_123__ap_done) begin
          C_drain_IO_L1_out_wrapper_123__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_123__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_123__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_123__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_123__ap_start = (C_drain_IO_L1_out_wrapper_123__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_124__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_124__is_done__q0 = (C_drain_IO_L1_out_wrapper_124__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_124__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_124__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_124__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_124__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_124__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_124__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_124__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_124__ap_done) begin
            C_drain_IO_L1_out_wrapper_124__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_124__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_124__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_124__ap_done) begin
          C_drain_IO_L1_out_wrapper_124__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_124__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_124__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_124__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_124__ap_start = (C_drain_IO_L1_out_wrapper_124__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_125__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_125__is_done__q0 = (C_drain_IO_L1_out_wrapper_125__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_125__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_125__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_125__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_125__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_125__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_125__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_125__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_125__ap_done) begin
            C_drain_IO_L1_out_wrapper_125__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_125__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_125__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_125__ap_done) begin
          C_drain_IO_L1_out_wrapper_125__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_125__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_125__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_125__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_125__ap_start = (C_drain_IO_L1_out_wrapper_125__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_126__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_126__is_done__q0 = (C_drain_IO_L1_out_wrapper_126__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_126__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_126__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_126__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_126__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_126__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_126__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_126__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_126__ap_done) begin
            C_drain_IO_L1_out_wrapper_126__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_126__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_126__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_126__ap_done) begin
          C_drain_IO_L1_out_wrapper_126__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_126__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_126__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_126__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_126__ap_start = (C_drain_IO_L1_out_wrapper_126__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_127__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_127__is_done__q0 = (C_drain_IO_L1_out_wrapper_127__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_127__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_127__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_127__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_127__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_127__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_127__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_127__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_127__ap_done) begin
            C_drain_IO_L1_out_wrapper_127__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_127__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_127__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_127__ap_done) begin
          C_drain_IO_L1_out_wrapper_127__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_127__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_127__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_127__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_127__ap_start = (C_drain_IO_L1_out_wrapper_127__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_128__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_128__is_done__q0 = (C_drain_IO_L1_out_wrapper_128__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_128__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_128__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_128__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_128__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_128__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_128__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_128__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_128__ap_done) begin
            C_drain_IO_L1_out_wrapper_128__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_128__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_128__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_128__ap_done) begin
          C_drain_IO_L1_out_wrapper_128__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_128__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_128__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_128__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_128__ap_start = (C_drain_IO_L1_out_wrapper_128__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_129__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_129__is_done__q0 = (C_drain_IO_L1_out_wrapper_129__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_129__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_129__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_129__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_129__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_129__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_129__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_129__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_129__ap_done) begin
            C_drain_IO_L1_out_wrapper_129__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_129__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_129__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_129__ap_done) begin
          C_drain_IO_L1_out_wrapper_129__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_129__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_129__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_129__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_129__ap_start = (C_drain_IO_L1_out_wrapper_129__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_130__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_130__is_done__q0 = (C_drain_IO_L1_out_wrapper_130__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_130__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_130__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_130__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_130__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_130__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_130__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_130__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_130__ap_done) begin
            C_drain_IO_L1_out_wrapper_130__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_130__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_130__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_130__ap_done) begin
          C_drain_IO_L1_out_wrapper_130__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_130__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_130__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_130__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_130__ap_start = (C_drain_IO_L1_out_wrapper_130__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_131__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_131__is_done__q0 = (C_drain_IO_L1_out_wrapper_131__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_131__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_131__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_131__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_131__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_131__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_131__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_131__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_131__ap_done) begin
            C_drain_IO_L1_out_wrapper_131__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_131__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_131__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_131__ap_done) begin
          C_drain_IO_L1_out_wrapper_131__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_131__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_131__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_131__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_131__ap_start = (C_drain_IO_L1_out_wrapper_131__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_132__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_132__is_done__q0 = (C_drain_IO_L1_out_wrapper_132__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_132__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_132__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_132__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_132__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_132__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_132__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_132__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_132__ap_done) begin
            C_drain_IO_L1_out_wrapper_132__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_132__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_132__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_132__ap_done) begin
          C_drain_IO_L1_out_wrapper_132__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_132__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_132__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_132__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_132__ap_start = (C_drain_IO_L1_out_wrapper_132__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_133__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_133__is_done__q0 = (C_drain_IO_L1_out_wrapper_133__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_133__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_133__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_133__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_133__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_133__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_133__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_133__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_133__ap_done) begin
            C_drain_IO_L1_out_wrapper_133__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_133__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_133__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_133__ap_done) begin
          C_drain_IO_L1_out_wrapper_133__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_133__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_133__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_133__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_133__ap_start = (C_drain_IO_L1_out_wrapper_133__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_134__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_134__is_done__q0 = (C_drain_IO_L1_out_wrapper_134__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_134__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_134__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_134__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_134__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_134__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_134__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_134__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_134__ap_done) begin
            C_drain_IO_L1_out_wrapper_134__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_134__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_134__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_134__ap_done) begin
          C_drain_IO_L1_out_wrapper_134__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_134__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_134__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_134__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_134__ap_start = (C_drain_IO_L1_out_wrapper_134__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_135__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_135__is_done__q0 = (C_drain_IO_L1_out_wrapper_135__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_135__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_135__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_135__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_135__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_135__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_135__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_135__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_135__ap_done) begin
            C_drain_IO_L1_out_wrapper_135__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_135__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_135__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_135__ap_done) begin
          C_drain_IO_L1_out_wrapper_135__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_135__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_135__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_135__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_135__ap_start = (C_drain_IO_L1_out_wrapper_135__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_136__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_136__is_done__q0 = (C_drain_IO_L1_out_wrapper_136__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_136__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_136__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_136__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_136__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_136__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_136__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_136__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_136__ap_done) begin
            C_drain_IO_L1_out_wrapper_136__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_136__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_136__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_136__ap_done) begin
          C_drain_IO_L1_out_wrapper_136__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_136__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_136__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_136__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_136__ap_start = (C_drain_IO_L1_out_wrapper_136__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_137__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_137__is_done__q0 = (C_drain_IO_L1_out_wrapper_137__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_137__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_137__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_137__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_137__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_137__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_137__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_137__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_137__ap_done) begin
            C_drain_IO_L1_out_wrapper_137__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_137__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_137__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_137__ap_done) begin
          C_drain_IO_L1_out_wrapper_137__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_137__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_137__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_137__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_137__ap_start = (C_drain_IO_L1_out_wrapper_137__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_138__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_138__is_done__q0 = (C_drain_IO_L1_out_wrapper_138__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_138__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_138__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_138__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_138__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_138__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_138__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_138__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_138__ap_done) begin
            C_drain_IO_L1_out_wrapper_138__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_138__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_138__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_138__ap_done) begin
          C_drain_IO_L1_out_wrapper_138__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_138__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_138__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_138__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_138__ap_start = (C_drain_IO_L1_out_wrapper_138__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_139__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_139__is_done__q0 = (C_drain_IO_L1_out_wrapper_139__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_139__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_139__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_139__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_139__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_139__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_139__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_139__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_139__ap_done) begin
            C_drain_IO_L1_out_wrapper_139__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_139__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_139__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_139__ap_done) begin
          C_drain_IO_L1_out_wrapper_139__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_139__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_139__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_139__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_139__ap_start = (C_drain_IO_L1_out_wrapper_139__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_140__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_140__is_done__q0 = (C_drain_IO_L1_out_wrapper_140__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_140__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_140__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_140__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_140__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_140__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_140__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_140__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_140__ap_done) begin
            C_drain_IO_L1_out_wrapper_140__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_140__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_140__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_140__ap_done) begin
          C_drain_IO_L1_out_wrapper_140__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_140__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_140__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_140__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_140__ap_start = (C_drain_IO_L1_out_wrapper_140__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_141__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_141__is_done__q0 = (C_drain_IO_L1_out_wrapper_141__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_141__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_141__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_141__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_141__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_141__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_141__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_141__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_141__ap_done) begin
            C_drain_IO_L1_out_wrapper_141__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_141__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_141__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_141__ap_done) begin
          C_drain_IO_L1_out_wrapper_141__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_141__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_141__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_141__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_141__ap_start = (C_drain_IO_L1_out_wrapper_141__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_142__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_142__is_done__q0 = (C_drain_IO_L1_out_wrapper_142__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_142__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_142__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_142__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_142__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_142__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_142__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_142__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_142__ap_done) begin
            C_drain_IO_L1_out_wrapper_142__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_142__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_142__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_142__ap_done) begin
          C_drain_IO_L1_out_wrapper_142__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_142__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_142__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_142__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_142__ap_start = (C_drain_IO_L1_out_wrapper_142__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_143__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_143__is_done__q0 = (C_drain_IO_L1_out_wrapper_143__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_143__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_143__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_143__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_143__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_143__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_143__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_143__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_143__ap_done) begin
            C_drain_IO_L1_out_wrapper_143__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_143__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_143__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_143__ap_done) begin
          C_drain_IO_L1_out_wrapper_143__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_143__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_143__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_143__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_143__ap_start = (C_drain_IO_L1_out_wrapper_143__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_144__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_144__is_done__q0 = (C_drain_IO_L1_out_wrapper_144__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_144__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_144__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_144__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_144__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_144__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_144__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_144__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_144__ap_done) begin
            C_drain_IO_L1_out_wrapper_144__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_144__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_144__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_144__ap_done) begin
          C_drain_IO_L1_out_wrapper_144__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_144__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_144__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_144__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_144__ap_start = (C_drain_IO_L1_out_wrapper_144__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_145__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_145__is_done__q0 = (C_drain_IO_L1_out_wrapper_145__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_145__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_145__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_145__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_145__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_145__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_145__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_145__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_145__ap_done) begin
            C_drain_IO_L1_out_wrapper_145__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_145__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_145__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_145__ap_done) begin
          C_drain_IO_L1_out_wrapper_145__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_145__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_145__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_145__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_145__ap_start = (C_drain_IO_L1_out_wrapper_145__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_146__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_146__is_done__q0 = (C_drain_IO_L1_out_wrapper_146__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_146__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_146__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_146__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_146__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_146__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_146__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_146__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_146__ap_done) begin
            C_drain_IO_L1_out_wrapper_146__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_146__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_146__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_146__ap_done) begin
          C_drain_IO_L1_out_wrapper_146__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_146__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_146__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_146__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_146__ap_start = (C_drain_IO_L1_out_wrapper_146__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_147__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_147__is_done__q0 = (C_drain_IO_L1_out_wrapper_147__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_147__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_147__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_147__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_147__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_147__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_147__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_147__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_147__ap_done) begin
            C_drain_IO_L1_out_wrapper_147__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_147__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_147__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_147__ap_done) begin
          C_drain_IO_L1_out_wrapper_147__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_147__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_147__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_147__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_147__ap_start = (C_drain_IO_L1_out_wrapper_147__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_148__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_148__is_done__q0 = (C_drain_IO_L1_out_wrapper_148__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_148__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_148__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_148__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_148__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_148__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_148__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_148__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_148__ap_done) begin
            C_drain_IO_L1_out_wrapper_148__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_148__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_148__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_148__ap_done) begin
          C_drain_IO_L1_out_wrapper_148__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_148__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_148__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_148__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_148__ap_start = (C_drain_IO_L1_out_wrapper_148__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_149__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_149__is_done__q0 = (C_drain_IO_L1_out_wrapper_149__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_149__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_149__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_149__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_149__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_149__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_149__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_149__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_149__ap_done) begin
            C_drain_IO_L1_out_wrapper_149__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_149__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_149__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_149__ap_done) begin
          C_drain_IO_L1_out_wrapper_149__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_149__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_149__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_149__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_149__ap_start = (C_drain_IO_L1_out_wrapper_149__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_150__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_150__is_done__q0 = (C_drain_IO_L1_out_wrapper_150__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_150__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_150__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_150__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_150__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_150__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_150__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_150__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_150__ap_done) begin
            C_drain_IO_L1_out_wrapper_150__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_150__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_150__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_150__ap_done) begin
          C_drain_IO_L1_out_wrapper_150__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_150__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_150__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_150__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_150__ap_start = (C_drain_IO_L1_out_wrapper_150__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_151__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_151__is_done__q0 = (C_drain_IO_L1_out_wrapper_151__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_151__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_151__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_151__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_151__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_151__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_151__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_151__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_151__ap_done) begin
            C_drain_IO_L1_out_wrapper_151__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_151__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_151__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_151__ap_done) begin
          C_drain_IO_L1_out_wrapper_151__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_151__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_151__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_151__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_151__ap_start = (C_drain_IO_L1_out_wrapper_151__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_152__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_152__is_done__q0 = (C_drain_IO_L1_out_wrapper_152__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_152__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_152__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_152__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_152__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_152__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_152__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_152__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_152__ap_done) begin
            C_drain_IO_L1_out_wrapper_152__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_152__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_152__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_152__ap_done) begin
          C_drain_IO_L1_out_wrapper_152__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_152__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_152__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_152__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_152__ap_start = (C_drain_IO_L1_out_wrapper_152__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_153__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_153__is_done__q0 = (C_drain_IO_L1_out_wrapper_153__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_153__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_153__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_153__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_153__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_153__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_153__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_153__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_153__ap_done) begin
            C_drain_IO_L1_out_wrapper_153__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_153__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_153__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_153__ap_done) begin
          C_drain_IO_L1_out_wrapper_153__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_153__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_153__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_153__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_153__ap_start = (C_drain_IO_L1_out_wrapper_153__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_154__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_154__is_done__q0 = (C_drain_IO_L1_out_wrapper_154__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_154__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_154__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_154__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_154__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_154__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_154__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_154__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_154__ap_done) begin
            C_drain_IO_L1_out_wrapper_154__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_154__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_154__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_154__ap_done) begin
          C_drain_IO_L1_out_wrapper_154__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_154__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_154__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_154__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_154__ap_start = (C_drain_IO_L1_out_wrapper_154__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_155__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_155__is_done__q0 = (C_drain_IO_L1_out_wrapper_155__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_155__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_155__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_155__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_155__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_155__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_155__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_155__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_155__ap_done) begin
            C_drain_IO_L1_out_wrapper_155__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_155__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_155__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_155__ap_done) begin
          C_drain_IO_L1_out_wrapper_155__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_155__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_155__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_155__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_155__ap_start = (C_drain_IO_L1_out_wrapper_155__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_156__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_156__is_done__q0 = (C_drain_IO_L1_out_wrapper_156__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_156__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_156__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_156__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_156__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_156__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_156__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_156__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_156__ap_done) begin
            C_drain_IO_L1_out_wrapper_156__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_156__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_156__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_156__ap_done) begin
          C_drain_IO_L1_out_wrapper_156__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_156__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_156__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_156__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_156__ap_start = (C_drain_IO_L1_out_wrapper_156__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_157__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_157__is_done__q0 = (C_drain_IO_L1_out_wrapper_157__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_157__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_157__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_157__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_157__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_157__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_157__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_157__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_157__ap_done) begin
            C_drain_IO_L1_out_wrapper_157__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_157__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_157__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_157__ap_done) begin
          C_drain_IO_L1_out_wrapper_157__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_157__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_157__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_157__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_157__ap_start = (C_drain_IO_L1_out_wrapper_157__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_158__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_158__is_done__q0 = (C_drain_IO_L1_out_wrapper_158__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_158__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_158__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_158__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_158__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_158__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_158__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_158__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_158__ap_done) begin
            C_drain_IO_L1_out_wrapper_158__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_158__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_158__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_158__ap_done) begin
          C_drain_IO_L1_out_wrapper_158__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_158__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_158__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_158__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_158__ap_start = (C_drain_IO_L1_out_wrapper_158__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_159__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_159__is_done__q0 = (C_drain_IO_L1_out_wrapper_159__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_159__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_159__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_159__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_159__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_159__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_159__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_159__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_159__ap_done) begin
            C_drain_IO_L1_out_wrapper_159__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_159__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_159__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_159__ap_done) begin
          C_drain_IO_L1_out_wrapper_159__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_159__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_159__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_159__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_159__ap_start = (C_drain_IO_L1_out_wrapper_159__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_160__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_160__is_done__q0 = (C_drain_IO_L1_out_wrapper_160__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_160__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_160__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_160__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_160__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_160__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_160__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_160__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_160__ap_done) begin
            C_drain_IO_L1_out_wrapper_160__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_160__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_160__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_160__ap_done) begin
          C_drain_IO_L1_out_wrapper_160__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_160__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_160__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_160__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_160__ap_start = (C_drain_IO_L1_out_wrapper_160__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_161__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_161__is_done__q0 = (C_drain_IO_L1_out_wrapper_161__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_161__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_161__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_161__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_161__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_161__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_161__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_161__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_161__ap_done) begin
            C_drain_IO_L1_out_wrapper_161__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_161__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_161__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_161__ap_done) begin
          C_drain_IO_L1_out_wrapper_161__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_161__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_161__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_161__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_161__ap_start = (C_drain_IO_L1_out_wrapper_161__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_162__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_162__is_done__q0 = (C_drain_IO_L1_out_wrapper_162__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_162__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_162__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_162__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_162__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_162__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_162__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_162__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_162__ap_done) begin
            C_drain_IO_L1_out_wrapper_162__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_162__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_162__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_162__ap_done) begin
          C_drain_IO_L1_out_wrapper_162__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_162__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_162__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_162__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_162__ap_start = (C_drain_IO_L1_out_wrapper_162__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_163__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_163__is_done__q0 = (C_drain_IO_L1_out_wrapper_163__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_163__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_163__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_163__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_163__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_163__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_163__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_163__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_163__ap_done) begin
            C_drain_IO_L1_out_wrapper_163__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_163__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_163__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_163__ap_done) begin
          C_drain_IO_L1_out_wrapper_163__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_163__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_163__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_163__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_163__ap_start = (C_drain_IO_L1_out_wrapper_163__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_164__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_164__is_done__q0 = (C_drain_IO_L1_out_wrapper_164__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_164__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_164__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_164__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_164__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_164__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_164__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_164__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_164__ap_done) begin
            C_drain_IO_L1_out_wrapper_164__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_164__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_164__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_164__ap_done) begin
          C_drain_IO_L1_out_wrapper_164__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_164__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_164__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_164__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_164__ap_start = (C_drain_IO_L1_out_wrapper_164__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_165__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_165__is_done__q0 = (C_drain_IO_L1_out_wrapper_165__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_165__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_165__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_165__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_165__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_165__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_165__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_165__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_165__ap_done) begin
            C_drain_IO_L1_out_wrapper_165__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_165__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_165__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_165__ap_done) begin
          C_drain_IO_L1_out_wrapper_165__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_165__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_165__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_165__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_165__ap_start = (C_drain_IO_L1_out_wrapper_165__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_166__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_166__is_done__q0 = (C_drain_IO_L1_out_wrapper_166__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_166__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_166__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_166__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_166__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_166__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_166__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_166__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_166__ap_done) begin
            C_drain_IO_L1_out_wrapper_166__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_166__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_166__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_166__ap_done) begin
          C_drain_IO_L1_out_wrapper_166__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_166__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_166__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_166__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_166__ap_start = (C_drain_IO_L1_out_wrapper_166__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_167__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_167__is_done__q0 = (C_drain_IO_L1_out_wrapper_167__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_167__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_167__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_167__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_167__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_167__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_167__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_167__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_167__ap_done) begin
            C_drain_IO_L1_out_wrapper_167__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_167__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_167__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_167__ap_done) begin
          C_drain_IO_L1_out_wrapper_167__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_167__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_167__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_167__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_167__ap_start = (C_drain_IO_L1_out_wrapper_167__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_168__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_168__is_done__q0 = (C_drain_IO_L1_out_wrapper_168__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_168__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_168__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_168__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_168__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_168__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_168__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_168__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_168__ap_done) begin
            C_drain_IO_L1_out_wrapper_168__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_168__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_168__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_168__ap_done) begin
          C_drain_IO_L1_out_wrapper_168__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_168__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_168__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_168__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_168__ap_start = (C_drain_IO_L1_out_wrapper_168__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_169__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_169__is_done__q0 = (C_drain_IO_L1_out_wrapper_169__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_169__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_169__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_169__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_169__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_169__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_169__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_169__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_169__ap_done) begin
            C_drain_IO_L1_out_wrapper_169__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_169__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_169__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_169__ap_done) begin
          C_drain_IO_L1_out_wrapper_169__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_169__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_169__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_169__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_169__ap_start = (C_drain_IO_L1_out_wrapper_169__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_170__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_170__is_done__q0 = (C_drain_IO_L1_out_wrapper_170__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_170__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_170__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_170__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_170__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_170__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_170__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_170__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_170__ap_done) begin
            C_drain_IO_L1_out_wrapper_170__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_170__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_170__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_170__ap_done) begin
          C_drain_IO_L1_out_wrapper_170__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_170__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_170__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_170__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_170__ap_start = (C_drain_IO_L1_out_wrapper_170__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_171__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_171__is_done__q0 = (C_drain_IO_L1_out_wrapper_171__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_171__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_171__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_171__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_171__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_171__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_171__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_171__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_171__ap_done) begin
            C_drain_IO_L1_out_wrapper_171__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_171__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_171__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_171__ap_done) begin
          C_drain_IO_L1_out_wrapper_171__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_171__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_171__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_171__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_171__ap_start = (C_drain_IO_L1_out_wrapper_171__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_172__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_172__is_done__q0 = (C_drain_IO_L1_out_wrapper_172__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_172__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_172__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_172__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_172__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_172__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_172__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_172__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_172__ap_done) begin
            C_drain_IO_L1_out_wrapper_172__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_172__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_172__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_172__ap_done) begin
          C_drain_IO_L1_out_wrapper_172__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_172__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_172__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_172__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_172__ap_start = (C_drain_IO_L1_out_wrapper_172__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_173__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_173__is_done__q0 = (C_drain_IO_L1_out_wrapper_173__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_173__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_173__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_173__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_173__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_173__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_173__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_173__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_173__ap_done) begin
            C_drain_IO_L1_out_wrapper_173__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_173__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_173__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_173__ap_done) begin
          C_drain_IO_L1_out_wrapper_173__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_173__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_173__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_173__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_173__ap_start = (C_drain_IO_L1_out_wrapper_173__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_174__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_174__is_done__q0 = (C_drain_IO_L1_out_wrapper_174__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_174__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_174__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_174__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_174__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_174__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_174__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_174__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_174__ap_done) begin
            C_drain_IO_L1_out_wrapper_174__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_174__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_174__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_174__ap_done) begin
          C_drain_IO_L1_out_wrapper_174__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_174__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_174__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_174__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_174__ap_start = (C_drain_IO_L1_out_wrapper_174__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_175__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_175__is_done__q0 = (C_drain_IO_L1_out_wrapper_175__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_175__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_175__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_175__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_175__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_175__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_175__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_175__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_175__ap_done) begin
            C_drain_IO_L1_out_wrapper_175__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_175__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_175__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_175__ap_done) begin
          C_drain_IO_L1_out_wrapper_175__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_175__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_175__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_175__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_175__ap_start = (C_drain_IO_L1_out_wrapper_175__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_176__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_176__is_done__q0 = (C_drain_IO_L1_out_wrapper_176__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_176__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_176__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_176__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_176__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_176__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_176__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_176__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_176__ap_done) begin
            C_drain_IO_L1_out_wrapper_176__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_176__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_176__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_176__ap_done) begin
          C_drain_IO_L1_out_wrapper_176__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_176__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_176__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_176__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_176__ap_start = (C_drain_IO_L1_out_wrapper_176__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_177__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_177__is_done__q0 = (C_drain_IO_L1_out_wrapper_177__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_177__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_177__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_177__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_177__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_177__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_177__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_177__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_177__ap_done) begin
            C_drain_IO_L1_out_wrapper_177__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_177__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_177__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_177__ap_done) begin
          C_drain_IO_L1_out_wrapper_177__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_177__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_177__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_177__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_177__ap_start = (C_drain_IO_L1_out_wrapper_177__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_178__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_178__is_done__q0 = (C_drain_IO_L1_out_wrapper_178__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_178__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_178__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_178__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_178__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_178__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_178__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_178__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_178__ap_done) begin
            C_drain_IO_L1_out_wrapper_178__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_178__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_178__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_178__ap_done) begin
          C_drain_IO_L1_out_wrapper_178__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_178__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_178__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_178__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_178__ap_start = (C_drain_IO_L1_out_wrapper_178__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_179__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_179__is_done__q0 = (C_drain_IO_L1_out_wrapper_179__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_179__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_179__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_179__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_179__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_179__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_179__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_179__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_179__ap_done) begin
            C_drain_IO_L1_out_wrapper_179__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_179__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_179__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_179__ap_done) begin
          C_drain_IO_L1_out_wrapper_179__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_179__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_179__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_179__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_179__ap_start = (C_drain_IO_L1_out_wrapper_179__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_180__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_180__is_done__q0 = (C_drain_IO_L1_out_wrapper_180__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_180__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_180__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_180__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_180__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_180__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_180__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_180__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_180__ap_done) begin
            C_drain_IO_L1_out_wrapper_180__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_180__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_180__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_180__ap_done) begin
          C_drain_IO_L1_out_wrapper_180__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_180__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_180__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_180__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_180__ap_start = (C_drain_IO_L1_out_wrapper_180__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_181__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_181__is_done__q0 = (C_drain_IO_L1_out_wrapper_181__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_181__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_181__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_181__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_181__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_181__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_181__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_181__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_181__ap_done) begin
            C_drain_IO_L1_out_wrapper_181__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_181__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_181__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_181__ap_done) begin
          C_drain_IO_L1_out_wrapper_181__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_181__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_181__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_181__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_181__ap_start = (C_drain_IO_L1_out_wrapper_181__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_182__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_182__is_done__q0 = (C_drain_IO_L1_out_wrapper_182__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_182__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_182__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_182__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_182__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_182__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_182__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_182__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_182__ap_done) begin
            C_drain_IO_L1_out_wrapper_182__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_182__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_182__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_182__ap_done) begin
          C_drain_IO_L1_out_wrapper_182__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_182__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_182__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_182__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_182__ap_start = (C_drain_IO_L1_out_wrapper_182__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_183__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_183__is_done__q0 = (C_drain_IO_L1_out_wrapper_183__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_183__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_183__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_183__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_183__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_183__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_183__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_183__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_183__ap_done) begin
            C_drain_IO_L1_out_wrapper_183__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_183__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_183__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_183__ap_done) begin
          C_drain_IO_L1_out_wrapper_183__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_183__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_183__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_183__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_183__ap_start = (C_drain_IO_L1_out_wrapper_183__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_184__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_184__is_done__q0 = (C_drain_IO_L1_out_wrapper_184__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_184__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_184__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_184__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_184__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_184__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_184__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_184__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_184__ap_done) begin
            C_drain_IO_L1_out_wrapper_184__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_184__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_184__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_184__ap_done) begin
          C_drain_IO_L1_out_wrapper_184__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_184__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_184__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_184__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_184__ap_start = (C_drain_IO_L1_out_wrapper_184__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_185__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_185__is_done__q0 = (C_drain_IO_L1_out_wrapper_185__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_185__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_185__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_185__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_185__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_185__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_185__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_185__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_185__ap_done) begin
            C_drain_IO_L1_out_wrapper_185__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_185__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_185__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_185__ap_done) begin
          C_drain_IO_L1_out_wrapper_185__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_185__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_185__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_185__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_185__ap_start = (C_drain_IO_L1_out_wrapper_185__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_186__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_186__is_done__q0 = (C_drain_IO_L1_out_wrapper_186__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_186__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_186__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_186__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_186__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_186__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_186__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_186__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_186__ap_done) begin
            C_drain_IO_L1_out_wrapper_186__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_186__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_186__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_186__ap_done) begin
          C_drain_IO_L1_out_wrapper_186__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_186__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_186__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_186__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_186__ap_start = (C_drain_IO_L1_out_wrapper_186__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_187__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_187__is_done__q0 = (C_drain_IO_L1_out_wrapper_187__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_187__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_187__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_187__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_187__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_187__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_187__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_187__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_187__ap_done) begin
            C_drain_IO_L1_out_wrapper_187__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_187__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_187__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_187__ap_done) begin
          C_drain_IO_L1_out_wrapper_187__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_187__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_187__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_187__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_187__ap_start = (C_drain_IO_L1_out_wrapper_187__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_188__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_188__is_done__q0 = (C_drain_IO_L1_out_wrapper_188__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_188__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_188__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_188__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_188__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_188__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_188__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_188__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_188__ap_done) begin
            C_drain_IO_L1_out_wrapper_188__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_188__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_188__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_188__ap_done) begin
          C_drain_IO_L1_out_wrapper_188__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_188__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_188__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_188__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_188__ap_start = (C_drain_IO_L1_out_wrapper_188__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_189__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_189__is_done__q0 = (C_drain_IO_L1_out_wrapper_189__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_189__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_189__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_189__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_189__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_189__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_189__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_189__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_189__ap_done) begin
            C_drain_IO_L1_out_wrapper_189__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_189__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_189__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_189__ap_done) begin
          C_drain_IO_L1_out_wrapper_189__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_189__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_189__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_189__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_189__ap_start = (C_drain_IO_L1_out_wrapper_189__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_190__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_190__is_done__q0 = (C_drain_IO_L1_out_wrapper_190__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_190__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_190__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_190__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_190__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_190__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_190__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_190__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_190__ap_done) begin
            C_drain_IO_L1_out_wrapper_190__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_190__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_190__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_190__ap_done) begin
          C_drain_IO_L1_out_wrapper_190__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_190__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_190__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_190__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_190__ap_start = (C_drain_IO_L1_out_wrapper_190__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_191__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_191__is_done__q0 = (C_drain_IO_L1_out_wrapper_191__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_191__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_191__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_191__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_191__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_191__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_191__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_191__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_191__ap_done) begin
            C_drain_IO_L1_out_wrapper_191__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_191__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_191__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_191__ap_done) begin
          C_drain_IO_L1_out_wrapper_191__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_191__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_191__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_191__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_191__ap_start = (C_drain_IO_L1_out_wrapper_191__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_192__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_192__is_done__q0 = (C_drain_IO_L1_out_wrapper_192__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_192__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_192__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_192__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_192__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_192__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_192__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_192__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_192__ap_done) begin
            C_drain_IO_L1_out_wrapper_192__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_192__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_192__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_192__ap_done) begin
          C_drain_IO_L1_out_wrapper_192__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_192__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_192__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_192__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_192__ap_start = (C_drain_IO_L1_out_wrapper_192__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_193__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_193__is_done__q0 = (C_drain_IO_L1_out_wrapper_193__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_193__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_193__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_193__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_193__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_193__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_193__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_193__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_193__ap_done) begin
            C_drain_IO_L1_out_wrapper_193__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_193__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_193__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_193__ap_done) begin
          C_drain_IO_L1_out_wrapper_193__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_193__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_193__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_193__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_193__ap_start = (C_drain_IO_L1_out_wrapper_193__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_194__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_194__is_done__q0 = (C_drain_IO_L1_out_wrapper_194__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_194__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_194__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_194__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_194__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_194__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_194__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_194__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_194__ap_done) begin
            C_drain_IO_L1_out_wrapper_194__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_194__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_194__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_194__ap_done) begin
          C_drain_IO_L1_out_wrapper_194__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_194__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_194__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_194__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_194__ap_start = (C_drain_IO_L1_out_wrapper_194__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_195__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_195__is_done__q0 = (C_drain_IO_L1_out_wrapper_195__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_195__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_195__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_195__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_195__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_195__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_195__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_195__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_195__ap_done) begin
            C_drain_IO_L1_out_wrapper_195__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_195__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_195__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_195__ap_done) begin
          C_drain_IO_L1_out_wrapper_195__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_195__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_195__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_195__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_195__ap_start = (C_drain_IO_L1_out_wrapper_195__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_196__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_196__is_done__q0 = (C_drain_IO_L1_out_wrapper_196__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_196__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_196__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_196__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_196__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_196__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_196__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_196__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_196__ap_done) begin
            C_drain_IO_L1_out_wrapper_196__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_196__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_196__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_196__ap_done) begin
          C_drain_IO_L1_out_wrapper_196__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_196__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_196__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_196__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_196__ap_start = (C_drain_IO_L1_out_wrapper_196__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_197__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_197__is_done__q0 = (C_drain_IO_L1_out_wrapper_197__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_197__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_197__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_197__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_197__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_197__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_197__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_197__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_197__ap_done) begin
            C_drain_IO_L1_out_wrapper_197__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_197__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_197__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_197__ap_done) begin
          C_drain_IO_L1_out_wrapper_197__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_197__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_197__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_197__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_197__ap_start = (C_drain_IO_L1_out_wrapper_197__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_198__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_198__is_done__q0 = (C_drain_IO_L1_out_wrapper_198__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_198__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_198__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_198__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_198__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_198__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_198__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_198__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_198__ap_done) begin
            C_drain_IO_L1_out_wrapper_198__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_198__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_198__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_198__ap_done) begin
          C_drain_IO_L1_out_wrapper_198__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_198__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_198__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_198__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_198__ap_start = (C_drain_IO_L1_out_wrapper_198__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_199__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_199__is_done__q0 = (C_drain_IO_L1_out_wrapper_199__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_199__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_199__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_199__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_199__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_199__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_199__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_199__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_199__ap_done) begin
            C_drain_IO_L1_out_wrapper_199__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_199__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_199__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_199__ap_done) begin
          C_drain_IO_L1_out_wrapper_199__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_199__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_199__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_199__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_199__ap_start = (C_drain_IO_L1_out_wrapper_199__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_200__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_200__is_done__q0 = (C_drain_IO_L1_out_wrapper_200__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_200__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_200__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_200__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_200__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_200__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_200__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_200__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_200__ap_done) begin
            C_drain_IO_L1_out_wrapper_200__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_200__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_200__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_200__ap_done) begin
          C_drain_IO_L1_out_wrapper_200__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_200__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_200__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_200__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_200__ap_start = (C_drain_IO_L1_out_wrapper_200__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_201__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_201__is_done__q0 = (C_drain_IO_L1_out_wrapper_201__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_201__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_201__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_201__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_201__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_201__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_201__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_201__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_201__ap_done) begin
            C_drain_IO_L1_out_wrapper_201__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_201__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_201__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_201__ap_done) begin
          C_drain_IO_L1_out_wrapper_201__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_201__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_201__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_201__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_201__ap_start = (C_drain_IO_L1_out_wrapper_201__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_202__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_202__is_done__q0 = (C_drain_IO_L1_out_wrapper_202__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_202__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_202__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_202__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_202__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_202__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_202__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_202__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_202__ap_done) begin
            C_drain_IO_L1_out_wrapper_202__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_202__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_202__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_202__ap_done) begin
          C_drain_IO_L1_out_wrapper_202__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_202__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_202__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_202__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_202__ap_start = (C_drain_IO_L1_out_wrapper_202__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_203__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_203__is_done__q0 = (C_drain_IO_L1_out_wrapper_203__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_203__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_203__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_203__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_203__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_203__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_203__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_203__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_203__ap_done) begin
            C_drain_IO_L1_out_wrapper_203__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_203__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_203__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_203__ap_done) begin
          C_drain_IO_L1_out_wrapper_203__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_203__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_203__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_203__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_203__ap_start = (C_drain_IO_L1_out_wrapper_203__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_204__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_204__is_done__q0 = (C_drain_IO_L1_out_wrapper_204__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_204__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_204__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_204__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_204__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_204__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_204__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_204__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_204__ap_done) begin
            C_drain_IO_L1_out_wrapper_204__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_204__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_204__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_204__ap_done) begin
          C_drain_IO_L1_out_wrapper_204__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_204__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_204__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_204__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_204__ap_start = (C_drain_IO_L1_out_wrapper_204__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_205__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_205__is_done__q0 = (C_drain_IO_L1_out_wrapper_205__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_205__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_205__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_205__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_205__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_205__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_205__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_205__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_205__ap_done) begin
            C_drain_IO_L1_out_wrapper_205__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_205__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_205__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_205__ap_done) begin
          C_drain_IO_L1_out_wrapper_205__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_205__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_205__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_205__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_205__ap_start = (C_drain_IO_L1_out_wrapper_205__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_206__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_206__is_done__q0 = (C_drain_IO_L1_out_wrapper_206__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_206__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_206__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_206__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_206__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_206__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_206__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_206__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_206__ap_done) begin
            C_drain_IO_L1_out_wrapper_206__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_206__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_206__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_206__ap_done) begin
          C_drain_IO_L1_out_wrapper_206__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_206__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_206__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_206__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_206__ap_start = (C_drain_IO_L1_out_wrapper_206__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_207__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_207__is_done__q0 = (C_drain_IO_L1_out_wrapper_207__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_207__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_207__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_207__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_207__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_207__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_207__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_207__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_207__ap_done) begin
            C_drain_IO_L1_out_wrapper_207__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_207__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_207__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_207__ap_done) begin
          C_drain_IO_L1_out_wrapper_207__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_207__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_207__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_207__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_207__ap_start = (C_drain_IO_L1_out_wrapper_207__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_208__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_208__is_done__q0 = (C_drain_IO_L1_out_wrapper_208__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_208__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_208__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_208__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_208__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_208__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_208__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_208__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_208__ap_done) begin
            C_drain_IO_L1_out_wrapper_208__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_208__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_208__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_208__ap_done) begin
          C_drain_IO_L1_out_wrapper_208__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_208__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_208__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_208__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_208__ap_start = (C_drain_IO_L1_out_wrapper_208__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_209__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_209__is_done__q0 = (C_drain_IO_L1_out_wrapper_209__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_209__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_209__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_209__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_209__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_209__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_209__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_209__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_209__ap_done) begin
            C_drain_IO_L1_out_wrapper_209__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_209__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_209__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_209__ap_done) begin
          C_drain_IO_L1_out_wrapper_209__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_209__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_209__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_209__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_209__ap_start = (C_drain_IO_L1_out_wrapper_209__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_210__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_210__is_done__q0 = (C_drain_IO_L1_out_wrapper_210__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_210__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_210__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_210__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_210__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_210__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_210__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_210__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_210__ap_done) begin
            C_drain_IO_L1_out_wrapper_210__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_210__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_210__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_210__ap_done) begin
          C_drain_IO_L1_out_wrapper_210__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_210__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_210__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_210__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_210__ap_start = (C_drain_IO_L1_out_wrapper_210__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_211__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_211__is_done__q0 = (C_drain_IO_L1_out_wrapper_211__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_211__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_211__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_211__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_211__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_211__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_211__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_211__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_211__ap_done) begin
            C_drain_IO_L1_out_wrapper_211__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_211__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_211__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_211__ap_done) begin
          C_drain_IO_L1_out_wrapper_211__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_211__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_211__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_211__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_211__ap_start = (C_drain_IO_L1_out_wrapper_211__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_212__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_212__is_done__q0 = (C_drain_IO_L1_out_wrapper_212__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_212__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_212__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_212__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_212__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_212__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_212__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_212__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_212__ap_done) begin
            C_drain_IO_L1_out_wrapper_212__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_212__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_212__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_212__ap_done) begin
          C_drain_IO_L1_out_wrapper_212__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_212__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_212__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_212__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_212__ap_start = (C_drain_IO_L1_out_wrapper_212__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_213__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_213__is_done__q0 = (C_drain_IO_L1_out_wrapper_213__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_213__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_213__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_213__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_213__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_213__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_213__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_213__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_213__ap_done) begin
            C_drain_IO_L1_out_wrapper_213__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_213__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_213__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_213__ap_done) begin
          C_drain_IO_L1_out_wrapper_213__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_213__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_213__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_213__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_213__ap_start = (C_drain_IO_L1_out_wrapper_213__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_214__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_214__is_done__q0 = (C_drain_IO_L1_out_wrapper_214__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_214__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_214__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_214__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_214__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_214__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_214__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_214__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_214__ap_done) begin
            C_drain_IO_L1_out_wrapper_214__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_214__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_214__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_214__ap_done) begin
          C_drain_IO_L1_out_wrapper_214__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_214__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_214__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_214__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_214__ap_start = (C_drain_IO_L1_out_wrapper_214__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_215__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_215__is_done__q0 = (C_drain_IO_L1_out_wrapper_215__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_215__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_215__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_215__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_215__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_215__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_215__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_215__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_215__ap_done) begin
            C_drain_IO_L1_out_wrapper_215__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_215__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_215__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_215__ap_done) begin
          C_drain_IO_L1_out_wrapper_215__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_215__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_215__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_215__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_215__ap_start = (C_drain_IO_L1_out_wrapper_215__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_216__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_216__is_done__q0 = (C_drain_IO_L1_out_wrapper_216__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_216__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_216__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_216__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_216__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_216__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_216__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_216__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_216__ap_done) begin
            C_drain_IO_L1_out_wrapper_216__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_216__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_216__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_216__ap_done) begin
          C_drain_IO_L1_out_wrapper_216__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_216__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_216__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_216__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_216__ap_start = (C_drain_IO_L1_out_wrapper_216__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_217__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_217__is_done__q0 = (C_drain_IO_L1_out_wrapper_217__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_217__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_217__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_217__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_217__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_217__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_217__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_217__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_217__ap_done) begin
            C_drain_IO_L1_out_wrapper_217__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_217__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_217__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_217__ap_done) begin
          C_drain_IO_L1_out_wrapper_217__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_217__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_217__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_217__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_217__ap_start = (C_drain_IO_L1_out_wrapper_217__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_218__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_218__is_done__q0 = (C_drain_IO_L1_out_wrapper_218__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_218__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_218__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_218__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_218__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_218__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_218__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_218__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_218__ap_done) begin
            C_drain_IO_L1_out_wrapper_218__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_218__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_218__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_218__ap_done) begin
          C_drain_IO_L1_out_wrapper_218__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_218__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_218__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_218__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_218__ap_start = (C_drain_IO_L1_out_wrapper_218__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_219__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_219__is_done__q0 = (C_drain_IO_L1_out_wrapper_219__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_219__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_219__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_219__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_219__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_219__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_219__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_219__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_219__ap_done) begin
            C_drain_IO_L1_out_wrapper_219__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_219__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_219__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_219__ap_done) begin
          C_drain_IO_L1_out_wrapper_219__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_219__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_219__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_219__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_219__ap_start = (C_drain_IO_L1_out_wrapper_219__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_220__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_220__is_done__q0 = (C_drain_IO_L1_out_wrapper_220__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_220__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_220__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_220__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_220__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_220__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_220__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_220__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_220__ap_done) begin
            C_drain_IO_L1_out_wrapper_220__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_220__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_220__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_220__ap_done) begin
          C_drain_IO_L1_out_wrapper_220__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_220__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_220__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_220__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_220__ap_start = (C_drain_IO_L1_out_wrapper_220__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_221__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_221__is_done__q0 = (C_drain_IO_L1_out_wrapper_221__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_221__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_221__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_221__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_221__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_221__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_221__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_221__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_221__ap_done) begin
            C_drain_IO_L1_out_wrapper_221__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_221__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_221__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_221__ap_done) begin
          C_drain_IO_L1_out_wrapper_221__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_221__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_221__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_221__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_221__ap_start = (C_drain_IO_L1_out_wrapper_221__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_222__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_222__is_done__q0 = (C_drain_IO_L1_out_wrapper_222__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_222__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_222__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_222__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_222__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_222__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_222__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_222__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_222__ap_done) begin
            C_drain_IO_L1_out_wrapper_222__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_222__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_222__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_222__ap_done) begin
          C_drain_IO_L1_out_wrapper_222__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_222__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_222__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_222__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_222__ap_start = (C_drain_IO_L1_out_wrapper_222__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_223__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_223__is_done__q0 = (C_drain_IO_L1_out_wrapper_223__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_223__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_223__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_223__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_223__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_223__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_223__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_223__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_223__ap_done) begin
            C_drain_IO_L1_out_wrapper_223__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_223__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_223__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_223__ap_done) begin
          C_drain_IO_L1_out_wrapper_223__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_223__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_223__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_223__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_223__ap_start = (C_drain_IO_L1_out_wrapper_223__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_224__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_224__is_done__q0 = (C_drain_IO_L1_out_wrapper_224__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_224__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_224__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_224__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_224__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_224__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_224__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_224__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_224__ap_done) begin
            C_drain_IO_L1_out_wrapper_224__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_224__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_224__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_224__ap_done) begin
          C_drain_IO_L1_out_wrapper_224__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_224__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_224__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_224__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_224__ap_start = (C_drain_IO_L1_out_wrapper_224__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_225__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_225__is_done__q0 = (C_drain_IO_L1_out_wrapper_225__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_225__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_225__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_225__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_225__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_225__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_225__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_225__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_225__ap_done) begin
            C_drain_IO_L1_out_wrapper_225__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_225__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_225__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_225__ap_done) begin
          C_drain_IO_L1_out_wrapper_225__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_225__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_225__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_225__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_225__ap_start = (C_drain_IO_L1_out_wrapper_225__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_226__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_226__is_done__q0 = (C_drain_IO_L1_out_wrapper_226__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_226__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_226__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_226__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_226__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_226__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_226__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_226__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_226__ap_done) begin
            C_drain_IO_L1_out_wrapper_226__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_226__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_226__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_226__ap_done) begin
          C_drain_IO_L1_out_wrapper_226__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_226__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_226__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_226__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_226__ap_start = (C_drain_IO_L1_out_wrapper_226__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_227__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_227__is_done__q0 = (C_drain_IO_L1_out_wrapper_227__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_227__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_227__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_227__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_227__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_227__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_227__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_227__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_227__ap_done) begin
            C_drain_IO_L1_out_wrapper_227__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_227__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_227__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_227__ap_done) begin
          C_drain_IO_L1_out_wrapper_227__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_227__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_227__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_227__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_227__ap_start = (C_drain_IO_L1_out_wrapper_227__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_228__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_228__is_done__q0 = (C_drain_IO_L1_out_wrapper_228__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_228__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_228__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_228__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_228__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_228__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_228__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_228__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_228__ap_done) begin
            C_drain_IO_L1_out_wrapper_228__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_228__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_228__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_228__ap_done) begin
          C_drain_IO_L1_out_wrapper_228__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_228__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_228__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_228__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_228__ap_start = (C_drain_IO_L1_out_wrapper_228__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_229__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_229__is_done__q0 = (C_drain_IO_L1_out_wrapper_229__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_229__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_229__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_229__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_229__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_229__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_229__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_229__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_229__ap_done) begin
            C_drain_IO_L1_out_wrapper_229__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_229__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_229__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_229__ap_done) begin
          C_drain_IO_L1_out_wrapper_229__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_229__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_229__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_229__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_229__ap_start = (C_drain_IO_L1_out_wrapper_229__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_230__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_230__is_done__q0 = (C_drain_IO_L1_out_wrapper_230__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_230__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_230__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_230__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_230__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_230__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_230__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_230__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_230__ap_done) begin
            C_drain_IO_L1_out_wrapper_230__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_230__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_230__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_230__ap_done) begin
          C_drain_IO_L1_out_wrapper_230__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_230__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_230__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_230__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_230__ap_start = (C_drain_IO_L1_out_wrapper_230__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_231__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_231__is_done__q0 = (C_drain_IO_L1_out_wrapper_231__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_231__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_231__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_231__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_231__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_231__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_231__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_231__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_231__ap_done) begin
            C_drain_IO_L1_out_wrapper_231__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_231__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_231__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_231__ap_done) begin
          C_drain_IO_L1_out_wrapper_231__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_231__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_231__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_231__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_231__ap_start = (C_drain_IO_L1_out_wrapper_231__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_232__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_232__is_done__q0 = (C_drain_IO_L1_out_wrapper_232__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_232__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_232__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_232__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_232__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_232__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_232__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_232__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_232__ap_done) begin
            C_drain_IO_L1_out_wrapper_232__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_232__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_232__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_232__ap_done) begin
          C_drain_IO_L1_out_wrapper_232__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_232__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_232__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_232__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_232__ap_start = (C_drain_IO_L1_out_wrapper_232__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_233__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_233__is_done__q0 = (C_drain_IO_L1_out_wrapper_233__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_233__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_233__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_233__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_233__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_233__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_233__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_233__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_233__ap_done) begin
            C_drain_IO_L1_out_wrapper_233__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_233__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_233__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_233__ap_done) begin
          C_drain_IO_L1_out_wrapper_233__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_233__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_233__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_233__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_233__ap_start = (C_drain_IO_L1_out_wrapper_233__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_234__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_234__is_done__q0 = (C_drain_IO_L1_out_wrapper_234__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_234__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_234__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_234__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_234__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_234__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_234__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_234__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_234__ap_done) begin
            C_drain_IO_L1_out_wrapper_234__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_234__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_234__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_234__ap_done) begin
          C_drain_IO_L1_out_wrapper_234__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_234__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_234__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_234__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_234__ap_start = (C_drain_IO_L1_out_wrapper_234__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_235__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_235__is_done__q0 = (C_drain_IO_L1_out_wrapper_235__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_235__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_235__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_235__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_235__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_235__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_235__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_235__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_235__ap_done) begin
            C_drain_IO_L1_out_wrapper_235__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_235__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_235__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_235__ap_done) begin
          C_drain_IO_L1_out_wrapper_235__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_235__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_235__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_235__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_235__ap_start = (C_drain_IO_L1_out_wrapper_235__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_236__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_236__is_done__q0 = (C_drain_IO_L1_out_wrapper_236__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_236__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_236__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_236__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_236__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_236__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_236__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_236__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_236__ap_done) begin
            C_drain_IO_L1_out_wrapper_236__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_236__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_236__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_236__ap_done) begin
          C_drain_IO_L1_out_wrapper_236__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_236__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_236__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_236__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_236__ap_start = (C_drain_IO_L1_out_wrapper_236__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_237__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_237__is_done__q0 = (C_drain_IO_L1_out_wrapper_237__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_237__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_237__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_237__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_237__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_237__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_237__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_237__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_237__ap_done) begin
            C_drain_IO_L1_out_wrapper_237__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_237__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_237__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_237__ap_done) begin
          C_drain_IO_L1_out_wrapper_237__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_237__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_237__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_237__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_237__ap_start = (C_drain_IO_L1_out_wrapper_237__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_238__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_238__is_done__q0 = (C_drain_IO_L1_out_wrapper_238__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_238__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_238__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_238__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_238__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_238__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_238__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_238__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_238__ap_done) begin
            C_drain_IO_L1_out_wrapper_238__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_238__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_238__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_238__ap_done) begin
          C_drain_IO_L1_out_wrapper_238__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_238__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_238__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_238__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_238__ap_start = (C_drain_IO_L1_out_wrapper_238__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_239__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_239__is_done__q0 = (C_drain_IO_L1_out_wrapper_239__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_239__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_239__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_239__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_239__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_239__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_239__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_239__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_239__ap_done) begin
            C_drain_IO_L1_out_wrapper_239__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_239__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_239__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_239__ap_done) begin
          C_drain_IO_L1_out_wrapper_239__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_239__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_239__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_239__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_239__ap_start = (C_drain_IO_L1_out_wrapper_239__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_240__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_240__is_done__q0 = (C_drain_IO_L1_out_wrapper_240__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_240__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_240__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_240__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_240__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_240__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_240__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_240__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_240__ap_done) begin
            C_drain_IO_L1_out_wrapper_240__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_240__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_240__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_240__ap_done) begin
          C_drain_IO_L1_out_wrapper_240__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_240__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_240__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_240__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_240__ap_start = (C_drain_IO_L1_out_wrapper_240__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_241__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_241__is_done__q0 = (C_drain_IO_L1_out_wrapper_241__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_241__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_241__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_241__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_241__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_241__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_241__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_241__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_241__ap_done) begin
            C_drain_IO_L1_out_wrapper_241__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_241__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_241__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_241__ap_done) begin
          C_drain_IO_L1_out_wrapper_241__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_241__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_241__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_241__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_241__ap_start = (C_drain_IO_L1_out_wrapper_241__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_242__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_242__is_done__q0 = (C_drain_IO_L1_out_wrapper_242__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_242__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_242__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_242__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_242__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_242__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_242__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_242__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_242__ap_done) begin
            C_drain_IO_L1_out_wrapper_242__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_242__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_242__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_242__ap_done) begin
          C_drain_IO_L1_out_wrapper_242__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_242__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_242__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_242__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_242__ap_start = (C_drain_IO_L1_out_wrapper_242__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_243__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_243__is_done__q0 = (C_drain_IO_L1_out_wrapper_243__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_243__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_243__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_243__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_243__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_243__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_243__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_243__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_243__ap_done) begin
            C_drain_IO_L1_out_wrapper_243__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_243__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_243__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_243__ap_done) begin
          C_drain_IO_L1_out_wrapper_243__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_243__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_243__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_243__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_243__ap_start = (C_drain_IO_L1_out_wrapper_243__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_244__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_244__is_done__q0 = (C_drain_IO_L1_out_wrapper_244__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_244__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_244__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_244__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_244__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_244__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_244__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_244__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_244__ap_done) begin
            C_drain_IO_L1_out_wrapper_244__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_244__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_244__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_244__ap_done) begin
          C_drain_IO_L1_out_wrapper_244__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_244__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_244__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_244__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_244__ap_start = (C_drain_IO_L1_out_wrapper_244__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_245__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_245__is_done__q0 = (C_drain_IO_L1_out_wrapper_245__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_245__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_245__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_245__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_245__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_245__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_245__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_245__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_245__ap_done) begin
            C_drain_IO_L1_out_wrapper_245__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_245__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_245__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_245__ap_done) begin
          C_drain_IO_L1_out_wrapper_245__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_245__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_245__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_245__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_245__ap_start = (C_drain_IO_L1_out_wrapper_245__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_246__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_246__is_done__q0 = (C_drain_IO_L1_out_wrapper_246__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_246__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_246__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_246__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_246__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_246__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_246__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_246__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_246__ap_done) begin
            C_drain_IO_L1_out_wrapper_246__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_246__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_246__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_246__ap_done) begin
          C_drain_IO_L1_out_wrapper_246__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_246__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_246__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_246__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_246__ap_start = (C_drain_IO_L1_out_wrapper_246__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_247__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_247__is_done__q0 = (C_drain_IO_L1_out_wrapper_247__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_247__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_247__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_247__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_247__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_247__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_247__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_247__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_247__ap_done) begin
            C_drain_IO_L1_out_wrapper_247__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_247__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_247__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_247__ap_done) begin
          C_drain_IO_L1_out_wrapper_247__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_247__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_247__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_247__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_247__ap_start = (C_drain_IO_L1_out_wrapper_247__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_248__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_248__is_done__q0 = (C_drain_IO_L1_out_wrapper_248__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_248__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_248__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_248__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_248__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_248__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_248__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_248__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_248__ap_done) begin
            C_drain_IO_L1_out_wrapper_248__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_248__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_248__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_248__ap_done) begin
          C_drain_IO_L1_out_wrapper_248__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_248__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_248__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_248__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_248__ap_start = (C_drain_IO_L1_out_wrapper_248__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_249__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_249__is_done__q0 = (C_drain_IO_L1_out_wrapper_249__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_249__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_249__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_249__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_249__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_249__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_249__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_249__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_249__ap_done) begin
            C_drain_IO_L1_out_wrapper_249__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_249__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_249__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_249__ap_done) begin
          C_drain_IO_L1_out_wrapper_249__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_249__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_249__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_249__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_249__ap_start = (C_drain_IO_L1_out_wrapper_249__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_250__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_250__is_done__q0 = (C_drain_IO_L1_out_wrapper_250__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_250__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_250__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_250__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_250__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_250__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_250__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_250__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_250__ap_done) begin
            C_drain_IO_L1_out_wrapper_250__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_250__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_250__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_250__ap_done) begin
          C_drain_IO_L1_out_wrapper_250__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_250__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_250__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_250__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_250__ap_start = (C_drain_IO_L1_out_wrapper_250__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_251__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_251__is_done__q0 = (C_drain_IO_L1_out_wrapper_251__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_251__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_251__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_251__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_251__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_251__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_251__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_251__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_251__ap_done) begin
            C_drain_IO_L1_out_wrapper_251__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_251__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_251__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_251__ap_done) begin
          C_drain_IO_L1_out_wrapper_251__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_251__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_251__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_251__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_251__ap_start = (C_drain_IO_L1_out_wrapper_251__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_252__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_252__is_done__q0 = (C_drain_IO_L1_out_wrapper_252__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_252__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_252__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_252__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_252__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_252__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_252__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_252__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_252__ap_done) begin
            C_drain_IO_L1_out_wrapper_252__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_252__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_252__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_252__ap_done) begin
          C_drain_IO_L1_out_wrapper_252__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_252__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_252__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_252__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_252__ap_start = (C_drain_IO_L1_out_wrapper_252__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_253__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_253__is_done__q0 = (C_drain_IO_L1_out_wrapper_253__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_253__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_253__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_253__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_253__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_253__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_253__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_253__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_253__ap_done) begin
            C_drain_IO_L1_out_wrapper_253__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_253__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_253__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_253__ap_done) begin
          C_drain_IO_L1_out_wrapper_253__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_253__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_253__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_253__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_253__ap_start = (C_drain_IO_L1_out_wrapper_253__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_254__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_254__is_done__q0 = (C_drain_IO_L1_out_wrapper_254__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_254__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_254__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_254__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_254__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_254__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_254__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_254__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_254__ap_done) begin
            C_drain_IO_L1_out_wrapper_254__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_254__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_254__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_254__ap_done) begin
          C_drain_IO_L1_out_wrapper_254__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_254__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_254__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_254__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_254__ap_start = (C_drain_IO_L1_out_wrapper_254__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_255__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_255__is_done__q0 = (C_drain_IO_L1_out_wrapper_255__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_255__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_255__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_255__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_255__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_255__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_255__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_255__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_255__ap_done) begin
            C_drain_IO_L1_out_wrapper_255__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_255__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_255__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_255__ap_done) begin
          C_drain_IO_L1_out_wrapper_255__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_255__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_255__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_255__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_255__ap_start = (C_drain_IO_L1_out_wrapper_255__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_256__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_256__is_done__q0 = (C_drain_IO_L1_out_wrapper_256__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_256__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_256__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_256__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_256__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_256__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_256__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_256__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_256__ap_done) begin
            C_drain_IO_L1_out_wrapper_256__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_256__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_256__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_256__ap_done) begin
          C_drain_IO_L1_out_wrapper_256__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_256__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_256__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_256__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_256__ap_start = (C_drain_IO_L1_out_wrapper_256__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_257__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_257__is_done__q0 = (C_drain_IO_L1_out_wrapper_257__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_257__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_257__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_257__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_257__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_257__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_257__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_257__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_257__ap_done) begin
            C_drain_IO_L1_out_wrapper_257__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_257__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_257__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_257__ap_done) begin
          C_drain_IO_L1_out_wrapper_257__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_257__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_257__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_257__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_257__ap_start = (C_drain_IO_L1_out_wrapper_257__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_258__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_258__is_done__q0 = (C_drain_IO_L1_out_wrapper_258__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_258__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_258__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_258__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_258__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_258__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_258__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_258__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_258__ap_done) begin
            C_drain_IO_L1_out_wrapper_258__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_258__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_258__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_258__ap_done) begin
          C_drain_IO_L1_out_wrapper_258__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_258__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_258__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_258__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_258__ap_start = (C_drain_IO_L1_out_wrapper_258__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_259__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_259__is_done__q0 = (C_drain_IO_L1_out_wrapper_259__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_259__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_259__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_259__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_259__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_259__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_259__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_259__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_259__ap_done) begin
            C_drain_IO_L1_out_wrapper_259__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_259__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_259__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_259__ap_done) begin
          C_drain_IO_L1_out_wrapper_259__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_259__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_259__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_259__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_259__ap_start = (C_drain_IO_L1_out_wrapper_259__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_260__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_260__is_done__q0 = (C_drain_IO_L1_out_wrapper_260__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_260__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_260__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_260__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_260__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_260__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_260__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_260__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_260__ap_done) begin
            C_drain_IO_L1_out_wrapper_260__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_260__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_260__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_260__ap_done) begin
          C_drain_IO_L1_out_wrapper_260__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_260__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_260__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_260__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_260__ap_start = (C_drain_IO_L1_out_wrapper_260__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_261__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_261__is_done__q0 = (C_drain_IO_L1_out_wrapper_261__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_261__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_261__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_261__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_261__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_261__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_261__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_261__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_261__ap_done) begin
            C_drain_IO_L1_out_wrapper_261__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_261__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_261__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_261__ap_done) begin
          C_drain_IO_L1_out_wrapper_261__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_261__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_261__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_261__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_261__ap_start = (C_drain_IO_L1_out_wrapper_261__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_262__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_262__is_done__q0 = (C_drain_IO_L1_out_wrapper_262__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_262__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_262__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_262__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_262__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_262__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_262__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_262__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_262__ap_done) begin
            C_drain_IO_L1_out_wrapper_262__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_262__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_262__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_262__ap_done) begin
          C_drain_IO_L1_out_wrapper_262__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_262__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_262__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_262__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_262__ap_start = (C_drain_IO_L1_out_wrapper_262__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_263__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_263__is_done__q0 = (C_drain_IO_L1_out_wrapper_263__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_263__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_263__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_263__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_263__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_263__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_263__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_263__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_263__ap_done) begin
            C_drain_IO_L1_out_wrapper_263__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_263__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_263__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_263__ap_done) begin
          C_drain_IO_L1_out_wrapper_263__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_263__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_263__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_263__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_263__ap_start = (C_drain_IO_L1_out_wrapper_263__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_264__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_264__is_done__q0 = (C_drain_IO_L1_out_wrapper_264__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_264__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_264__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_264__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_264__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_264__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_264__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_264__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_264__ap_done) begin
            C_drain_IO_L1_out_wrapper_264__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_264__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_264__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_264__ap_done) begin
          C_drain_IO_L1_out_wrapper_264__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_264__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_264__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_264__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_264__ap_start = (C_drain_IO_L1_out_wrapper_264__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_265__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_265__is_done__q0 = (C_drain_IO_L1_out_wrapper_265__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_265__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_265__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_265__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_265__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_265__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_265__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_265__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_265__ap_done) begin
            C_drain_IO_L1_out_wrapper_265__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_265__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_265__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_265__ap_done) begin
          C_drain_IO_L1_out_wrapper_265__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_265__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_265__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_265__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_265__ap_start = (C_drain_IO_L1_out_wrapper_265__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_266__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_266__is_done__q0 = (C_drain_IO_L1_out_wrapper_266__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_266__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_266__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_266__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_266__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_266__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_266__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_266__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_266__ap_done) begin
            C_drain_IO_L1_out_wrapper_266__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_266__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_266__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_266__ap_done) begin
          C_drain_IO_L1_out_wrapper_266__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_266__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_266__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_266__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_266__ap_start = (C_drain_IO_L1_out_wrapper_266__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_267__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_267__is_done__q0 = (C_drain_IO_L1_out_wrapper_267__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_267__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_267__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_267__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_267__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_267__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_267__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_267__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_267__ap_done) begin
            C_drain_IO_L1_out_wrapper_267__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_267__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_267__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_267__ap_done) begin
          C_drain_IO_L1_out_wrapper_267__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_267__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_267__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_267__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_267__ap_start = (C_drain_IO_L1_out_wrapper_267__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_268__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_268__is_done__q0 = (C_drain_IO_L1_out_wrapper_268__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_268__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_268__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_268__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_268__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_268__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_268__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_268__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_268__ap_done) begin
            C_drain_IO_L1_out_wrapper_268__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_268__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_268__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_268__ap_done) begin
          C_drain_IO_L1_out_wrapper_268__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_268__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_268__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_268__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_268__ap_start = (C_drain_IO_L1_out_wrapper_268__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_269__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_269__is_done__q0 = (C_drain_IO_L1_out_wrapper_269__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_269__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_269__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_269__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_269__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_269__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_269__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_269__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_269__ap_done) begin
            C_drain_IO_L1_out_wrapper_269__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_269__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_269__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_269__ap_done) begin
          C_drain_IO_L1_out_wrapper_269__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_269__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_269__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_269__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_269__ap_start = (C_drain_IO_L1_out_wrapper_269__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_270__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_270__is_done__q0 = (C_drain_IO_L1_out_wrapper_270__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_270__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_270__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_270__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_270__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_270__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_270__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_270__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_270__ap_done) begin
            C_drain_IO_L1_out_wrapper_270__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_270__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_270__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_270__ap_done) begin
          C_drain_IO_L1_out_wrapper_270__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_270__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_270__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_270__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_270__ap_start = (C_drain_IO_L1_out_wrapper_270__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_271__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_271__is_done__q0 = (C_drain_IO_L1_out_wrapper_271__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_271__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_271__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_271__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_271__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_271__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_271__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_271__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_271__ap_done) begin
            C_drain_IO_L1_out_wrapper_271__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_271__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_271__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_271__ap_done) begin
          C_drain_IO_L1_out_wrapper_271__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_271__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_271__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_271__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_271__ap_start = (C_drain_IO_L1_out_wrapper_271__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_272__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_272__is_done__q0 = (C_drain_IO_L1_out_wrapper_272__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_272__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_272__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_272__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_272__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_272__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_272__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_272__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_272__ap_done) begin
            C_drain_IO_L1_out_wrapper_272__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_272__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_272__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_272__ap_done) begin
          C_drain_IO_L1_out_wrapper_272__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_272__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_272__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_272__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_272__ap_start = (C_drain_IO_L1_out_wrapper_272__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_273__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_273__is_done__q0 = (C_drain_IO_L1_out_wrapper_273__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_273__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_273__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_273__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_273__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_273__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_273__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_273__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_273__ap_done) begin
            C_drain_IO_L1_out_wrapper_273__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_273__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_273__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_273__ap_done) begin
          C_drain_IO_L1_out_wrapper_273__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_273__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_273__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_273__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_273__ap_start = (C_drain_IO_L1_out_wrapper_273__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_274__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_274__is_done__q0 = (C_drain_IO_L1_out_wrapper_274__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_274__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_274__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_274__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_274__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_274__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_274__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_274__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_274__ap_done) begin
            C_drain_IO_L1_out_wrapper_274__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_274__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_274__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_274__ap_done) begin
          C_drain_IO_L1_out_wrapper_274__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_274__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_274__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_274__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_274__ap_start = (C_drain_IO_L1_out_wrapper_274__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_275__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_275__is_done__q0 = (C_drain_IO_L1_out_wrapper_275__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_275__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_275__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_275__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_275__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_275__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_275__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_275__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_275__ap_done) begin
            C_drain_IO_L1_out_wrapper_275__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_275__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_275__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_275__ap_done) begin
          C_drain_IO_L1_out_wrapper_275__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_275__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_275__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_275__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_275__ap_start = (C_drain_IO_L1_out_wrapper_275__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_276__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_276__is_done__q0 = (C_drain_IO_L1_out_wrapper_276__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_276__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_276__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_276__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_276__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_276__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_276__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_276__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_276__ap_done) begin
            C_drain_IO_L1_out_wrapper_276__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_276__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_276__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_276__ap_done) begin
          C_drain_IO_L1_out_wrapper_276__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_276__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_276__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_276__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_276__ap_start = (C_drain_IO_L1_out_wrapper_276__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_277__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_277__is_done__q0 = (C_drain_IO_L1_out_wrapper_277__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_277__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_277__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_277__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_277__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_277__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_277__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_277__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_277__ap_done) begin
            C_drain_IO_L1_out_wrapper_277__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_277__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_277__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_277__ap_done) begin
          C_drain_IO_L1_out_wrapper_277__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_277__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_277__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_277__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_277__ap_start = (C_drain_IO_L1_out_wrapper_277__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_278__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_278__is_done__q0 = (C_drain_IO_L1_out_wrapper_278__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_278__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_278__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_278__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_278__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_278__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_278__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_278__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_278__ap_done) begin
            C_drain_IO_L1_out_wrapper_278__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_278__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_278__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_278__ap_done) begin
          C_drain_IO_L1_out_wrapper_278__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_278__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_278__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_278__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_278__ap_start = (C_drain_IO_L1_out_wrapper_278__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_279__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_279__is_done__q0 = (C_drain_IO_L1_out_wrapper_279__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_279__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_279__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_279__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_279__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_279__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_279__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_279__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_279__ap_done) begin
            C_drain_IO_L1_out_wrapper_279__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_279__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_279__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_279__ap_done) begin
          C_drain_IO_L1_out_wrapper_279__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_279__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_279__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_279__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_279__ap_start = (C_drain_IO_L1_out_wrapper_279__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_280__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_280__is_done__q0 = (C_drain_IO_L1_out_wrapper_280__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_280__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_280__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_280__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_280__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_280__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_280__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_280__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_280__ap_done) begin
            C_drain_IO_L1_out_wrapper_280__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_280__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_280__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_280__ap_done) begin
          C_drain_IO_L1_out_wrapper_280__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_280__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_280__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_280__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_280__ap_start = (C_drain_IO_L1_out_wrapper_280__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_281__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_281__is_done__q0 = (C_drain_IO_L1_out_wrapper_281__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_281__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_281__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_281__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_281__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_281__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_281__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_281__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_281__ap_done) begin
            C_drain_IO_L1_out_wrapper_281__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_281__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_281__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_281__ap_done) begin
          C_drain_IO_L1_out_wrapper_281__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_281__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_281__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_281__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_281__ap_start = (C_drain_IO_L1_out_wrapper_281__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_282__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_282__is_done__q0 = (C_drain_IO_L1_out_wrapper_282__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_282__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_282__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_282__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_282__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_282__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_282__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_282__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_282__ap_done) begin
            C_drain_IO_L1_out_wrapper_282__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_282__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_282__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_282__ap_done) begin
          C_drain_IO_L1_out_wrapper_282__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_282__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_282__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_282__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_282__ap_start = (C_drain_IO_L1_out_wrapper_282__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_283__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_283__is_done__q0 = (C_drain_IO_L1_out_wrapper_283__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_283__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_283__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_283__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_283__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_283__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_283__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_283__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_283__ap_done) begin
            C_drain_IO_L1_out_wrapper_283__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_283__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_283__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_283__ap_done) begin
          C_drain_IO_L1_out_wrapper_283__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_283__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_283__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_283__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_283__ap_start = (C_drain_IO_L1_out_wrapper_283__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_284__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_284__is_done__q0 = (C_drain_IO_L1_out_wrapper_284__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_284__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_284__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_284__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_284__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_284__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_284__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_284__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_284__ap_done) begin
            C_drain_IO_L1_out_wrapper_284__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_284__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_284__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_284__ap_done) begin
          C_drain_IO_L1_out_wrapper_284__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_284__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_284__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_284__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_284__ap_start = (C_drain_IO_L1_out_wrapper_284__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_285__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_285__is_done__q0 = (C_drain_IO_L1_out_wrapper_285__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_285__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_285__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_285__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_285__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_285__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_285__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_285__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_285__ap_done) begin
            C_drain_IO_L1_out_wrapper_285__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_285__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_285__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_285__ap_done) begin
          C_drain_IO_L1_out_wrapper_285__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_285__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_285__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_285__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_285__ap_start = (C_drain_IO_L1_out_wrapper_285__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_286__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_286__is_done__q0 = (C_drain_IO_L1_out_wrapper_286__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_286__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_286__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_286__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_286__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_286__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_286__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_286__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_286__ap_done) begin
            C_drain_IO_L1_out_wrapper_286__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_286__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_286__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_286__ap_done) begin
          C_drain_IO_L1_out_wrapper_286__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_286__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_286__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_286__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_286__ap_start = (C_drain_IO_L1_out_wrapper_286__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_287__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_287__is_done__q0 = (C_drain_IO_L1_out_wrapper_287__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_287__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_287__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_287__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_287__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_287__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_287__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_287__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_287__ap_done) begin
            C_drain_IO_L1_out_wrapper_287__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_287__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_287__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_287__ap_done) begin
          C_drain_IO_L1_out_wrapper_287__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_287__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_287__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_287__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_287__ap_start = (C_drain_IO_L1_out_wrapper_287__state == 2'b01);
  assign C_drain_IO_L1_out_wrapper_288__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L1_out_wrapper_288__is_done__q0 = (C_drain_IO_L1_out_wrapper_288__state == 2'b10);
  assign C_drain_IO_L1_out_wrapper_288__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L1_out_wrapper_288__state <= 2'b00;
    end else begin
      if(C_drain_IO_L1_out_wrapper_288__state == 2'b00) begin
        if(C_drain_IO_L1_out_wrapper_288__ap_start_global__q0) begin
          C_drain_IO_L1_out_wrapper_288__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_288__state == 2'b01) begin
        if(C_drain_IO_L1_out_wrapper_288__ap_ready) begin
          if(C_drain_IO_L1_out_wrapper_288__ap_done) begin
            C_drain_IO_L1_out_wrapper_288__state <= 2'b10;
          end else begin
            C_drain_IO_L1_out_wrapper_288__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_288__state == 2'b11) begin
        if(C_drain_IO_L1_out_wrapper_288__ap_done) begin
          C_drain_IO_L1_out_wrapper_288__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L1_out_wrapper_288__state == 2'b10) begin
        if(C_drain_IO_L1_out_wrapper_288__ap_done_global__q0) begin
          C_drain_IO_L1_out_wrapper_288__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L1_out_wrapper_288__ap_start = (C_drain_IO_L1_out_wrapper_288__state == 2'b01);
  assign C_drain_IO_L2_out_0__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L2_out_0__is_done__q0 = (C_drain_IO_L2_out_0__state == 2'b10);
  assign C_drain_IO_L2_out_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L2_out_0__state <= 2'b00;
    end else begin
      if(C_drain_IO_L2_out_0__state == 2'b00) begin
        if(C_drain_IO_L2_out_0__ap_start_global__q0) begin
          C_drain_IO_L2_out_0__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L2_out_0__state == 2'b01) begin
        if(C_drain_IO_L2_out_0__ap_ready) begin
          if(C_drain_IO_L2_out_0__ap_done) begin
            C_drain_IO_L2_out_0__state <= 2'b10;
          end else begin
            C_drain_IO_L2_out_0__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L2_out_0__state == 2'b11) begin
        if(C_drain_IO_L2_out_0__ap_done) begin
          C_drain_IO_L2_out_0__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L2_out_0__state == 2'b10) begin
        if(C_drain_IO_L2_out_0__ap_done_global__q0) begin
          C_drain_IO_L2_out_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L2_out_0__ap_start = (C_drain_IO_L2_out_0__state == 2'b01);
  assign C_drain_IO_L2_out_1__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L2_out_1__is_done__q0 = (C_drain_IO_L2_out_1__state == 2'b10);
  assign C_drain_IO_L2_out_1__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L2_out_1__state <= 2'b00;
    end else begin
      if(C_drain_IO_L2_out_1__state == 2'b00) begin
        if(C_drain_IO_L2_out_1__ap_start_global__q0) begin
          C_drain_IO_L2_out_1__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L2_out_1__state == 2'b01) begin
        if(C_drain_IO_L2_out_1__ap_ready) begin
          if(C_drain_IO_L2_out_1__ap_done) begin
            C_drain_IO_L2_out_1__state <= 2'b10;
          end else begin
            C_drain_IO_L2_out_1__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L2_out_1__state == 2'b11) begin
        if(C_drain_IO_L2_out_1__ap_done) begin
          C_drain_IO_L2_out_1__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L2_out_1__state == 2'b10) begin
        if(C_drain_IO_L2_out_1__ap_done_global__q0) begin
          C_drain_IO_L2_out_1__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L2_out_1__ap_start = (C_drain_IO_L2_out_1__state == 2'b01);
  assign C_drain_IO_L2_out_2__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L2_out_2__is_done__q0 = (C_drain_IO_L2_out_2__state == 2'b10);
  assign C_drain_IO_L2_out_2__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L2_out_2__state <= 2'b00;
    end else begin
      if(C_drain_IO_L2_out_2__state == 2'b00) begin
        if(C_drain_IO_L2_out_2__ap_start_global__q0) begin
          C_drain_IO_L2_out_2__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L2_out_2__state == 2'b01) begin
        if(C_drain_IO_L2_out_2__ap_ready) begin
          if(C_drain_IO_L2_out_2__ap_done) begin
            C_drain_IO_L2_out_2__state <= 2'b10;
          end else begin
            C_drain_IO_L2_out_2__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L2_out_2__state == 2'b11) begin
        if(C_drain_IO_L2_out_2__ap_done) begin
          C_drain_IO_L2_out_2__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L2_out_2__state == 2'b10) begin
        if(C_drain_IO_L2_out_2__ap_done_global__q0) begin
          C_drain_IO_L2_out_2__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L2_out_2__ap_start = (C_drain_IO_L2_out_2__state == 2'b01);
  assign C_drain_IO_L2_out_3__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L2_out_3__is_done__q0 = (C_drain_IO_L2_out_3__state == 2'b10);
  assign C_drain_IO_L2_out_3__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L2_out_3__state <= 2'b00;
    end else begin
      if(C_drain_IO_L2_out_3__state == 2'b00) begin
        if(C_drain_IO_L2_out_3__ap_start_global__q0) begin
          C_drain_IO_L2_out_3__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L2_out_3__state == 2'b01) begin
        if(C_drain_IO_L2_out_3__ap_ready) begin
          if(C_drain_IO_L2_out_3__ap_done) begin
            C_drain_IO_L2_out_3__state <= 2'b10;
          end else begin
            C_drain_IO_L2_out_3__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L2_out_3__state == 2'b11) begin
        if(C_drain_IO_L2_out_3__ap_done) begin
          C_drain_IO_L2_out_3__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L2_out_3__state == 2'b10) begin
        if(C_drain_IO_L2_out_3__ap_done_global__q0) begin
          C_drain_IO_L2_out_3__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L2_out_3__ap_start = (C_drain_IO_L2_out_3__state == 2'b01);
  assign C_drain_IO_L2_out_4__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L2_out_4__is_done__q0 = (C_drain_IO_L2_out_4__state == 2'b10);
  assign C_drain_IO_L2_out_4__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L2_out_4__state <= 2'b00;
    end else begin
      if(C_drain_IO_L2_out_4__state == 2'b00) begin
        if(C_drain_IO_L2_out_4__ap_start_global__q0) begin
          C_drain_IO_L2_out_4__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L2_out_4__state == 2'b01) begin
        if(C_drain_IO_L2_out_4__ap_ready) begin
          if(C_drain_IO_L2_out_4__ap_done) begin
            C_drain_IO_L2_out_4__state <= 2'b10;
          end else begin
            C_drain_IO_L2_out_4__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L2_out_4__state == 2'b11) begin
        if(C_drain_IO_L2_out_4__ap_done) begin
          C_drain_IO_L2_out_4__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L2_out_4__state == 2'b10) begin
        if(C_drain_IO_L2_out_4__ap_done_global__q0) begin
          C_drain_IO_L2_out_4__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L2_out_4__ap_start = (C_drain_IO_L2_out_4__state == 2'b01);
  assign C_drain_IO_L2_out_5__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L2_out_5__is_done__q0 = (C_drain_IO_L2_out_5__state == 2'b10);
  assign C_drain_IO_L2_out_5__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L2_out_5__state <= 2'b00;
    end else begin
      if(C_drain_IO_L2_out_5__state == 2'b00) begin
        if(C_drain_IO_L2_out_5__ap_start_global__q0) begin
          C_drain_IO_L2_out_5__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L2_out_5__state == 2'b01) begin
        if(C_drain_IO_L2_out_5__ap_ready) begin
          if(C_drain_IO_L2_out_5__ap_done) begin
            C_drain_IO_L2_out_5__state <= 2'b10;
          end else begin
            C_drain_IO_L2_out_5__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L2_out_5__state == 2'b11) begin
        if(C_drain_IO_L2_out_5__ap_done) begin
          C_drain_IO_L2_out_5__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L2_out_5__state == 2'b10) begin
        if(C_drain_IO_L2_out_5__ap_done_global__q0) begin
          C_drain_IO_L2_out_5__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L2_out_5__ap_start = (C_drain_IO_L2_out_5__state == 2'b01);
  assign C_drain_IO_L2_out_6__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L2_out_6__is_done__q0 = (C_drain_IO_L2_out_6__state == 2'b10);
  assign C_drain_IO_L2_out_6__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L2_out_6__state <= 2'b00;
    end else begin
      if(C_drain_IO_L2_out_6__state == 2'b00) begin
        if(C_drain_IO_L2_out_6__ap_start_global__q0) begin
          C_drain_IO_L2_out_6__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L2_out_6__state == 2'b01) begin
        if(C_drain_IO_L2_out_6__ap_ready) begin
          if(C_drain_IO_L2_out_6__ap_done) begin
            C_drain_IO_L2_out_6__state <= 2'b10;
          end else begin
            C_drain_IO_L2_out_6__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L2_out_6__state == 2'b11) begin
        if(C_drain_IO_L2_out_6__ap_done) begin
          C_drain_IO_L2_out_6__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L2_out_6__state == 2'b10) begin
        if(C_drain_IO_L2_out_6__ap_done_global__q0) begin
          C_drain_IO_L2_out_6__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L2_out_6__ap_start = (C_drain_IO_L2_out_6__state == 2'b01);
  assign C_drain_IO_L2_out_7__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L2_out_7__is_done__q0 = (C_drain_IO_L2_out_7__state == 2'b10);
  assign C_drain_IO_L2_out_7__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L2_out_7__state <= 2'b00;
    end else begin
      if(C_drain_IO_L2_out_7__state == 2'b00) begin
        if(C_drain_IO_L2_out_7__ap_start_global__q0) begin
          C_drain_IO_L2_out_7__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L2_out_7__state == 2'b01) begin
        if(C_drain_IO_L2_out_7__ap_ready) begin
          if(C_drain_IO_L2_out_7__ap_done) begin
            C_drain_IO_L2_out_7__state <= 2'b10;
          end else begin
            C_drain_IO_L2_out_7__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L2_out_7__state == 2'b11) begin
        if(C_drain_IO_L2_out_7__ap_done) begin
          C_drain_IO_L2_out_7__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L2_out_7__state == 2'b10) begin
        if(C_drain_IO_L2_out_7__ap_done_global__q0) begin
          C_drain_IO_L2_out_7__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L2_out_7__ap_start = (C_drain_IO_L2_out_7__state == 2'b01);
  assign C_drain_IO_L2_out_8__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L2_out_8__is_done__q0 = (C_drain_IO_L2_out_8__state == 2'b10);
  assign C_drain_IO_L2_out_8__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L2_out_8__state <= 2'b00;
    end else begin
      if(C_drain_IO_L2_out_8__state == 2'b00) begin
        if(C_drain_IO_L2_out_8__ap_start_global__q0) begin
          C_drain_IO_L2_out_8__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L2_out_8__state == 2'b01) begin
        if(C_drain_IO_L2_out_8__ap_ready) begin
          if(C_drain_IO_L2_out_8__ap_done) begin
            C_drain_IO_L2_out_8__state <= 2'b10;
          end else begin
            C_drain_IO_L2_out_8__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L2_out_8__state == 2'b11) begin
        if(C_drain_IO_L2_out_8__ap_done) begin
          C_drain_IO_L2_out_8__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L2_out_8__state == 2'b10) begin
        if(C_drain_IO_L2_out_8__ap_done_global__q0) begin
          C_drain_IO_L2_out_8__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L2_out_8__ap_start = (C_drain_IO_L2_out_8__state == 2'b01);
  assign C_drain_IO_L2_out_9__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L2_out_9__is_done__q0 = (C_drain_IO_L2_out_9__state == 2'b10);
  assign C_drain_IO_L2_out_9__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L2_out_9__state <= 2'b00;
    end else begin
      if(C_drain_IO_L2_out_9__state == 2'b00) begin
        if(C_drain_IO_L2_out_9__ap_start_global__q0) begin
          C_drain_IO_L2_out_9__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L2_out_9__state == 2'b01) begin
        if(C_drain_IO_L2_out_9__ap_ready) begin
          if(C_drain_IO_L2_out_9__ap_done) begin
            C_drain_IO_L2_out_9__state <= 2'b10;
          end else begin
            C_drain_IO_L2_out_9__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L2_out_9__state == 2'b11) begin
        if(C_drain_IO_L2_out_9__ap_done) begin
          C_drain_IO_L2_out_9__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L2_out_9__state == 2'b10) begin
        if(C_drain_IO_L2_out_9__ap_done_global__q0) begin
          C_drain_IO_L2_out_9__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L2_out_9__ap_start = (C_drain_IO_L2_out_9__state == 2'b01);
  assign C_drain_IO_L2_out_10__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L2_out_10__is_done__q0 = (C_drain_IO_L2_out_10__state == 2'b10);
  assign C_drain_IO_L2_out_10__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L2_out_10__state <= 2'b00;
    end else begin
      if(C_drain_IO_L2_out_10__state == 2'b00) begin
        if(C_drain_IO_L2_out_10__ap_start_global__q0) begin
          C_drain_IO_L2_out_10__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L2_out_10__state == 2'b01) begin
        if(C_drain_IO_L2_out_10__ap_ready) begin
          if(C_drain_IO_L2_out_10__ap_done) begin
            C_drain_IO_L2_out_10__state <= 2'b10;
          end else begin
            C_drain_IO_L2_out_10__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L2_out_10__state == 2'b11) begin
        if(C_drain_IO_L2_out_10__ap_done) begin
          C_drain_IO_L2_out_10__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L2_out_10__state == 2'b10) begin
        if(C_drain_IO_L2_out_10__ap_done_global__q0) begin
          C_drain_IO_L2_out_10__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L2_out_10__ap_start = (C_drain_IO_L2_out_10__state == 2'b01);
  assign C_drain_IO_L2_out_11__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L2_out_11__is_done__q0 = (C_drain_IO_L2_out_11__state == 2'b10);
  assign C_drain_IO_L2_out_11__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L2_out_11__state <= 2'b00;
    end else begin
      if(C_drain_IO_L2_out_11__state == 2'b00) begin
        if(C_drain_IO_L2_out_11__ap_start_global__q0) begin
          C_drain_IO_L2_out_11__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L2_out_11__state == 2'b01) begin
        if(C_drain_IO_L2_out_11__ap_ready) begin
          if(C_drain_IO_L2_out_11__ap_done) begin
            C_drain_IO_L2_out_11__state <= 2'b10;
          end else begin
            C_drain_IO_L2_out_11__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L2_out_11__state == 2'b11) begin
        if(C_drain_IO_L2_out_11__ap_done) begin
          C_drain_IO_L2_out_11__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L2_out_11__state == 2'b10) begin
        if(C_drain_IO_L2_out_11__ap_done_global__q0) begin
          C_drain_IO_L2_out_11__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L2_out_11__ap_start = (C_drain_IO_L2_out_11__state == 2'b01);
  assign C_drain_IO_L2_out_12__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L2_out_12__is_done__q0 = (C_drain_IO_L2_out_12__state == 2'b10);
  assign C_drain_IO_L2_out_12__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L2_out_12__state <= 2'b00;
    end else begin
      if(C_drain_IO_L2_out_12__state == 2'b00) begin
        if(C_drain_IO_L2_out_12__ap_start_global__q0) begin
          C_drain_IO_L2_out_12__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L2_out_12__state == 2'b01) begin
        if(C_drain_IO_L2_out_12__ap_ready) begin
          if(C_drain_IO_L2_out_12__ap_done) begin
            C_drain_IO_L2_out_12__state <= 2'b10;
          end else begin
            C_drain_IO_L2_out_12__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L2_out_12__state == 2'b11) begin
        if(C_drain_IO_L2_out_12__ap_done) begin
          C_drain_IO_L2_out_12__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L2_out_12__state == 2'b10) begin
        if(C_drain_IO_L2_out_12__ap_done_global__q0) begin
          C_drain_IO_L2_out_12__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L2_out_12__ap_start = (C_drain_IO_L2_out_12__state == 2'b01);
  assign C_drain_IO_L2_out_13__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L2_out_13__is_done__q0 = (C_drain_IO_L2_out_13__state == 2'b10);
  assign C_drain_IO_L2_out_13__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L2_out_13__state <= 2'b00;
    end else begin
      if(C_drain_IO_L2_out_13__state == 2'b00) begin
        if(C_drain_IO_L2_out_13__ap_start_global__q0) begin
          C_drain_IO_L2_out_13__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L2_out_13__state == 2'b01) begin
        if(C_drain_IO_L2_out_13__ap_ready) begin
          if(C_drain_IO_L2_out_13__ap_done) begin
            C_drain_IO_L2_out_13__state <= 2'b10;
          end else begin
            C_drain_IO_L2_out_13__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L2_out_13__state == 2'b11) begin
        if(C_drain_IO_L2_out_13__ap_done) begin
          C_drain_IO_L2_out_13__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L2_out_13__state == 2'b10) begin
        if(C_drain_IO_L2_out_13__ap_done_global__q0) begin
          C_drain_IO_L2_out_13__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L2_out_13__ap_start = (C_drain_IO_L2_out_13__state == 2'b01);
  assign C_drain_IO_L2_out_14__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L2_out_14__is_done__q0 = (C_drain_IO_L2_out_14__state == 2'b10);
  assign C_drain_IO_L2_out_14__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L2_out_14__state <= 2'b00;
    end else begin
      if(C_drain_IO_L2_out_14__state == 2'b00) begin
        if(C_drain_IO_L2_out_14__ap_start_global__q0) begin
          C_drain_IO_L2_out_14__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L2_out_14__state == 2'b01) begin
        if(C_drain_IO_L2_out_14__ap_ready) begin
          if(C_drain_IO_L2_out_14__ap_done) begin
            C_drain_IO_L2_out_14__state <= 2'b10;
          end else begin
            C_drain_IO_L2_out_14__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L2_out_14__state == 2'b11) begin
        if(C_drain_IO_L2_out_14__ap_done) begin
          C_drain_IO_L2_out_14__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L2_out_14__state == 2'b10) begin
        if(C_drain_IO_L2_out_14__ap_done_global__q0) begin
          C_drain_IO_L2_out_14__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L2_out_14__ap_start = (C_drain_IO_L2_out_14__state == 2'b01);
  assign C_drain_IO_L2_out_15__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L2_out_15__is_done__q0 = (C_drain_IO_L2_out_15__state == 2'b10);
  assign C_drain_IO_L2_out_15__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L2_out_15__state <= 2'b00;
    end else begin
      if(C_drain_IO_L2_out_15__state == 2'b00) begin
        if(C_drain_IO_L2_out_15__ap_start_global__q0) begin
          C_drain_IO_L2_out_15__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L2_out_15__state == 2'b01) begin
        if(C_drain_IO_L2_out_15__ap_ready) begin
          if(C_drain_IO_L2_out_15__ap_done) begin
            C_drain_IO_L2_out_15__state <= 2'b10;
          end else begin
            C_drain_IO_L2_out_15__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L2_out_15__state == 2'b11) begin
        if(C_drain_IO_L2_out_15__ap_done) begin
          C_drain_IO_L2_out_15__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L2_out_15__state == 2'b10) begin
        if(C_drain_IO_L2_out_15__ap_done_global__q0) begin
          C_drain_IO_L2_out_15__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L2_out_15__ap_start = (C_drain_IO_L2_out_15__state == 2'b01);
  assign C_drain_IO_L2_out_boundary_0__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L2_out_boundary_0__is_done__q0 = (C_drain_IO_L2_out_boundary_0__state == 2'b10);
  assign C_drain_IO_L2_out_boundary_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L2_out_boundary_0__state <= 2'b00;
    end else begin
      if(C_drain_IO_L2_out_boundary_0__state == 2'b00) begin
        if(C_drain_IO_L2_out_boundary_0__ap_start_global__q0) begin
          C_drain_IO_L2_out_boundary_0__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L2_out_boundary_0__state == 2'b01) begin
        if(C_drain_IO_L2_out_boundary_0__ap_ready) begin
          if(C_drain_IO_L2_out_boundary_0__ap_done) begin
            C_drain_IO_L2_out_boundary_0__state <= 2'b10;
          end else begin
            C_drain_IO_L2_out_boundary_0__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L2_out_boundary_0__state == 2'b11) begin
        if(C_drain_IO_L2_out_boundary_0__ap_done) begin
          C_drain_IO_L2_out_boundary_0__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L2_out_boundary_0__state == 2'b10) begin
        if(C_drain_IO_L2_out_boundary_0__ap_done_global__q0) begin
          C_drain_IO_L2_out_boundary_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L2_out_boundary_0__ap_start = (C_drain_IO_L2_out_boundary_0__state == 2'b01);
  assign C_drain_IO_L3_out_0__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L3_out_0__is_done__q0 = (C_drain_IO_L3_out_0__state == 2'b10);
  assign C_drain_IO_L3_out_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L3_out_0__state <= 2'b00;
    end else begin
      if(C_drain_IO_L3_out_0__state == 2'b00) begin
        if(C_drain_IO_L3_out_0__ap_start_global__q0) begin
          C_drain_IO_L3_out_0__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L3_out_0__state == 2'b01) begin
        if(C_drain_IO_L3_out_0__ap_ready) begin
          if(C_drain_IO_L3_out_0__ap_done) begin
            C_drain_IO_L3_out_0__state <= 2'b10;
          end else begin
            C_drain_IO_L3_out_0__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L3_out_0__state == 2'b11) begin
        if(C_drain_IO_L3_out_0__ap_done) begin
          C_drain_IO_L3_out_0__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L3_out_0__state == 2'b10) begin
        if(C_drain_IO_L3_out_0__ap_done_global__q0) begin
          C_drain_IO_L3_out_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L3_out_0__ap_start = (C_drain_IO_L3_out_0__state == 2'b01);
  assign C_drain_IO_L3_out_serialize_0___C__q0 = C;
  assign C_drain_IO_L3_out_serialize_0__ap_start_global__q0 = ap_start__q0;
  assign C_drain_IO_L3_out_serialize_0__is_done__q0 = (C_drain_IO_L3_out_serialize_0__state == 2'b10);
  assign C_drain_IO_L3_out_serialize_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      C_drain_IO_L3_out_serialize_0__state <= 2'b00;
    end else begin
      if(C_drain_IO_L3_out_serialize_0__state == 2'b00) begin
        if(C_drain_IO_L3_out_serialize_0__ap_start_global__q0) begin
          C_drain_IO_L3_out_serialize_0__state <= 2'b01;
        end 
      end 
      if(C_drain_IO_L3_out_serialize_0__state == 2'b01) begin
        if(C_drain_IO_L3_out_serialize_0__ap_ready) begin
          if(C_drain_IO_L3_out_serialize_0__ap_done) begin
            C_drain_IO_L3_out_serialize_0__state <= 2'b10;
          end else begin
            C_drain_IO_L3_out_serialize_0__state <= 2'b11;
          end
        end 
      end 
      if(C_drain_IO_L3_out_serialize_0__state == 2'b11) begin
        if(C_drain_IO_L3_out_serialize_0__ap_done) begin
          C_drain_IO_L3_out_serialize_0__state <= 2'b10;
        end 
      end 
      if(C_drain_IO_L3_out_serialize_0__state == 2'b10) begin
        if(C_drain_IO_L3_out_serialize_0__ap_done_global__q0) begin
          C_drain_IO_L3_out_serialize_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign C_drain_IO_L3_out_serialize_0__ap_start = (C_drain_IO_L3_out_serialize_0__state == 2'b01);
  assign PE_wrapper_0__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_0__is_done__q0 = (PE_wrapper_0__state == 2'b10);
  assign PE_wrapper_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_0__state <= 2'b00;
    end else begin
      if(PE_wrapper_0__state == 2'b00) begin
        if(PE_wrapper_0__ap_start_global__q0) begin
          PE_wrapper_0__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_0__state == 2'b01) begin
        if(PE_wrapper_0__ap_ready) begin
          if(PE_wrapper_0__ap_done) begin
            PE_wrapper_0__state <= 2'b10;
          end else begin
            PE_wrapper_0__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_0__state == 2'b11) begin
        if(PE_wrapper_0__ap_done) begin
          PE_wrapper_0__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_0__state == 2'b10) begin
        if(PE_wrapper_0__ap_done_global__q0) begin
          PE_wrapper_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_0__ap_start = (PE_wrapper_0__state == 2'b01);
  assign PE_wrapper_1__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_1__is_done__q0 = (PE_wrapper_1__state == 2'b10);
  assign PE_wrapper_1__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_1__state <= 2'b00;
    end else begin
      if(PE_wrapper_1__state == 2'b00) begin
        if(PE_wrapper_1__ap_start_global__q0) begin
          PE_wrapper_1__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_1__state == 2'b01) begin
        if(PE_wrapper_1__ap_ready) begin
          if(PE_wrapper_1__ap_done) begin
            PE_wrapper_1__state <= 2'b10;
          end else begin
            PE_wrapper_1__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_1__state == 2'b11) begin
        if(PE_wrapper_1__ap_done) begin
          PE_wrapper_1__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_1__state == 2'b10) begin
        if(PE_wrapper_1__ap_done_global__q0) begin
          PE_wrapper_1__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_1__ap_start = (PE_wrapper_1__state == 2'b01);
  assign PE_wrapper_2__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_2__is_done__q0 = (PE_wrapper_2__state == 2'b10);
  assign PE_wrapper_2__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_2__state <= 2'b00;
    end else begin
      if(PE_wrapper_2__state == 2'b00) begin
        if(PE_wrapper_2__ap_start_global__q0) begin
          PE_wrapper_2__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_2__state == 2'b01) begin
        if(PE_wrapper_2__ap_ready) begin
          if(PE_wrapper_2__ap_done) begin
            PE_wrapper_2__state <= 2'b10;
          end else begin
            PE_wrapper_2__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_2__state == 2'b11) begin
        if(PE_wrapper_2__ap_done) begin
          PE_wrapper_2__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_2__state == 2'b10) begin
        if(PE_wrapper_2__ap_done_global__q0) begin
          PE_wrapper_2__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_2__ap_start = (PE_wrapper_2__state == 2'b01);
  assign PE_wrapper_3__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_3__is_done__q0 = (PE_wrapper_3__state == 2'b10);
  assign PE_wrapper_3__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_3__state <= 2'b00;
    end else begin
      if(PE_wrapper_3__state == 2'b00) begin
        if(PE_wrapper_3__ap_start_global__q0) begin
          PE_wrapper_3__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_3__state == 2'b01) begin
        if(PE_wrapper_3__ap_ready) begin
          if(PE_wrapper_3__ap_done) begin
            PE_wrapper_3__state <= 2'b10;
          end else begin
            PE_wrapper_3__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_3__state == 2'b11) begin
        if(PE_wrapper_3__ap_done) begin
          PE_wrapper_3__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_3__state == 2'b10) begin
        if(PE_wrapper_3__ap_done_global__q0) begin
          PE_wrapper_3__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_3__ap_start = (PE_wrapper_3__state == 2'b01);
  assign PE_wrapper_4__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_4__is_done__q0 = (PE_wrapper_4__state == 2'b10);
  assign PE_wrapper_4__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_4__state <= 2'b00;
    end else begin
      if(PE_wrapper_4__state == 2'b00) begin
        if(PE_wrapper_4__ap_start_global__q0) begin
          PE_wrapper_4__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_4__state == 2'b01) begin
        if(PE_wrapper_4__ap_ready) begin
          if(PE_wrapper_4__ap_done) begin
            PE_wrapper_4__state <= 2'b10;
          end else begin
            PE_wrapper_4__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_4__state == 2'b11) begin
        if(PE_wrapper_4__ap_done) begin
          PE_wrapper_4__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_4__state == 2'b10) begin
        if(PE_wrapper_4__ap_done_global__q0) begin
          PE_wrapper_4__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_4__ap_start = (PE_wrapper_4__state == 2'b01);
  assign PE_wrapper_5__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_5__is_done__q0 = (PE_wrapper_5__state == 2'b10);
  assign PE_wrapper_5__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_5__state <= 2'b00;
    end else begin
      if(PE_wrapper_5__state == 2'b00) begin
        if(PE_wrapper_5__ap_start_global__q0) begin
          PE_wrapper_5__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_5__state == 2'b01) begin
        if(PE_wrapper_5__ap_ready) begin
          if(PE_wrapper_5__ap_done) begin
            PE_wrapper_5__state <= 2'b10;
          end else begin
            PE_wrapper_5__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_5__state == 2'b11) begin
        if(PE_wrapper_5__ap_done) begin
          PE_wrapper_5__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_5__state == 2'b10) begin
        if(PE_wrapper_5__ap_done_global__q0) begin
          PE_wrapper_5__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_5__ap_start = (PE_wrapper_5__state == 2'b01);
  assign PE_wrapper_6__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_6__is_done__q0 = (PE_wrapper_6__state == 2'b10);
  assign PE_wrapper_6__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_6__state <= 2'b00;
    end else begin
      if(PE_wrapper_6__state == 2'b00) begin
        if(PE_wrapper_6__ap_start_global__q0) begin
          PE_wrapper_6__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_6__state == 2'b01) begin
        if(PE_wrapper_6__ap_ready) begin
          if(PE_wrapper_6__ap_done) begin
            PE_wrapper_6__state <= 2'b10;
          end else begin
            PE_wrapper_6__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_6__state == 2'b11) begin
        if(PE_wrapper_6__ap_done) begin
          PE_wrapper_6__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_6__state == 2'b10) begin
        if(PE_wrapper_6__ap_done_global__q0) begin
          PE_wrapper_6__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_6__ap_start = (PE_wrapper_6__state == 2'b01);
  assign PE_wrapper_7__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_7__is_done__q0 = (PE_wrapper_7__state == 2'b10);
  assign PE_wrapper_7__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_7__state <= 2'b00;
    end else begin
      if(PE_wrapper_7__state == 2'b00) begin
        if(PE_wrapper_7__ap_start_global__q0) begin
          PE_wrapper_7__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_7__state == 2'b01) begin
        if(PE_wrapper_7__ap_ready) begin
          if(PE_wrapper_7__ap_done) begin
            PE_wrapper_7__state <= 2'b10;
          end else begin
            PE_wrapper_7__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_7__state == 2'b11) begin
        if(PE_wrapper_7__ap_done) begin
          PE_wrapper_7__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_7__state == 2'b10) begin
        if(PE_wrapper_7__ap_done_global__q0) begin
          PE_wrapper_7__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_7__ap_start = (PE_wrapper_7__state == 2'b01);
  assign PE_wrapper_8__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_8__is_done__q0 = (PE_wrapper_8__state == 2'b10);
  assign PE_wrapper_8__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_8__state <= 2'b00;
    end else begin
      if(PE_wrapper_8__state == 2'b00) begin
        if(PE_wrapper_8__ap_start_global__q0) begin
          PE_wrapper_8__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_8__state == 2'b01) begin
        if(PE_wrapper_8__ap_ready) begin
          if(PE_wrapper_8__ap_done) begin
            PE_wrapper_8__state <= 2'b10;
          end else begin
            PE_wrapper_8__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_8__state == 2'b11) begin
        if(PE_wrapper_8__ap_done) begin
          PE_wrapper_8__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_8__state == 2'b10) begin
        if(PE_wrapper_8__ap_done_global__q0) begin
          PE_wrapper_8__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_8__ap_start = (PE_wrapper_8__state == 2'b01);
  assign PE_wrapper_9__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_9__is_done__q0 = (PE_wrapper_9__state == 2'b10);
  assign PE_wrapper_9__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_9__state <= 2'b00;
    end else begin
      if(PE_wrapper_9__state == 2'b00) begin
        if(PE_wrapper_9__ap_start_global__q0) begin
          PE_wrapper_9__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_9__state == 2'b01) begin
        if(PE_wrapper_9__ap_ready) begin
          if(PE_wrapper_9__ap_done) begin
            PE_wrapper_9__state <= 2'b10;
          end else begin
            PE_wrapper_9__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_9__state == 2'b11) begin
        if(PE_wrapper_9__ap_done) begin
          PE_wrapper_9__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_9__state == 2'b10) begin
        if(PE_wrapper_9__ap_done_global__q0) begin
          PE_wrapper_9__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_9__ap_start = (PE_wrapper_9__state == 2'b01);
  assign PE_wrapper_10__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_10__is_done__q0 = (PE_wrapper_10__state == 2'b10);
  assign PE_wrapper_10__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_10__state <= 2'b00;
    end else begin
      if(PE_wrapper_10__state == 2'b00) begin
        if(PE_wrapper_10__ap_start_global__q0) begin
          PE_wrapper_10__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_10__state == 2'b01) begin
        if(PE_wrapper_10__ap_ready) begin
          if(PE_wrapper_10__ap_done) begin
            PE_wrapper_10__state <= 2'b10;
          end else begin
            PE_wrapper_10__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_10__state == 2'b11) begin
        if(PE_wrapper_10__ap_done) begin
          PE_wrapper_10__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_10__state == 2'b10) begin
        if(PE_wrapper_10__ap_done_global__q0) begin
          PE_wrapper_10__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_10__ap_start = (PE_wrapper_10__state == 2'b01);
  assign PE_wrapper_11__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_11__is_done__q0 = (PE_wrapper_11__state == 2'b10);
  assign PE_wrapper_11__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_11__state <= 2'b00;
    end else begin
      if(PE_wrapper_11__state == 2'b00) begin
        if(PE_wrapper_11__ap_start_global__q0) begin
          PE_wrapper_11__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_11__state == 2'b01) begin
        if(PE_wrapper_11__ap_ready) begin
          if(PE_wrapper_11__ap_done) begin
            PE_wrapper_11__state <= 2'b10;
          end else begin
            PE_wrapper_11__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_11__state == 2'b11) begin
        if(PE_wrapper_11__ap_done) begin
          PE_wrapper_11__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_11__state == 2'b10) begin
        if(PE_wrapper_11__ap_done_global__q0) begin
          PE_wrapper_11__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_11__ap_start = (PE_wrapper_11__state == 2'b01);
  assign PE_wrapper_12__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_12__is_done__q0 = (PE_wrapper_12__state == 2'b10);
  assign PE_wrapper_12__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_12__state <= 2'b00;
    end else begin
      if(PE_wrapper_12__state == 2'b00) begin
        if(PE_wrapper_12__ap_start_global__q0) begin
          PE_wrapper_12__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_12__state == 2'b01) begin
        if(PE_wrapper_12__ap_ready) begin
          if(PE_wrapper_12__ap_done) begin
            PE_wrapper_12__state <= 2'b10;
          end else begin
            PE_wrapper_12__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_12__state == 2'b11) begin
        if(PE_wrapper_12__ap_done) begin
          PE_wrapper_12__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_12__state == 2'b10) begin
        if(PE_wrapper_12__ap_done_global__q0) begin
          PE_wrapper_12__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_12__ap_start = (PE_wrapper_12__state == 2'b01);
  assign PE_wrapper_13__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_13__is_done__q0 = (PE_wrapper_13__state == 2'b10);
  assign PE_wrapper_13__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_13__state <= 2'b00;
    end else begin
      if(PE_wrapper_13__state == 2'b00) begin
        if(PE_wrapper_13__ap_start_global__q0) begin
          PE_wrapper_13__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_13__state == 2'b01) begin
        if(PE_wrapper_13__ap_ready) begin
          if(PE_wrapper_13__ap_done) begin
            PE_wrapper_13__state <= 2'b10;
          end else begin
            PE_wrapper_13__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_13__state == 2'b11) begin
        if(PE_wrapper_13__ap_done) begin
          PE_wrapper_13__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_13__state == 2'b10) begin
        if(PE_wrapper_13__ap_done_global__q0) begin
          PE_wrapper_13__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_13__ap_start = (PE_wrapper_13__state == 2'b01);
  assign PE_wrapper_14__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_14__is_done__q0 = (PE_wrapper_14__state == 2'b10);
  assign PE_wrapper_14__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_14__state <= 2'b00;
    end else begin
      if(PE_wrapper_14__state == 2'b00) begin
        if(PE_wrapper_14__ap_start_global__q0) begin
          PE_wrapper_14__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_14__state == 2'b01) begin
        if(PE_wrapper_14__ap_ready) begin
          if(PE_wrapper_14__ap_done) begin
            PE_wrapper_14__state <= 2'b10;
          end else begin
            PE_wrapper_14__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_14__state == 2'b11) begin
        if(PE_wrapper_14__ap_done) begin
          PE_wrapper_14__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_14__state == 2'b10) begin
        if(PE_wrapper_14__ap_done_global__q0) begin
          PE_wrapper_14__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_14__ap_start = (PE_wrapper_14__state == 2'b01);
  assign PE_wrapper_15__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_15__is_done__q0 = (PE_wrapper_15__state == 2'b10);
  assign PE_wrapper_15__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_15__state <= 2'b00;
    end else begin
      if(PE_wrapper_15__state == 2'b00) begin
        if(PE_wrapper_15__ap_start_global__q0) begin
          PE_wrapper_15__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_15__state == 2'b01) begin
        if(PE_wrapper_15__ap_ready) begin
          if(PE_wrapper_15__ap_done) begin
            PE_wrapper_15__state <= 2'b10;
          end else begin
            PE_wrapper_15__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_15__state == 2'b11) begin
        if(PE_wrapper_15__ap_done) begin
          PE_wrapper_15__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_15__state == 2'b10) begin
        if(PE_wrapper_15__ap_done_global__q0) begin
          PE_wrapper_15__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_15__ap_start = (PE_wrapper_15__state == 2'b01);
  assign PE_wrapper_16__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_16__is_done__q0 = (PE_wrapper_16__state == 2'b10);
  assign PE_wrapper_16__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_16__state <= 2'b00;
    end else begin
      if(PE_wrapper_16__state == 2'b00) begin
        if(PE_wrapper_16__ap_start_global__q0) begin
          PE_wrapper_16__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_16__state == 2'b01) begin
        if(PE_wrapper_16__ap_ready) begin
          if(PE_wrapper_16__ap_done) begin
            PE_wrapper_16__state <= 2'b10;
          end else begin
            PE_wrapper_16__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_16__state == 2'b11) begin
        if(PE_wrapper_16__ap_done) begin
          PE_wrapper_16__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_16__state == 2'b10) begin
        if(PE_wrapper_16__ap_done_global__q0) begin
          PE_wrapper_16__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_16__ap_start = (PE_wrapper_16__state == 2'b01);
  assign PE_wrapper_17__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_17__is_done__q0 = (PE_wrapper_17__state == 2'b10);
  assign PE_wrapper_17__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_17__state <= 2'b00;
    end else begin
      if(PE_wrapper_17__state == 2'b00) begin
        if(PE_wrapper_17__ap_start_global__q0) begin
          PE_wrapper_17__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_17__state == 2'b01) begin
        if(PE_wrapper_17__ap_ready) begin
          if(PE_wrapper_17__ap_done) begin
            PE_wrapper_17__state <= 2'b10;
          end else begin
            PE_wrapper_17__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_17__state == 2'b11) begin
        if(PE_wrapper_17__ap_done) begin
          PE_wrapper_17__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_17__state == 2'b10) begin
        if(PE_wrapper_17__ap_done_global__q0) begin
          PE_wrapper_17__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_17__ap_start = (PE_wrapper_17__state == 2'b01);
  assign PE_wrapper_18__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_18__is_done__q0 = (PE_wrapper_18__state == 2'b10);
  assign PE_wrapper_18__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_18__state <= 2'b00;
    end else begin
      if(PE_wrapper_18__state == 2'b00) begin
        if(PE_wrapper_18__ap_start_global__q0) begin
          PE_wrapper_18__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_18__state == 2'b01) begin
        if(PE_wrapper_18__ap_ready) begin
          if(PE_wrapper_18__ap_done) begin
            PE_wrapper_18__state <= 2'b10;
          end else begin
            PE_wrapper_18__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_18__state == 2'b11) begin
        if(PE_wrapper_18__ap_done) begin
          PE_wrapper_18__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_18__state == 2'b10) begin
        if(PE_wrapper_18__ap_done_global__q0) begin
          PE_wrapper_18__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_18__ap_start = (PE_wrapper_18__state == 2'b01);
  assign PE_wrapper_19__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_19__is_done__q0 = (PE_wrapper_19__state == 2'b10);
  assign PE_wrapper_19__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_19__state <= 2'b00;
    end else begin
      if(PE_wrapper_19__state == 2'b00) begin
        if(PE_wrapper_19__ap_start_global__q0) begin
          PE_wrapper_19__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_19__state == 2'b01) begin
        if(PE_wrapper_19__ap_ready) begin
          if(PE_wrapper_19__ap_done) begin
            PE_wrapper_19__state <= 2'b10;
          end else begin
            PE_wrapper_19__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_19__state == 2'b11) begin
        if(PE_wrapper_19__ap_done) begin
          PE_wrapper_19__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_19__state == 2'b10) begin
        if(PE_wrapper_19__ap_done_global__q0) begin
          PE_wrapper_19__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_19__ap_start = (PE_wrapper_19__state == 2'b01);
  assign PE_wrapper_20__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_20__is_done__q0 = (PE_wrapper_20__state == 2'b10);
  assign PE_wrapper_20__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_20__state <= 2'b00;
    end else begin
      if(PE_wrapper_20__state == 2'b00) begin
        if(PE_wrapper_20__ap_start_global__q0) begin
          PE_wrapper_20__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_20__state == 2'b01) begin
        if(PE_wrapper_20__ap_ready) begin
          if(PE_wrapper_20__ap_done) begin
            PE_wrapper_20__state <= 2'b10;
          end else begin
            PE_wrapper_20__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_20__state == 2'b11) begin
        if(PE_wrapper_20__ap_done) begin
          PE_wrapper_20__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_20__state == 2'b10) begin
        if(PE_wrapper_20__ap_done_global__q0) begin
          PE_wrapper_20__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_20__ap_start = (PE_wrapper_20__state == 2'b01);
  assign PE_wrapper_21__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_21__is_done__q0 = (PE_wrapper_21__state == 2'b10);
  assign PE_wrapper_21__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_21__state <= 2'b00;
    end else begin
      if(PE_wrapper_21__state == 2'b00) begin
        if(PE_wrapper_21__ap_start_global__q0) begin
          PE_wrapper_21__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_21__state == 2'b01) begin
        if(PE_wrapper_21__ap_ready) begin
          if(PE_wrapper_21__ap_done) begin
            PE_wrapper_21__state <= 2'b10;
          end else begin
            PE_wrapper_21__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_21__state == 2'b11) begin
        if(PE_wrapper_21__ap_done) begin
          PE_wrapper_21__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_21__state == 2'b10) begin
        if(PE_wrapper_21__ap_done_global__q0) begin
          PE_wrapper_21__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_21__ap_start = (PE_wrapper_21__state == 2'b01);
  assign PE_wrapper_22__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_22__is_done__q0 = (PE_wrapper_22__state == 2'b10);
  assign PE_wrapper_22__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_22__state <= 2'b00;
    end else begin
      if(PE_wrapper_22__state == 2'b00) begin
        if(PE_wrapper_22__ap_start_global__q0) begin
          PE_wrapper_22__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_22__state == 2'b01) begin
        if(PE_wrapper_22__ap_ready) begin
          if(PE_wrapper_22__ap_done) begin
            PE_wrapper_22__state <= 2'b10;
          end else begin
            PE_wrapper_22__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_22__state == 2'b11) begin
        if(PE_wrapper_22__ap_done) begin
          PE_wrapper_22__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_22__state == 2'b10) begin
        if(PE_wrapper_22__ap_done_global__q0) begin
          PE_wrapper_22__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_22__ap_start = (PE_wrapper_22__state == 2'b01);
  assign PE_wrapper_23__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_23__is_done__q0 = (PE_wrapper_23__state == 2'b10);
  assign PE_wrapper_23__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_23__state <= 2'b00;
    end else begin
      if(PE_wrapper_23__state == 2'b00) begin
        if(PE_wrapper_23__ap_start_global__q0) begin
          PE_wrapper_23__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_23__state == 2'b01) begin
        if(PE_wrapper_23__ap_ready) begin
          if(PE_wrapper_23__ap_done) begin
            PE_wrapper_23__state <= 2'b10;
          end else begin
            PE_wrapper_23__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_23__state == 2'b11) begin
        if(PE_wrapper_23__ap_done) begin
          PE_wrapper_23__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_23__state == 2'b10) begin
        if(PE_wrapper_23__ap_done_global__q0) begin
          PE_wrapper_23__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_23__ap_start = (PE_wrapper_23__state == 2'b01);
  assign PE_wrapper_24__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_24__is_done__q0 = (PE_wrapper_24__state == 2'b10);
  assign PE_wrapper_24__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_24__state <= 2'b00;
    end else begin
      if(PE_wrapper_24__state == 2'b00) begin
        if(PE_wrapper_24__ap_start_global__q0) begin
          PE_wrapper_24__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_24__state == 2'b01) begin
        if(PE_wrapper_24__ap_ready) begin
          if(PE_wrapper_24__ap_done) begin
            PE_wrapper_24__state <= 2'b10;
          end else begin
            PE_wrapper_24__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_24__state == 2'b11) begin
        if(PE_wrapper_24__ap_done) begin
          PE_wrapper_24__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_24__state == 2'b10) begin
        if(PE_wrapper_24__ap_done_global__q0) begin
          PE_wrapper_24__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_24__ap_start = (PE_wrapper_24__state == 2'b01);
  assign PE_wrapper_25__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_25__is_done__q0 = (PE_wrapper_25__state == 2'b10);
  assign PE_wrapper_25__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_25__state <= 2'b00;
    end else begin
      if(PE_wrapper_25__state == 2'b00) begin
        if(PE_wrapper_25__ap_start_global__q0) begin
          PE_wrapper_25__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_25__state == 2'b01) begin
        if(PE_wrapper_25__ap_ready) begin
          if(PE_wrapper_25__ap_done) begin
            PE_wrapper_25__state <= 2'b10;
          end else begin
            PE_wrapper_25__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_25__state == 2'b11) begin
        if(PE_wrapper_25__ap_done) begin
          PE_wrapper_25__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_25__state == 2'b10) begin
        if(PE_wrapper_25__ap_done_global__q0) begin
          PE_wrapper_25__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_25__ap_start = (PE_wrapper_25__state == 2'b01);
  assign PE_wrapper_26__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_26__is_done__q0 = (PE_wrapper_26__state == 2'b10);
  assign PE_wrapper_26__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_26__state <= 2'b00;
    end else begin
      if(PE_wrapper_26__state == 2'b00) begin
        if(PE_wrapper_26__ap_start_global__q0) begin
          PE_wrapper_26__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_26__state == 2'b01) begin
        if(PE_wrapper_26__ap_ready) begin
          if(PE_wrapper_26__ap_done) begin
            PE_wrapper_26__state <= 2'b10;
          end else begin
            PE_wrapper_26__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_26__state == 2'b11) begin
        if(PE_wrapper_26__ap_done) begin
          PE_wrapper_26__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_26__state == 2'b10) begin
        if(PE_wrapper_26__ap_done_global__q0) begin
          PE_wrapper_26__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_26__ap_start = (PE_wrapper_26__state == 2'b01);
  assign PE_wrapper_27__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_27__is_done__q0 = (PE_wrapper_27__state == 2'b10);
  assign PE_wrapper_27__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_27__state <= 2'b00;
    end else begin
      if(PE_wrapper_27__state == 2'b00) begin
        if(PE_wrapper_27__ap_start_global__q0) begin
          PE_wrapper_27__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_27__state == 2'b01) begin
        if(PE_wrapper_27__ap_ready) begin
          if(PE_wrapper_27__ap_done) begin
            PE_wrapper_27__state <= 2'b10;
          end else begin
            PE_wrapper_27__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_27__state == 2'b11) begin
        if(PE_wrapper_27__ap_done) begin
          PE_wrapper_27__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_27__state == 2'b10) begin
        if(PE_wrapper_27__ap_done_global__q0) begin
          PE_wrapper_27__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_27__ap_start = (PE_wrapper_27__state == 2'b01);
  assign PE_wrapper_28__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_28__is_done__q0 = (PE_wrapper_28__state == 2'b10);
  assign PE_wrapper_28__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_28__state <= 2'b00;
    end else begin
      if(PE_wrapper_28__state == 2'b00) begin
        if(PE_wrapper_28__ap_start_global__q0) begin
          PE_wrapper_28__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_28__state == 2'b01) begin
        if(PE_wrapper_28__ap_ready) begin
          if(PE_wrapper_28__ap_done) begin
            PE_wrapper_28__state <= 2'b10;
          end else begin
            PE_wrapper_28__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_28__state == 2'b11) begin
        if(PE_wrapper_28__ap_done) begin
          PE_wrapper_28__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_28__state == 2'b10) begin
        if(PE_wrapper_28__ap_done_global__q0) begin
          PE_wrapper_28__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_28__ap_start = (PE_wrapper_28__state == 2'b01);
  assign PE_wrapper_29__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_29__is_done__q0 = (PE_wrapper_29__state == 2'b10);
  assign PE_wrapper_29__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_29__state <= 2'b00;
    end else begin
      if(PE_wrapper_29__state == 2'b00) begin
        if(PE_wrapper_29__ap_start_global__q0) begin
          PE_wrapper_29__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_29__state == 2'b01) begin
        if(PE_wrapper_29__ap_ready) begin
          if(PE_wrapper_29__ap_done) begin
            PE_wrapper_29__state <= 2'b10;
          end else begin
            PE_wrapper_29__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_29__state == 2'b11) begin
        if(PE_wrapper_29__ap_done) begin
          PE_wrapper_29__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_29__state == 2'b10) begin
        if(PE_wrapper_29__ap_done_global__q0) begin
          PE_wrapper_29__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_29__ap_start = (PE_wrapper_29__state == 2'b01);
  assign PE_wrapper_30__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_30__is_done__q0 = (PE_wrapper_30__state == 2'b10);
  assign PE_wrapper_30__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_30__state <= 2'b00;
    end else begin
      if(PE_wrapper_30__state == 2'b00) begin
        if(PE_wrapper_30__ap_start_global__q0) begin
          PE_wrapper_30__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_30__state == 2'b01) begin
        if(PE_wrapper_30__ap_ready) begin
          if(PE_wrapper_30__ap_done) begin
            PE_wrapper_30__state <= 2'b10;
          end else begin
            PE_wrapper_30__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_30__state == 2'b11) begin
        if(PE_wrapper_30__ap_done) begin
          PE_wrapper_30__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_30__state == 2'b10) begin
        if(PE_wrapper_30__ap_done_global__q0) begin
          PE_wrapper_30__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_30__ap_start = (PE_wrapper_30__state == 2'b01);
  assign PE_wrapper_31__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_31__is_done__q0 = (PE_wrapper_31__state == 2'b10);
  assign PE_wrapper_31__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_31__state <= 2'b00;
    end else begin
      if(PE_wrapper_31__state == 2'b00) begin
        if(PE_wrapper_31__ap_start_global__q0) begin
          PE_wrapper_31__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_31__state == 2'b01) begin
        if(PE_wrapper_31__ap_ready) begin
          if(PE_wrapper_31__ap_done) begin
            PE_wrapper_31__state <= 2'b10;
          end else begin
            PE_wrapper_31__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_31__state == 2'b11) begin
        if(PE_wrapper_31__ap_done) begin
          PE_wrapper_31__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_31__state == 2'b10) begin
        if(PE_wrapper_31__ap_done_global__q0) begin
          PE_wrapper_31__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_31__ap_start = (PE_wrapper_31__state == 2'b01);
  assign PE_wrapper_32__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_32__is_done__q0 = (PE_wrapper_32__state == 2'b10);
  assign PE_wrapper_32__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_32__state <= 2'b00;
    end else begin
      if(PE_wrapper_32__state == 2'b00) begin
        if(PE_wrapper_32__ap_start_global__q0) begin
          PE_wrapper_32__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_32__state == 2'b01) begin
        if(PE_wrapper_32__ap_ready) begin
          if(PE_wrapper_32__ap_done) begin
            PE_wrapper_32__state <= 2'b10;
          end else begin
            PE_wrapper_32__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_32__state == 2'b11) begin
        if(PE_wrapper_32__ap_done) begin
          PE_wrapper_32__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_32__state == 2'b10) begin
        if(PE_wrapper_32__ap_done_global__q0) begin
          PE_wrapper_32__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_32__ap_start = (PE_wrapper_32__state == 2'b01);
  assign PE_wrapper_33__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_33__is_done__q0 = (PE_wrapper_33__state == 2'b10);
  assign PE_wrapper_33__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_33__state <= 2'b00;
    end else begin
      if(PE_wrapper_33__state == 2'b00) begin
        if(PE_wrapper_33__ap_start_global__q0) begin
          PE_wrapper_33__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_33__state == 2'b01) begin
        if(PE_wrapper_33__ap_ready) begin
          if(PE_wrapper_33__ap_done) begin
            PE_wrapper_33__state <= 2'b10;
          end else begin
            PE_wrapper_33__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_33__state == 2'b11) begin
        if(PE_wrapper_33__ap_done) begin
          PE_wrapper_33__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_33__state == 2'b10) begin
        if(PE_wrapper_33__ap_done_global__q0) begin
          PE_wrapper_33__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_33__ap_start = (PE_wrapper_33__state == 2'b01);
  assign PE_wrapper_34__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_34__is_done__q0 = (PE_wrapper_34__state == 2'b10);
  assign PE_wrapper_34__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_34__state <= 2'b00;
    end else begin
      if(PE_wrapper_34__state == 2'b00) begin
        if(PE_wrapper_34__ap_start_global__q0) begin
          PE_wrapper_34__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_34__state == 2'b01) begin
        if(PE_wrapper_34__ap_ready) begin
          if(PE_wrapper_34__ap_done) begin
            PE_wrapper_34__state <= 2'b10;
          end else begin
            PE_wrapper_34__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_34__state == 2'b11) begin
        if(PE_wrapper_34__ap_done) begin
          PE_wrapper_34__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_34__state == 2'b10) begin
        if(PE_wrapper_34__ap_done_global__q0) begin
          PE_wrapper_34__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_34__ap_start = (PE_wrapper_34__state == 2'b01);
  assign PE_wrapper_35__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_35__is_done__q0 = (PE_wrapper_35__state == 2'b10);
  assign PE_wrapper_35__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_35__state <= 2'b00;
    end else begin
      if(PE_wrapper_35__state == 2'b00) begin
        if(PE_wrapper_35__ap_start_global__q0) begin
          PE_wrapper_35__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_35__state == 2'b01) begin
        if(PE_wrapper_35__ap_ready) begin
          if(PE_wrapper_35__ap_done) begin
            PE_wrapper_35__state <= 2'b10;
          end else begin
            PE_wrapper_35__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_35__state == 2'b11) begin
        if(PE_wrapper_35__ap_done) begin
          PE_wrapper_35__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_35__state == 2'b10) begin
        if(PE_wrapper_35__ap_done_global__q0) begin
          PE_wrapper_35__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_35__ap_start = (PE_wrapper_35__state == 2'b01);
  assign PE_wrapper_36__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_36__is_done__q0 = (PE_wrapper_36__state == 2'b10);
  assign PE_wrapper_36__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_36__state <= 2'b00;
    end else begin
      if(PE_wrapper_36__state == 2'b00) begin
        if(PE_wrapper_36__ap_start_global__q0) begin
          PE_wrapper_36__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_36__state == 2'b01) begin
        if(PE_wrapper_36__ap_ready) begin
          if(PE_wrapper_36__ap_done) begin
            PE_wrapper_36__state <= 2'b10;
          end else begin
            PE_wrapper_36__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_36__state == 2'b11) begin
        if(PE_wrapper_36__ap_done) begin
          PE_wrapper_36__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_36__state == 2'b10) begin
        if(PE_wrapper_36__ap_done_global__q0) begin
          PE_wrapper_36__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_36__ap_start = (PE_wrapper_36__state == 2'b01);
  assign PE_wrapper_37__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_37__is_done__q0 = (PE_wrapper_37__state == 2'b10);
  assign PE_wrapper_37__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_37__state <= 2'b00;
    end else begin
      if(PE_wrapper_37__state == 2'b00) begin
        if(PE_wrapper_37__ap_start_global__q0) begin
          PE_wrapper_37__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_37__state == 2'b01) begin
        if(PE_wrapper_37__ap_ready) begin
          if(PE_wrapper_37__ap_done) begin
            PE_wrapper_37__state <= 2'b10;
          end else begin
            PE_wrapper_37__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_37__state == 2'b11) begin
        if(PE_wrapper_37__ap_done) begin
          PE_wrapper_37__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_37__state == 2'b10) begin
        if(PE_wrapper_37__ap_done_global__q0) begin
          PE_wrapper_37__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_37__ap_start = (PE_wrapper_37__state == 2'b01);
  assign PE_wrapper_38__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_38__is_done__q0 = (PE_wrapper_38__state == 2'b10);
  assign PE_wrapper_38__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_38__state <= 2'b00;
    end else begin
      if(PE_wrapper_38__state == 2'b00) begin
        if(PE_wrapper_38__ap_start_global__q0) begin
          PE_wrapper_38__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_38__state == 2'b01) begin
        if(PE_wrapper_38__ap_ready) begin
          if(PE_wrapper_38__ap_done) begin
            PE_wrapper_38__state <= 2'b10;
          end else begin
            PE_wrapper_38__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_38__state == 2'b11) begin
        if(PE_wrapper_38__ap_done) begin
          PE_wrapper_38__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_38__state == 2'b10) begin
        if(PE_wrapper_38__ap_done_global__q0) begin
          PE_wrapper_38__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_38__ap_start = (PE_wrapper_38__state == 2'b01);
  assign PE_wrapper_39__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_39__is_done__q0 = (PE_wrapper_39__state == 2'b10);
  assign PE_wrapper_39__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_39__state <= 2'b00;
    end else begin
      if(PE_wrapper_39__state == 2'b00) begin
        if(PE_wrapper_39__ap_start_global__q0) begin
          PE_wrapper_39__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_39__state == 2'b01) begin
        if(PE_wrapper_39__ap_ready) begin
          if(PE_wrapper_39__ap_done) begin
            PE_wrapper_39__state <= 2'b10;
          end else begin
            PE_wrapper_39__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_39__state == 2'b11) begin
        if(PE_wrapper_39__ap_done) begin
          PE_wrapper_39__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_39__state == 2'b10) begin
        if(PE_wrapper_39__ap_done_global__q0) begin
          PE_wrapper_39__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_39__ap_start = (PE_wrapper_39__state == 2'b01);
  assign PE_wrapper_40__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_40__is_done__q0 = (PE_wrapper_40__state == 2'b10);
  assign PE_wrapper_40__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_40__state <= 2'b00;
    end else begin
      if(PE_wrapper_40__state == 2'b00) begin
        if(PE_wrapper_40__ap_start_global__q0) begin
          PE_wrapper_40__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_40__state == 2'b01) begin
        if(PE_wrapper_40__ap_ready) begin
          if(PE_wrapper_40__ap_done) begin
            PE_wrapper_40__state <= 2'b10;
          end else begin
            PE_wrapper_40__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_40__state == 2'b11) begin
        if(PE_wrapper_40__ap_done) begin
          PE_wrapper_40__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_40__state == 2'b10) begin
        if(PE_wrapper_40__ap_done_global__q0) begin
          PE_wrapper_40__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_40__ap_start = (PE_wrapper_40__state == 2'b01);
  assign PE_wrapper_41__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_41__is_done__q0 = (PE_wrapper_41__state == 2'b10);
  assign PE_wrapper_41__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_41__state <= 2'b00;
    end else begin
      if(PE_wrapper_41__state == 2'b00) begin
        if(PE_wrapper_41__ap_start_global__q0) begin
          PE_wrapper_41__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_41__state == 2'b01) begin
        if(PE_wrapper_41__ap_ready) begin
          if(PE_wrapper_41__ap_done) begin
            PE_wrapper_41__state <= 2'b10;
          end else begin
            PE_wrapper_41__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_41__state == 2'b11) begin
        if(PE_wrapper_41__ap_done) begin
          PE_wrapper_41__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_41__state == 2'b10) begin
        if(PE_wrapper_41__ap_done_global__q0) begin
          PE_wrapper_41__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_41__ap_start = (PE_wrapper_41__state == 2'b01);
  assign PE_wrapper_42__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_42__is_done__q0 = (PE_wrapper_42__state == 2'b10);
  assign PE_wrapper_42__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_42__state <= 2'b00;
    end else begin
      if(PE_wrapper_42__state == 2'b00) begin
        if(PE_wrapper_42__ap_start_global__q0) begin
          PE_wrapper_42__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_42__state == 2'b01) begin
        if(PE_wrapper_42__ap_ready) begin
          if(PE_wrapper_42__ap_done) begin
            PE_wrapper_42__state <= 2'b10;
          end else begin
            PE_wrapper_42__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_42__state == 2'b11) begin
        if(PE_wrapper_42__ap_done) begin
          PE_wrapper_42__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_42__state == 2'b10) begin
        if(PE_wrapper_42__ap_done_global__q0) begin
          PE_wrapper_42__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_42__ap_start = (PE_wrapper_42__state == 2'b01);
  assign PE_wrapper_43__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_43__is_done__q0 = (PE_wrapper_43__state == 2'b10);
  assign PE_wrapper_43__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_43__state <= 2'b00;
    end else begin
      if(PE_wrapper_43__state == 2'b00) begin
        if(PE_wrapper_43__ap_start_global__q0) begin
          PE_wrapper_43__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_43__state == 2'b01) begin
        if(PE_wrapper_43__ap_ready) begin
          if(PE_wrapper_43__ap_done) begin
            PE_wrapper_43__state <= 2'b10;
          end else begin
            PE_wrapper_43__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_43__state == 2'b11) begin
        if(PE_wrapper_43__ap_done) begin
          PE_wrapper_43__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_43__state == 2'b10) begin
        if(PE_wrapper_43__ap_done_global__q0) begin
          PE_wrapper_43__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_43__ap_start = (PE_wrapper_43__state == 2'b01);
  assign PE_wrapper_44__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_44__is_done__q0 = (PE_wrapper_44__state == 2'b10);
  assign PE_wrapper_44__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_44__state <= 2'b00;
    end else begin
      if(PE_wrapper_44__state == 2'b00) begin
        if(PE_wrapper_44__ap_start_global__q0) begin
          PE_wrapper_44__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_44__state == 2'b01) begin
        if(PE_wrapper_44__ap_ready) begin
          if(PE_wrapper_44__ap_done) begin
            PE_wrapper_44__state <= 2'b10;
          end else begin
            PE_wrapper_44__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_44__state == 2'b11) begin
        if(PE_wrapper_44__ap_done) begin
          PE_wrapper_44__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_44__state == 2'b10) begin
        if(PE_wrapper_44__ap_done_global__q0) begin
          PE_wrapper_44__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_44__ap_start = (PE_wrapper_44__state == 2'b01);
  assign PE_wrapper_45__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_45__is_done__q0 = (PE_wrapper_45__state == 2'b10);
  assign PE_wrapper_45__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_45__state <= 2'b00;
    end else begin
      if(PE_wrapper_45__state == 2'b00) begin
        if(PE_wrapper_45__ap_start_global__q0) begin
          PE_wrapper_45__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_45__state == 2'b01) begin
        if(PE_wrapper_45__ap_ready) begin
          if(PE_wrapper_45__ap_done) begin
            PE_wrapper_45__state <= 2'b10;
          end else begin
            PE_wrapper_45__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_45__state == 2'b11) begin
        if(PE_wrapper_45__ap_done) begin
          PE_wrapper_45__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_45__state == 2'b10) begin
        if(PE_wrapper_45__ap_done_global__q0) begin
          PE_wrapper_45__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_45__ap_start = (PE_wrapper_45__state == 2'b01);
  assign PE_wrapper_46__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_46__is_done__q0 = (PE_wrapper_46__state == 2'b10);
  assign PE_wrapper_46__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_46__state <= 2'b00;
    end else begin
      if(PE_wrapper_46__state == 2'b00) begin
        if(PE_wrapper_46__ap_start_global__q0) begin
          PE_wrapper_46__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_46__state == 2'b01) begin
        if(PE_wrapper_46__ap_ready) begin
          if(PE_wrapper_46__ap_done) begin
            PE_wrapper_46__state <= 2'b10;
          end else begin
            PE_wrapper_46__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_46__state == 2'b11) begin
        if(PE_wrapper_46__ap_done) begin
          PE_wrapper_46__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_46__state == 2'b10) begin
        if(PE_wrapper_46__ap_done_global__q0) begin
          PE_wrapper_46__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_46__ap_start = (PE_wrapper_46__state == 2'b01);
  assign PE_wrapper_47__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_47__is_done__q0 = (PE_wrapper_47__state == 2'b10);
  assign PE_wrapper_47__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_47__state <= 2'b00;
    end else begin
      if(PE_wrapper_47__state == 2'b00) begin
        if(PE_wrapper_47__ap_start_global__q0) begin
          PE_wrapper_47__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_47__state == 2'b01) begin
        if(PE_wrapper_47__ap_ready) begin
          if(PE_wrapper_47__ap_done) begin
            PE_wrapper_47__state <= 2'b10;
          end else begin
            PE_wrapper_47__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_47__state == 2'b11) begin
        if(PE_wrapper_47__ap_done) begin
          PE_wrapper_47__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_47__state == 2'b10) begin
        if(PE_wrapper_47__ap_done_global__q0) begin
          PE_wrapper_47__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_47__ap_start = (PE_wrapper_47__state == 2'b01);
  assign PE_wrapper_48__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_48__is_done__q0 = (PE_wrapper_48__state == 2'b10);
  assign PE_wrapper_48__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_48__state <= 2'b00;
    end else begin
      if(PE_wrapper_48__state == 2'b00) begin
        if(PE_wrapper_48__ap_start_global__q0) begin
          PE_wrapper_48__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_48__state == 2'b01) begin
        if(PE_wrapper_48__ap_ready) begin
          if(PE_wrapper_48__ap_done) begin
            PE_wrapper_48__state <= 2'b10;
          end else begin
            PE_wrapper_48__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_48__state == 2'b11) begin
        if(PE_wrapper_48__ap_done) begin
          PE_wrapper_48__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_48__state == 2'b10) begin
        if(PE_wrapper_48__ap_done_global__q0) begin
          PE_wrapper_48__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_48__ap_start = (PE_wrapper_48__state == 2'b01);
  assign PE_wrapper_49__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_49__is_done__q0 = (PE_wrapper_49__state == 2'b10);
  assign PE_wrapper_49__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_49__state <= 2'b00;
    end else begin
      if(PE_wrapper_49__state == 2'b00) begin
        if(PE_wrapper_49__ap_start_global__q0) begin
          PE_wrapper_49__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_49__state == 2'b01) begin
        if(PE_wrapper_49__ap_ready) begin
          if(PE_wrapper_49__ap_done) begin
            PE_wrapper_49__state <= 2'b10;
          end else begin
            PE_wrapper_49__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_49__state == 2'b11) begin
        if(PE_wrapper_49__ap_done) begin
          PE_wrapper_49__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_49__state == 2'b10) begin
        if(PE_wrapper_49__ap_done_global__q0) begin
          PE_wrapper_49__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_49__ap_start = (PE_wrapper_49__state == 2'b01);
  assign PE_wrapper_50__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_50__is_done__q0 = (PE_wrapper_50__state == 2'b10);
  assign PE_wrapper_50__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_50__state <= 2'b00;
    end else begin
      if(PE_wrapper_50__state == 2'b00) begin
        if(PE_wrapper_50__ap_start_global__q0) begin
          PE_wrapper_50__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_50__state == 2'b01) begin
        if(PE_wrapper_50__ap_ready) begin
          if(PE_wrapper_50__ap_done) begin
            PE_wrapper_50__state <= 2'b10;
          end else begin
            PE_wrapper_50__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_50__state == 2'b11) begin
        if(PE_wrapper_50__ap_done) begin
          PE_wrapper_50__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_50__state == 2'b10) begin
        if(PE_wrapper_50__ap_done_global__q0) begin
          PE_wrapper_50__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_50__ap_start = (PE_wrapper_50__state == 2'b01);
  assign PE_wrapper_51__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_51__is_done__q0 = (PE_wrapper_51__state == 2'b10);
  assign PE_wrapper_51__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_51__state <= 2'b00;
    end else begin
      if(PE_wrapper_51__state == 2'b00) begin
        if(PE_wrapper_51__ap_start_global__q0) begin
          PE_wrapper_51__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_51__state == 2'b01) begin
        if(PE_wrapper_51__ap_ready) begin
          if(PE_wrapper_51__ap_done) begin
            PE_wrapper_51__state <= 2'b10;
          end else begin
            PE_wrapper_51__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_51__state == 2'b11) begin
        if(PE_wrapper_51__ap_done) begin
          PE_wrapper_51__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_51__state == 2'b10) begin
        if(PE_wrapper_51__ap_done_global__q0) begin
          PE_wrapper_51__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_51__ap_start = (PE_wrapper_51__state == 2'b01);
  assign PE_wrapper_52__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_52__is_done__q0 = (PE_wrapper_52__state == 2'b10);
  assign PE_wrapper_52__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_52__state <= 2'b00;
    end else begin
      if(PE_wrapper_52__state == 2'b00) begin
        if(PE_wrapper_52__ap_start_global__q0) begin
          PE_wrapper_52__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_52__state == 2'b01) begin
        if(PE_wrapper_52__ap_ready) begin
          if(PE_wrapper_52__ap_done) begin
            PE_wrapper_52__state <= 2'b10;
          end else begin
            PE_wrapper_52__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_52__state == 2'b11) begin
        if(PE_wrapper_52__ap_done) begin
          PE_wrapper_52__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_52__state == 2'b10) begin
        if(PE_wrapper_52__ap_done_global__q0) begin
          PE_wrapper_52__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_52__ap_start = (PE_wrapper_52__state == 2'b01);
  assign PE_wrapper_53__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_53__is_done__q0 = (PE_wrapper_53__state == 2'b10);
  assign PE_wrapper_53__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_53__state <= 2'b00;
    end else begin
      if(PE_wrapper_53__state == 2'b00) begin
        if(PE_wrapper_53__ap_start_global__q0) begin
          PE_wrapper_53__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_53__state == 2'b01) begin
        if(PE_wrapper_53__ap_ready) begin
          if(PE_wrapper_53__ap_done) begin
            PE_wrapper_53__state <= 2'b10;
          end else begin
            PE_wrapper_53__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_53__state == 2'b11) begin
        if(PE_wrapper_53__ap_done) begin
          PE_wrapper_53__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_53__state == 2'b10) begin
        if(PE_wrapper_53__ap_done_global__q0) begin
          PE_wrapper_53__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_53__ap_start = (PE_wrapper_53__state == 2'b01);
  assign PE_wrapper_54__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_54__is_done__q0 = (PE_wrapper_54__state == 2'b10);
  assign PE_wrapper_54__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_54__state <= 2'b00;
    end else begin
      if(PE_wrapper_54__state == 2'b00) begin
        if(PE_wrapper_54__ap_start_global__q0) begin
          PE_wrapper_54__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_54__state == 2'b01) begin
        if(PE_wrapper_54__ap_ready) begin
          if(PE_wrapper_54__ap_done) begin
            PE_wrapper_54__state <= 2'b10;
          end else begin
            PE_wrapper_54__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_54__state == 2'b11) begin
        if(PE_wrapper_54__ap_done) begin
          PE_wrapper_54__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_54__state == 2'b10) begin
        if(PE_wrapper_54__ap_done_global__q0) begin
          PE_wrapper_54__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_54__ap_start = (PE_wrapper_54__state == 2'b01);
  assign PE_wrapper_55__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_55__is_done__q0 = (PE_wrapper_55__state == 2'b10);
  assign PE_wrapper_55__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_55__state <= 2'b00;
    end else begin
      if(PE_wrapper_55__state == 2'b00) begin
        if(PE_wrapper_55__ap_start_global__q0) begin
          PE_wrapper_55__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_55__state == 2'b01) begin
        if(PE_wrapper_55__ap_ready) begin
          if(PE_wrapper_55__ap_done) begin
            PE_wrapper_55__state <= 2'b10;
          end else begin
            PE_wrapper_55__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_55__state == 2'b11) begin
        if(PE_wrapper_55__ap_done) begin
          PE_wrapper_55__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_55__state == 2'b10) begin
        if(PE_wrapper_55__ap_done_global__q0) begin
          PE_wrapper_55__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_55__ap_start = (PE_wrapper_55__state == 2'b01);
  assign PE_wrapper_56__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_56__is_done__q0 = (PE_wrapper_56__state == 2'b10);
  assign PE_wrapper_56__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_56__state <= 2'b00;
    end else begin
      if(PE_wrapper_56__state == 2'b00) begin
        if(PE_wrapper_56__ap_start_global__q0) begin
          PE_wrapper_56__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_56__state == 2'b01) begin
        if(PE_wrapper_56__ap_ready) begin
          if(PE_wrapper_56__ap_done) begin
            PE_wrapper_56__state <= 2'b10;
          end else begin
            PE_wrapper_56__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_56__state == 2'b11) begin
        if(PE_wrapper_56__ap_done) begin
          PE_wrapper_56__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_56__state == 2'b10) begin
        if(PE_wrapper_56__ap_done_global__q0) begin
          PE_wrapper_56__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_56__ap_start = (PE_wrapper_56__state == 2'b01);
  assign PE_wrapper_57__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_57__is_done__q0 = (PE_wrapper_57__state == 2'b10);
  assign PE_wrapper_57__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_57__state <= 2'b00;
    end else begin
      if(PE_wrapper_57__state == 2'b00) begin
        if(PE_wrapper_57__ap_start_global__q0) begin
          PE_wrapper_57__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_57__state == 2'b01) begin
        if(PE_wrapper_57__ap_ready) begin
          if(PE_wrapper_57__ap_done) begin
            PE_wrapper_57__state <= 2'b10;
          end else begin
            PE_wrapper_57__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_57__state == 2'b11) begin
        if(PE_wrapper_57__ap_done) begin
          PE_wrapper_57__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_57__state == 2'b10) begin
        if(PE_wrapper_57__ap_done_global__q0) begin
          PE_wrapper_57__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_57__ap_start = (PE_wrapper_57__state == 2'b01);
  assign PE_wrapper_58__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_58__is_done__q0 = (PE_wrapper_58__state == 2'b10);
  assign PE_wrapper_58__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_58__state <= 2'b00;
    end else begin
      if(PE_wrapper_58__state == 2'b00) begin
        if(PE_wrapper_58__ap_start_global__q0) begin
          PE_wrapper_58__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_58__state == 2'b01) begin
        if(PE_wrapper_58__ap_ready) begin
          if(PE_wrapper_58__ap_done) begin
            PE_wrapper_58__state <= 2'b10;
          end else begin
            PE_wrapper_58__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_58__state == 2'b11) begin
        if(PE_wrapper_58__ap_done) begin
          PE_wrapper_58__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_58__state == 2'b10) begin
        if(PE_wrapper_58__ap_done_global__q0) begin
          PE_wrapper_58__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_58__ap_start = (PE_wrapper_58__state == 2'b01);
  assign PE_wrapper_59__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_59__is_done__q0 = (PE_wrapper_59__state == 2'b10);
  assign PE_wrapper_59__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_59__state <= 2'b00;
    end else begin
      if(PE_wrapper_59__state == 2'b00) begin
        if(PE_wrapper_59__ap_start_global__q0) begin
          PE_wrapper_59__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_59__state == 2'b01) begin
        if(PE_wrapper_59__ap_ready) begin
          if(PE_wrapper_59__ap_done) begin
            PE_wrapper_59__state <= 2'b10;
          end else begin
            PE_wrapper_59__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_59__state == 2'b11) begin
        if(PE_wrapper_59__ap_done) begin
          PE_wrapper_59__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_59__state == 2'b10) begin
        if(PE_wrapper_59__ap_done_global__q0) begin
          PE_wrapper_59__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_59__ap_start = (PE_wrapper_59__state == 2'b01);
  assign PE_wrapper_60__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_60__is_done__q0 = (PE_wrapper_60__state == 2'b10);
  assign PE_wrapper_60__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_60__state <= 2'b00;
    end else begin
      if(PE_wrapper_60__state == 2'b00) begin
        if(PE_wrapper_60__ap_start_global__q0) begin
          PE_wrapper_60__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_60__state == 2'b01) begin
        if(PE_wrapper_60__ap_ready) begin
          if(PE_wrapper_60__ap_done) begin
            PE_wrapper_60__state <= 2'b10;
          end else begin
            PE_wrapper_60__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_60__state == 2'b11) begin
        if(PE_wrapper_60__ap_done) begin
          PE_wrapper_60__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_60__state == 2'b10) begin
        if(PE_wrapper_60__ap_done_global__q0) begin
          PE_wrapper_60__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_60__ap_start = (PE_wrapper_60__state == 2'b01);
  assign PE_wrapper_61__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_61__is_done__q0 = (PE_wrapper_61__state == 2'b10);
  assign PE_wrapper_61__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_61__state <= 2'b00;
    end else begin
      if(PE_wrapper_61__state == 2'b00) begin
        if(PE_wrapper_61__ap_start_global__q0) begin
          PE_wrapper_61__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_61__state == 2'b01) begin
        if(PE_wrapper_61__ap_ready) begin
          if(PE_wrapper_61__ap_done) begin
            PE_wrapper_61__state <= 2'b10;
          end else begin
            PE_wrapper_61__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_61__state == 2'b11) begin
        if(PE_wrapper_61__ap_done) begin
          PE_wrapper_61__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_61__state == 2'b10) begin
        if(PE_wrapper_61__ap_done_global__q0) begin
          PE_wrapper_61__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_61__ap_start = (PE_wrapper_61__state == 2'b01);
  assign PE_wrapper_62__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_62__is_done__q0 = (PE_wrapper_62__state == 2'b10);
  assign PE_wrapper_62__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_62__state <= 2'b00;
    end else begin
      if(PE_wrapper_62__state == 2'b00) begin
        if(PE_wrapper_62__ap_start_global__q0) begin
          PE_wrapper_62__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_62__state == 2'b01) begin
        if(PE_wrapper_62__ap_ready) begin
          if(PE_wrapper_62__ap_done) begin
            PE_wrapper_62__state <= 2'b10;
          end else begin
            PE_wrapper_62__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_62__state == 2'b11) begin
        if(PE_wrapper_62__ap_done) begin
          PE_wrapper_62__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_62__state == 2'b10) begin
        if(PE_wrapper_62__ap_done_global__q0) begin
          PE_wrapper_62__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_62__ap_start = (PE_wrapper_62__state == 2'b01);
  assign PE_wrapper_63__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_63__is_done__q0 = (PE_wrapper_63__state == 2'b10);
  assign PE_wrapper_63__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_63__state <= 2'b00;
    end else begin
      if(PE_wrapper_63__state == 2'b00) begin
        if(PE_wrapper_63__ap_start_global__q0) begin
          PE_wrapper_63__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_63__state == 2'b01) begin
        if(PE_wrapper_63__ap_ready) begin
          if(PE_wrapper_63__ap_done) begin
            PE_wrapper_63__state <= 2'b10;
          end else begin
            PE_wrapper_63__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_63__state == 2'b11) begin
        if(PE_wrapper_63__ap_done) begin
          PE_wrapper_63__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_63__state == 2'b10) begin
        if(PE_wrapper_63__ap_done_global__q0) begin
          PE_wrapper_63__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_63__ap_start = (PE_wrapper_63__state == 2'b01);
  assign PE_wrapper_64__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_64__is_done__q0 = (PE_wrapper_64__state == 2'b10);
  assign PE_wrapper_64__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_64__state <= 2'b00;
    end else begin
      if(PE_wrapper_64__state == 2'b00) begin
        if(PE_wrapper_64__ap_start_global__q0) begin
          PE_wrapper_64__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_64__state == 2'b01) begin
        if(PE_wrapper_64__ap_ready) begin
          if(PE_wrapper_64__ap_done) begin
            PE_wrapper_64__state <= 2'b10;
          end else begin
            PE_wrapper_64__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_64__state == 2'b11) begin
        if(PE_wrapper_64__ap_done) begin
          PE_wrapper_64__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_64__state == 2'b10) begin
        if(PE_wrapper_64__ap_done_global__q0) begin
          PE_wrapper_64__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_64__ap_start = (PE_wrapper_64__state == 2'b01);
  assign PE_wrapper_65__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_65__is_done__q0 = (PE_wrapper_65__state == 2'b10);
  assign PE_wrapper_65__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_65__state <= 2'b00;
    end else begin
      if(PE_wrapper_65__state == 2'b00) begin
        if(PE_wrapper_65__ap_start_global__q0) begin
          PE_wrapper_65__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_65__state == 2'b01) begin
        if(PE_wrapper_65__ap_ready) begin
          if(PE_wrapper_65__ap_done) begin
            PE_wrapper_65__state <= 2'b10;
          end else begin
            PE_wrapper_65__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_65__state == 2'b11) begin
        if(PE_wrapper_65__ap_done) begin
          PE_wrapper_65__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_65__state == 2'b10) begin
        if(PE_wrapper_65__ap_done_global__q0) begin
          PE_wrapper_65__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_65__ap_start = (PE_wrapper_65__state == 2'b01);
  assign PE_wrapper_66__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_66__is_done__q0 = (PE_wrapper_66__state == 2'b10);
  assign PE_wrapper_66__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_66__state <= 2'b00;
    end else begin
      if(PE_wrapper_66__state == 2'b00) begin
        if(PE_wrapper_66__ap_start_global__q0) begin
          PE_wrapper_66__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_66__state == 2'b01) begin
        if(PE_wrapper_66__ap_ready) begin
          if(PE_wrapper_66__ap_done) begin
            PE_wrapper_66__state <= 2'b10;
          end else begin
            PE_wrapper_66__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_66__state == 2'b11) begin
        if(PE_wrapper_66__ap_done) begin
          PE_wrapper_66__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_66__state == 2'b10) begin
        if(PE_wrapper_66__ap_done_global__q0) begin
          PE_wrapper_66__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_66__ap_start = (PE_wrapper_66__state == 2'b01);
  assign PE_wrapper_67__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_67__is_done__q0 = (PE_wrapper_67__state == 2'b10);
  assign PE_wrapper_67__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_67__state <= 2'b00;
    end else begin
      if(PE_wrapper_67__state == 2'b00) begin
        if(PE_wrapper_67__ap_start_global__q0) begin
          PE_wrapper_67__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_67__state == 2'b01) begin
        if(PE_wrapper_67__ap_ready) begin
          if(PE_wrapper_67__ap_done) begin
            PE_wrapper_67__state <= 2'b10;
          end else begin
            PE_wrapper_67__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_67__state == 2'b11) begin
        if(PE_wrapper_67__ap_done) begin
          PE_wrapper_67__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_67__state == 2'b10) begin
        if(PE_wrapper_67__ap_done_global__q0) begin
          PE_wrapper_67__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_67__ap_start = (PE_wrapper_67__state == 2'b01);
  assign PE_wrapper_68__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_68__is_done__q0 = (PE_wrapper_68__state == 2'b10);
  assign PE_wrapper_68__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_68__state <= 2'b00;
    end else begin
      if(PE_wrapper_68__state == 2'b00) begin
        if(PE_wrapper_68__ap_start_global__q0) begin
          PE_wrapper_68__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_68__state == 2'b01) begin
        if(PE_wrapper_68__ap_ready) begin
          if(PE_wrapper_68__ap_done) begin
            PE_wrapper_68__state <= 2'b10;
          end else begin
            PE_wrapper_68__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_68__state == 2'b11) begin
        if(PE_wrapper_68__ap_done) begin
          PE_wrapper_68__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_68__state == 2'b10) begin
        if(PE_wrapper_68__ap_done_global__q0) begin
          PE_wrapper_68__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_68__ap_start = (PE_wrapper_68__state == 2'b01);
  assign PE_wrapper_69__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_69__is_done__q0 = (PE_wrapper_69__state == 2'b10);
  assign PE_wrapper_69__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_69__state <= 2'b00;
    end else begin
      if(PE_wrapper_69__state == 2'b00) begin
        if(PE_wrapper_69__ap_start_global__q0) begin
          PE_wrapper_69__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_69__state == 2'b01) begin
        if(PE_wrapper_69__ap_ready) begin
          if(PE_wrapper_69__ap_done) begin
            PE_wrapper_69__state <= 2'b10;
          end else begin
            PE_wrapper_69__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_69__state == 2'b11) begin
        if(PE_wrapper_69__ap_done) begin
          PE_wrapper_69__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_69__state == 2'b10) begin
        if(PE_wrapper_69__ap_done_global__q0) begin
          PE_wrapper_69__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_69__ap_start = (PE_wrapper_69__state == 2'b01);
  assign PE_wrapper_70__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_70__is_done__q0 = (PE_wrapper_70__state == 2'b10);
  assign PE_wrapper_70__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_70__state <= 2'b00;
    end else begin
      if(PE_wrapper_70__state == 2'b00) begin
        if(PE_wrapper_70__ap_start_global__q0) begin
          PE_wrapper_70__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_70__state == 2'b01) begin
        if(PE_wrapper_70__ap_ready) begin
          if(PE_wrapper_70__ap_done) begin
            PE_wrapper_70__state <= 2'b10;
          end else begin
            PE_wrapper_70__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_70__state == 2'b11) begin
        if(PE_wrapper_70__ap_done) begin
          PE_wrapper_70__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_70__state == 2'b10) begin
        if(PE_wrapper_70__ap_done_global__q0) begin
          PE_wrapper_70__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_70__ap_start = (PE_wrapper_70__state == 2'b01);
  assign PE_wrapper_71__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_71__is_done__q0 = (PE_wrapper_71__state == 2'b10);
  assign PE_wrapper_71__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_71__state <= 2'b00;
    end else begin
      if(PE_wrapper_71__state == 2'b00) begin
        if(PE_wrapper_71__ap_start_global__q0) begin
          PE_wrapper_71__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_71__state == 2'b01) begin
        if(PE_wrapper_71__ap_ready) begin
          if(PE_wrapper_71__ap_done) begin
            PE_wrapper_71__state <= 2'b10;
          end else begin
            PE_wrapper_71__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_71__state == 2'b11) begin
        if(PE_wrapper_71__ap_done) begin
          PE_wrapper_71__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_71__state == 2'b10) begin
        if(PE_wrapper_71__ap_done_global__q0) begin
          PE_wrapper_71__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_71__ap_start = (PE_wrapper_71__state == 2'b01);
  assign PE_wrapper_72__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_72__is_done__q0 = (PE_wrapper_72__state == 2'b10);
  assign PE_wrapper_72__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_72__state <= 2'b00;
    end else begin
      if(PE_wrapper_72__state == 2'b00) begin
        if(PE_wrapper_72__ap_start_global__q0) begin
          PE_wrapper_72__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_72__state == 2'b01) begin
        if(PE_wrapper_72__ap_ready) begin
          if(PE_wrapper_72__ap_done) begin
            PE_wrapper_72__state <= 2'b10;
          end else begin
            PE_wrapper_72__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_72__state == 2'b11) begin
        if(PE_wrapper_72__ap_done) begin
          PE_wrapper_72__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_72__state == 2'b10) begin
        if(PE_wrapper_72__ap_done_global__q0) begin
          PE_wrapper_72__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_72__ap_start = (PE_wrapper_72__state == 2'b01);
  assign PE_wrapper_73__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_73__is_done__q0 = (PE_wrapper_73__state == 2'b10);
  assign PE_wrapper_73__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_73__state <= 2'b00;
    end else begin
      if(PE_wrapper_73__state == 2'b00) begin
        if(PE_wrapper_73__ap_start_global__q0) begin
          PE_wrapper_73__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_73__state == 2'b01) begin
        if(PE_wrapper_73__ap_ready) begin
          if(PE_wrapper_73__ap_done) begin
            PE_wrapper_73__state <= 2'b10;
          end else begin
            PE_wrapper_73__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_73__state == 2'b11) begin
        if(PE_wrapper_73__ap_done) begin
          PE_wrapper_73__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_73__state == 2'b10) begin
        if(PE_wrapper_73__ap_done_global__q0) begin
          PE_wrapper_73__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_73__ap_start = (PE_wrapper_73__state == 2'b01);
  assign PE_wrapper_74__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_74__is_done__q0 = (PE_wrapper_74__state == 2'b10);
  assign PE_wrapper_74__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_74__state <= 2'b00;
    end else begin
      if(PE_wrapper_74__state == 2'b00) begin
        if(PE_wrapper_74__ap_start_global__q0) begin
          PE_wrapper_74__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_74__state == 2'b01) begin
        if(PE_wrapper_74__ap_ready) begin
          if(PE_wrapper_74__ap_done) begin
            PE_wrapper_74__state <= 2'b10;
          end else begin
            PE_wrapper_74__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_74__state == 2'b11) begin
        if(PE_wrapper_74__ap_done) begin
          PE_wrapper_74__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_74__state == 2'b10) begin
        if(PE_wrapper_74__ap_done_global__q0) begin
          PE_wrapper_74__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_74__ap_start = (PE_wrapper_74__state == 2'b01);
  assign PE_wrapper_75__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_75__is_done__q0 = (PE_wrapper_75__state == 2'b10);
  assign PE_wrapper_75__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_75__state <= 2'b00;
    end else begin
      if(PE_wrapper_75__state == 2'b00) begin
        if(PE_wrapper_75__ap_start_global__q0) begin
          PE_wrapper_75__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_75__state == 2'b01) begin
        if(PE_wrapper_75__ap_ready) begin
          if(PE_wrapper_75__ap_done) begin
            PE_wrapper_75__state <= 2'b10;
          end else begin
            PE_wrapper_75__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_75__state == 2'b11) begin
        if(PE_wrapper_75__ap_done) begin
          PE_wrapper_75__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_75__state == 2'b10) begin
        if(PE_wrapper_75__ap_done_global__q0) begin
          PE_wrapper_75__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_75__ap_start = (PE_wrapper_75__state == 2'b01);
  assign PE_wrapper_76__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_76__is_done__q0 = (PE_wrapper_76__state == 2'b10);
  assign PE_wrapper_76__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_76__state <= 2'b00;
    end else begin
      if(PE_wrapper_76__state == 2'b00) begin
        if(PE_wrapper_76__ap_start_global__q0) begin
          PE_wrapper_76__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_76__state == 2'b01) begin
        if(PE_wrapper_76__ap_ready) begin
          if(PE_wrapper_76__ap_done) begin
            PE_wrapper_76__state <= 2'b10;
          end else begin
            PE_wrapper_76__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_76__state == 2'b11) begin
        if(PE_wrapper_76__ap_done) begin
          PE_wrapper_76__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_76__state == 2'b10) begin
        if(PE_wrapper_76__ap_done_global__q0) begin
          PE_wrapper_76__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_76__ap_start = (PE_wrapper_76__state == 2'b01);
  assign PE_wrapper_77__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_77__is_done__q0 = (PE_wrapper_77__state == 2'b10);
  assign PE_wrapper_77__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_77__state <= 2'b00;
    end else begin
      if(PE_wrapper_77__state == 2'b00) begin
        if(PE_wrapper_77__ap_start_global__q0) begin
          PE_wrapper_77__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_77__state == 2'b01) begin
        if(PE_wrapper_77__ap_ready) begin
          if(PE_wrapper_77__ap_done) begin
            PE_wrapper_77__state <= 2'b10;
          end else begin
            PE_wrapper_77__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_77__state == 2'b11) begin
        if(PE_wrapper_77__ap_done) begin
          PE_wrapper_77__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_77__state == 2'b10) begin
        if(PE_wrapper_77__ap_done_global__q0) begin
          PE_wrapper_77__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_77__ap_start = (PE_wrapper_77__state == 2'b01);
  assign PE_wrapper_78__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_78__is_done__q0 = (PE_wrapper_78__state == 2'b10);
  assign PE_wrapper_78__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_78__state <= 2'b00;
    end else begin
      if(PE_wrapper_78__state == 2'b00) begin
        if(PE_wrapper_78__ap_start_global__q0) begin
          PE_wrapper_78__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_78__state == 2'b01) begin
        if(PE_wrapper_78__ap_ready) begin
          if(PE_wrapper_78__ap_done) begin
            PE_wrapper_78__state <= 2'b10;
          end else begin
            PE_wrapper_78__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_78__state == 2'b11) begin
        if(PE_wrapper_78__ap_done) begin
          PE_wrapper_78__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_78__state == 2'b10) begin
        if(PE_wrapper_78__ap_done_global__q0) begin
          PE_wrapper_78__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_78__ap_start = (PE_wrapper_78__state == 2'b01);
  assign PE_wrapper_79__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_79__is_done__q0 = (PE_wrapper_79__state == 2'b10);
  assign PE_wrapper_79__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_79__state <= 2'b00;
    end else begin
      if(PE_wrapper_79__state == 2'b00) begin
        if(PE_wrapper_79__ap_start_global__q0) begin
          PE_wrapper_79__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_79__state == 2'b01) begin
        if(PE_wrapper_79__ap_ready) begin
          if(PE_wrapper_79__ap_done) begin
            PE_wrapper_79__state <= 2'b10;
          end else begin
            PE_wrapper_79__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_79__state == 2'b11) begin
        if(PE_wrapper_79__ap_done) begin
          PE_wrapper_79__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_79__state == 2'b10) begin
        if(PE_wrapper_79__ap_done_global__q0) begin
          PE_wrapper_79__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_79__ap_start = (PE_wrapper_79__state == 2'b01);
  assign PE_wrapper_80__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_80__is_done__q0 = (PE_wrapper_80__state == 2'b10);
  assign PE_wrapper_80__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_80__state <= 2'b00;
    end else begin
      if(PE_wrapper_80__state == 2'b00) begin
        if(PE_wrapper_80__ap_start_global__q0) begin
          PE_wrapper_80__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_80__state == 2'b01) begin
        if(PE_wrapper_80__ap_ready) begin
          if(PE_wrapper_80__ap_done) begin
            PE_wrapper_80__state <= 2'b10;
          end else begin
            PE_wrapper_80__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_80__state == 2'b11) begin
        if(PE_wrapper_80__ap_done) begin
          PE_wrapper_80__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_80__state == 2'b10) begin
        if(PE_wrapper_80__ap_done_global__q0) begin
          PE_wrapper_80__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_80__ap_start = (PE_wrapper_80__state == 2'b01);
  assign PE_wrapper_81__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_81__is_done__q0 = (PE_wrapper_81__state == 2'b10);
  assign PE_wrapper_81__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_81__state <= 2'b00;
    end else begin
      if(PE_wrapper_81__state == 2'b00) begin
        if(PE_wrapper_81__ap_start_global__q0) begin
          PE_wrapper_81__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_81__state == 2'b01) begin
        if(PE_wrapper_81__ap_ready) begin
          if(PE_wrapper_81__ap_done) begin
            PE_wrapper_81__state <= 2'b10;
          end else begin
            PE_wrapper_81__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_81__state == 2'b11) begin
        if(PE_wrapper_81__ap_done) begin
          PE_wrapper_81__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_81__state == 2'b10) begin
        if(PE_wrapper_81__ap_done_global__q0) begin
          PE_wrapper_81__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_81__ap_start = (PE_wrapper_81__state == 2'b01);
  assign PE_wrapper_82__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_82__is_done__q0 = (PE_wrapper_82__state == 2'b10);
  assign PE_wrapper_82__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_82__state <= 2'b00;
    end else begin
      if(PE_wrapper_82__state == 2'b00) begin
        if(PE_wrapper_82__ap_start_global__q0) begin
          PE_wrapper_82__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_82__state == 2'b01) begin
        if(PE_wrapper_82__ap_ready) begin
          if(PE_wrapper_82__ap_done) begin
            PE_wrapper_82__state <= 2'b10;
          end else begin
            PE_wrapper_82__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_82__state == 2'b11) begin
        if(PE_wrapper_82__ap_done) begin
          PE_wrapper_82__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_82__state == 2'b10) begin
        if(PE_wrapper_82__ap_done_global__q0) begin
          PE_wrapper_82__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_82__ap_start = (PE_wrapper_82__state == 2'b01);
  assign PE_wrapper_83__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_83__is_done__q0 = (PE_wrapper_83__state == 2'b10);
  assign PE_wrapper_83__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_83__state <= 2'b00;
    end else begin
      if(PE_wrapper_83__state == 2'b00) begin
        if(PE_wrapper_83__ap_start_global__q0) begin
          PE_wrapper_83__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_83__state == 2'b01) begin
        if(PE_wrapper_83__ap_ready) begin
          if(PE_wrapper_83__ap_done) begin
            PE_wrapper_83__state <= 2'b10;
          end else begin
            PE_wrapper_83__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_83__state == 2'b11) begin
        if(PE_wrapper_83__ap_done) begin
          PE_wrapper_83__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_83__state == 2'b10) begin
        if(PE_wrapper_83__ap_done_global__q0) begin
          PE_wrapper_83__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_83__ap_start = (PE_wrapper_83__state == 2'b01);
  assign PE_wrapper_84__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_84__is_done__q0 = (PE_wrapper_84__state == 2'b10);
  assign PE_wrapper_84__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_84__state <= 2'b00;
    end else begin
      if(PE_wrapper_84__state == 2'b00) begin
        if(PE_wrapper_84__ap_start_global__q0) begin
          PE_wrapper_84__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_84__state == 2'b01) begin
        if(PE_wrapper_84__ap_ready) begin
          if(PE_wrapper_84__ap_done) begin
            PE_wrapper_84__state <= 2'b10;
          end else begin
            PE_wrapper_84__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_84__state == 2'b11) begin
        if(PE_wrapper_84__ap_done) begin
          PE_wrapper_84__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_84__state == 2'b10) begin
        if(PE_wrapper_84__ap_done_global__q0) begin
          PE_wrapper_84__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_84__ap_start = (PE_wrapper_84__state == 2'b01);
  assign PE_wrapper_85__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_85__is_done__q0 = (PE_wrapper_85__state == 2'b10);
  assign PE_wrapper_85__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_85__state <= 2'b00;
    end else begin
      if(PE_wrapper_85__state == 2'b00) begin
        if(PE_wrapper_85__ap_start_global__q0) begin
          PE_wrapper_85__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_85__state == 2'b01) begin
        if(PE_wrapper_85__ap_ready) begin
          if(PE_wrapper_85__ap_done) begin
            PE_wrapper_85__state <= 2'b10;
          end else begin
            PE_wrapper_85__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_85__state == 2'b11) begin
        if(PE_wrapper_85__ap_done) begin
          PE_wrapper_85__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_85__state == 2'b10) begin
        if(PE_wrapper_85__ap_done_global__q0) begin
          PE_wrapper_85__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_85__ap_start = (PE_wrapper_85__state == 2'b01);
  assign PE_wrapper_86__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_86__is_done__q0 = (PE_wrapper_86__state == 2'b10);
  assign PE_wrapper_86__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_86__state <= 2'b00;
    end else begin
      if(PE_wrapper_86__state == 2'b00) begin
        if(PE_wrapper_86__ap_start_global__q0) begin
          PE_wrapper_86__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_86__state == 2'b01) begin
        if(PE_wrapper_86__ap_ready) begin
          if(PE_wrapper_86__ap_done) begin
            PE_wrapper_86__state <= 2'b10;
          end else begin
            PE_wrapper_86__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_86__state == 2'b11) begin
        if(PE_wrapper_86__ap_done) begin
          PE_wrapper_86__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_86__state == 2'b10) begin
        if(PE_wrapper_86__ap_done_global__q0) begin
          PE_wrapper_86__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_86__ap_start = (PE_wrapper_86__state == 2'b01);
  assign PE_wrapper_87__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_87__is_done__q0 = (PE_wrapper_87__state == 2'b10);
  assign PE_wrapper_87__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_87__state <= 2'b00;
    end else begin
      if(PE_wrapper_87__state == 2'b00) begin
        if(PE_wrapper_87__ap_start_global__q0) begin
          PE_wrapper_87__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_87__state == 2'b01) begin
        if(PE_wrapper_87__ap_ready) begin
          if(PE_wrapper_87__ap_done) begin
            PE_wrapper_87__state <= 2'b10;
          end else begin
            PE_wrapper_87__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_87__state == 2'b11) begin
        if(PE_wrapper_87__ap_done) begin
          PE_wrapper_87__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_87__state == 2'b10) begin
        if(PE_wrapper_87__ap_done_global__q0) begin
          PE_wrapper_87__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_87__ap_start = (PE_wrapper_87__state == 2'b01);
  assign PE_wrapper_88__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_88__is_done__q0 = (PE_wrapper_88__state == 2'b10);
  assign PE_wrapper_88__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_88__state <= 2'b00;
    end else begin
      if(PE_wrapper_88__state == 2'b00) begin
        if(PE_wrapper_88__ap_start_global__q0) begin
          PE_wrapper_88__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_88__state == 2'b01) begin
        if(PE_wrapper_88__ap_ready) begin
          if(PE_wrapper_88__ap_done) begin
            PE_wrapper_88__state <= 2'b10;
          end else begin
            PE_wrapper_88__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_88__state == 2'b11) begin
        if(PE_wrapper_88__ap_done) begin
          PE_wrapper_88__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_88__state == 2'b10) begin
        if(PE_wrapper_88__ap_done_global__q0) begin
          PE_wrapper_88__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_88__ap_start = (PE_wrapper_88__state == 2'b01);
  assign PE_wrapper_89__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_89__is_done__q0 = (PE_wrapper_89__state == 2'b10);
  assign PE_wrapper_89__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_89__state <= 2'b00;
    end else begin
      if(PE_wrapper_89__state == 2'b00) begin
        if(PE_wrapper_89__ap_start_global__q0) begin
          PE_wrapper_89__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_89__state == 2'b01) begin
        if(PE_wrapper_89__ap_ready) begin
          if(PE_wrapper_89__ap_done) begin
            PE_wrapper_89__state <= 2'b10;
          end else begin
            PE_wrapper_89__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_89__state == 2'b11) begin
        if(PE_wrapper_89__ap_done) begin
          PE_wrapper_89__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_89__state == 2'b10) begin
        if(PE_wrapper_89__ap_done_global__q0) begin
          PE_wrapper_89__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_89__ap_start = (PE_wrapper_89__state == 2'b01);
  assign PE_wrapper_90__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_90__is_done__q0 = (PE_wrapper_90__state == 2'b10);
  assign PE_wrapper_90__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_90__state <= 2'b00;
    end else begin
      if(PE_wrapper_90__state == 2'b00) begin
        if(PE_wrapper_90__ap_start_global__q0) begin
          PE_wrapper_90__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_90__state == 2'b01) begin
        if(PE_wrapper_90__ap_ready) begin
          if(PE_wrapper_90__ap_done) begin
            PE_wrapper_90__state <= 2'b10;
          end else begin
            PE_wrapper_90__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_90__state == 2'b11) begin
        if(PE_wrapper_90__ap_done) begin
          PE_wrapper_90__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_90__state == 2'b10) begin
        if(PE_wrapper_90__ap_done_global__q0) begin
          PE_wrapper_90__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_90__ap_start = (PE_wrapper_90__state == 2'b01);
  assign PE_wrapper_91__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_91__is_done__q0 = (PE_wrapper_91__state == 2'b10);
  assign PE_wrapper_91__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_91__state <= 2'b00;
    end else begin
      if(PE_wrapper_91__state == 2'b00) begin
        if(PE_wrapper_91__ap_start_global__q0) begin
          PE_wrapper_91__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_91__state == 2'b01) begin
        if(PE_wrapper_91__ap_ready) begin
          if(PE_wrapper_91__ap_done) begin
            PE_wrapper_91__state <= 2'b10;
          end else begin
            PE_wrapper_91__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_91__state == 2'b11) begin
        if(PE_wrapper_91__ap_done) begin
          PE_wrapper_91__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_91__state == 2'b10) begin
        if(PE_wrapper_91__ap_done_global__q0) begin
          PE_wrapper_91__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_91__ap_start = (PE_wrapper_91__state == 2'b01);
  assign PE_wrapper_92__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_92__is_done__q0 = (PE_wrapper_92__state == 2'b10);
  assign PE_wrapper_92__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_92__state <= 2'b00;
    end else begin
      if(PE_wrapper_92__state == 2'b00) begin
        if(PE_wrapper_92__ap_start_global__q0) begin
          PE_wrapper_92__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_92__state == 2'b01) begin
        if(PE_wrapper_92__ap_ready) begin
          if(PE_wrapper_92__ap_done) begin
            PE_wrapper_92__state <= 2'b10;
          end else begin
            PE_wrapper_92__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_92__state == 2'b11) begin
        if(PE_wrapper_92__ap_done) begin
          PE_wrapper_92__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_92__state == 2'b10) begin
        if(PE_wrapper_92__ap_done_global__q0) begin
          PE_wrapper_92__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_92__ap_start = (PE_wrapper_92__state == 2'b01);
  assign PE_wrapper_93__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_93__is_done__q0 = (PE_wrapper_93__state == 2'b10);
  assign PE_wrapper_93__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_93__state <= 2'b00;
    end else begin
      if(PE_wrapper_93__state == 2'b00) begin
        if(PE_wrapper_93__ap_start_global__q0) begin
          PE_wrapper_93__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_93__state == 2'b01) begin
        if(PE_wrapper_93__ap_ready) begin
          if(PE_wrapper_93__ap_done) begin
            PE_wrapper_93__state <= 2'b10;
          end else begin
            PE_wrapper_93__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_93__state == 2'b11) begin
        if(PE_wrapper_93__ap_done) begin
          PE_wrapper_93__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_93__state == 2'b10) begin
        if(PE_wrapper_93__ap_done_global__q0) begin
          PE_wrapper_93__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_93__ap_start = (PE_wrapper_93__state == 2'b01);
  assign PE_wrapper_94__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_94__is_done__q0 = (PE_wrapper_94__state == 2'b10);
  assign PE_wrapper_94__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_94__state <= 2'b00;
    end else begin
      if(PE_wrapper_94__state == 2'b00) begin
        if(PE_wrapper_94__ap_start_global__q0) begin
          PE_wrapper_94__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_94__state == 2'b01) begin
        if(PE_wrapper_94__ap_ready) begin
          if(PE_wrapper_94__ap_done) begin
            PE_wrapper_94__state <= 2'b10;
          end else begin
            PE_wrapper_94__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_94__state == 2'b11) begin
        if(PE_wrapper_94__ap_done) begin
          PE_wrapper_94__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_94__state == 2'b10) begin
        if(PE_wrapper_94__ap_done_global__q0) begin
          PE_wrapper_94__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_94__ap_start = (PE_wrapper_94__state == 2'b01);
  assign PE_wrapper_95__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_95__is_done__q0 = (PE_wrapper_95__state == 2'b10);
  assign PE_wrapper_95__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_95__state <= 2'b00;
    end else begin
      if(PE_wrapper_95__state == 2'b00) begin
        if(PE_wrapper_95__ap_start_global__q0) begin
          PE_wrapper_95__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_95__state == 2'b01) begin
        if(PE_wrapper_95__ap_ready) begin
          if(PE_wrapper_95__ap_done) begin
            PE_wrapper_95__state <= 2'b10;
          end else begin
            PE_wrapper_95__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_95__state == 2'b11) begin
        if(PE_wrapper_95__ap_done) begin
          PE_wrapper_95__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_95__state == 2'b10) begin
        if(PE_wrapper_95__ap_done_global__q0) begin
          PE_wrapper_95__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_95__ap_start = (PE_wrapper_95__state == 2'b01);
  assign PE_wrapper_96__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_96__is_done__q0 = (PE_wrapper_96__state == 2'b10);
  assign PE_wrapper_96__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_96__state <= 2'b00;
    end else begin
      if(PE_wrapper_96__state == 2'b00) begin
        if(PE_wrapper_96__ap_start_global__q0) begin
          PE_wrapper_96__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_96__state == 2'b01) begin
        if(PE_wrapper_96__ap_ready) begin
          if(PE_wrapper_96__ap_done) begin
            PE_wrapper_96__state <= 2'b10;
          end else begin
            PE_wrapper_96__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_96__state == 2'b11) begin
        if(PE_wrapper_96__ap_done) begin
          PE_wrapper_96__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_96__state == 2'b10) begin
        if(PE_wrapper_96__ap_done_global__q0) begin
          PE_wrapper_96__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_96__ap_start = (PE_wrapper_96__state == 2'b01);
  assign PE_wrapper_97__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_97__is_done__q0 = (PE_wrapper_97__state == 2'b10);
  assign PE_wrapper_97__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_97__state <= 2'b00;
    end else begin
      if(PE_wrapper_97__state == 2'b00) begin
        if(PE_wrapper_97__ap_start_global__q0) begin
          PE_wrapper_97__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_97__state == 2'b01) begin
        if(PE_wrapper_97__ap_ready) begin
          if(PE_wrapper_97__ap_done) begin
            PE_wrapper_97__state <= 2'b10;
          end else begin
            PE_wrapper_97__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_97__state == 2'b11) begin
        if(PE_wrapper_97__ap_done) begin
          PE_wrapper_97__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_97__state == 2'b10) begin
        if(PE_wrapper_97__ap_done_global__q0) begin
          PE_wrapper_97__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_97__ap_start = (PE_wrapper_97__state == 2'b01);
  assign PE_wrapper_98__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_98__is_done__q0 = (PE_wrapper_98__state == 2'b10);
  assign PE_wrapper_98__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_98__state <= 2'b00;
    end else begin
      if(PE_wrapper_98__state == 2'b00) begin
        if(PE_wrapper_98__ap_start_global__q0) begin
          PE_wrapper_98__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_98__state == 2'b01) begin
        if(PE_wrapper_98__ap_ready) begin
          if(PE_wrapper_98__ap_done) begin
            PE_wrapper_98__state <= 2'b10;
          end else begin
            PE_wrapper_98__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_98__state == 2'b11) begin
        if(PE_wrapper_98__ap_done) begin
          PE_wrapper_98__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_98__state == 2'b10) begin
        if(PE_wrapper_98__ap_done_global__q0) begin
          PE_wrapper_98__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_98__ap_start = (PE_wrapper_98__state == 2'b01);
  assign PE_wrapper_99__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_99__is_done__q0 = (PE_wrapper_99__state == 2'b10);
  assign PE_wrapper_99__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_99__state <= 2'b00;
    end else begin
      if(PE_wrapper_99__state == 2'b00) begin
        if(PE_wrapper_99__ap_start_global__q0) begin
          PE_wrapper_99__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_99__state == 2'b01) begin
        if(PE_wrapper_99__ap_ready) begin
          if(PE_wrapper_99__ap_done) begin
            PE_wrapper_99__state <= 2'b10;
          end else begin
            PE_wrapper_99__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_99__state == 2'b11) begin
        if(PE_wrapper_99__ap_done) begin
          PE_wrapper_99__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_99__state == 2'b10) begin
        if(PE_wrapper_99__ap_done_global__q0) begin
          PE_wrapper_99__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_99__ap_start = (PE_wrapper_99__state == 2'b01);
  assign PE_wrapper_100__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_100__is_done__q0 = (PE_wrapper_100__state == 2'b10);
  assign PE_wrapper_100__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_100__state <= 2'b00;
    end else begin
      if(PE_wrapper_100__state == 2'b00) begin
        if(PE_wrapper_100__ap_start_global__q0) begin
          PE_wrapper_100__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_100__state == 2'b01) begin
        if(PE_wrapper_100__ap_ready) begin
          if(PE_wrapper_100__ap_done) begin
            PE_wrapper_100__state <= 2'b10;
          end else begin
            PE_wrapper_100__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_100__state == 2'b11) begin
        if(PE_wrapper_100__ap_done) begin
          PE_wrapper_100__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_100__state == 2'b10) begin
        if(PE_wrapper_100__ap_done_global__q0) begin
          PE_wrapper_100__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_100__ap_start = (PE_wrapper_100__state == 2'b01);
  assign PE_wrapper_101__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_101__is_done__q0 = (PE_wrapper_101__state == 2'b10);
  assign PE_wrapper_101__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_101__state <= 2'b00;
    end else begin
      if(PE_wrapper_101__state == 2'b00) begin
        if(PE_wrapper_101__ap_start_global__q0) begin
          PE_wrapper_101__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_101__state == 2'b01) begin
        if(PE_wrapper_101__ap_ready) begin
          if(PE_wrapper_101__ap_done) begin
            PE_wrapper_101__state <= 2'b10;
          end else begin
            PE_wrapper_101__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_101__state == 2'b11) begin
        if(PE_wrapper_101__ap_done) begin
          PE_wrapper_101__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_101__state == 2'b10) begin
        if(PE_wrapper_101__ap_done_global__q0) begin
          PE_wrapper_101__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_101__ap_start = (PE_wrapper_101__state == 2'b01);
  assign PE_wrapper_102__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_102__is_done__q0 = (PE_wrapper_102__state == 2'b10);
  assign PE_wrapper_102__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_102__state <= 2'b00;
    end else begin
      if(PE_wrapper_102__state == 2'b00) begin
        if(PE_wrapper_102__ap_start_global__q0) begin
          PE_wrapper_102__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_102__state == 2'b01) begin
        if(PE_wrapper_102__ap_ready) begin
          if(PE_wrapper_102__ap_done) begin
            PE_wrapper_102__state <= 2'b10;
          end else begin
            PE_wrapper_102__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_102__state == 2'b11) begin
        if(PE_wrapper_102__ap_done) begin
          PE_wrapper_102__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_102__state == 2'b10) begin
        if(PE_wrapper_102__ap_done_global__q0) begin
          PE_wrapper_102__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_102__ap_start = (PE_wrapper_102__state == 2'b01);
  assign PE_wrapper_103__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_103__is_done__q0 = (PE_wrapper_103__state == 2'b10);
  assign PE_wrapper_103__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_103__state <= 2'b00;
    end else begin
      if(PE_wrapper_103__state == 2'b00) begin
        if(PE_wrapper_103__ap_start_global__q0) begin
          PE_wrapper_103__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_103__state == 2'b01) begin
        if(PE_wrapper_103__ap_ready) begin
          if(PE_wrapper_103__ap_done) begin
            PE_wrapper_103__state <= 2'b10;
          end else begin
            PE_wrapper_103__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_103__state == 2'b11) begin
        if(PE_wrapper_103__ap_done) begin
          PE_wrapper_103__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_103__state == 2'b10) begin
        if(PE_wrapper_103__ap_done_global__q0) begin
          PE_wrapper_103__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_103__ap_start = (PE_wrapper_103__state == 2'b01);
  assign PE_wrapper_104__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_104__is_done__q0 = (PE_wrapper_104__state == 2'b10);
  assign PE_wrapper_104__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_104__state <= 2'b00;
    end else begin
      if(PE_wrapper_104__state == 2'b00) begin
        if(PE_wrapper_104__ap_start_global__q0) begin
          PE_wrapper_104__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_104__state == 2'b01) begin
        if(PE_wrapper_104__ap_ready) begin
          if(PE_wrapper_104__ap_done) begin
            PE_wrapper_104__state <= 2'b10;
          end else begin
            PE_wrapper_104__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_104__state == 2'b11) begin
        if(PE_wrapper_104__ap_done) begin
          PE_wrapper_104__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_104__state == 2'b10) begin
        if(PE_wrapper_104__ap_done_global__q0) begin
          PE_wrapper_104__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_104__ap_start = (PE_wrapper_104__state == 2'b01);
  assign PE_wrapper_105__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_105__is_done__q0 = (PE_wrapper_105__state == 2'b10);
  assign PE_wrapper_105__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_105__state <= 2'b00;
    end else begin
      if(PE_wrapper_105__state == 2'b00) begin
        if(PE_wrapper_105__ap_start_global__q0) begin
          PE_wrapper_105__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_105__state == 2'b01) begin
        if(PE_wrapper_105__ap_ready) begin
          if(PE_wrapper_105__ap_done) begin
            PE_wrapper_105__state <= 2'b10;
          end else begin
            PE_wrapper_105__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_105__state == 2'b11) begin
        if(PE_wrapper_105__ap_done) begin
          PE_wrapper_105__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_105__state == 2'b10) begin
        if(PE_wrapper_105__ap_done_global__q0) begin
          PE_wrapper_105__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_105__ap_start = (PE_wrapper_105__state == 2'b01);
  assign PE_wrapper_106__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_106__is_done__q0 = (PE_wrapper_106__state == 2'b10);
  assign PE_wrapper_106__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_106__state <= 2'b00;
    end else begin
      if(PE_wrapper_106__state == 2'b00) begin
        if(PE_wrapper_106__ap_start_global__q0) begin
          PE_wrapper_106__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_106__state == 2'b01) begin
        if(PE_wrapper_106__ap_ready) begin
          if(PE_wrapper_106__ap_done) begin
            PE_wrapper_106__state <= 2'b10;
          end else begin
            PE_wrapper_106__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_106__state == 2'b11) begin
        if(PE_wrapper_106__ap_done) begin
          PE_wrapper_106__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_106__state == 2'b10) begin
        if(PE_wrapper_106__ap_done_global__q0) begin
          PE_wrapper_106__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_106__ap_start = (PE_wrapper_106__state == 2'b01);
  assign PE_wrapper_107__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_107__is_done__q0 = (PE_wrapper_107__state == 2'b10);
  assign PE_wrapper_107__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_107__state <= 2'b00;
    end else begin
      if(PE_wrapper_107__state == 2'b00) begin
        if(PE_wrapper_107__ap_start_global__q0) begin
          PE_wrapper_107__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_107__state == 2'b01) begin
        if(PE_wrapper_107__ap_ready) begin
          if(PE_wrapper_107__ap_done) begin
            PE_wrapper_107__state <= 2'b10;
          end else begin
            PE_wrapper_107__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_107__state == 2'b11) begin
        if(PE_wrapper_107__ap_done) begin
          PE_wrapper_107__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_107__state == 2'b10) begin
        if(PE_wrapper_107__ap_done_global__q0) begin
          PE_wrapper_107__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_107__ap_start = (PE_wrapper_107__state == 2'b01);
  assign PE_wrapper_108__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_108__is_done__q0 = (PE_wrapper_108__state == 2'b10);
  assign PE_wrapper_108__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_108__state <= 2'b00;
    end else begin
      if(PE_wrapper_108__state == 2'b00) begin
        if(PE_wrapper_108__ap_start_global__q0) begin
          PE_wrapper_108__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_108__state == 2'b01) begin
        if(PE_wrapper_108__ap_ready) begin
          if(PE_wrapper_108__ap_done) begin
            PE_wrapper_108__state <= 2'b10;
          end else begin
            PE_wrapper_108__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_108__state == 2'b11) begin
        if(PE_wrapper_108__ap_done) begin
          PE_wrapper_108__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_108__state == 2'b10) begin
        if(PE_wrapper_108__ap_done_global__q0) begin
          PE_wrapper_108__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_108__ap_start = (PE_wrapper_108__state == 2'b01);
  assign PE_wrapper_109__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_109__is_done__q0 = (PE_wrapper_109__state == 2'b10);
  assign PE_wrapper_109__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_109__state <= 2'b00;
    end else begin
      if(PE_wrapper_109__state == 2'b00) begin
        if(PE_wrapper_109__ap_start_global__q0) begin
          PE_wrapper_109__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_109__state == 2'b01) begin
        if(PE_wrapper_109__ap_ready) begin
          if(PE_wrapper_109__ap_done) begin
            PE_wrapper_109__state <= 2'b10;
          end else begin
            PE_wrapper_109__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_109__state == 2'b11) begin
        if(PE_wrapper_109__ap_done) begin
          PE_wrapper_109__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_109__state == 2'b10) begin
        if(PE_wrapper_109__ap_done_global__q0) begin
          PE_wrapper_109__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_109__ap_start = (PE_wrapper_109__state == 2'b01);
  assign PE_wrapper_110__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_110__is_done__q0 = (PE_wrapper_110__state == 2'b10);
  assign PE_wrapper_110__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_110__state <= 2'b00;
    end else begin
      if(PE_wrapper_110__state == 2'b00) begin
        if(PE_wrapper_110__ap_start_global__q0) begin
          PE_wrapper_110__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_110__state == 2'b01) begin
        if(PE_wrapper_110__ap_ready) begin
          if(PE_wrapper_110__ap_done) begin
            PE_wrapper_110__state <= 2'b10;
          end else begin
            PE_wrapper_110__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_110__state == 2'b11) begin
        if(PE_wrapper_110__ap_done) begin
          PE_wrapper_110__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_110__state == 2'b10) begin
        if(PE_wrapper_110__ap_done_global__q0) begin
          PE_wrapper_110__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_110__ap_start = (PE_wrapper_110__state == 2'b01);
  assign PE_wrapper_111__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_111__is_done__q0 = (PE_wrapper_111__state == 2'b10);
  assign PE_wrapper_111__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_111__state <= 2'b00;
    end else begin
      if(PE_wrapper_111__state == 2'b00) begin
        if(PE_wrapper_111__ap_start_global__q0) begin
          PE_wrapper_111__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_111__state == 2'b01) begin
        if(PE_wrapper_111__ap_ready) begin
          if(PE_wrapper_111__ap_done) begin
            PE_wrapper_111__state <= 2'b10;
          end else begin
            PE_wrapper_111__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_111__state == 2'b11) begin
        if(PE_wrapper_111__ap_done) begin
          PE_wrapper_111__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_111__state == 2'b10) begin
        if(PE_wrapper_111__ap_done_global__q0) begin
          PE_wrapper_111__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_111__ap_start = (PE_wrapper_111__state == 2'b01);
  assign PE_wrapper_112__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_112__is_done__q0 = (PE_wrapper_112__state == 2'b10);
  assign PE_wrapper_112__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_112__state <= 2'b00;
    end else begin
      if(PE_wrapper_112__state == 2'b00) begin
        if(PE_wrapper_112__ap_start_global__q0) begin
          PE_wrapper_112__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_112__state == 2'b01) begin
        if(PE_wrapper_112__ap_ready) begin
          if(PE_wrapper_112__ap_done) begin
            PE_wrapper_112__state <= 2'b10;
          end else begin
            PE_wrapper_112__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_112__state == 2'b11) begin
        if(PE_wrapper_112__ap_done) begin
          PE_wrapper_112__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_112__state == 2'b10) begin
        if(PE_wrapper_112__ap_done_global__q0) begin
          PE_wrapper_112__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_112__ap_start = (PE_wrapper_112__state == 2'b01);
  assign PE_wrapper_113__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_113__is_done__q0 = (PE_wrapper_113__state == 2'b10);
  assign PE_wrapper_113__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_113__state <= 2'b00;
    end else begin
      if(PE_wrapper_113__state == 2'b00) begin
        if(PE_wrapper_113__ap_start_global__q0) begin
          PE_wrapper_113__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_113__state == 2'b01) begin
        if(PE_wrapper_113__ap_ready) begin
          if(PE_wrapper_113__ap_done) begin
            PE_wrapper_113__state <= 2'b10;
          end else begin
            PE_wrapper_113__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_113__state == 2'b11) begin
        if(PE_wrapper_113__ap_done) begin
          PE_wrapper_113__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_113__state == 2'b10) begin
        if(PE_wrapper_113__ap_done_global__q0) begin
          PE_wrapper_113__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_113__ap_start = (PE_wrapper_113__state == 2'b01);
  assign PE_wrapper_114__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_114__is_done__q0 = (PE_wrapper_114__state == 2'b10);
  assign PE_wrapper_114__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_114__state <= 2'b00;
    end else begin
      if(PE_wrapper_114__state == 2'b00) begin
        if(PE_wrapper_114__ap_start_global__q0) begin
          PE_wrapper_114__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_114__state == 2'b01) begin
        if(PE_wrapper_114__ap_ready) begin
          if(PE_wrapper_114__ap_done) begin
            PE_wrapper_114__state <= 2'b10;
          end else begin
            PE_wrapper_114__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_114__state == 2'b11) begin
        if(PE_wrapper_114__ap_done) begin
          PE_wrapper_114__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_114__state == 2'b10) begin
        if(PE_wrapper_114__ap_done_global__q0) begin
          PE_wrapper_114__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_114__ap_start = (PE_wrapper_114__state == 2'b01);
  assign PE_wrapper_115__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_115__is_done__q0 = (PE_wrapper_115__state == 2'b10);
  assign PE_wrapper_115__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_115__state <= 2'b00;
    end else begin
      if(PE_wrapper_115__state == 2'b00) begin
        if(PE_wrapper_115__ap_start_global__q0) begin
          PE_wrapper_115__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_115__state == 2'b01) begin
        if(PE_wrapper_115__ap_ready) begin
          if(PE_wrapper_115__ap_done) begin
            PE_wrapper_115__state <= 2'b10;
          end else begin
            PE_wrapper_115__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_115__state == 2'b11) begin
        if(PE_wrapper_115__ap_done) begin
          PE_wrapper_115__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_115__state == 2'b10) begin
        if(PE_wrapper_115__ap_done_global__q0) begin
          PE_wrapper_115__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_115__ap_start = (PE_wrapper_115__state == 2'b01);
  assign PE_wrapper_116__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_116__is_done__q0 = (PE_wrapper_116__state == 2'b10);
  assign PE_wrapper_116__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_116__state <= 2'b00;
    end else begin
      if(PE_wrapper_116__state == 2'b00) begin
        if(PE_wrapper_116__ap_start_global__q0) begin
          PE_wrapper_116__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_116__state == 2'b01) begin
        if(PE_wrapper_116__ap_ready) begin
          if(PE_wrapper_116__ap_done) begin
            PE_wrapper_116__state <= 2'b10;
          end else begin
            PE_wrapper_116__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_116__state == 2'b11) begin
        if(PE_wrapper_116__ap_done) begin
          PE_wrapper_116__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_116__state == 2'b10) begin
        if(PE_wrapper_116__ap_done_global__q0) begin
          PE_wrapper_116__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_116__ap_start = (PE_wrapper_116__state == 2'b01);
  assign PE_wrapper_117__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_117__is_done__q0 = (PE_wrapper_117__state == 2'b10);
  assign PE_wrapper_117__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_117__state <= 2'b00;
    end else begin
      if(PE_wrapper_117__state == 2'b00) begin
        if(PE_wrapper_117__ap_start_global__q0) begin
          PE_wrapper_117__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_117__state == 2'b01) begin
        if(PE_wrapper_117__ap_ready) begin
          if(PE_wrapper_117__ap_done) begin
            PE_wrapper_117__state <= 2'b10;
          end else begin
            PE_wrapper_117__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_117__state == 2'b11) begin
        if(PE_wrapper_117__ap_done) begin
          PE_wrapper_117__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_117__state == 2'b10) begin
        if(PE_wrapper_117__ap_done_global__q0) begin
          PE_wrapper_117__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_117__ap_start = (PE_wrapper_117__state == 2'b01);
  assign PE_wrapper_118__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_118__is_done__q0 = (PE_wrapper_118__state == 2'b10);
  assign PE_wrapper_118__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_118__state <= 2'b00;
    end else begin
      if(PE_wrapper_118__state == 2'b00) begin
        if(PE_wrapper_118__ap_start_global__q0) begin
          PE_wrapper_118__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_118__state == 2'b01) begin
        if(PE_wrapper_118__ap_ready) begin
          if(PE_wrapper_118__ap_done) begin
            PE_wrapper_118__state <= 2'b10;
          end else begin
            PE_wrapper_118__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_118__state == 2'b11) begin
        if(PE_wrapper_118__ap_done) begin
          PE_wrapper_118__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_118__state == 2'b10) begin
        if(PE_wrapper_118__ap_done_global__q0) begin
          PE_wrapper_118__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_118__ap_start = (PE_wrapper_118__state == 2'b01);
  assign PE_wrapper_119__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_119__is_done__q0 = (PE_wrapper_119__state == 2'b10);
  assign PE_wrapper_119__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_119__state <= 2'b00;
    end else begin
      if(PE_wrapper_119__state == 2'b00) begin
        if(PE_wrapper_119__ap_start_global__q0) begin
          PE_wrapper_119__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_119__state == 2'b01) begin
        if(PE_wrapper_119__ap_ready) begin
          if(PE_wrapper_119__ap_done) begin
            PE_wrapper_119__state <= 2'b10;
          end else begin
            PE_wrapper_119__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_119__state == 2'b11) begin
        if(PE_wrapper_119__ap_done) begin
          PE_wrapper_119__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_119__state == 2'b10) begin
        if(PE_wrapper_119__ap_done_global__q0) begin
          PE_wrapper_119__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_119__ap_start = (PE_wrapper_119__state == 2'b01);
  assign PE_wrapper_120__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_120__is_done__q0 = (PE_wrapper_120__state == 2'b10);
  assign PE_wrapper_120__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_120__state <= 2'b00;
    end else begin
      if(PE_wrapper_120__state == 2'b00) begin
        if(PE_wrapper_120__ap_start_global__q0) begin
          PE_wrapper_120__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_120__state == 2'b01) begin
        if(PE_wrapper_120__ap_ready) begin
          if(PE_wrapper_120__ap_done) begin
            PE_wrapper_120__state <= 2'b10;
          end else begin
            PE_wrapper_120__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_120__state == 2'b11) begin
        if(PE_wrapper_120__ap_done) begin
          PE_wrapper_120__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_120__state == 2'b10) begin
        if(PE_wrapper_120__ap_done_global__q0) begin
          PE_wrapper_120__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_120__ap_start = (PE_wrapper_120__state == 2'b01);
  assign PE_wrapper_121__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_121__is_done__q0 = (PE_wrapper_121__state == 2'b10);
  assign PE_wrapper_121__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_121__state <= 2'b00;
    end else begin
      if(PE_wrapper_121__state == 2'b00) begin
        if(PE_wrapper_121__ap_start_global__q0) begin
          PE_wrapper_121__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_121__state == 2'b01) begin
        if(PE_wrapper_121__ap_ready) begin
          if(PE_wrapper_121__ap_done) begin
            PE_wrapper_121__state <= 2'b10;
          end else begin
            PE_wrapper_121__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_121__state == 2'b11) begin
        if(PE_wrapper_121__ap_done) begin
          PE_wrapper_121__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_121__state == 2'b10) begin
        if(PE_wrapper_121__ap_done_global__q0) begin
          PE_wrapper_121__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_121__ap_start = (PE_wrapper_121__state == 2'b01);
  assign PE_wrapper_122__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_122__is_done__q0 = (PE_wrapper_122__state == 2'b10);
  assign PE_wrapper_122__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_122__state <= 2'b00;
    end else begin
      if(PE_wrapper_122__state == 2'b00) begin
        if(PE_wrapper_122__ap_start_global__q0) begin
          PE_wrapper_122__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_122__state == 2'b01) begin
        if(PE_wrapper_122__ap_ready) begin
          if(PE_wrapper_122__ap_done) begin
            PE_wrapper_122__state <= 2'b10;
          end else begin
            PE_wrapper_122__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_122__state == 2'b11) begin
        if(PE_wrapper_122__ap_done) begin
          PE_wrapper_122__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_122__state == 2'b10) begin
        if(PE_wrapper_122__ap_done_global__q0) begin
          PE_wrapper_122__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_122__ap_start = (PE_wrapper_122__state == 2'b01);
  assign PE_wrapper_123__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_123__is_done__q0 = (PE_wrapper_123__state == 2'b10);
  assign PE_wrapper_123__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_123__state <= 2'b00;
    end else begin
      if(PE_wrapper_123__state == 2'b00) begin
        if(PE_wrapper_123__ap_start_global__q0) begin
          PE_wrapper_123__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_123__state == 2'b01) begin
        if(PE_wrapper_123__ap_ready) begin
          if(PE_wrapper_123__ap_done) begin
            PE_wrapper_123__state <= 2'b10;
          end else begin
            PE_wrapper_123__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_123__state == 2'b11) begin
        if(PE_wrapper_123__ap_done) begin
          PE_wrapper_123__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_123__state == 2'b10) begin
        if(PE_wrapper_123__ap_done_global__q0) begin
          PE_wrapper_123__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_123__ap_start = (PE_wrapper_123__state == 2'b01);
  assign PE_wrapper_124__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_124__is_done__q0 = (PE_wrapper_124__state == 2'b10);
  assign PE_wrapper_124__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_124__state <= 2'b00;
    end else begin
      if(PE_wrapper_124__state == 2'b00) begin
        if(PE_wrapper_124__ap_start_global__q0) begin
          PE_wrapper_124__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_124__state == 2'b01) begin
        if(PE_wrapper_124__ap_ready) begin
          if(PE_wrapper_124__ap_done) begin
            PE_wrapper_124__state <= 2'b10;
          end else begin
            PE_wrapper_124__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_124__state == 2'b11) begin
        if(PE_wrapper_124__ap_done) begin
          PE_wrapper_124__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_124__state == 2'b10) begin
        if(PE_wrapper_124__ap_done_global__q0) begin
          PE_wrapper_124__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_124__ap_start = (PE_wrapper_124__state == 2'b01);
  assign PE_wrapper_125__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_125__is_done__q0 = (PE_wrapper_125__state == 2'b10);
  assign PE_wrapper_125__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_125__state <= 2'b00;
    end else begin
      if(PE_wrapper_125__state == 2'b00) begin
        if(PE_wrapper_125__ap_start_global__q0) begin
          PE_wrapper_125__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_125__state == 2'b01) begin
        if(PE_wrapper_125__ap_ready) begin
          if(PE_wrapper_125__ap_done) begin
            PE_wrapper_125__state <= 2'b10;
          end else begin
            PE_wrapper_125__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_125__state == 2'b11) begin
        if(PE_wrapper_125__ap_done) begin
          PE_wrapper_125__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_125__state == 2'b10) begin
        if(PE_wrapper_125__ap_done_global__q0) begin
          PE_wrapper_125__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_125__ap_start = (PE_wrapper_125__state == 2'b01);
  assign PE_wrapper_126__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_126__is_done__q0 = (PE_wrapper_126__state == 2'b10);
  assign PE_wrapper_126__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_126__state <= 2'b00;
    end else begin
      if(PE_wrapper_126__state == 2'b00) begin
        if(PE_wrapper_126__ap_start_global__q0) begin
          PE_wrapper_126__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_126__state == 2'b01) begin
        if(PE_wrapper_126__ap_ready) begin
          if(PE_wrapper_126__ap_done) begin
            PE_wrapper_126__state <= 2'b10;
          end else begin
            PE_wrapper_126__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_126__state == 2'b11) begin
        if(PE_wrapper_126__ap_done) begin
          PE_wrapper_126__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_126__state == 2'b10) begin
        if(PE_wrapper_126__ap_done_global__q0) begin
          PE_wrapper_126__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_126__ap_start = (PE_wrapper_126__state == 2'b01);
  assign PE_wrapper_127__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_127__is_done__q0 = (PE_wrapper_127__state == 2'b10);
  assign PE_wrapper_127__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_127__state <= 2'b00;
    end else begin
      if(PE_wrapper_127__state == 2'b00) begin
        if(PE_wrapper_127__ap_start_global__q0) begin
          PE_wrapper_127__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_127__state == 2'b01) begin
        if(PE_wrapper_127__ap_ready) begin
          if(PE_wrapper_127__ap_done) begin
            PE_wrapper_127__state <= 2'b10;
          end else begin
            PE_wrapper_127__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_127__state == 2'b11) begin
        if(PE_wrapper_127__ap_done) begin
          PE_wrapper_127__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_127__state == 2'b10) begin
        if(PE_wrapper_127__ap_done_global__q0) begin
          PE_wrapper_127__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_127__ap_start = (PE_wrapper_127__state == 2'b01);
  assign PE_wrapper_128__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_128__is_done__q0 = (PE_wrapper_128__state == 2'b10);
  assign PE_wrapper_128__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_128__state <= 2'b00;
    end else begin
      if(PE_wrapper_128__state == 2'b00) begin
        if(PE_wrapper_128__ap_start_global__q0) begin
          PE_wrapper_128__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_128__state == 2'b01) begin
        if(PE_wrapper_128__ap_ready) begin
          if(PE_wrapper_128__ap_done) begin
            PE_wrapper_128__state <= 2'b10;
          end else begin
            PE_wrapper_128__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_128__state == 2'b11) begin
        if(PE_wrapper_128__ap_done) begin
          PE_wrapper_128__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_128__state == 2'b10) begin
        if(PE_wrapper_128__ap_done_global__q0) begin
          PE_wrapper_128__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_128__ap_start = (PE_wrapper_128__state == 2'b01);
  assign PE_wrapper_129__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_129__is_done__q0 = (PE_wrapper_129__state == 2'b10);
  assign PE_wrapper_129__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_129__state <= 2'b00;
    end else begin
      if(PE_wrapper_129__state == 2'b00) begin
        if(PE_wrapper_129__ap_start_global__q0) begin
          PE_wrapper_129__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_129__state == 2'b01) begin
        if(PE_wrapper_129__ap_ready) begin
          if(PE_wrapper_129__ap_done) begin
            PE_wrapper_129__state <= 2'b10;
          end else begin
            PE_wrapper_129__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_129__state == 2'b11) begin
        if(PE_wrapper_129__ap_done) begin
          PE_wrapper_129__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_129__state == 2'b10) begin
        if(PE_wrapper_129__ap_done_global__q0) begin
          PE_wrapper_129__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_129__ap_start = (PE_wrapper_129__state == 2'b01);
  assign PE_wrapper_130__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_130__is_done__q0 = (PE_wrapper_130__state == 2'b10);
  assign PE_wrapper_130__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_130__state <= 2'b00;
    end else begin
      if(PE_wrapper_130__state == 2'b00) begin
        if(PE_wrapper_130__ap_start_global__q0) begin
          PE_wrapper_130__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_130__state == 2'b01) begin
        if(PE_wrapper_130__ap_ready) begin
          if(PE_wrapper_130__ap_done) begin
            PE_wrapper_130__state <= 2'b10;
          end else begin
            PE_wrapper_130__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_130__state == 2'b11) begin
        if(PE_wrapper_130__ap_done) begin
          PE_wrapper_130__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_130__state == 2'b10) begin
        if(PE_wrapper_130__ap_done_global__q0) begin
          PE_wrapper_130__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_130__ap_start = (PE_wrapper_130__state == 2'b01);
  assign PE_wrapper_131__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_131__is_done__q0 = (PE_wrapper_131__state == 2'b10);
  assign PE_wrapper_131__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_131__state <= 2'b00;
    end else begin
      if(PE_wrapper_131__state == 2'b00) begin
        if(PE_wrapper_131__ap_start_global__q0) begin
          PE_wrapper_131__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_131__state == 2'b01) begin
        if(PE_wrapper_131__ap_ready) begin
          if(PE_wrapper_131__ap_done) begin
            PE_wrapper_131__state <= 2'b10;
          end else begin
            PE_wrapper_131__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_131__state == 2'b11) begin
        if(PE_wrapper_131__ap_done) begin
          PE_wrapper_131__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_131__state == 2'b10) begin
        if(PE_wrapper_131__ap_done_global__q0) begin
          PE_wrapper_131__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_131__ap_start = (PE_wrapper_131__state == 2'b01);
  assign PE_wrapper_132__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_132__is_done__q0 = (PE_wrapper_132__state == 2'b10);
  assign PE_wrapper_132__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_132__state <= 2'b00;
    end else begin
      if(PE_wrapper_132__state == 2'b00) begin
        if(PE_wrapper_132__ap_start_global__q0) begin
          PE_wrapper_132__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_132__state == 2'b01) begin
        if(PE_wrapper_132__ap_ready) begin
          if(PE_wrapper_132__ap_done) begin
            PE_wrapper_132__state <= 2'b10;
          end else begin
            PE_wrapper_132__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_132__state == 2'b11) begin
        if(PE_wrapper_132__ap_done) begin
          PE_wrapper_132__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_132__state == 2'b10) begin
        if(PE_wrapper_132__ap_done_global__q0) begin
          PE_wrapper_132__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_132__ap_start = (PE_wrapper_132__state == 2'b01);
  assign PE_wrapper_133__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_133__is_done__q0 = (PE_wrapper_133__state == 2'b10);
  assign PE_wrapper_133__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_133__state <= 2'b00;
    end else begin
      if(PE_wrapper_133__state == 2'b00) begin
        if(PE_wrapper_133__ap_start_global__q0) begin
          PE_wrapper_133__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_133__state == 2'b01) begin
        if(PE_wrapper_133__ap_ready) begin
          if(PE_wrapper_133__ap_done) begin
            PE_wrapper_133__state <= 2'b10;
          end else begin
            PE_wrapper_133__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_133__state == 2'b11) begin
        if(PE_wrapper_133__ap_done) begin
          PE_wrapper_133__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_133__state == 2'b10) begin
        if(PE_wrapper_133__ap_done_global__q0) begin
          PE_wrapper_133__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_133__ap_start = (PE_wrapper_133__state == 2'b01);
  assign PE_wrapper_134__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_134__is_done__q0 = (PE_wrapper_134__state == 2'b10);
  assign PE_wrapper_134__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_134__state <= 2'b00;
    end else begin
      if(PE_wrapper_134__state == 2'b00) begin
        if(PE_wrapper_134__ap_start_global__q0) begin
          PE_wrapper_134__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_134__state == 2'b01) begin
        if(PE_wrapper_134__ap_ready) begin
          if(PE_wrapper_134__ap_done) begin
            PE_wrapper_134__state <= 2'b10;
          end else begin
            PE_wrapper_134__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_134__state == 2'b11) begin
        if(PE_wrapper_134__ap_done) begin
          PE_wrapper_134__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_134__state == 2'b10) begin
        if(PE_wrapper_134__ap_done_global__q0) begin
          PE_wrapper_134__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_134__ap_start = (PE_wrapper_134__state == 2'b01);
  assign PE_wrapper_135__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_135__is_done__q0 = (PE_wrapper_135__state == 2'b10);
  assign PE_wrapper_135__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_135__state <= 2'b00;
    end else begin
      if(PE_wrapper_135__state == 2'b00) begin
        if(PE_wrapper_135__ap_start_global__q0) begin
          PE_wrapper_135__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_135__state == 2'b01) begin
        if(PE_wrapper_135__ap_ready) begin
          if(PE_wrapper_135__ap_done) begin
            PE_wrapper_135__state <= 2'b10;
          end else begin
            PE_wrapper_135__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_135__state == 2'b11) begin
        if(PE_wrapper_135__ap_done) begin
          PE_wrapper_135__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_135__state == 2'b10) begin
        if(PE_wrapper_135__ap_done_global__q0) begin
          PE_wrapper_135__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_135__ap_start = (PE_wrapper_135__state == 2'b01);
  assign PE_wrapper_136__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_136__is_done__q0 = (PE_wrapper_136__state == 2'b10);
  assign PE_wrapper_136__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_136__state <= 2'b00;
    end else begin
      if(PE_wrapper_136__state == 2'b00) begin
        if(PE_wrapper_136__ap_start_global__q0) begin
          PE_wrapper_136__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_136__state == 2'b01) begin
        if(PE_wrapper_136__ap_ready) begin
          if(PE_wrapper_136__ap_done) begin
            PE_wrapper_136__state <= 2'b10;
          end else begin
            PE_wrapper_136__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_136__state == 2'b11) begin
        if(PE_wrapper_136__ap_done) begin
          PE_wrapper_136__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_136__state == 2'b10) begin
        if(PE_wrapper_136__ap_done_global__q0) begin
          PE_wrapper_136__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_136__ap_start = (PE_wrapper_136__state == 2'b01);
  assign PE_wrapper_137__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_137__is_done__q0 = (PE_wrapper_137__state == 2'b10);
  assign PE_wrapper_137__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_137__state <= 2'b00;
    end else begin
      if(PE_wrapper_137__state == 2'b00) begin
        if(PE_wrapper_137__ap_start_global__q0) begin
          PE_wrapper_137__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_137__state == 2'b01) begin
        if(PE_wrapper_137__ap_ready) begin
          if(PE_wrapper_137__ap_done) begin
            PE_wrapper_137__state <= 2'b10;
          end else begin
            PE_wrapper_137__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_137__state == 2'b11) begin
        if(PE_wrapper_137__ap_done) begin
          PE_wrapper_137__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_137__state == 2'b10) begin
        if(PE_wrapper_137__ap_done_global__q0) begin
          PE_wrapper_137__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_137__ap_start = (PE_wrapper_137__state == 2'b01);
  assign PE_wrapper_138__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_138__is_done__q0 = (PE_wrapper_138__state == 2'b10);
  assign PE_wrapper_138__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_138__state <= 2'b00;
    end else begin
      if(PE_wrapper_138__state == 2'b00) begin
        if(PE_wrapper_138__ap_start_global__q0) begin
          PE_wrapper_138__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_138__state == 2'b01) begin
        if(PE_wrapper_138__ap_ready) begin
          if(PE_wrapper_138__ap_done) begin
            PE_wrapper_138__state <= 2'b10;
          end else begin
            PE_wrapper_138__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_138__state == 2'b11) begin
        if(PE_wrapper_138__ap_done) begin
          PE_wrapper_138__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_138__state == 2'b10) begin
        if(PE_wrapper_138__ap_done_global__q0) begin
          PE_wrapper_138__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_138__ap_start = (PE_wrapper_138__state == 2'b01);
  assign PE_wrapper_139__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_139__is_done__q0 = (PE_wrapper_139__state == 2'b10);
  assign PE_wrapper_139__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_139__state <= 2'b00;
    end else begin
      if(PE_wrapper_139__state == 2'b00) begin
        if(PE_wrapper_139__ap_start_global__q0) begin
          PE_wrapper_139__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_139__state == 2'b01) begin
        if(PE_wrapper_139__ap_ready) begin
          if(PE_wrapper_139__ap_done) begin
            PE_wrapper_139__state <= 2'b10;
          end else begin
            PE_wrapper_139__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_139__state == 2'b11) begin
        if(PE_wrapper_139__ap_done) begin
          PE_wrapper_139__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_139__state == 2'b10) begin
        if(PE_wrapper_139__ap_done_global__q0) begin
          PE_wrapper_139__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_139__ap_start = (PE_wrapper_139__state == 2'b01);
  assign PE_wrapper_140__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_140__is_done__q0 = (PE_wrapper_140__state == 2'b10);
  assign PE_wrapper_140__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_140__state <= 2'b00;
    end else begin
      if(PE_wrapper_140__state == 2'b00) begin
        if(PE_wrapper_140__ap_start_global__q0) begin
          PE_wrapper_140__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_140__state == 2'b01) begin
        if(PE_wrapper_140__ap_ready) begin
          if(PE_wrapper_140__ap_done) begin
            PE_wrapper_140__state <= 2'b10;
          end else begin
            PE_wrapper_140__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_140__state == 2'b11) begin
        if(PE_wrapper_140__ap_done) begin
          PE_wrapper_140__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_140__state == 2'b10) begin
        if(PE_wrapper_140__ap_done_global__q0) begin
          PE_wrapper_140__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_140__ap_start = (PE_wrapper_140__state == 2'b01);
  assign PE_wrapper_141__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_141__is_done__q0 = (PE_wrapper_141__state == 2'b10);
  assign PE_wrapper_141__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_141__state <= 2'b00;
    end else begin
      if(PE_wrapper_141__state == 2'b00) begin
        if(PE_wrapper_141__ap_start_global__q0) begin
          PE_wrapper_141__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_141__state == 2'b01) begin
        if(PE_wrapper_141__ap_ready) begin
          if(PE_wrapper_141__ap_done) begin
            PE_wrapper_141__state <= 2'b10;
          end else begin
            PE_wrapper_141__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_141__state == 2'b11) begin
        if(PE_wrapper_141__ap_done) begin
          PE_wrapper_141__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_141__state == 2'b10) begin
        if(PE_wrapper_141__ap_done_global__q0) begin
          PE_wrapper_141__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_141__ap_start = (PE_wrapper_141__state == 2'b01);
  assign PE_wrapper_142__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_142__is_done__q0 = (PE_wrapper_142__state == 2'b10);
  assign PE_wrapper_142__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_142__state <= 2'b00;
    end else begin
      if(PE_wrapper_142__state == 2'b00) begin
        if(PE_wrapper_142__ap_start_global__q0) begin
          PE_wrapper_142__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_142__state == 2'b01) begin
        if(PE_wrapper_142__ap_ready) begin
          if(PE_wrapper_142__ap_done) begin
            PE_wrapper_142__state <= 2'b10;
          end else begin
            PE_wrapper_142__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_142__state == 2'b11) begin
        if(PE_wrapper_142__ap_done) begin
          PE_wrapper_142__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_142__state == 2'b10) begin
        if(PE_wrapper_142__ap_done_global__q0) begin
          PE_wrapper_142__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_142__ap_start = (PE_wrapper_142__state == 2'b01);
  assign PE_wrapper_143__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_143__is_done__q0 = (PE_wrapper_143__state == 2'b10);
  assign PE_wrapper_143__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_143__state <= 2'b00;
    end else begin
      if(PE_wrapper_143__state == 2'b00) begin
        if(PE_wrapper_143__ap_start_global__q0) begin
          PE_wrapper_143__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_143__state == 2'b01) begin
        if(PE_wrapper_143__ap_ready) begin
          if(PE_wrapper_143__ap_done) begin
            PE_wrapper_143__state <= 2'b10;
          end else begin
            PE_wrapper_143__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_143__state == 2'b11) begin
        if(PE_wrapper_143__ap_done) begin
          PE_wrapper_143__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_143__state == 2'b10) begin
        if(PE_wrapper_143__ap_done_global__q0) begin
          PE_wrapper_143__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_143__ap_start = (PE_wrapper_143__state == 2'b01);
  assign PE_wrapper_144__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_144__is_done__q0 = (PE_wrapper_144__state == 2'b10);
  assign PE_wrapper_144__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_144__state <= 2'b00;
    end else begin
      if(PE_wrapper_144__state == 2'b00) begin
        if(PE_wrapper_144__ap_start_global__q0) begin
          PE_wrapper_144__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_144__state == 2'b01) begin
        if(PE_wrapper_144__ap_ready) begin
          if(PE_wrapper_144__ap_done) begin
            PE_wrapper_144__state <= 2'b10;
          end else begin
            PE_wrapper_144__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_144__state == 2'b11) begin
        if(PE_wrapper_144__ap_done) begin
          PE_wrapper_144__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_144__state == 2'b10) begin
        if(PE_wrapper_144__ap_done_global__q0) begin
          PE_wrapper_144__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_144__ap_start = (PE_wrapper_144__state == 2'b01);
  assign PE_wrapper_145__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_145__is_done__q0 = (PE_wrapper_145__state == 2'b10);
  assign PE_wrapper_145__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_145__state <= 2'b00;
    end else begin
      if(PE_wrapper_145__state == 2'b00) begin
        if(PE_wrapper_145__ap_start_global__q0) begin
          PE_wrapper_145__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_145__state == 2'b01) begin
        if(PE_wrapper_145__ap_ready) begin
          if(PE_wrapper_145__ap_done) begin
            PE_wrapper_145__state <= 2'b10;
          end else begin
            PE_wrapper_145__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_145__state == 2'b11) begin
        if(PE_wrapper_145__ap_done) begin
          PE_wrapper_145__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_145__state == 2'b10) begin
        if(PE_wrapper_145__ap_done_global__q0) begin
          PE_wrapper_145__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_145__ap_start = (PE_wrapper_145__state == 2'b01);
  assign PE_wrapper_146__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_146__is_done__q0 = (PE_wrapper_146__state == 2'b10);
  assign PE_wrapper_146__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_146__state <= 2'b00;
    end else begin
      if(PE_wrapper_146__state == 2'b00) begin
        if(PE_wrapper_146__ap_start_global__q0) begin
          PE_wrapper_146__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_146__state == 2'b01) begin
        if(PE_wrapper_146__ap_ready) begin
          if(PE_wrapper_146__ap_done) begin
            PE_wrapper_146__state <= 2'b10;
          end else begin
            PE_wrapper_146__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_146__state == 2'b11) begin
        if(PE_wrapper_146__ap_done) begin
          PE_wrapper_146__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_146__state == 2'b10) begin
        if(PE_wrapper_146__ap_done_global__q0) begin
          PE_wrapper_146__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_146__ap_start = (PE_wrapper_146__state == 2'b01);
  assign PE_wrapper_147__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_147__is_done__q0 = (PE_wrapper_147__state == 2'b10);
  assign PE_wrapper_147__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_147__state <= 2'b00;
    end else begin
      if(PE_wrapper_147__state == 2'b00) begin
        if(PE_wrapper_147__ap_start_global__q0) begin
          PE_wrapper_147__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_147__state == 2'b01) begin
        if(PE_wrapper_147__ap_ready) begin
          if(PE_wrapper_147__ap_done) begin
            PE_wrapper_147__state <= 2'b10;
          end else begin
            PE_wrapper_147__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_147__state == 2'b11) begin
        if(PE_wrapper_147__ap_done) begin
          PE_wrapper_147__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_147__state == 2'b10) begin
        if(PE_wrapper_147__ap_done_global__q0) begin
          PE_wrapper_147__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_147__ap_start = (PE_wrapper_147__state == 2'b01);
  assign PE_wrapper_148__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_148__is_done__q0 = (PE_wrapper_148__state == 2'b10);
  assign PE_wrapper_148__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_148__state <= 2'b00;
    end else begin
      if(PE_wrapper_148__state == 2'b00) begin
        if(PE_wrapper_148__ap_start_global__q0) begin
          PE_wrapper_148__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_148__state == 2'b01) begin
        if(PE_wrapper_148__ap_ready) begin
          if(PE_wrapper_148__ap_done) begin
            PE_wrapper_148__state <= 2'b10;
          end else begin
            PE_wrapper_148__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_148__state == 2'b11) begin
        if(PE_wrapper_148__ap_done) begin
          PE_wrapper_148__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_148__state == 2'b10) begin
        if(PE_wrapper_148__ap_done_global__q0) begin
          PE_wrapper_148__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_148__ap_start = (PE_wrapper_148__state == 2'b01);
  assign PE_wrapper_149__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_149__is_done__q0 = (PE_wrapper_149__state == 2'b10);
  assign PE_wrapper_149__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_149__state <= 2'b00;
    end else begin
      if(PE_wrapper_149__state == 2'b00) begin
        if(PE_wrapper_149__ap_start_global__q0) begin
          PE_wrapper_149__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_149__state == 2'b01) begin
        if(PE_wrapper_149__ap_ready) begin
          if(PE_wrapper_149__ap_done) begin
            PE_wrapper_149__state <= 2'b10;
          end else begin
            PE_wrapper_149__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_149__state == 2'b11) begin
        if(PE_wrapper_149__ap_done) begin
          PE_wrapper_149__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_149__state == 2'b10) begin
        if(PE_wrapper_149__ap_done_global__q0) begin
          PE_wrapper_149__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_149__ap_start = (PE_wrapper_149__state == 2'b01);
  assign PE_wrapper_150__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_150__is_done__q0 = (PE_wrapper_150__state == 2'b10);
  assign PE_wrapper_150__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_150__state <= 2'b00;
    end else begin
      if(PE_wrapper_150__state == 2'b00) begin
        if(PE_wrapper_150__ap_start_global__q0) begin
          PE_wrapper_150__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_150__state == 2'b01) begin
        if(PE_wrapper_150__ap_ready) begin
          if(PE_wrapper_150__ap_done) begin
            PE_wrapper_150__state <= 2'b10;
          end else begin
            PE_wrapper_150__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_150__state == 2'b11) begin
        if(PE_wrapper_150__ap_done) begin
          PE_wrapper_150__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_150__state == 2'b10) begin
        if(PE_wrapper_150__ap_done_global__q0) begin
          PE_wrapper_150__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_150__ap_start = (PE_wrapper_150__state == 2'b01);
  assign PE_wrapper_151__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_151__is_done__q0 = (PE_wrapper_151__state == 2'b10);
  assign PE_wrapper_151__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_151__state <= 2'b00;
    end else begin
      if(PE_wrapper_151__state == 2'b00) begin
        if(PE_wrapper_151__ap_start_global__q0) begin
          PE_wrapper_151__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_151__state == 2'b01) begin
        if(PE_wrapper_151__ap_ready) begin
          if(PE_wrapper_151__ap_done) begin
            PE_wrapper_151__state <= 2'b10;
          end else begin
            PE_wrapper_151__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_151__state == 2'b11) begin
        if(PE_wrapper_151__ap_done) begin
          PE_wrapper_151__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_151__state == 2'b10) begin
        if(PE_wrapper_151__ap_done_global__q0) begin
          PE_wrapper_151__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_151__ap_start = (PE_wrapper_151__state == 2'b01);
  assign PE_wrapper_152__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_152__is_done__q0 = (PE_wrapper_152__state == 2'b10);
  assign PE_wrapper_152__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_152__state <= 2'b00;
    end else begin
      if(PE_wrapper_152__state == 2'b00) begin
        if(PE_wrapper_152__ap_start_global__q0) begin
          PE_wrapper_152__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_152__state == 2'b01) begin
        if(PE_wrapper_152__ap_ready) begin
          if(PE_wrapper_152__ap_done) begin
            PE_wrapper_152__state <= 2'b10;
          end else begin
            PE_wrapper_152__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_152__state == 2'b11) begin
        if(PE_wrapper_152__ap_done) begin
          PE_wrapper_152__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_152__state == 2'b10) begin
        if(PE_wrapper_152__ap_done_global__q0) begin
          PE_wrapper_152__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_152__ap_start = (PE_wrapper_152__state == 2'b01);
  assign PE_wrapper_153__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_153__is_done__q0 = (PE_wrapper_153__state == 2'b10);
  assign PE_wrapper_153__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_153__state <= 2'b00;
    end else begin
      if(PE_wrapper_153__state == 2'b00) begin
        if(PE_wrapper_153__ap_start_global__q0) begin
          PE_wrapper_153__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_153__state == 2'b01) begin
        if(PE_wrapper_153__ap_ready) begin
          if(PE_wrapper_153__ap_done) begin
            PE_wrapper_153__state <= 2'b10;
          end else begin
            PE_wrapper_153__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_153__state == 2'b11) begin
        if(PE_wrapper_153__ap_done) begin
          PE_wrapper_153__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_153__state == 2'b10) begin
        if(PE_wrapper_153__ap_done_global__q0) begin
          PE_wrapper_153__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_153__ap_start = (PE_wrapper_153__state == 2'b01);
  assign PE_wrapper_154__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_154__is_done__q0 = (PE_wrapper_154__state == 2'b10);
  assign PE_wrapper_154__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_154__state <= 2'b00;
    end else begin
      if(PE_wrapper_154__state == 2'b00) begin
        if(PE_wrapper_154__ap_start_global__q0) begin
          PE_wrapper_154__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_154__state == 2'b01) begin
        if(PE_wrapper_154__ap_ready) begin
          if(PE_wrapper_154__ap_done) begin
            PE_wrapper_154__state <= 2'b10;
          end else begin
            PE_wrapper_154__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_154__state == 2'b11) begin
        if(PE_wrapper_154__ap_done) begin
          PE_wrapper_154__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_154__state == 2'b10) begin
        if(PE_wrapper_154__ap_done_global__q0) begin
          PE_wrapper_154__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_154__ap_start = (PE_wrapper_154__state == 2'b01);
  assign PE_wrapper_155__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_155__is_done__q0 = (PE_wrapper_155__state == 2'b10);
  assign PE_wrapper_155__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_155__state <= 2'b00;
    end else begin
      if(PE_wrapper_155__state == 2'b00) begin
        if(PE_wrapper_155__ap_start_global__q0) begin
          PE_wrapper_155__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_155__state == 2'b01) begin
        if(PE_wrapper_155__ap_ready) begin
          if(PE_wrapper_155__ap_done) begin
            PE_wrapper_155__state <= 2'b10;
          end else begin
            PE_wrapper_155__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_155__state == 2'b11) begin
        if(PE_wrapper_155__ap_done) begin
          PE_wrapper_155__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_155__state == 2'b10) begin
        if(PE_wrapper_155__ap_done_global__q0) begin
          PE_wrapper_155__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_155__ap_start = (PE_wrapper_155__state == 2'b01);
  assign PE_wrapper_156__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_156__is_done__q0 = (PE_wrapper_156__state == 2'b10);
  assign PE_wrapper_156__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_156__state <= 2'b00;
    end else begin
      if(PE_wrapper_156__state == 2'b00) begin
        if(PE_wrapper_156__ap_start_global__q0) begin
          PE_wrapper_156__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_156__state == 2'b01) begin
        if(PE_wrapper_156__ap_ready) begin
          if(PE_wrapper_156__ap_done) begin
            PE_wrapper_156__state <= 2'b10;
          end else begin
            PE_wrapper_156__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_156__state == 2'b11) begin
        if(PE_wrapper_156__ap_done) begin
          PE_wrapper_156__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_156__state == 2'b10) begin
        if(PE_wrapper_156__ap_done_global__q0) begin
          PE_wrapper_156__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_156__ap_start = (PE_wrapper_156__state == 2'b01);
  assign PE_wrapper_157__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_157__is_done__q0 = (PE_wrapper_157__state == 2'b10);
  assign PE_wrapper_157__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_157__state <= 2'b00;
    end else begin
      if(PE_wrapper_157__state == 2'b00) begin
        if(PE_wrapper_157__ap_start_global__q0) begin
          PE_wrapper_157__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_157__state == 2'b01) begin
        if(PE_wrapper_157__ap_ready) begin
          if(PE_wrapper_157__ap_done) begin
            PE_wrapper_157__state <= 2'b10;
          end else begin
            PE_wrapper_157__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_157__state == 2'b11) begin
        if(PE_wrapper_157__ap_done) begin
          PE_wrapper_157__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_157__state == 2'b10) begin
        if(PE_wrapper_157__ap_done_global__q0) begin
          PE_wrapper_157__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_157__ap_start = (PE_wrapper_157__state == 2'b01);
  assign PE_wrapper_158__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_158__is_done__q0 = (PE_wrapper_158__state == 2'b10);
  assign PE_wrapper_158__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_158__state <= 2'b00;
    end else begin
      if(PE_wrapper_158__state == 2'b00) begin
        if(PE_wrapper_158__ap_start_global__q0) begin
          PE_wrapper_158__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_158__state == 2'b01) begin
        if(PE_wrapper_158__ap_ready) begin
          if(PE_wrapper_158__ap_done) begin
            PE_wrapper_158__state <= 2'b10;
          end else begin
            PE_wrapper_158__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_158__state == 2'b11) begin
        if(PE_wrapper_158__ap_done) begin
          PE_wrapper_158__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_158__state == 2'b10) begin
        if(PE_wrapper_158__ap_done_global__q0) begin
          PE_wrapper_158__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_158__ap_start = (PE_wrapper_158__state == 2'b01);
  assign PE_wrapper_159__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_159__is_done__q0 = (PE_wrapper_159__state == 2'b10);
  assign PE_wrapper_159__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_159__state <= 2'b00;
    end else begin
      if(PE_wrapper_159__state == 2'b00) begin
        if(PE_wrapper_159__ap_start_global__q0) begin
          PE_wrapper_159__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_159__state == 2'b01) begin
        if(PE_wrapper_159__ap_ready) begin
          if(PE_wrapper_159__ap_done) begin
            PE_wrapper_159__state <= 2'b10;
          end else begin
            PE_wrapper_159__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_159__state == 2'b11) begin
        if(PE_wrapper_159__ap_done) begin
          PE_wrapper_159__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_159__state == 2'b10) begin
        if(PE_wrapper_159__ap_done_global__q0) begin
          PE_wrapper_159__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_159__ap_start = (PE_wrapper_159__state == 2'b01);
  assign PE_wrapper_160__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_160__is_done__q0 = (PE_wrapper_160__state == 2'b10);
  assign PE_wrapper_160__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_160__state <= 2'b00;
    end else begin
      if(PE_wrapper_160__state == 2'b00) begin
        if(PE_wrapper_160__ap_start_global__q0) begin
          PE_wrapper_160__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_160__state == 2'b01) begin
        if(PE_wrapper_160__ap_ready) begin
          if(PE_wrapper_160__ap_done) begin
            PE_wrapper_160__state <= 2'b10;
          end else begin
            PE_wrapper_160__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_160__state == 2'b11) begin
        if(PE_wrapper_160__ap_done) begin
          PE_wrapper_160__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_160__state == 2'b10) begin
        if(PE_wrapper_160__ap_done_global__q0) begin
          PE_wrapper_160__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_160__ap_start = (PE_wrapper_160__state == 2'b01);
  assign PE_wrapper_161__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_161__is_done__q0 = (PE_wrapper_161__state == 2'b10);
  assign PE_wrapper_161__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_161__state <= 2'b00;
    end else begin
      if(PE_wrapper_161__state == 2'b00) begin
        if(PE_wrapper_161__ap_start_global__q0) begin
          PE_wrapper_161__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_161__state == 2'b01) begin
        if(PE_wrapper_161__ap_ready) begin
          if(PE_wrapper_161__ap_done) begin
            PE_wrapper_161__state <= 2'b10;
          end else begin
            PE_wrapper_161__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_161__state == 2'b11) begin
        if(PE_wrapper_161__ap_done) begin
          PE_wrapper_161__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_161__state == 2'b10) begin
        if(PE_wrapper_161__ap_done_global__q0) begin
          PE_wrapper_161__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_161__ap_start = (PE_wrapper_161__state == 2'b01);
  assign PE_wrapper_162__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_162__is_done__q0 = (PE_wrapper_162__state == 2'b10);
  assign PE_wrapper_162__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_162__state <= 2'b00;
    end else begin
      if(PE_wrapper_162__state == 2'b00) begin
        if(PE_wrapper_162__ap_start_global__q0) begin
          PE_wrapper_162__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_162__state == 2'b01) begin
        if(PE_wrapper_162__ap_ready) begin
          if(PE_wrapper_162__ap_done) begin
            PE_wrapper_162__state <= 2'b10;
          end else begin
            PE_wrapper_162__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_162__state == 2'b11) begin
        if(PE_wrapper_162__ap_done) begin
          PE_wrapper_162__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_162__state == 2'b10) begin
        if(PE_wrapper_162__ap_done_global__q0) begin
          PE_wrapper_162__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_162__ap_start = (PE_wrapper_162__state == 2'b01);
  assign PE_wrapper_163__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_163__is_done__q0 = (PE_wrapper_163__state == 2'b10);
  assign PE_wrapper_163__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_163__state <= 2'b00;
    end else begin
      if(PE_wrapper_163__state == 2'b00) begin
        if(PE_wrapper_163__ap_start_global__q0) begin
          PE_wrapper_163__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_163__state == 2'b01) begin
        if(PE_wrapper_163__ap_ready) begin
          if(PE_wrapper_163__ap_done) begin
            PE_wrapper_163__state <= 2'b10;
          end else begin
            PE_wrapper_163__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_163__state == 2'b11) begin
        if(PE_wrapper_163__ap_done) begin
          PE_wrapper_163__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_163__state == 2'b10) begin
        if(PE_wrapper_163__ap_done_global__q0) begin
          PE_wrapper_163__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_163__ap_start = (PE_wrapper_163__state == 2'b01);
  assign PE_wrapper_164__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_164__is_done__q0 = (PE_wrapper_164__state == 2'b10);
  assign PE_wrapper_164__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_164__state <= 2'b00;
    end else begin
      if(PE_wrapper_164__state == 2'b00) begin
        if(PE_wrapper_164__ap_start_global__q0) begin
          PE_wrapper_164__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_164__state == 2'b01) begin
        if(PE_wrapper_164__ap_ready) begin
          if(PE_wrapper_164__ap_done) begin
            PE_wrapper_164__state <= 2'b10;
          end else begin
            PE_wrapper_164__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_164__state == 2'b11) begin
        if(PE_wrapper_164__ap_done) begin
          PE_wrapper_164__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_164__state == 2'b10) begin
        if(PE_wrapper_164__ap_done_global__q0) begin
          PE_wrapper_164__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_164__ap_start = (PE_wrapper_164__state == 2'b01);
  assign PE_wrapper_165__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_165__is_done__q0 = (PE_wrapper_165__state == 2'b10);
  assign PE_wrapper_165__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_165__state <= 2'b00;
    end else begin
      if(PE_wrapper_165__state == 2'b00) begin
        if(PE_wrapper_165__ap_start_global__q0) begin
          PE_wrapper_165__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_165__state == 2'b01) begin
        if(PE_wrapper_165__ap_ready) begin
          if(PE_wrapper_165__ap_done) begin
            PE_wrapper_165__state <= 2'b10;
          end else begin
            PE_wrapper_165__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_165__state == 2'b11) begin
        if(PE_wrapper_165__ap_done) begin
          PE_wrapper_165__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_165__state == 2'b10) begin
        if(PE_wrapper_165__ap_done_global__q0) begin
          PE_wrapper_165__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_165__ap_start = (PE_wrapper_165__state == 2'b01);
  assign PE_wrapper_166__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_166__is_done__q0 = (PE_wrapper_166__state == 2'b10);
  assign PE_wrapper_166__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_166__state <= 2'b00;
    end else begin
      if(PE_wrapper_166__state == 2'b00) begin
        if(PE_wrapper_166__ap_start_global__q0) begin
          PE_wrapper_166__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_166__state == 2'b01) begin
        if(PE_wrapper_166__ap_ready) begin
          if(PE_wrapper_166__ap_done) begin
            PE_wrapper_166__state <= 2'b10;
          end else begin
            PE_wrapper_166__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_166__state == 2'b11) begin
        if(PE_wrapper_166__ap_done) begin
          PE_wrapper_166__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_166__state == 2'b10) begin
        if(PE_wrapper_166__ap_done_global__q0) begin
          PE_wrapper_166__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_166__ap_start = (PE_wrapper_166__state == 2'b01);
  assign PE_wrapper_167__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_167__is_done__q0 = (PE_wrapper_167__state == 2'b10);
  assign PE_wrapper_167__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_167__state <= 2'b00;
    end else begin
      if(PE_wrapper_167__state == 2'b00) begin
        if(PE_wrapper_167__ap_start_global__q0) begin
          PE_wrapper_167__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_167__state == 2'b01) begin
        if(PE_wrapper_167__ap_ready) begin
          if(PE_wrapper_167__ap_done) begin
            PE_wrapper_167__state <= 2'b10;
          end else begin
            PE_wrapper_167__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_167__state == 2'b11) begin
        if(PE_wrapper_167__ap_done) begin
          PE_wrapper_167__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_167__state == 2'b10) begin
        if(PE_wrapper_167__ap_done_global__q0) begin
          PE_wrapper_167__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_167__ap_start = (PE_wrapper_167__state == 2'b01);
  assign PE_wrapper_168__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_168__is_done__q0 = (PE_wrapper_168__state == 2'b10);
  assign PE_wrapper_168__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_168__state <= 2'b00;
    end else begin
      if(PE_wrapper_168__state == 2'b00) begin
        if(PE_wrapper_168__ap_start_global__q0) begin
          PE_wrapper_168__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_168__state == 2'b01) begin
        if(PE_wrapper_168__ap_ready) begin
          if(PE_wrapper_168__ap_done) begin
            PE_wrapper_168__state <= 2'b10;
          end else begin
            PE_wrapper_168__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_168__state == 2'b11) begin
        if(PE_wrapper_168__ap_done) begin
          PE_wrapper_168__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_168__state == 2'b10) begin
        if(PE_wrapper_168__ap_done_global__q0) begin
          PE_wrapper_168__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_168__ap_start = (PE_wrapper_168__state == 2'b01);
  assign PE_wrapper_169__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_169__is_done__q0 = (PE_wrapper_169__state == 2'b10);
  assign PE_wrapper_169__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_169__state <= 2'b00;
    end else begin
      if(PE_wrapper_169__state == 2'b00) begin
        if(PE_wrapper_169__ap_start_global__q0) begin
          PE_wrapper_169__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_169__state == 2'b01) begin
        if(PE_wrapper_169__ap_ready) begin
          if(PE_wrapper_169__ap_done) begin
            PE_wrapper_169__state <= 2'b10;
          end else begin
            PE_wrapper_169__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_169__state == 2'b11) begin
        if(PE_wrapper_169__ap_done) begin
          PE_wrapper_169__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_169__state == 2'b10) begin
        if(PE_wrapper_169__ap_done_global__q0) begin
          PE_wrapper_169__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_169__ap_start = (PE_wrapper_169__state == 2'b01);
  assign PE_wrapper_170__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_170__is_done__q0 = (PE_wrapper_170__state == 2'b10);
  assign PE_wrapper_170__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_170__state <= 2'b00;
    end else begin
      if(PE_wrapper_170__state == 2'b00) begin
        if(PE_wrapper_170__ap_start_global__q0) begin
          PE_wrapper_170__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_170__state == 2'b01) begin
        if(PE_wrapper_170__ap_ready) begin
          if(PE_wrapper_170__ap_done) begin
            PE_wrapper_170__state <= 2'b10;
          end else begin
            PE_wrapper_170__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_170__state == 2'b11) begin
        if(PE_wrapper_170__ap_done) begin
          PE_wrapper_170__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_170__state == 2'b10) begin
        if(PE_wrapper_170__ap_done_global__q0) begin
          PE_wrapper_170__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_170__ap_start = (PE_wrapper_170__state == 2'b01);
  assign PE_wrapper_171__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_171__is_done__q0 = (PE_wrapper_171__state == 2'b10);
  assign PE_wrapper_171__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_171__state <= 2'b00;
    end else begin
      if(PE_wrapper_171__state == 2'b00) begin
        if(PE_wrapper_171__ap_start_global__q0) begin
          PE_wrapper_171__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_171__state == 2'b01) begin
        if(PE_wrapper_171__ap_ready) begin
          if(PE_wrapper_171__ap_done) begin
            PE_wrapper_171__state <= 2'b10;
          end else begin
            PE_wrapper_171__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_171__state == 2'b11) begin
        if(PE_wrapper_171__ap_done) begin
          PE_wrapper_171__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_171__state == 2'b10) begin
        if(PE_wrapper_171__ap_done_global__q0) begin
          PE_wrapper_171__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_171__ap_start = (PE_wrapper_171__state == 2'b01);
  assign PE_wrapper_172__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_172__is_done__q0 = (PE_wrapper_172__state == 2'b10);
  assign PE_wrapper_172__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_172__state <= 2'b00;
    end else begin
      if(PE_wrapper_172__state == 2'b00) begin
        if(PE_wrapper_172__ap_start_global__q0) begin
          PE_wrapper_172__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_172__state == 2'b01) begin
        if(PE_wrapper_172__ap_ready) begin
          if(PE_wrapper_172__ap_done) begin
            PE_wrapper_172__state <= 2'b10;
          end else begin
            PE_wrapper_172__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_172__state == 2'b11) begin
        if(PE_wrapper_172__ap_done) begin
          PE_wrapper_172__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_172__state == 2'b10) begin
        if(PE_wrapper_172__ap_done_global__q0) begin
          PE_wrapper_172__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_172__ap_start = (PE_wrapper_172__state == 2'b01);
  assign PE_wrapper_173__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_173__is_done__q0 = (PE_wrapper_173__state == 2'b10);
  assign PE_wrapper_173__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_173__state <= 2'b00;
    end else begin
      if(PE_wrapper_173__state == 2'b00) begin
        if(PE_wrapper_173__ap_start_global__q0) begin
          PE_wrapper_173__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_173__state == 2'b01) begin
        if(PE_wrapper_173__ap_ready) begin
          if(PE_wrapper_173__ap_done) begin
            PE_wrapper_173__state <= 2'b10;
          end else begin
            PE_wrapper_173__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_173__state == 2'b11) begin
        if(PE_wrapper_173__ap_done) begin
          PE_wrapper_173__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_173__state == 2'b10) begin
        if(PE_wrapper_173__ap_done_global__q0) begin
          PE_wrapper_173__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_173__ap_start = (PE_wrapper_173__state == 2'b01);
  assign PE_wrapper_174__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_174__is_done__q0 = (PE_wrapper_174__state == 2'b10);
  assign PE_wrapper_174__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_174__state <= 2'b00;
    end else begin
      if(PE_wrapper_174__state == 2'b00) begin
        if(PE_wrapper_174__ap_start_global__q0) begin
          PE_wrapper_174__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_174__state == 2'b01) begin
        if(PE_wrapper_174__ap_ready) begin
          if(PE_wrapper_174__ap_done) begin
            PE_wrapper_174__state <= 2'b10;
          end else begin
            PE_wrapper_174__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_174__state == 2'b11) begin
        if(PE_wrapper_174__ap_done) begin
          PE_wrapper_174__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_174__state == 2'b10) begin
        if(PE_wrapper_174__ap_done_global__q0) begin
          PE_wrapper_174__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_174__ap_start = (PE_wrapper_174__state == 2'b01);
  assign PE_wrapper_175__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_175__is_done__q0 = (PE_wrapper_175__state == 2'b10);
  assign PE_wrapper_175__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_175__state <= 2'b00;
    end else begin
      if(PE_wrapper_175__state == 2'b00) begin
        if(PE_wrapper_175__ap_start_global__q0) begin
          PE_wrapper_175__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_175__state == 2'b01) begin
        if(PE_wrapper_175__ap_ready) begin
          if(PE_wrapper_175__ap_done) begin
            PE_wrapper_175__state <= 2'b10;
          end else begin
            PE_wrapper_175__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_175__state == 2'b11) begin
        if(PE_wrapper_175__ap_done) begin
          PE_wrapper_175__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_175__state == 2'b10) begin
        if(PE_wrapper_175__ap_done_global__q0) begin
          PE_wrapper_175__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_175__ap_start = (PE_wrapper_175__state == 2'b01);
  assign PE_wrapper_176__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_176__is_done__q0 = (PE_wrapper_176__state == 2'b10);
  assign PE_wrapper_176__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_176__state <= 2'b00;
    end else begin
      if(PE_wrapper_176__state == 2'b00) begin
        if(PE_wrapper_176__ap_start_global__q0) begin
          PE_wrapper_176__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_176__state == 2'b01) begin
        if(PE_wrapper_176__ap_ready) begin
          if(PE_wrapper_176__ap_done) begin
            PE_wrapper_176__state <= 2'b10;
          end else begin
            PE_wrapper_176__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_176__state == 2'b11) begin
        if(PE_wrapper_176__ap_done) begin
          PE_wrapper_176__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_176__state == 2'b10) begin
        if(PE_wrapper_176__ap_done_global__q0) begin
          PE_wrapper_176__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_176__ap_start = (PE_wrapper_176__state == 2'b01);
  assign PE_wrapper_177__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_177__is_done__q0 = (PE_wrapper_177__state == 2'b10);
  assign PE_wrapper_177__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_177__state <= 2'b00;
    end else begin
      if(PE_wrapper_177__state == 2'b00) begin
        if(PE_wrapper_177__ap_start_global__q0) begin
          PE_wrapper_177__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_177__state == 2'b01) begin
        if(PE_wrapper_177__ap_ready) begin
          if(PE_wrapper_177__ap_done) begin
            PE_wrapper_177__state <= 2'b10;
          end else begin
            PE_wrapper_177__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_177__state == 2'b11) begin
        if(PE_wrapper_177__ap_done) begin
          PE_wrapper_177__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_177__state == 2'b10) begin
        if(PE_wrapper_177__ap_done_global__q0) begin
          PE_wrapper_177__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_177__ap_start = (PE_wrapper_177__state == 2'b01);
  assign PE_wrapper_178__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_178__is_done__q0 = (PE_wrapper_178__state == 2'b10);
  assign PE_wrapper_178__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_178__state <= 2'b00;
    end else begin
      if(PE_wrapper_178__state == 2'b00) begin
        if(PE_wrapper_178__ap_start_global__q0) begin
          PE_wrapper_178__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_178__state == 2'b01) begin
        if(PE_wrapper_178__ap_ready) begin
          if(PE_wrapper_178__ap_done) begin
            PE_wrapper_178__state <= 2'b10;
          end else begin
            PE_wrapper_178__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_178__state == 2'b11) begin
        if(PE_wrapper_178__ap_done) begin
          PE_wrapper_178__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_178__state == 2'b10) begin
        if(PE_wrapper_178__ap_done_global__q0) begin
          PE_wrapper_178__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_178__ap_start = (PE_wrapper_178__state == 2'b01);
  assign PE_wrapper_179__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_179__is_done__q0 = (PE_wrapper_179__state == 2'b10);
  assign PE_wrapper_179__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_179__state <= 2'b00;
    end else begin
      if(PE_wrapper_179__state == 2'b00) begin
        if(PE_wrapper_179__ap_start_global__q0) begin
          PE_wrapper_179__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_179__state == 2'b01) begin
        if(PE_wrapper_179__ap_ready) begin
          if(PE_wrapper_179__ap_done) begin
            PE_wrapper_179__state <= 2'b10;
          end else begin
            PE_wrapper_179__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_179__state == 2'b11) begin
        if(PE_wrapper_179__ap_done) begin
          PE_wrapper_179__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_179__state == 2'b10) begin
        if(PE_wrapper_179__ap_done_global__q0) begin
          PE_wrapper_179__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_179__ap_start = (PE_wrapper_179__state == 2'b01);
  assign PE_wrapper_180__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_180__is_done__q0 = (PE_wrapper_180__state == 2'b10);
  assign PE_wrapper_180__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_180__state <= 2'b00;
    end else begin
      if(PE_wrapper_180__state == 2'b00) begin
        if(PE_wrapper_180__ap_start_global__q0) begin
          PE_wrapper_180__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_180__state == 2'b01) begin
        if(PE_wrapper_180__ap_ready) begin
          if(PE_wrapper_180__ap_done) begin
            PE_wrapper_180__state <= 2'b10;
          end else begin
            PE_wrapper_180__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_180__state == 2'b11) begin
        if(PE_wrapper_180__ap_done) begin
          PE_wrapper_180__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_180__state == 2'b10) begin
        if(PE_wrapper_180__ap_done_global__q0) begin
          PE_wrapper_180__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_180__ap_start = (PE_wrapper_180__state == 2'b01);
  assign PE_wrapper_181__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_181__is_done__q0 = (PE_wrapper_181__state == 2'b10);
  assign PE_wrapper_181__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_181__state <= 2'b00;
    end else begin
      if(PE_wrapper_181__state == 2'b00) begin
        if(PE_wrapper_181__ap_start_global__q0) begin
          PE_wrapper_181__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_181__state == 2'b01) begin
        if(PE_wrapper_181__ap_ready) begin
          if(PE_wrapper_181__ap_done) begin
            PE_wrapper_181__state <= 2'b10;
          end else begin
            PE_wrapper_181__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_181__state == 2'b11) begin
        if(PE_wrapper_181__ap_done) begin
          PE_wrapper_181__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_181__state == 2'b10) begin
        if(PE_wrapper_181__ap_done_global__q0) begin
          PE_wrapper_181__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_181__ap_start = (PE_wrapper_181__state == 2'b01);
  assign PE_wrapper_182__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_182__is_done__q0 = (PE_wrapper_182__state == 2'b10);
  assign PE_wrapper_182__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_182__state <= 2'b00;
    end else begin
      if(PE_wrapper_182__state == 2'b00) begin
        if(PE_wrapper_182__ap_start_global__q0) begin
          PE_wrapper_182__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_182__state == 2'b01) begin
        if(PE_wrapper_182__ap_ready) begin
          if(PE_wrapper_182__ap_done) begin
            PE_wrapper_182__state <= 2'b10;
          end else begin
            PE_wrapper_182__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_182__state == 2'b11) begin
        if(PE_wrapper_182__ap_done) begin
          PE_wrapper_182__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_182__state == 2'b10) begin
        if(PE_wrapper_182__ap_done_global__q0) begin
          PE_wrapper_182__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_182__ap_start = (PE_wrapper_182__state == 2'b01);
  assign PE_wrapper_183__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_183__is_done__q0 = (PE_wrapper_183__state == 2'b10);
  assign PE_wrapper_183__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_183__state <= 2'b00;
    end else begin
      if(PE_wrapper_183__state == 2'b00) begin
        if(PE_wrapper_183__ap_start_global__q0) begin
          PE_wrapper_183__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_183__state == 2'b01) begin
        if(PE_wrapper_183__ap_ready) begin
          if(PE_wrapper_183__ap_done) begin
            PE_wrapper_183__state <= 2'b10;
          end else begin
            PE_wrapper_183__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_183__state == 2'b11) begin
        if(PE_wrapper_183__ap_done) begin
          PE_wrapper_183__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_183__state == 2'b10) begin
        if(PE_wrapper_183__ap_done_global__q0) begin
          PE_wrapper_183__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_183__ap_start = (PE_wrapper_183__state == 2'b01);
  assign PE_wrapper_184__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_184__is_done__q0 = (PE_wrapper_184__state == 2'b10);
  assign PE_wrapper_184__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_184__state <= 2'b00;
    end else begin
      if(PE_wrapper_184__state == 2'b00) begin
        if(PE_wrapper_184__ap_start_global__q0) begin
          PE_wrapper_184__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_184__state == 2'b01) begin
        if(PE_wrapper_184__ap_ready) begin
          if(PE_wrapper_184__ap_done) begin
            PE_wrapper_184__state <= 2'b10;
          end else begin
            PE_wrapper_184__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_184__state == 2'b11) begin
        if(PE_wrapper_184__ap_done) begin
          PE_wrapper_184__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_184__state == 2'b10) begin
        if(PE_wrapper_184__ap_done_global__q0) begin
          PE_wrapper_184__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_184__ap_start = (PE_wrapper_184__state == 2'b01);
  assign PE_wrapper_185__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_185__is_done__q0 = (PE_wrapper_185__state == 2'b10);
  assign PE_wrapper_185__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_185__state <= 2'b00;
    end else begin
      if(PE_wrapper_185__state == 2'b00) begin
        if(PE_wrapper_185__ap_start_global__q0) begin
          PE_wrapper_185__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_185__state == 2'b01) begin
        if(PE_wrapper_185__ap_ready) begin
          if(PE_wrapper_185__ap_done) begin
            PE_wrapper_185__state <= 2'b10;
          end else begin
            PE_wrapper_185__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_185__state == 2'b11) begin
        if(PE_wrapper_185__ap_done) begin
          PE_wrapper_185__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_185__state == 2'b10) begin
        if(PE_wrapper_185__ap_done_global__q0) begin
          PE_wrapper_185__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_185__ap_start = (PE_wrapper_185__state == 2'b01);
  assign PE_wrapper_186__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_186__is_done__q0 = (PE_wrapper_186__state == 2'b10);
  assign PE_wrapper_186__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_186__state <= 2'b00;
    end else begin
      if(PE_wrapper_186__state == 2'b00) begin
        if(PE_wrapper_186__ap_start_global__q0) begin
          PE_wrapper_186__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_186__state == 2'b01) begin
        if(PE_wrapper_186__ap_ready) begin
          if(PE_wrapper_186__ap_done) begin
            PE_wrapper_186__state <= 2'b10;
          end else begin
            PE_wrapper_186__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_186__state == 2'b11) begin
        if(PE_wrapper_186__ap_done) begin
          PE_wrapper_186__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_186__state == 2'b10) begin
        if(PE_wrapper_186__ap_done_global__q0) begin
          PE_wrapper_186__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_186__ap_start = (PE_wrapper_186__state == 2'b01);
  assign PE_wrapper_187__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_187__is_done__q0 = (PE_wrapper_187__state == 2'b10);
  assign PE_wrapper_187__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_187__state <= 2'b00;
    end else begin
      if(PE_wrapper_187__state == 2'b00) begin
        if(PE_wrapper_187__ap_start_global__q0) begin
          PE_wrapper_187__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_187__state == 2'b01) begin
        if(PE_wrapper_187__ap_ready) begin
          if(PE_wrapper_187__ap_done) begin
            PE_wrapper_187__state <= 2'b10;
          end else begin
            PE_wrapper_187__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_187__state == 2'b11) begin
        if(PE_wrapper_187__ap_done) begin
          PE_wrapper_187__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_187__state == 2'b10) begin
        if(PE_wrapper_187__ap_done_global__q0) begin
          PE_wrapper_187__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_187__ap_start = (PE_wrapper_187__state == 2'b01);
  assign PE_wrapper_188__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_188__is_done__q0 = (PE_wrapper_188__state == 2'b10);
  assign PE_wrapper_188__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_188__state <= 2'b00;
    end else begin
      if(PE_wrapper_188__state == 2'b00) begin
        if(PE_wrapper_188__ap_start_global__q0) begin
          PE_wrapper_188__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_188__state == 2'b01) begin
        if(PE_wrapper_188__ap_ready) begin
          if(PE_wrapper_188__ap_done) begin
            PE_wrapper_188__state <= 2'b10;
          end else begin
            PE_wrapper_188__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_188__state == 2'b11) begin
        if(PE_wrapper_188__ap_done) begin
          PE_wrapper_188__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_188__state == 2'b10) begin
        if(PE_wrapper_188__ap_done_global__q0) begin
          PE_wrapper_188__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_188__ap_start = (PE_wrapper_188__state == 2'b01);
  assign PE_wrapper_189__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_189__is_done__q0 = (PE_wrapper_189__state == 2'b10);
  assign PE_wrapper_189__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_189__state <= 2'b00;
    end else begin
      if(PE_wrapper_189__state == 2'b00) begin
        if(PE_wrapper_189__ap_start_global__q0) begin
          PE_wrapper_189__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_189__state == 2'b01) begin
        if(PE_wrapper_189__ap_ready) begin
          if(PE_wrapper_189__ap_done) begin
            PE_wrapper_189__state <= 2'b10;
          end else begin
            PE_wrapper_189__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_189__state == 2'b11) begin
        if(PE_wrapper_189__ap_done) begin
          PE_wrapper_189__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_189__state == 2'b10) begin
        if(PE_wrapper_189__ap_done_global__q0) begin
          PE_wrapper_189__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_189__ap_start = (PE_wrapper_189__state == 2'b01);
  assign PE_wrapper_190__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_190__is_done__q0 = (PE_wrapper_190__state == 2'b10);
  assign PE_wrapper_190__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_190__state <= 2'b00;
    end else begin
      if(PE_wrapper_190__state == 2'b00) begin
        if(PE_wrapper_190__ap_start_global__q0) begin
          PE_wrapper_190__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_190__state == 2'b01) begin
        if(PE_wrapper_190__ap_ready) begin
          if(PE_wrapper_190__ap_done) begin
            PE_wrapper_190__state <= 2'b10;
          end else begin
            PE_wrapper_190__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_190__state == 2'b11) begin
        if(PE_wrapper_190__ap_done) begin
          PE_wrapper_190__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_190__state == 2'b10) begin
        if(PE_wrapper_190__ap_done_global__q0) begin
          PE_wrapper_190__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_190__ap_start = (PE_wrapper_190__state == 2'b01);
  assign PE_wrapper_191__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_191__is_done__q0 = (PE_wrapper_191__state == 2'b10);
  assign PE_wrapper_191__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_191__state <= 2'b00;
    end else begin
      if(PE_wrapper_191__state == 2'b00) begin
        if(PE_wrapper_191__ap_start_global__q0) begin
          PE_wrapper_191__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_191__state == 2'b01) begin
        if(PE_wrapper_191__ap_ready) begin
          if(PE_wrapper_191__ap_done) begin
            PE_wrapper_191__state <= 2'b10;
          end else begin
            PE_wrapper_191__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_191__state == 2'b11) begin
        if(PE_wrapper_191__ap_done) begin
          PE_wrapper_191__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_191__state == 2'b10) begin
        if(PE_wrapper_191__ap_done_global__q0) begin
          PE_wrapper_191__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_191__ap_start = (PE_wrapper_191__state == 2'b01);
  assign PE_wrapper_192__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_192__is_done__q0 = (PE_wrapper_192__state == 2'b10);
  assign PE_wrapper_192__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_192__state <= 2'b00;
    end else begin
      if(PE_wrapper_192__state == 2'b00) begin
        if(PE_wrapper_192__ap_start_global__q0) begin
          PE_wrapper_192__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_192__state == 2'b01) begin
        if(PE_wrapper_192__ap_ready) begin
          if(PE_wrapper_192__ap_done) begin
            PE_wrapper_192__state <= 2'b10;
          end else begin
            PE_wrapper_192__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_192__state == 2'b11) begin
        if(PE_wrapper_192__ap_done) begin
          PE_wrapper_192__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_192__state == 2'b10) begin
        if(PE_wrapper_192__ap_done_global__q0) begin
          PE_wrapper_192__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_192__ap_start = (PE_wrapper_192__state == 2'b01);
  assign PE_wrapper_193__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_193__is_done__q0 = (PE_wrapper_193__state == 2'b10);
  assign PE_wrapper_193__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_193__state <= 2'b00;
    end else begin
      if(PE_wrapper_193__state == 2'b00) begin
        if(PE_wrapper_193__ap_start_global__q0) begin
          PE_wrapper_193__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_193__state == 2'b01) begin
        if(PE_wrapper_193__ap_ready) begin
          if(PE_wrapper_193__ap_done) begin
            PE_wrapper_193__state <= 2'b10;
          end else begin
            PE_wrapper_193__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_193__state == 2'b11) begin
        if(PE_wrapper_193__ap_done) begin
          PE_wrapper_193__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_193__state == 2'b10) begin
        if(PE_wrapper_193__ap_done_global__q0) begin
          PE_wrapper_193__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_193__ap_start = (PE_wrapper_193__state == 2'b01);
  assign PE_wrapper_194__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_194__is_done__q0 = (PE_wrapper_194__state == 2'b10);
  assign PE_wrapper_194__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_194__state <= 2'b00;
    end else begin
      if(PE_wrapper_194__state == 2'b00) begin
        if(PE_wrapper_194__ap_start_global__q0) begin
          PE_wrapper_194__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_194__state == 2'b01) begin
        if(PE_wrapper_194__ap_ready) begin
          if(PE_wrapper_194__ap_done) begin
            PE_wrapper_194__state <= 2'b10;
          end else begin
            PE_wrapper_194__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_194__state == 2'b11) begin
        if(PE_wrapper_194__ap_done) begin
          PE_wrapper_194__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_194__state == 2'b10) begin
        if(PE_wrapper_194__ap_done_global__q0) begin
          PE_wrapper_194__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_194__ap_start = (PE_wrapper_194__state == 2'b01);
  assign PE_wrapper_195__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_195__is_done__q0 = (PE_wrapper_195__state == 2'b10);
  assign PE_wrapper_195__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_195__state <= 2'b00;
    end else begin
      if(PE_wrapper_195__state == 2'b00) begin
        if(PE_wrapper_195__ap_start_global__q0) begin
          PE_wrapper_195__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_195__state == 2'b01) begin
        if(PE_wrapper_195__ap_ready) begin
          if(PE_wrapper_195__ap_done) begin
            PE_wrapper_195__state <= 2'b10;
          end else begin
            PE_wrapper_195__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_195__state == 2'b11) begin
        if(PE_wrapper_195__ap_done) begin
          PE_wrapper_195__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_195__state == 2'b10) begin
        if(PE_wrapper_195__ap_done_global__q0) begin
          PE_wrapper_195__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_195__ap_start = (PE_wrapper_195__state == 2'b01);
  assign PE_wrapper_196__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_196__is_done__q0 = (PE_wrapper_196__state == 2'b10);
  assign PE_wrapper_196__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_196__state <= 2'b00;
    end else begin
      if(PE_wrapper_196__state == 2'b00) begin
        if(PE_wrapper_196__ap_start_global__q0) begin
          PE_wrapper_196__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_196__state == 2'b01) begin
        if(PE_wrapper_196__ap_ready) begin
          if(PE_wrapper_196__ap_done) begin
            PE_wrapper_196__state <= 2'b10;
          end else begin
            PE_wrapper_196__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_196__state == 2'b11) begin
        if(PE_wrapper_196__ap_done) begin
          PE_wrapper_196__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_196__state == 2'b10) begin
        if(PE_wrapper_196__ap_done_global__q0) begin
          PE_wrapper_196__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_196__ap_start = (PE_wrapper_196__state == 2'b01);
  assign PE_wrapper_197__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_197__is_done__q0 = (PE_wrapper_197__state == 2'b10);
  assign PE_wrapper_197__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_197__state <= 2'b00;
    end else begin
      if(PE_wrapper_197__state == 2'b00) begin
        if(PE_wrapper_197__ap_start_global__q0) begin
          PE_wrapper_197__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_197__state == 2'b01) begin
        if(PE_wrapper_197__ap_ready) begin
          if(PE_wrapper_197__ap_done) begin
            PE_wrapper_197__state <= 2'b10;
          end else begin
            PE_wrapper_197__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_197__state == 2'b11) begin
        if(PE_wrapper_197__ap_done) begin
          PE_wrapper_197__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_197__state == 2'b10) begin
        if(PE_wrapper_197__ap_done_global__q0) begin
          PE_wrapper_197__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_197__ap_start = (PE_wrapper_197__state == 2'b01);
  assign PE_wrapper_198__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_198__is_done__q0 = (PE_wrapper_198__state == 2'b10);
  assign PE_wrapper_198__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_198__state <= 2'b00;
    end else begin
      if(PE_wrapper_198__state == 2'b00) begin
        if(PE_wrapper_198__ap_start_global__q0) begin
          PE_wrapper_198__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_198__state == 2'b01) begin
        if(PE_wrapper_198__ap_ready) begin
          if(PE_wrapper_198__ap_done) begin
            PE_wrapper_198__state <= 2'b10;
          end else begin
            PE_wrapper_198__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_198__state == 2'b11) begin
        if(PE_wrapper_198__ap_done) begin
          PE_wrapper_198__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_198__state == 2'b10) begin
        if(PE_wrapper_198__ap_done_global__q0) begin
          PE_wrapper_198__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_198__ap_start = (PE_wrapper_198__state == 2'b01);
  assign PE_wrapper_199__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_199__is_done__q0 = (PE_wrapper_199__state == 2'b10);
  assign PE_wrapper_199__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_199__state <= 2'b00;
    end else begin
      if(PE_wrapper_199__state == 2'b00) begin
        if(PE_wrapper_199__ap_start_global__q0) begin
          PE_wrapper_199__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_199__state == 2'b01) begin
        if(PE_wrapper_199__ap_ready) begin
          if(PE_wrapper_199__ap_done) begin
            PE_wrapper_199__state <= 2'b10;
          end else begin
            PE_wrapper_199__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_199__state == 2'b11) begin
        if(PE_wrapper_199__ap_done) begin
          PE_wrapper_199__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_199__state == 2'b10) begin
        if(PE_wrapper_199__ap_done_global__q0) begin
          PE_wrapper_199__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_199__ap_start = (PE_wrapper_199__state == 2'b01);
  assign PE_wrapper_200__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_200__is_done__q0 = (PE_wrapper_200__state == 2'b10);
  assign PE_wrapper_200__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_200__state <= 2'b00;
    end else begin
      if(PE_wrapper_200__state == 2'b00) begin
        if(PE_wrapper_200__ap_start_global__q0) begin
          PE_wrapper_200__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_200__state == 2'b01) begin
        if(PE_wrapper_200__ap_ready) begin
          if(PE_wrapper_200__ap_done) begin
            PE_wrapper_200__state <= 2'b10;
          end else begin
            PE_wrapper_200__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_200__state == 2'b11) begin
        if(PE_wrapper_200__ap_done) begin
          PE_wrapper_200__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_200__state == 2'b10) begin
        if(PE_wrapper_200__ap_done_global__q0) begin
          PE_wrapper_200__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_200__ap_start = (PE_wrapper_200__state == 2'b01);
  assign PE_wrapper_201__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_201__is_done__q0 = (PE_wrapper_201__state == 2'b10);
  assign PE_wrapper_201__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_201__state <= 2'b00;
    end else begin
      if(PE_wrapper_201__state == 2'b00) begin
        if(PE_wrapper_201__ap_start_global__q0) begin
          PE_wrapper_201__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_201__state == 2'b01) begin
        if(PE_wrapper_201__ap_ready) begin
          if(PE_wrapper_201__ap_done) begin
            PE_wrapper_201__state <= 2'b10;
          end else begin
            PE_wrapper_201__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_201__state == 2'b11) begin
        if(PE_wrapper_201__ap_done) begin
          PE_wrapper_201__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_201__state == 2'b10) begin
        if(PE_wrapper_201__ap_done_global__q0) begin
          PE_wrapper_201__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_201__ap_start = (PE_wrapper_201__state == 2'b01);
  assign PE_wrapper_202__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_202__is_done__q0 = (PE_wrapper_202__state == 2'b10);
  assign PE_wrapper_202__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_202__state <= 2'b00;
    end else begin
      if(PE_wrapper_202__state == 2'b00) begin
        if(PE_wrapper_202__ap_start_global__q0) begin
          PE_wrapper_202__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_202__state == 2'b01) begin
        if(PE_wrapper_202__ap_ready) begin
          if(PE_wrapper_202__ap_done) begin
            PE_wrapper_202__state <= 2'b10;
          end else begin
            PE_wrapper_202__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_202__state == 2'b11) begin
        if(PE_wrapper_202__ap_done) begin
          PE_wrapper_202__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_202__state == 2'b10) begin
        if(PE_wrapper_202__ap_done_global__q0) begin
          PE_wrapper_202__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_202__ap_start = (PE_wrapper_202__state == 2'b01);
  assign PE_wrapper_203__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_203__is_done__q0 = (PE_wrapper_203__state == 2'b10);
  assign PE_wrapper_203__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_203__state <= 2'b00;
    end else begin
      if(PE_wrapper_203__state == 2'b00) begin
        if(PE_wrapper_203__ap_start_global__q0) begin
          PE_wrapper_203__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_203__state == 2'b01) begin
        if(PE_wrapper_203__ap_ready) begin
          if(PE_wrapper_203__ap_done) begin
            PE_wrapper_203__state <= 2'b10;
          end else begin
            PE_wrapper_203__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_203__state == 2'b11) begin
        if(PE_wrapper_203__ap_done) begin
          PE_wrapper_203__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_203__state == 2'b10) begin
        if(PE_wrapper_203__ap_done_global__q0) begin
          PE_wrapper_203__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_203__ap_start = (PE_wrapper_203__state == 2'b01);
  assign PE_wrapper_204__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_204__is_done__q0 = (PE_wrapper_204__state == 2'b10);
  assign PE_wrapper_204__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_204__state <= 2'b00;
    end else begin
      if(PE_wrapper_204__state == 2'b00) begin
        if(PE_wrapper_204__ap_start_global__q0) begin
          PE_wrapper_204__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_204__state == 2'b01) begin
        if(PE_wrapper_204__ap_ready) begin
          if(PE_wrapper_204__ap_done) begin
            PE_wrapper_204__state <= 2'b10;
          end else begin
            PE_wrapper_204__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_204__state == 2'b11) begin
        if(PE_wrapper_204__ap_done) begin
          PE_wrapper_204__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_204__state == 2'b10) begin
        if(PE_wrapper_204__ap_done_global__q0) begin
          PE_wrapper_204__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_204__ap_start = (PE_wrapper_204__state == 2'b01);
  assign PE_wrapper_205__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_205__is_done__q0 = (PE_wrapper_205__state == 2'b10);
  assign PE_wrapper_205__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_205__state <= 2'b00;
    end else begin
      if(PE_wrapper_205__state == 2'b00) begin
        if(PE_wrapper_205__ap_start_global__q0) begin
          PE_wrapper_205__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_205__state == 2'b01) begin
        if(PE_wrapper_205__ap_ready) begin
          if(PE_wrapper_205__ap_done) begin
            PE_wrapper_205__state <= 2'b10;
          end else begin
            PE_wrapper_205__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_205__state == 2'b11) begin
        if(PE_wrapper_205__ap_done) begin
          PE_wrapper_205__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_205__state == 2'b10) begin
        if(PE_wrapper_205__ap_done_global__q0) begin
          PE_wrapper_205__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_205__ap_start = (PE_wrapper_205__state == 2'b01);
  assign PE_wrapper_206__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_206__is_done__q0 = (PE_wrapper_206__state == 2'b10);
  assign PE_wrapper_206__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_206__state <= 2'b00;
    end else begin
      if(PE_wrapper_206__state == 2'b00) begin
        if(PE_wrapper_206__ap_start_global__q0) begin
          PE_wrapper_206__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_206__state == 2'b01) begin
        if(PE_wrapper_206__ap_ready) begin
          if(PE_wrapper_206__ap_done) begin
            PE_wrapper_206__state <= 2'b10;
          end else begin
            PE_wrapper_206__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_206__state == 2'b11) begin
        if(PE_wrapper_206__ap_done) begin
          PE_wrapper_206__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_206__state == 2'b10) begin
        if(PE_wrapper_206__ap_done_global__q0) begin
          PE_wrapper_206__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_206__ap_start = (PE_wrapper_206__state == 2'b01);
  assign PE_wrapper_207__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_207__is_done__q0 = (PE_wrapper_207__state == 2'b10);
  assign PE_wrapper_207__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_207__state <= 2'b00;
    end else begin
      if(PE_wrapper_207__state == 2'b00) begin
        if(PE_wrapper_207__ap_start_global__q0) begin
          PE_wrapper_207__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_207__state == 2'b01) begin
        if(PE_wrapper_207__ap_ready) begin
          if(PE_wrapper_207__ap_done) begin
            PE_wrapper_207__state <= 2'b10;
          end else begin
            PE_wrapper_207__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_207__state == 2'b11) begin
        if(PE_wrapper_207__ap_done) begin
          PE_wrapper_207__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_207__state == 2'b10) begin
        if(PE_wrapper_207__ap_done_global__q0) begin
          PE_wrapper_207__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_207__ap_start = (PE_wrapper_207__state == 2'b01);
  assign PE_wrapper_208__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_208__is_done__q0 = (PE_wrapper_208__state == 2'b10);
  assign PE_wrapper_208__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_208__state <= 2'b00;
    end else begin
      if(PE_wrapper_208__state == 2'b00) begin
        if(PE_wrapper_208__ap_start_global__q0) begin
          PE_wrapper_208__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_208__state == 2'b01) begin
        if(PE_wrapper_208__ap_ready) begin
          if(PE_wrapper_208__ap_done) begin
            PE_wrapper_208__state <= 2'b10;
          end else begin
            PE_wrapper_208__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_208__state == 2'b11) begin
        if(PE_wrapper_208__ap_done) begin
          PE_wrapper_208__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_208__state == 2'b10) begin
        if(PE_wrapper_208__ap_done_global__q0) begin
          PE_wrapper_208__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_208__ap_start = (PE_wrapper_208__state == 2'b01);
  assign PE_wrapper_209__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_209__is_done__q0 = (PE_wrapper_209__state == 2'b10);
  assign PE_wrapper_209__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_209__state <= 2'b00;
    end else begin
      if(PE_wrapper_209__state == 2'b00) begin
        if(PE_wrapper_209__ap_start_global__q0) begin
          PE_wrapper_209__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_209__state == 2'b01) begin
        if(PE_wrapper_209__ap_ready) begin
          if(PE_wrapper_209__ap_done) begin
            PE_wrapper_209__state <= 2'b10;
          end else begin
            PE_wrapper_209__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_209__state == 2'b11) begin
        if(PE_wrapper_209__ap_done) begin
          PE_wrapper_209__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_209__state == 2'b10) begin
        if(PE_wrapper_209__ap_done_global__q0) begin
          PE_wrapper_209__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_209__ap_start = (PE_wrapper_209__state == 2'b01);
  assign PE_wrapper_210__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_210__is_done__q0 = (PE_wrapper_210__state == 2'b10);
  assign PE_wrapper_210__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_210__state <= 2'b00;
    end else begin
      if(PE_wrapper_210__state == 2'b00) begin
        if(PE_wrapper_210__ap_start_global__q0) begin
          PE_wrapper_210__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_210__state == 2'b01) begin
        if(PE_wrapper_210__ap_ready) begin
          if(PE_wrapper_210__ap_done) begin
            PE_wrapper_210__state <= 2'b10;
          end else begin
            PE_wrapper_210__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_210__state == 2'b11) begin
        if(PE_wrapper_210__ap_done) begin
          PE_wrapper_210__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_210__state == 2'b10) begin
        if(PE_wrapper_210__ap_done_global__q0) begin
          PE_wrapper_210__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_210__ap_start = (PE_wrapper_210__state == 2'b01);
  assign PE_wrapper_211__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_211__is_done__q0 = (PE_wrapper_211__state == 2'b10);
  assign PE_wrapper_211__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_211__state <= 2'b00;
    end else begin
      if(PE_wrapper_211__state == 2'b00) begin
        if(PE_wrapper_211__ap_start_global__q0) begin
          PE_wrapper_211__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_211__state == 2'b01) begin
        if(PE_wrapper_211__ap_ready) begin
          if(PE_wrapper_211__ap_done) begin
            PE_wrapper_211__state <= 2'b10;
          end else begin
            PE_wrapper_211__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_211__state == 2'b11) begin
        if(PE_wrapper_211__ap_done) begin
          PE_wrapper_211__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_211__state == 2'b10) begin
        if(PE_wrapper_211__ap_done_global__q0) begin
          PE_wrapper_211__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_211__ap_start = (PE_wrapper_211__state == 2'b01);
  assign PE_wrapper_212__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_212__is_done__q0 = (PE_wrapper_212__state == 2'b10);
  assign PE_wrapper_212__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_212__state <= 2'b00;
    end else begin
      if(PE_wrapper_212__state == 2'b00) begin
        if(PE_wrapper_212__ap_start_global__q0) begin
          PE_wrapper_212__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_212__state == 2'b01) begin
        if(PE_wrapper_212__ap_ready) begin
          if(PE_wrapper_212__ap_done) begin
            PE_wrapper_212__state <= 2'b10;
          end else begin
            PE_wrapper_212__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_212__state == 2'b11) begin
        if(PE_wrapper_212__ap_done) begin
          PE_wrapper_212__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_212__state == 2'b10) begin
        if(PE_wrapper_212__ap_done_global__q0) begin
          PE_wrapper_212__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_212__ap_start = (PE_wrapper_212__state == 2'b01);
  assign PE_wrapper_213__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_213__is_done__q0 = (PE_wrapper_213__state == 2'b10);
  assign PE_wrapper_213__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_213__state <= 2'b00;
    end else begin
      if(PE_wrapper_213__state == 2'b00) begin
        if(PE_wrapper_213__ap_start_global__q0) begin
          PE_wrapper_213__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_213__state == 2'b01) begin
        if(PE_wrapper_213__ap_ready) begin
          if(PE_wrapper_213__ap_done) begin
            PE_wrapper_213__state <= 2'b10;
          end else begin
            PE_wrapper_213__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_213__state == 2'b11) begin
        if(PE_wrapper_213__ap_done) begin
          PE_wrapper_213__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_213__state == 2'b10) begin
        if(PE_wrapper_213__ap_done_global__q0) begin
          PE_wrapper_213__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_213__ap_start = (PE_wrapper_213__state == 2'b01);
  assign PE_wrapper_214__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_214__is_done__q0 = (PE_wrapper_214__state == 2'b10);
  assign PE_wrapper_214__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_214__state <= 2'b00;
    end else begin
      if(PE_wrapper_214__state == 2'b00) begin
        if(PE_wrapper_214__ap_start_global__q0) begin
          PE_wrapper_214__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_214__state == 2'b01) begin
        if(PE_wrapper_214__ap_ready) begin
          if(PE_wrapper_214__ap_done) begin
            PE_wrapper_214__state <= 2'b10;
          end else begin
            PE_wrapper_214__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_214__state == 2'b11) begin
        if(PE_wrapper_214__ap_done) begin
          PE_wrapper_214__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_214__state == 2'b10) begin
        if(PE_wrapper_214__ap_done_global__q0) begin
          PE_wrapper_214__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_214__ap_start = (PE_wrapper_214__state == 2'b01);
  assign PE_wrapper_215__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_215__is_done__q0 = (PE_wrapper_215__state == 2'b10);
  assign PE_wrapper_215__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_215__state <= 2'b00;
    end else begin
      if(PE_wrapper_215__state == 2'b00) begin
        if(PE_wrapper_215__ap_start_global__q0) begin
          PE_wrapper_215__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_215__state == 2'b01) begin
        if(PE_wrapper_215__ap_ready) begin
          if(PE_wrapper_215__ap_done) begin
            PE_wrapper_215__state <= 2'b10;
          end else begin
            PE_wrapper_215__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_215__state == 2'b11) begin
        if(PE_wrapper_215__ap_done) begin
          PE_wrapper_215__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_215__state == 2'b10) begin
        if(PE_wrapper_215__ap_done_global__q0) begin
          PE_wrapper_215__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_215__ap_start = (PE_wrapper_215__state == 2'b01);
  assign PE_wrapper_216__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_216__is_done__q0 = (PE_wrapper_216__state == 2'b10);
  assign PE_wrapper_216__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_216__state <= 2'b00;
    end else begin
      if(PE_wrapper_216__state == 2'b00) begin
        if(PE_wrapper_216__ap_start_global__q0) begin
          PE_wrapper_216__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_216__state == 2'b01) begin
        if(PE_wrapper_216__ap_ready) begin
          if(PE_wrapper_216__ap_done) begin
            PE_wrapper_216__state <= 2'b10;
          end else begin
            PE_wrapper_216__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_216__state == 2'b11) begin
        if(PE_wrapper_216__ap_done) begin
          PE_wrapper_216__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_216__state == 2'b10) begin
        if(PE_wrapper_216__ap_done_global__q0) begin
          PE_wrapper_216__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_216__ap_start = (PE_wrapper_216__state == 2'b01);
  assign PE_wrapper_217__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_217__is_done__q0 = (PE_wrapper_217__state == 2'b10);
  assign PE_wrapper_217__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_217__state <= 2'b00;
    end else begin
      if(PE_wrapper_217__state == 2'b00) begin
        if(PE_wrapper_217__ap_start_global__q0) begin
          PE_wrapper_217__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_217__state == 2'b01) begin
        if(PE_wrapper_217__ap_ready) begin
          if(PE_wrapper_217__ap_done) begin
            PE_wrapper_217__state <= 2'b10;
          end else begin
            PE_wrapper_217__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_217__state == 2'b11) begin
        if(PE_wrapper_217__ap_done) begin
          PE_wrapper_217__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_217__state == 2'b10) begin
        if(PE_wrapper_217__ap_done_global__q0) begin
          PE_wrapper_217__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_217__ap_start = (PE_wrapper_217__state == 2'b01);
  assign PE_wrapper_218__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_218__is_done__q0 = (PE_wrapper_218__state == 2'b10);
  assign PE_wrapper_218__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_218__state <= 2'b00;
    end else begin
      if(PE_wrapper_218__state == 2'b00) begin
        if(PE_wrapper_218__ap_start_global__q0) begin
          PE_wrapper_218__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_218__state == 2'b01) begin
        if(PE_wrapper_218__ap_ready) begin
          if(PE_wrapper_218__ap_done) begin
            PE_wrapper_218__state <= 2'b10;
          end else begin
            PE_wrapper_218__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_218__state == 2'b11) begin
        if(PE_wrapper_218__ap_done) begin
          PE_wrapper_218__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_218__state == 2'b10) begin
        if(PE_wrapper_218__ap_done_global__q0) begin
          PE_wrapper_218__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_218__ap_start = (PE_wrapper_218__state == 2'b01);
  assign PE_wrapper_219__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_219__is_done__q0 = (PE_wrapper_219__state == 2'b10);
  assign PE_wrapper_219__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_219__state <= 2'b00;
    end else begin
      if(PE_wrapper_219__state == 2'b00) begin
        if(PE_wrapper_219__ap_start_global__q0) begin
          PE_wrapper_219__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_219__state == 2'b01) begin
        if(PE_wrapper_219__ap_ready) begin
          if(PE_wrapper_219__ap_done) begin
            PE_wrapper_219__state <= 2'b10;
          end else begin
            PE_wrapper_219__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_219__state == 2'b11) begin
        if(PE_wrapper_219__ap_done) begin
          PE_wrapper_219__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_219__state == 2'b10) begin
        if(PE_wrapper_219__ap_done_global__q0) begin
          PE_wrapper_219__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_219__ap_start = (PE_wrapper_219__state == 2'b01);
  assign PE_wrapper_220__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_220__is_done__q0 = (PE_wrapper_220__state == 2'b10);
  assign PE_wrapper_220__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_220__state <= 2'b00;
    end else begin
      if(PE_wrapper_220__state == 2'b00) begin
        if(PE_wrapper_220__ap_start_global__q0) begin
          PE_wrapper_220__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_220__state == 2'b01) begin
        if(PE_wrapper_220__ap_ready) begin
          if(PE_wrapper_220__ap_done) begin
            PE_wrapper_220__state <= 2'b10;
          end else begin
            PE_wrapper_220__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_220__state == 2'b11) begin
        if(PE_wrapper_220__ap_done) begin
          PE_wrapper_220__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_220__state == 2'b10) begin
        if(PE_wrapper_220__ap_done_global__q0) begin
          PE_wrapper_220__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_220__ap_start = (PE_wrapper_220__state == 2'b01);
  assign PE_wrapper_221__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_221__is_done__q0 = (PE_wrapper_221__state == 2'b10);
  assign PE_wrapper_221__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_221__state <= 2'b00;
    end else begin
      if(PE_wrapper_221__state == 2'b00) begin
        if(PE_wrapper_221__ap_start_global__q0) begin
          PE_wrapper_221__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_221__state == 2'b01) begin
        if(PE_wrapper_221__ap_ready) begin
          if(PE_wrapper_221__ap_done) begin
            PE_wrapper_221__state <= 2'b10;
          end else begin
            PE_wrapper_221__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_221__state == 2'b11) begin
        if(PE_wrapper_221__ap_done) begin
          PE_wrapper_221__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_221__state == 2'b10) begin
        if(PE_wrapper_221__ap_done_global__q0) begin
          PE_wrapper_221__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_221__ap_start = (PE_wrapper_221__state == 2'b01);
  assign PE_wrapper_222__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_222__is_done__q0 = (PE_wrapper_222__state == 2'b10);
  assign PE_wrapper_222__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_222__state <= 2'b00;
    end else begin
      if(PE_wrapper_222__state == 2'b00) begin
        if(PE_wrapper_222__ap_start_global__q0) begin
          PE_wrapper_222__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_222__state == 2'b01) begin
        if(PE_wrapper_222__ap_ready) begin
          if(PE_wrapper_222__ap_done) begin
            PE_wrapper_222__state <= 2'b10;
          end else begin
            PE_wrapper_222__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_222__state == 2'b11) begin
        if(PE_wrapper_222__ap_done) begin
          PE_wrapper_222__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_222__state == 2'b10) begin
        if(PE_wrapper_222__ap_done_global__q0) begin
          PE_wrapper_222__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_222__ap_start = (PE_wrapper_222__state == 2'b01);
  assign PE_wrapper_223__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_223__is_done__q0 = (PE_wrapper_223__state == 2'b10);
  assign PE_wrapper_223__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_223__state <= 2'b00;
    end else begin
      if(PE_wrapper_223__state == 2'b00) begin
        if(PE_wrapper_223__ap_start_global__q0) begin
          PE_wrapper_223__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_223__state == 2'b01) begin
        if(PE_wrapper_223__ap_ready) begin
          if(PE_wrapper_223__ap_done) begin
            PE_wrapper_223__state <= 2'b10;
          end else begin
            PE_wrapper_223__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_223__state == 2'b11) begin
        if(PE_wrapper_223__ap_done) begin
          PE_wrapper_223__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_223__state == 2'b10) begin
        if(PE_wrapper_223__ap_done_global__q0) begin
          PE_wrapper_223__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_223__ap_start = (PE_wrapper_223__state == 2'b01);
  assign PE_wrapper_224__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_224__is_done__q0 = (PE_wrapper_224__state == 2'b10);
  assign PE_wrapper_224__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_224__state <= 2'b00;
    end else begin
      if(PE_wrapper_224__state == 2'b00) begin
        if(PE_wrapper_224__ap_start_global__q0) begin
          PE_wrapper_224__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_224__state == 2'b01) begin
        if(PE_wrapper_224__ap_ready) begin
          if(PE_wrapper_224__ap_done) begin
            PE_wrapper_224__state <= 2'b10;
          end else begin
            PE_wrapper_224__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_224__state == 2'b11) begin
        if(PE_wrapper_224__ap_done) begin
          PE_wrapper_224__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_224__state == 2'b10) begin
        if(PE_wrapper_224__ap_done_global__q0) begin
          PE_wrapper_224__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_224__ap_start = (PE_wrapper_224__state == 2'b01);
  assign PE_wrapper_225__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_225__is_done__q0 = (PE_wrapper_225__state == 2'b10);
  assign PE_wrapper_225__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_225__state <= 2'b00;
    end else begin
      if(PE_wrapper_225__state == 2'b00) begin
        if(PE_wrapper_225__ap_start_global__q0) begin
          PE_wrapper_225__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_225__state == 2'b01) begin
        if(PE_wrapper_225__ap_ready) begin
          if(PE_wrapper_225__ap_done) begin
            PE_wrapper_225__state <= 2'b10;
          end else begin
            PE_wrapper_225__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_225__state == 2'b11) begin
        if(PE_wrapper_225__ap_done) begin
          PE_wrapper_225__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_225__state == 2'b10) begin
        if(PE_wrapper_225__ap_done_global__q0) begin
          PE_wrapper_225__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_225__ap_start = (PE_wrapper_225__state == 2'b01);
  assign PE_wrapper_226__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_226__is_done__q0 = (PE_wrapper_226__state == 2'b10);
  assign PE_wrapper_226__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_226__state <= 2'b00;
    end else begin
      if(PE_wrapper_226__state == 2'b00) begin
        if(PE_wrapper_226__ap_start_global__q0) begin
          PE_wrapper_226__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_226__state == 2'b01) begin
        if(PE_wrapper_226__ap_ready) begin
          if(PE_wrapper_226__ap_done) begin
            PE_wrapper_226__state <= 2'b10;
          end else begin
            PE_wrapper_226__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_226__state == 2'b11) begin
        if(PE_wrapper_226__ap_done) begin
          PE_wrapper_226__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_226__state == 2'b10) begin
        if(PE_wrapper_226__ap_done_global__q0) begin
          PE_wrapper_226__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_226__ap_start = (PE_wrapper_226__state == 2'b01);
  assign PE_wrapper_227__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_227__is_done__q0 = (PE_wrapper_227__state == 2'b10);
  assign PE_wrapper_227__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_227__state <= 2'b00;
    end else begin
      if(PE_wrapper_227__state == 2'b00) begin
        if(PE_wrapper_227__ap_start_global__q0) begin
          PE_wrapper_227__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_227__state == 2'b01) begin
        if(PE_wrapper_227__ap_ready) begin
          if(PE_wrapper_227__ap_done) begin
            PE_wrapper_227__state <= 2'b10;
          end else begin
            PE_wrapper_227__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_227__state == 2'b11) begin
        if(PE_wrapper_227__ap_done) begin
          PE_wrapper_227__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_227__state == 2'b10) begin
        if(PE_wrapper_227__ap_done_global__q0) begin
          PE_wrapper_227__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_227__ap_start = (PE_wrapper_227__state == 2'b01);
  assign PE_wrapper_228__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_228__is_done__q0 = (PE_wrapper_228__state == 2'b10);
  assign PE_wrapper_228__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_228__state <= 2'b00;
    end else begin
      if(PE_wrapper_228__state == 2'b00) begin
        if(PE_wrapper_228__ap_start_global__q0) begin
          PE_wrapper_228__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_228__state == 2'b01) begin
        if(PE_wrapper_228__ap_ready) begin
          if(PE_wrapper_228__ap_done) begin
            PE_wrapper_228__state <= 2'b10;
          end else begin
            PE_wrapper_228__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_228__state == 2'b11) begin
        if(PE_wrapper_228__ap_done) begin
          PE_wrapper_228__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_228__state == 2'b10) begin
        if(PE_wrapper_228__ap_done_global__q0) begin
          PE_wrapper_228__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_228__ap_start = (PE_wrapper_228__state == 2'b01);
  assign PE_wrapper_229__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_229__is_done__q0 = (PE_wrapper_229__state == 2'b10);
  assign PE_wrapper_229__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_229__state <= 2'b00;
    end else begin
      if(PE_wrapper_229__state == 2'b00) begin
        if(PE_wrapper_229__ap_start_global__q0) begin
          PE_wrapper_229__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_229__state == 2'b01) begin
        if(PE_wrapper_229__ap_ready) begin
          if(PE_wrapper_229__ap_done) begin
            PE_wrapper_229__state <= 2'b10;
          end else begin
            PE_wrapper_229__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_229__state == 2'b11) begin
        if(PE_wrapper_229__ap_done) begin
          PE_wrapper_229__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_229__state == 2'b10) begin
        if(PE_wrapper_229__ap_done_global__q0) begin
          PE_wrapper_229__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_229__ap_start = (PE_wrapper_229__state == 2'b01);
  assign PE_wrapper_230__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_230__is_done__q0 = (PE_wrapper_230__state == 2'b10);
  assign PE_wrapper_230__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_230__state <= 2'b00;
    end else begin
      if(PE_wrapper_230__state == 2'b00) begin
        if(PE_wrapper_230__ap_start_global__q0) begin
          PE_wrapper_230__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_230__state == 2'b01) begin
        if(PE_wrapper_230__ap_ready) begin
          if(PE_wrapper_230__ap_done) begin
            PE_wrapper_230__state <= 2'b10;
          end else begin
            PE_wrapper_230__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_230__state == 2'b11) begin
        if(PE_wrapper_230__ap_done) begin
          PE_wrapper_230__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_230__state == 2'b10) begin
        if(PE_wrapper_230__ap_done_global__q0) begin
          PE_wrapper_230__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_230__ap_start = (PE_wrapper_230__state == 2'b01);
  assign PE_wrapper_231__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_231__is_done__q0 = (PE_wrapper_231__state == 2'b10);
  assign PE_wrapper_231__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_231__state <= 2'b00;
    end else begin
      if(PE_wrapper_231__state == 2'b00) begin
        if(PE_wrapper_231__ap_start_global__q0) begin
          PE_wrapper_231__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_231__state == 2'b01) begin
        if(PE_wrapper_231__ap_ready) begin
          if(PE_wrapper_231__ap_done) begin
            PE_wrapper_231__state <= 2'b10;
          end else begin
            PE_wrapper_231__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_231__state == 2'b11) begin
        if(PE_wrapper_231__ap_done) begin
          PE_wrapper_231__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_231__state == 2'b10) begin
        if(PE_wrapper_231__ap_done_global__q0) begin
          PE_wrapper_231__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_231__ap_start = (PE_wrapper_231__state == 2'b01);
  assign PE_wrapper_232__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_232__is_done__q0 = (PE_wrapper_232__state == 2'b10);
  assign PE_wrapper_232__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_232__state <= 2'b00;
    end else begin
      if(PE_wrapper_232__state == 2'b00) begin
        if(PE_wrapper_232__ap_start_global__q0) begin
          PE_wrapper_232__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_232__state == 2'b01) begin
        if(PE_wrapper_232__ap_ready) begin
          if(PE_wrapper_232__ap_done) begin
            PE_wrapper_232__state <= 2'b10;
          end else begin
            PE_wrapper_232__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_232__state == 2'b11) begin
        if(PE_wrapper_232__ap_done) begin
          PE_wrapper_232__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_232__state == 2'b10) begin
        if(PE_wrapper_232__ap_done_global__q0) begin
          PE_wrapper_232__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_232__ap_start = (PE_wrapper_232__state == 2'b01);
  assign PE_wrapper_233__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_233__is_done__q0 = (PE_wrapper_233__state == 2'b10);
  assign PE_wrapper_233__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_233__state <= 2'b00;
    end else begin
      if(PE_wrapper_233__state == 2'b00) begin
        if(PE_wrapper_233__ap_start_global__q0) begin
          PE_wrapper_233__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_233__state == 2'b01) begin
        if(PE_wrapper_233__ap_ready) begin
          if(PE_wrapper_233__ap_done) begin
            PE_wrapper_233__state <= 2'b10;
          end else begin
            PE_wrapper_233__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_233__state == 2'b11) begin
        if(PE_wrapper_233__ap_done) begin
          PE_wrapper_233__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_233__state == 2'b10) begin
        if(PE_wrapper_233__ap_done_global__q0) begin
          PE_wrapper_233__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_233__ap_start = (PE_wrapper_233__state == 2'b01);
  assign PE_wrapper_234__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_234__is_done__q0 = (PE_wrapper_234__state == 2'b10);
  assign PE_wrapper_234__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_234__state <= 2'b00;
    end else begin
      if(PE_wrapper_234__state == 2'b00) begin
        if(PE_wrapper_234__ap_start_global__q0) begin
          PE_wrapper_234__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_234__state == 2'b01) begin
        if(PE_wrapper_234__ap_ready) begin
          if(PE_wrapper_234__ap_done) begin
            PE_wrapper_234__state <= 2'b10;
          end else begin
            PE_wrapper_234__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_234__state == 2'b11) begin
        if(PE_wrapper_234__ap_done) begin
          PE_wrapper_234__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_234__state == 2'b10) begin
        if(PE_wrapper_234__ap_done_global__q0) begin
          PE_wrapper_234__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_234__ap_start = (PE_wrapper_234__state == 2'b01);
  assign PE_wrapper_235__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_235__is_done__q0 = (PE_wrapper_235__state == 2'b10);
  assign PE_wrapper_235__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_235__state <= 2'b00;
    end else begin
      if(PE_wrapper_235__state == 2'b00) begin
        if(PE_wrapper_235__ap_start_global__q0) begin
          PE_wrapper_235__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_235__state == 2'b01) begin
        if(PE_wrapper_235__ap_ready) begin
          if(PE_wrapper_235__ap_done) begin
            PE_wrapper_235__state <= 2'b10;
          end else begin
            PE_wrapper_235__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_235__state == 2'b11) begin
        if(PE_wrapper_235__ap_done) begin
          PE_wrapper_235__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_235__state == 2'b10) begin
        if(PE_wrapper_235__ap_done_global__q0) begin
          PE_wrapper_235__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_235__ap_start = (PE_wrapper_235__state == 2'b01);
  assign PE_wrapper_236__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_236__is_done__q0 = (PE_wrapper_236__state == 2'b10);
  assign PE_wrapper_236__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_236__state <= 2'b00;
    end else begin
      if(PE_wrapper_236__state == 2'b00) begin
        if(PE_wrapper_236__ap_start_global__q0) begin
          PE_wrapper_236__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_236__state == 2'b01) begin
        if(PE_wrapper_236__ap_ready) begin
          if(PE_wrapper_236__ap_done) begin
            PE_wrapper_236__state <= 2'b10;
          end else begin
            PE_wrapper_236__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_236__state == 2'b11) begin
        if(PE_wrapper_236__ap_done) begin
          PE_wrapper_236__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_236__state == 2'b10) begin
        if(PE_wrapper_236__ap_done_global__q0) begin
          PE_wrapper_236__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_236__ap_start = (PE_wrapper_236__state == 2'b01);
  assign PE_wrapper_237__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_237__is_done__q0 = (PE_wrapper_237__state == 2'b10);
  assign PE_wrapper_237__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_237__state <= 2'b00;
    end else begin
      if(PE_wrapper_237__state == 2'b00) begin
        if(PE_wrapper_237__ap_start_global__q0) begin
          PE_wrapper_237__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_237__state == 2'b01) begin
        if(PE_wrapper_237__ap_ready) begin
          if(PE_wrapper_237__ap_done) begin
            PE_wrapper_237__state <= 2'b10;
          end else begin
            PE_wrapper_237__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_237__state == 2'b11) begin
        if(PE_wrapper_237__ap_done) begin
          PE_wrapper_237__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_237__state == 2'b10) begin
        if(PE_wrapper_237__ap_done_global__q0) begin
          PE_wrapper_237__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_237__ap_start = (PE_wrapper_237__state == 2'b01);
  assign PE_wrapper_238__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_238__is_done__q0 = (PE_wrapper_238__state == 2'b10);
  assign PE_wrapper_238__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_238__state <= 2'b00;
    end else begin
      if(PE_wrapper_238__state == 2'b00) begin
        if(PE_wrapper_238__ap_start_global__q0) begin
          PE_wrapper_238__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_238__state == 2'b01) begin
        if(PE_wrapper_238__ap_ready) begin
          if(PE_wrapper_238__ap_done) begin
            PE_wrapper_238__state <= 2'b10;
          end else begin
            PE_wrapper_238__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_238__state == 2'b11) begin
        if(PE_wrapper_238__ap_done) begin
          PE_wrapper_238__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_238__state == 2'b10) begin
        if(PE_wrapper_238__ap_done_global__q0) begin
          PE_wrapper_238__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_238__ap_start = (PE_wrapper_238__state == 2'b01);
  assign PE_wrapper_239__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_239__is_done__q0 = (PE_wrapper_239__state == 2'b10);
  assign PE_wrapper_239__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_239__state <= 2'b00;
    end else begin
      if(PE_wrapper_239__state == 2'b00) begin
        if(PE_wrapper_239__ap_start_global__q0) begin
          PE_wrapper_239__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_239__state == 2'b01) begin
        if(PE_wrapper_239__ap_ready) begin
          if(PE_wrapper_239__ap_done) begin
            PE_wrapper_239__state <= 2'b10;
          end else begin
            PE_wrapper_239__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_239__state == 2'b11) begin
        if(PE_wrapper_239__ap_done) begin
          PE_wrapper_239__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_239__state == 2'b10) begin
        if(PE_wrapper_239__ap_done_global__q0) begin
          PE_wrapper_239__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_239__ap_start = (PE_wrapper_239__state == 2'b01);
  assign PE_wrapper_240__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_240__is_done__q0 = (PE_wrapper_240__state == 2'b10);
  assign PE_wrapper_240__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_240__state <= 2'b00;
    end else begin
      if(PE_wrapper_240__state == 2'b00) begin
        if(PE_wrapper_240__ap_start_global__q0) begin
          PE_wrapper_240__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_240__state == 2'b01) begin
        if(PE_wrapper_240__ap_ready) begin
          if(PE_wrapper_240__ap_done) begin
            PE_wrapper_240__state <= 2'b10;
          end else begin
            PE_wrapper_240__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_240__state == 2'b11) begin
        if(PE_wrapper_240__ap_done) begin
          PE_wrapper_240__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_240__state == 2'b10) begin
        if(PE_wrapper_240__ap_done_global__q0) begin
          PE_wrapper_240__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_240__ap_start = (PE_wrapper_240__state == 2'b01);
  assign PE_wrapper_241__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_241__is_done__q0 = (PE_wrapper_241__state == 2'b10);
  assign PE_wrapper_241__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_241__state <= 2'b00;
    end else begin
      if(PE_wrapper_241__state == 2'b00) begin
        if(PE_wrapper_241__ap_start_global__q0) begin
          PE_wrapper_241__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_241__state == 2'b01) begin
        if(PE_wrapper_241__ap_ready) begin
          if(PE_wrapper_241__ap_done) begin
            PE_wrapper_241__state <= 2'b10;
          end else begin
            PE_wrapper_241__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_241__state == 2'b11) begin
        if(PE_wrapper_241__ap_done) begin
          PE_wrapper_241__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_241__state == 2'b10) begin
        if(PE_wrapper_241__ap_done_global__q0) begin
          PE_wrapper_241__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_241__ap_start = (PE_wrapper_241__state == 2'b01);
  assign PE_wrapper_242__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_242__is_done__q0 = (PE_wrapper_242__state == 2'b10);
  assign PE_wrapper_242__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_242__state <= 2'b00;
    end else begin
      if(PE_wrapper_242__state == 2'b00) begin
        if(PE_wrapper_242__ap_start_global__q0) begin
          PE_wrapper_242__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_242__state == 2'b01) begin
        if(PE_wrapper_242__ap_ready) begin
          if(PE_wrapper_242__ap_done) begin
            PE_wrapper_242__state <= 2'b10;
          end else begin
            PE_wrapper_242__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_242__state == 2'b11) begin
        if(PE_wrapper_242__ap_done) begin
          PE_wrapper_242__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_242__state == 2'b10) begin
        if(PE_wrapper_242__ap_done_global__q0) begin
          PE_wrapper_242__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_242__ap_start = (PE_wrapper_242__state == 2'b01);
  assign PE_wrapper_243__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_243__is_done__q0 = (PE_wrapper_243__state == 2'b10);
  assign PE_wrapper_243__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_243__state <= 2'b00;
    end else begin
      if(PE_wrapper_243__state == 2'b00) begin
        if(PE_wrapper_243__ap_start_global__q0) begin
          PE_wrapper_243__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_243__state == 2'b01) begin
        if(PE_wrapper_243__ap_ready) begin
          if(PE_wrapper_243__ap_done) begin
            PE_wrapper_243__state <= 2'b10;
          end else begin
            PE_wrapper_243__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_243__state == 2'b11) begin
        if(PE_wrapper_243__ap_done) begin
          PE_wrapper_243__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_243__state == 2'b10) begin
        if(PE_wrapper_243__ap_done_global__q0) begin
          PE_wrapper_243__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_243__ap_start = (PE_wrapper_243__state == 2'b01);
  assign PE_wrapper_244__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_244__is_done__q0 = (PE_wrapper_244__state == 2'b10);
  assign PE_wrapper_244__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_244__state <= 2'b00;
    end else begin
      if(PE_wrapper_244__state == 2'b00) begin
        if(PE_wrapper_244__ap_start_global__q0) begin
          PE_wrapper_244__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_244__state == 2'b01) begin
        if(PE_wrapper_244__ap_ready) begin
          if(PE_wrapper_244__ap_done) begin
            PE_wrapper_244__state <= 2'b10;
          end else begin
            PE_wrapper_244__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_244__state == 2'b11) begin
        if(PE_wrapper_244__ap_done) begin
          PE_wrapper_244__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_244__state == 2'b10) begin
        if(PE_wrapper_244__ap_done_global__q0) begin
          PE_wrapper_244__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_244__ap_start = (PE_wrapper_244__state == 2'b01);
  assign PE_wrapper_245__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_245__is_done__q0 = (PE_wrapper_245__state == 2'b10);
  assign PE_wrapper_245__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_245__state <= 2'b00;
    end else begin
      if(PE_wrapper_245__state == 2'b00) begin
        if(PE_wrapper_245__ap_start_global__q0) begin
          PE_wrapper_245__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_245__state == 2'b01) begin
        if(PE_wrapper_245__ap_ready) begin
          if(PE_wrapper_245__ap_done) begin
            PE_wrapper_245__state <= 2'b10;
          end else begin
            PE_wrapper_245__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_245__state == 2'b11) begin
        if(PE_wrapper_245__ap_done) begin
          PE_wrapper_245__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_245__state == 2'b10) begin
        if(PE_wrapper_245__ap_done_global__q0) begin
          PE_wrapper_245__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_245__ap_start = (PE_wrapper_245__state == 2'b01);
  assign PE_wrapper_246__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_246__is_done__q0 = (PE_wrapper_246__state == 2'b10);
  assign PE_wrapper_246__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_246__state <= 2'b00;
    end else begin
      if(PE_wrapper_246__state == 2'b00) begin
        if(PE_wrapper_246__ap_start_global__q0) begin
          PE_wrapper_246__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_246__state == 2'b01) begin
        if(PE_wrapper_246__ap_ready) begin
          if(PE_wrapper_246__ap_done) begin
            PE_wrapper_246__state <= 2'b10;
          end else begin
            PE_wrapper_246__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_246__state == 2'b11) begin
        if(PE_wrapper_246__ap_done) begin
          PE_wrapper_246__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_246__state == 2'b10) begin
        if(PE_wrapper_246__ap_done_global__q0) begin
          PE_wrapper_246__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_246__ap_start = (PE_wrapper_246__state == 2'b01);
  assign PE_wrapper_247__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_247__is_done__q0 = (PE_wrapper_247__state == 2'b10);
  assign PE_wrapper_247__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_247__state <= 2'b00;
    end else begin
      if(PE_wrapper_247__state == 2'b00) begin
        if(PE_wrapper_247__ap_start_global__q0) begin
          PE_wrapper_247__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_247__state == 2'b01) begin
        if(PE_wrapper_247__ap_ready) begin
          if(PE_wrapper_247__ap_done) begin
            PE_wrapper_247__state <= 2'b10;
          end else begin
            PE_wrapper_247__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_247__state == 2'b11) begin
        if(PE_wrapper_247__ap_done) begin
          PE_wrapper_247__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_247__state == 2'b10) begin
        if(PE_wrapper_247__ap_done_global__q0) begin
          PE_wrapper_247__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_247__ap_start = (PE_wrapper_247__state == 2'b01);
  assign PE_wrapper_248__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_248__is_done__q0 = (PE_wrapper_248__state == 2'b10);
  assign PE_wrapper_248__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_248__state <= 2'b00;
    end else begin
      if(PE_wrapper_248__state == 2'b00) begin
        if(PE_wrapper_248__ap_start_global__q0) begin
          PE_wrapper_248__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_248__state == 2'b01) begin
        if(PE_wrapper_248__ap_ready) begin
          if(PE_wrapper_248__ap_done) begin
            PE_wrapper_248__state <= 2'b10;
          end else begin
            PE_wrapper_248__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_248__state == 2'b11) begin
        if(PE_wrapper_248__ap_done) begin
          PE_wrapper_248__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_248__state == 2'b10) begin
        if(PE_wrapper_248__ap_done_global__q0) begin
          PE_wrapper_248__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_248__ap_start = (PE_wrapper_248__state == 2'b01);
  assign PE_wrapper_249__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_249__is_done__q0 = (PE_wrapper_249__state == 2'b10);
  assign PE_wrapper_249__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_249__state <= 2'b00;
    end else begin
      if(PE_wrapper_249__state == 2'b00) begin
        if(PE_wrapper_249__ap_start_global__q0) begin
          PE_wrapper_249__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_249__state == 2'b01) begin
        if(PE_wrapper_249__ap_ready) begin
          if(PE_wrapper_249__ap_done) begin
            PE_wrapper_249__state <= 2'b10;
          end else begin
            PE_wrapper_249__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_249__state == 2'b11) begin
        if(PE_wrapper_249__ap_done) begin
          PE_wrapper_249__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_249__state == 2'b10) begin
        if(PE_wrapper_249__ap_done_global__q0) begin
          PE_wrapper_249__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_249__ap_start = (PE_wrapper_249__state == 2'b01);
  assign PE_wrapper_250__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_250__is_done__q0 = (PE_wrapper_250__state == 2'b10);
  assign PE_wrapper_250__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_250__state <= 2'b00;
    end else begin
      if(PE_wrapper_250__state == 2'b00) begin
        if(PE_wrapper_250__ap_start_global__q0) begin
          PE_wrapper_250__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_250__state == 2'b01) begin
        if(PE_wrapper_250__ap_ready) begin
          if(PE_wrapper_250__ap_done) begin
            PE_wrapper_250__state <= 2'b10;
          end else begin
            PE_wrapper_250__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_250__state == 2'b11) begin
        if(PE_wrapper_250__ap_done) begin
          PE_wrapper_250__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_250__state == 2'b10) begin
        if(PE_wrapper_250__ap_done_global__q0) begin
          PE_wrapper_250__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_250__ap_start = (PE_wrapper_250__state == 2'b01);
  assign PE_wrapper_251__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_251__is_done__q0 = (PE_wrapper_251__state == 2'b10);
  assign PE_wrapper_251__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_251__state <= 2'b00;
    end else begin
      if(PE_wrapper_251__state == 2'b00) begin
        if(PE_wrapper_251__ap_start_global__q0) begin
          PE_wrapper_251__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_251__state == 2'b01) begin
        if(PE_wrapper_251__ap_ready) begin
          if(PE_wrapper_251__ap_done) begin
            PE_wrapper_251__state <= 2'b10;
          end else begin
            PE_wrapper_251__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_251__state == 2'b11) begin
        if(PE_wrapper_251__ap_done) begin
          PE_wrapper_251__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_251__state == 2'b10) begin
        if(PE_wrapper_251__ap_done_global__q0) begin
          PE_wrapper_251__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_251__ap_start = (PE_wrapper_251__state == 2'b01);
  assign PE_wrapper_252__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_252__is_done__q0 = (PE_wrapper_252__state == 2'b10);
  assign PE_wrapper_252__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_252__state <= 2'b00;
    end else begin
      if(PE_wrapper_252__state == 2'b00) begin
        if(PE_wrapper_252__ap_start_global__q0) begin
          PE_wrapper_252__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_252__state == 2'b01) begin
        if(PE_wrapper_252__ap_ready) begin
          if(PE_wrapper_252__ap_done) begin
            PE_wrapper_252__state <= 2'b10;
          end else begin
            PE_wrapper_252__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_252__state == 2'b11) begin
        if(PE_wrapper_252__ap_done) begin
          PE_wrapper_252__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_252__state == 2'b10) begin
        if(PE_wrapper_252__ap_done_global__q0) begin
          PE_wrapper_252__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_252__ap_start = (PE_wrapper_252__state == 2'b01);
  assign PE_wrapper_253__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_253__is_done__q0 = (PE_wrapper_253__state == 2'b10);
  assign PE_wrapper_253__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_253__state <= 2'b00;
    end else begin
      if(PE_wrapper_253__state == 2'b00) begin
        if(PE_wrapper_253__ap_start_global__q0) begin
          PE_wrapper_253__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_253__state == 2'b01) begin
        if(PE_wrapper_253__ap_ready) begin
          if(PE_wrapper_253__ap_done) begin
            PE_wrapper_253__state <= 2'b10;
          end else begin
            PE_wrapper_253__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_253__state == 2'b11) begin
        if(PE_wrapper_253__ap_done) begin
          PE_wrapper_253__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_253__state == 2'b10) begin
        if(PE_wrapper_253__ap_done_global__q0) begin
          PE_wrapper_253__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_253__ap_start = (PE_wrapper_253__state == 2'b01);
  assign PE_wrapper_254__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_254__is_done__q0 = (PE_wrapper_254__state == 2'b10);
  assign PE_wrapper_254__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_254__state <= 2'b00;
    end else begin
      if(PE_wrapper_254__state == 2'b00) begin
        if(PE_wrapper_254__ap_start_global__q0) begin
          PE_wrapper_254__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_254__state == 2'b01) begin
        if(PE_wrapper_254__ap_ready) begin
          if(PE_wrapper_254__ap_done) begin
            PE_wrapper_254__state <= 2'b10;
          end else begin
            PE_wrapper_254__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_254__state == 2'b11) begin
        if(PE_wrapper_254__ap_done) begin
          PE_wrapper_254__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_254__state == 2'b10) begin
        if(PE_wrapper_254__ap_done_global__q0) begin
          PE_wrapper_254__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_254__ap_start = (PE_wrapper_254__state == 2'b01);
  assign PE_wrapper_255__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_255__is_done__q0 = (PE_wrapper_255__state == 2'b10);
  assign PE_wrapper_255__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_255__state <= 2'b00;
    end else begin
      if(PE_wrapper_255__state == 2'b00) begin
        if(PE_wrapper_255__ap_start_global__q0) begin
          PE_wrapper_255__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_255__state == 2'b01) begin
        if(PE_wrapper_255__ap_ready) begin
          if(PE_wrapper_255__ap_done) begin
            PE_wrapper_255__state <= 2'b10;
          end else begin
            PE_wrapper_255__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_255__state == 2'b11) begin
        if(PE_wrapper_255__ap_done) begin
          PE_wrapper_255__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_255__state == 2'b10) begin
        if(PE_wrapper_255__ap_done_global__q0) begin
          PE_wrapper_255__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_255__ap_start = (PE_wrapper_255__state == 2'b01);
  assign PE_wrapper_256__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_256__is_done__q0 = (PE_wrapper_256__state == 2'b10);
  assign PE_wrapper_256__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_256__state <= 2'b00;
    end else begin
      if(PE_wrapper_256__state == 2'b00) begin
        if(PE_wrapper_256__ap_start_global__q0) begin
          PE_wrapper_256__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_256__state == 2'b01) begin
        if(PE_wrapper_256__ap_ready) begin
          if(PE_wrapper_256__ap_done) begin
            PE_wrapper_256__state <= 2'b10;
          end else begin
            PE_wrapper_256__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_256__state == 2'b11) begin
        if(PE_wrapper_256__ap_done) begin
          PE_wrapper_256__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_256__state == 2'b10) begin
        if(PE_wrapper_256__ap_done_global__q0) begin
          PE_wrapper_256__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_256__ap_start = (PE_wrapper_256__state == 2'b01);
  assign PE_wrapper_257__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_257__is_done__q0 = (PE_wrapper_257__state == 2'b10);
  assign PE_wrapper_257__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_257__state <= 2'b00;
    end else begin
      if(PE_wrapper_257__state == 2'b00) begin
        if(PE_wrapper_257__ap_start_global__q0) begin
          PE_wrapper_257__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_257__state == 2'b01) begin
        if(PE_wrapper_257__ap_ready) begin
          if(PE_wrapper_257__ap_done) begin
            PE_wrapper_257__state <= 2'b10;
          end else begin
            PE_wrapper_257__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_257__state == 2'b11) begin
        if(PE_wrapper_257__ap_done) begin
          PE_wrapper_257__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_257__state == 2'b10) begin
        if(PE_wrapper_257__ap_done_global__q0) begin
          PE_wrapper_257__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_257__ap_start = (PE_wrapper_257__state == 2'b01);
  assign PE_wrapper_258__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_258__is_done__q0 = (PE_wrapper_258__state == 2'b10);
  assign PE_wrapper_258__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_258__state <= 2'b00;
    end else begin
      if(PE_wrapper_258__state == 2'b00) begin
        if(PE_wrapper_258__ap_start_global__q0) begin
          PE_wrapper_258__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_258__state == 2'b01) begin
        if(PE_wrapper_258__ap_ready) begin
          if(PE_wrapper_258__ap_done) begin
            PE_wrapper_258__state <= 2'b10;
          end else begin
            PE_wrapper_258__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_258__state == 2'b11) begin
        if(PE_wrapper_258__ap_done) begin
          PE_wrapper_258__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_258__state == 2'b10) begin
        if(PE_wrapper_258__ap_done_global__q0) begin
          PE_wrapper_258__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_258__ap_start = (PE_wrapper_258__state == 2'b01);
  assign PE_wrapper_259__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_259__is_done__q0 = (PE_wrapper_259__state == 2'b10);
  assign PE_wrapper_259__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_259__state <= 2'b00;
    end else begin
      if(PE_wrapper_259__state == 2'b00) begin
        if(PE_wrapper_259__ap_start_global__q0) begin
          PE_wrapper_259__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_259__state == 2'b01) begin
        if(PE_wrapper_259__ap_ready) begin
          if(PE_wrapper_259__ap_done) begin
            PE_wrapper_259__state <= 2'b10;
          end else begin
            PE_wrapper_259__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_259__state == 2'b11) begin
        if(PE_wrapper_259__ap_done) begin
          PE_wrapper_259__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_259__state == 2'b10) begin
        if(PE_wrapper_259__ap_done_global__q0) begin
          PE_wrapper_259__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_259__ap_start = (PE_wrapper_259__state == 2'b01);
  assign PE_wrapper_260__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_260__is_done__q0 = (PE_wrapper_260__state == 2'b10);
  assign PE_wrapper_260__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_260__state <= 2'b00;
    end else begin
      if(PE_wrapper_260__state == 2'b00) begin
        if(PE_wrapper_260__ap_start_global__q0) begin
          PE_wrapper_260__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_260__state == 2'b01) begin
        if(PE_wrapper_260__ap_ready) begin
          if(PE_wrapper_260__ap_done) begin
            PE_wrapper_260__state <= 2'b10;
          end else begin
            PE_wrapper_260__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_260__state == 2'b11) begin
        if(PE_wrapper_260__ap_done) begin
          PE_wrapper_260__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_260__state == 2'b10) begin
        if(PE_wrapper_260__ap_done_global__q0) begin
          PE_wrapper_260__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_260__ap_start = (PE_wrapper_260__state == 2'b01);
  assign PE_wrapper_261__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_261__is_done__q0 = (PE_wrapper_261__state == 2'b10);
  assign PE_wrapper_261__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_261__state <= 2'b00;
    end else begin
      if(PE_wrapper_261__state == 2'b00) begin
        if(PE_wrapper_261__ap_start_global__q0) begin
          PE_wrapper_261__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_261__state == 2'b01) begin
        if(PE_wrapper_261__ap_ready) begin
          if(PE_wrapper_261__ap_done) begin
            PE_wrapper_261__state <= 2'b10;
          end else begin
            PE_wrapper_261__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_261__state == 2'b11) begin
        if(PE_wrapper_261__ap_done) begin
          PE_wrapper_261__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_261__state == 2'b10) begin
        if(PE_wrapper_261__ap_done_global__q0) begin
          PE_wrapper_261__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_261__ap_start = (PE_wrapper_261__state == 2'b01);
  assign PE_wrapper_262__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_262__is_done__q0 = (PE_wrapper_262__state == 2'b10);
  assign PE_wrapper_262__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_262__state <= 2'b00;
    end else begin
      if(PE_wrapper_262__state == 2'b00) begin
        if(PE_wrapper_262__ap_start_global__q0) begin
          PE_wrapper_262__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_262__state == 2'b01) begin
        if(PE_wrapper_262__ap_ready) begin
          if(PE_wrapper_262__ap_done) begin
            PE_wrapper_262__state <= 2'b10;
          end else begin
            PE_wrapper_262__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_262__state == 2'b11) begin
        if(PE_wrapper_262__ap_done) begin
          PE_wrapper_262__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_262__state == 2'b10) begin
        if(PE_wrapper_262__ap_done_global__q0) begin
          PE_wrapper_262__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_262__ap_start = (PE_wrapper_262__state == 2'b01);
  assign PE_wrapper_263__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_263__is_done__q0 = (PE_wrapper_263__state == 2'b10);
  assign PE_wrapper_263__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_263__state <= 2'b00;
    end else begin
      if(PE_wrapper_263__state == 2'b00) begin
        if(PE_wrapper_263__ap_start_global__q0) begin
          PE_wrapper_263__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_263__state == 2'b01) begin
        if(PE_wrapper_263__ap_ready) begin
          if(PE_wrapper_263__ap_done) begin
            PE_wrapper_263__state <= 2'b10;
          end else begin
            PE_wrapper_263__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_263__state == 2'b11) begin
        if(PE_wrapper_263__ap_done) begin
          PE_wrapper_263__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_263__state == 2'b10) begin
        if(PE_wrapper_263__ap_done_global__q0) begin
          PE_wrapper_263__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_263__ap_start = (PE_wrapper_263__state == 2'b01);
  assign PE_wrapper_264__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_264__is_done__q0 = (PE_wrapper_264__state == 2'b10);
  assign PE_wrapper_264__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_264__state <= 2'b00;
    end else begin
      if(PE_wrapper_264__state == 2'b00) begin
        if(PE_wrapper_264__ap_start_global__q0) begin
          PE_wrapper_264__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_264__state == 2'b01) begin
        if(PE_wrapper_264__ap_ready) begin
          if(PE_wrapper_264__ap_done) begin
            PE_wrapper_264__state <= 2'b10;
          end else begin
            PE_wrapper_264__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_264__state == 2'b11) begin
        if(PE_wrapper_264__ap_done) begin
          PE_wrapper_264__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_264__state == 2'b10) begin
        if(PE_wrapper_264__ap_done_global__q0) begin
          PE_wrapper_264__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_264__ap_start = (PE_wrapper_264__state == 2'b01);
  assign PE_wrapper_265__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_265__is_done__q0 = (PE_wrapper_265__state == 2'b10);
  assign PE_wrapper_265__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_265__state <= 2'b00;
    end else begin
      if(PE_wrapper_265__state == 2'b00) begin
        if(PE_wrapper_265__ap_start_global__q0) begin
          PE_wrapper_265__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_265__state == 2'b01) begin
        if(PE_wrapper_265__ap_ready) begin
          if(PE_wrapper_265__ap_done) begin
            PE_wrapper_265__state <= 2'b10;
          end else begin
            PE_wrapper_265__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_265__state == 2'b11) begin
        if(PE_wrapper_265__ap_done) begin
          PE_wrapper_265__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_265__state == 2'b10) begin
        if(PE_wrapper_265__ap_done_global__q0) begin
          PE_wrapper_265__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_265__ap_start = (PE_wrapper_265__state == 2'b01);
  assign PE_wrapper_266__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_266__is_done__q0 = (PE_wrapper_266__state == 2'b10);
  assign PE_wrapper_266__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_266__state <= 2'b00;
    end else begin
      if(PE_wrapper_266__state == 2'b00) begin
        if(PE_wrapper_266__ap_start_global__q0) begin
          PE_wrapper_266__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_266__state == 2'b01) begin
        if(PE_wrapper_266__ap_ready) begin
          if(PE_wrapper_266__ap_done) begin
            PE_wrapper_266__state <= 2'b10;
          end else begin
            PE_wrapper_266__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_266__state == 2'b11) begin
        if(PE_wrapper_266__ap_done) begin
          PE_wrapper_266__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_266__state == 2'b10) begin
        if(PE_wrapper_266__ap_done_global__q0) begin
          PE_wrapper_266__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_266__ap_start = (PE_wrapper_266__state == 2'b01);
  assign PE_wrapper_267__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_267__is_done__q0 = (PE_wrapper_267__state == 2'b10);
  assign PE_wrapper_267__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_267__state <= 2'b00;
    end else begin
      if(PE_wrapper_267__state == 2'b00) begin
        if(PE_wrapper_267__ap_start_global__q0) begin
          PE_wrapper_267__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_267__state == 2'b01) begin
        if(PE_wrapper_267__ap_ready) begin
          if(PE_wrapper_267__ap_done) begin
            PE_wrapper_267__state <= 2'b10;
          end else begin
            PE_wrapper_267__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_267__state == 2'b11) begin
        if(PE_wrapper_267__ap_done) begin
          PE_wrapper_267__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_267__state == 2'b10) begin
        if(PE_wrapper_267__ap_done_global__q0) begin
          PE_wrapper_267__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_267__ap_start = (PE_wrapper_267__state == 2'b01);
  assign PE_wrapper_268__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_268__is_done__q0 = (PE_wrapper_268__state == 2'b10);
  assign PE_wrapper_268__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_268__state <= 2'b00;
    end else begin
      if(PE_wrapper_268__state == 2'b00) begin
        if(PE_wrapper_268__ap_start_global__q0) begin
          PE_wrapper_268__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_268__state == 2'b01) begin
        if(PE_wrapper_268__ap_ready) begin
          if(PE_wrapper_268__ap_done) begin
            PE_wrapper_268__state <= 2'b10;
          end else begin
            PE_wrapper_268__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_268__state == 2'b11) begin
        if(PE_wrapper_268__ap_done) begin
          PE_wrapper_268__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_268__state == 2'b10) begin
        if(PE_wrapper_268__ap_done_global__q0) begin
          PE_wrapper_268__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_268__ap_start = (PE_wrapper_268__state == 2'b01);
  assign PE_wrapper_269__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_269__is_done__q0 = (PE_wrapper_269__state == 2'b10);
  assign PE_wrapper_269__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_269__state <= 2'b00;
    end else begin
      if(PE_wrapper_269__state == 2'b00) begin
        if(PE_wrapper_269__ap_start_global__q0) begin
          PE_wrapper_269__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_269__state == 2'b01) begin
        if(PE_wrapper_269__ap_ready) begin
          if(PE_wrapper_269__ap_done) begin
            PE_wrapper_269__state <= 2'b10;
          end else begin
            PE_wrapper_269__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_269__state == 2'b11) begin
        if(PE_wrapper_269__ap_done) begin
          PE_wrapper_269__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_269__state == 2'b10) begin
        if(PE_wrapper_269__ap_done_global__q0) begin
          PE_wrapper_269__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_269__ap_start = (PE_wrapper_269__state == 2'b01);
  assign PE_wrapper_270__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_270__is_done__q0 = (PE_wrapper_270__state == 2'b10);
  assign PE_wrapper_270__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_270__state <= 2'b00;
    end else begin
      if(PE_wrapper_270__state == 2'b00) begin
        if(PE_wrapper_270__ap_start_global__q0) begin
          PE_wrapper_270__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_270__state == 2'b01) begin
        if(PE_wrapper_270__ap_ready) begin
          if(PE_wrapper_270__ap_done) begin
            PE_wrapper_270__state <= 2'b10;
          end else begin
            PE_wrapper_270__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_270__state == 2'b11) begin
        if(PE_wrapper_270__ap_done) begin
          PE_wrapper_270__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_270__state == 2'b10) begin
        if(PE_wrapper_270__ap_done_global__q0) begin
          PE_wrapper_270__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_270__ap_start = (PE_wrapper_270__state == 2'b01);
  assign PE_wrapper_271__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_271__is_done__q0 = (PE_wrapper_271__state == 2'b10);
  assign PE_wrapper_271__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_271__state <= 2'b00;
    end else begin
      if(PE_wrapper_271__state == 2'b00) begin
        if(PE_wrapper_271__ap_start_global__q0) begin
          PE_wrapper_271__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_271__state == 2'b01) begin
        if(PE_wrapper_271__ap_ready) begin
          if(PE_wrapper_271__ap_done) begin
            PE_wrapper_271__state <= 2'b10;
          end else begin
            PE_wrapper_271__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_271__state == 2'b11) begin
        if(PE_wrapper_271__ap_done) begin
          PE_wrapper_271__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_271__state == 2'b10) begin
        if(PE_wrapper_271__ap_done_global__q0) begin
          PE_wrapper_271__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_271__ap_start = (PE_wrapper_271__state == 2'b01);
  assign PE_wrapper_272__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_272__is_done__q0 = (PE_wrapper_272__state == 2'b10);
  assign PE_wrapper_272__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_272__state <= 2'b00;
    end else begin
      if(PE_wrapper_272__state == 2'b00) begin
        if(PE_wrapper_272__ap_start_global__q0) begin
          PE_wrapper_272__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_272__state == 2'b01) begin
        if(PE_wrapper_272__ap_ready) begin
          if(PE_wrapper_272__ap_done) begin
            PE_wrapper_272__state <= 2'b10;
          end else begin
            PE_wrapper_272__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_272__state == 2'b11) begin
        if(PE_wrapper_272__ap_done) begin
          PE_wrapper_272__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_272__state == 2'b10) begin
        if(PE_wrapper_272__ap_done_global__q0) begin
          PE_wrapper_272__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_272__ap_start = (PE_wrapper_272__state == 2'b01);
  assign PE_wrapper_273__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_273__is_done__q0 = (PE_wrapper_273__state == 2'b10);
  assign PE_wrapper_273__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_273__state <= 2'b00;
    end else begin
      if(PE_wrapper_273__state == 2'b00) begin
        if(PE_wrapper_273__ap_start_global__q0) begin
          PE_wrapper_273__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_273__state == 2'b01) begin
        if(PE_wrapper_273__ap_ready) begin
          if(PE_wrapper_273__ap_done) begin
            PE_wrapper_273__state <= 2'b10;
          end else begin
            PE_wrapper_273__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_273__state == 2'b11) begin
        if(PE_wrapper_273__ap_done) begin
          PE_wrapper_273__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_273__state == 2'b10) begin
        if(PE_wrapper_273__ap_done_global__q0) begin
          PE_wrapper_273__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_273__ap_start = (PE_wrapper_273__state == 2'b01);
  assign PE_wrapper_274__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_274__is_done__q0 = (PE_wrapper_274__state == 2'b10);
  assign PE_wrapper_274__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_274__state <= 2'b00;
    end else begin
      if(PE_wrapper_274__state == 2'b00) begin
        if(PE_wrapper_274__ap_start_global__q0) begin
          PE_wrapper_274__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_274__state == 2'b01) begin
        if(PE_wrapper_274__ap_ready) begin
          if(PE_wrapper_274__ap_done) begin
            PE_wrapper_274__state <= 2'b10;
          end else begin
            PE_wrapper_274__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_274__state == 2'b11) begin
        if(PE_wrapper_274__ap_done) begin
          PE_wrapper_274__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_274__state == 2'b10) begin
        if(PE_wrapper_274__ap_done_global__q0) begin
          PE_wrapper_274__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_274__ap_start = (PE_wrapper_274__state == 2'b01);
  assign PE_wrapper_275__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_275__is_done__q0 = (PE_wrapper_275__state == 2'b10);
  assign PE_wrapper_275__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_275__state <= 2'b00;
    end else begin
      if(PE_wrapper_275__state == 2'b00) begin
        if(PE_wrapper_275__ap_start_global__q0) begin
          PE_wrapper_275__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_275__state == 2'b01) begin
        if(PE_wrapper_275__ap_ready) begin
          if(PE_wrapper_275__ap_done) begin
            PE_wrapper_275__state <= 2'b10;
          end else begin
            PE_wrapper_275__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_275__state == 2'b11) begin
        if(PE_wrapper_275__ap_done) begin
          PE_wrapper_275__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_275__state == 2'b10) begin
        if(PE_wrapper_275__ap_done_global__q0) begin
          PE_wrapper_275__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_275__ap_start = (PE_wrapper_275__state == 2'b01);
  assign PE_wrapper_276__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_276__is_done__q0 = (PE_wrapper_276__state == 2'b10);
  assign PE_wrapper_276__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_276__state <= 2'b00;
    end else begin
      if(PE_wrapper_276__state == 2'b00) begin
        if(PE_wrapper_276__ap_start_global__q0) begin
          PE_wrapper_276__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_276__state == 2'b01) begin
        if(PE_wrapper_276__ap_ready) begin
          if(PE_wrapper_276__ap_done) begin
            PE_wrapper_276__state <= 2'b10;
          end else begin
            PE_wrapper_276__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_276__state == 2'b11) begin
        if(PE_wrapper_276__ap_done) begin
          PE_wrapper_276__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_276__state == 2'b10) begin
        if(PE_wrapper_276__ap_done_global__q0) begin
          PE_wrapper_276__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_276__ap_start = (PE_wrapper_276__state == 2'b01);
  assign PE_wrapper_277__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_277__is_done__q0 = (PE_wrapper_277__state == 2'b10);
  assign PE_wrapper_277__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_277__state <= 2'b00;
    end else begin
      if(PE_wrapper_277__state == 2'b00) begin
        if(PE_wrapper_277__ap_start_global__q0) begin
          PE_wrapper_277__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_277__state == 2'b01) begin
        if(PE_wrapper_277__ap_ready) begin
          if(PE_wrapper_277__ap_done) begin
            PE_wrapper_277__state <= 2'b10;
          end else begin
            PE_wrapper_277__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_277__state == 2'b11) begin
        if(PE_wrapper_277__ap_done) begin
          PE_wrapper_277__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_277__state == 2'b10) begin
        if(PE_wrapper_277__ap_done_global__q0) begin
          PE_wrapper_277__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_277__ap_start = (PE_wrapper_277__state == 2'b01);
  assign PE_wrapper_278__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_278__is_done__q0 = (PE_wrapper_278__state == 2'b10);
  assign PE_wrapper_278__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_278__state <= 2'b00;
    end else begin
      if(PE_wrapper_278__state == 2'b00) begin
        if(PE_wrapper_278__ap_start_global__q0) begin
          PE_wrapper_278__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_278__state == 2'b01) begin
        if(PE_wrapper_278__ap_ready) begin
          if(PE_wrapper_278__ap_done) begin
            PE_wrapper_278__state <= 2'b10;
          end else begin
            PE_wrapper_278__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_278__state == 2'b11) begin
        if(PE_wrapper_278__ap_done) begin
          PE_wrapper_278__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_278__state == 2'b10) begin
        if(PE_wrapper_278__ap_done_global__q0) begin
          PE_wrapper_278__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_278__ap_start = (PE_wrapper_278__state == 2'b01);
  assign PE_wrapper_279__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_279__is_done__q0 = (PE_wrapper_279__state == 2'b10);
  assign PE_wrapper_279__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_279__state <= 2'b00;
    end else begin
      if(PE_wrapper_279__state == 2'b00) begin
        if(PE_wrapper_279__ap_start_global__q0) begin
          PE_wrapper_279__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_279__state == 2'b01) begin
        if(PE_wrapper_279__ap_ready) begin
          if(PE_wrapper_279__ap_done) begin
            PE_wrapper_279__state <= 2'b10;
          end else begin
            PE_wrapper_279__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_279__state == 2'b11) begin
        if(PE_wrapper_279__ap_done) begin
          PE_wrapper_279__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_279__state == 2'b10) begin
        if(PE_wrapper_279__ap_done_global__q0) begin
          PE_wrapper_279__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_279__ap_start = (PE_wrapper_279__state == 2'b01);
  assign PE_wrapper_280__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_280__is_done__q0 = (PE_wrapper_280__state == 2'b10);
  assign PE_wrapper_280__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_280__state <= 2'b00;
    end else begin
      if(PE_wrapper_280__state == 2'b00) begin
        if(PE_wrapper_280__ap_start_global__q0) begin
          PE_wrapper_280__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_280__state == 2'b01) begin
        if(PE_wrapper_280__ap_ready) begin
          if(PE_wrapper_280__ap_done) begin
            PE_wrapper_280__state <= 2'b10;
          end else begin
            PE_wrapper_280__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_280__state == 2'b11) begin
        if(PE_wrapper_280__ap_done) begin
          PE_wrapper_280__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_280__state == 2'b10) begin
        if(PE_wrapper_280__ap_done_global__q0) begin
          PE_wrapper_280__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_280__ap_start = (PE_wrapper_280__state == 2'b01);
  assign PE_wrapper_281__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_281__is_done__q0 = (PE_wrapper_281__state == 2'b10);
  assign PE_wrapper_281__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_281__state <= 2'b00;
    end else begin
      if(PE_wrapper_281__state == 2'b00) begin
        if(PE_wrapper_281__ap_start_global__q0) begin
          PE_wrapper_281__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_281__state == 2'b01) begin
        if(PE_wrapper_281__ap_ready) begin
          if(PE_wrapper_281__ap_done) begin
            PE_wrapper_281__state <= 2'b10;
          end else begin
            PE_wrapper_281__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_281__state == 2'b11) begin
        if(PE_wrapper_281__ap_done) begin
          PE_wrapper_281__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_281__state == 2'b10) begin
        if(PE_wrapper_281__ap_done_global__q0) begin
          PE_wrapper_281__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_281__ap_start = (PE_wrapper_281__state == 2'b01);
  assign PE_wrapper_282__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_282__is_done__q0 = (PE_wrapper_282__state == 2'b10);
  assign PE_wrapper_282__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_282__state <= 2'b00;
    end else begin
      if(PE_wrapper_282__state == 2'b00) begin
        if(PE_wrapper_282__ap_start_global__q0) begin
          PE_wrapper_282__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_282__state == 2'b01) begin
        if(PE_wrapper_282__ap_ready) begin
          if(PE_wrapper_282__ap_done) begin
            PE_wrapper_282__state <= 2'b10;
          end else begin
            PE_wrapper_282__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_282__state == 2'b11) begin
        if(PE_wrapper_282__ap_done) begin
          PE_wrapper_282__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_282__state == 2'b10) begin
        if(PE_wrapper_282__ap_done_global__q0) begin
          PE_wrapper_282__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_282__ap_start = (PE_wrapper_282__state == 2'b01);
  assign PE_wrapper_283__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_283__is_done__q0 = (PE_wrapper_283__state == 2'b10);
  assign PE_wrapper_283__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_283__state <= 2'b00;
    end else begin
      if(PE_wrapper_283__state == 2'b00) begin
        if(PE_wrapper_283__ap_start_global__q0) begin
          PE_wrapper_283__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_283__state == 2'b01) begin
        if(PE_wrapper_283__ap_ready) begin
          if(PE_wrapper_283__ap_done) begin
            PE_wrapper_283__state <= 2'b10;
          end else begin
            PE_wrapper_283__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_283__state == 2'b11) begin
        if(PE_wrapper_283__ap_done) begin
          PE_wrapper_283__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_283__state == 2'b10) begin
        if(PE_wrapper_283__ap_done_global__q0) begin
          PE_wrapper_283__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_283__ap_start = (PE_wrapper_283__state == 2'b01);
  assign PE_wrapper_284__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_284__is_done__q0 = (PE_wrapper_284__state == 2'b10);
  assign PE_wrapper_284__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_284__state <= 2'b00;
    end else begin
      if(PE_wrapper_284__state == 2'b00) begin
        if(PE_wrapper_284__ap_start_global__q0) begin
          PE_wrapper_284__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_284__state == 2'b01) begin
        if(PE_wrapper_284__ap_ready) begin
          if(PE_wrapper_284__ap_done) begin
            PE_wrapper_284__state <= 2'b10;
          end else begin
            PE_wrapper_284__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_284__state == 2'b11) begin
        if(PE_wrapper_284__ap_done) begin
          PE_wrapper_284__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_284__state == 2'b10) begin
        if(PE_wrapper_284__ap_done_global__q0) begin
          PE_wrapper_284__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_284__ap_start = (PE_wrapper_284__state == 2'b01);
  assign PE_wrapper_285__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_285__is_done__q0 = (PE_wrapper_285__state == 2'b10);
  assign PE_wrapper_285__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_285__state <= 2'b00;
    end else begin
      if(PE_wrapper_285__state == 2'b00) begin
        if(PE_wrapper_285__ap_start_global__q0) begin
          PE_wrapper_285__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_285__state == 2'b01) begin
        if(PE_wrapper_285__ap_ready) begin
          if(PE_wrapper_285__ap_done) begin
            PE_wrapper_285__state <= 2'b10;
          end else begin
            PE_wrapper_285__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_285__state == 2'b11) begin
        if(PE_wrapper_285__ap_done) begin
          PE_wrapper_285__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_285__state == 2'b10) begin
        if(PE_wrapper_285__ap_done_global__q0) begin
          PE_wrapper_285__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_285__ap_start = (PE_wrapper_285__state == 2'b01);
  assign PE_wrapper_286__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_286__is_done__q0 = (PE_wrapper_286__state == 2'b10);
  assign PE_wrapper_286__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_286__state <= 2'b00;
    end else begin
      if(PE_wrapper_286__state == 2'b00) begin
        if(PE_wrapper_286__ap_start_global__q0) begin
          PE_wrapper_286__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_286__state == 2'b01) begin
        if(PE_wrapper_286__ap_ready) begin
          if(PE_wrapper_286__ap_done) begin
            PE_wrapper_286__state <= 2'b10;
          end else begin
            PE_wrapper_286__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_286__state == 2'b11) begin
        if(PE_wrapper_286__ap_done) begin
          PE_wrapper_286__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_286__state == 2'b10) begin
        if(PE_wrapper_286__ap_done_global__q0) begin
          PE_wrapper_286__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_286__ap_start = (PE_wrapper_286__state == 2'b01);
  assign PE_wrapper_287__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_287__is_done__q0 = (PE_wrapper_287__state == 2'b10);
  assign PE_wrapper_287__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_287__state <= 2'b00;
    end else begin
      if(PE_wrapper_287__state == 2'b00) begin
        if(PE_wrapper_287__ap_start_global__q0) begin
          PE_wrapper_287__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_287__state == 2'b01) begin
        if(PE_wrapper_287__ap_ready) begin
          if(PE_wrapper_287__ap_done) begin
            PE_wrapper_287__state <= 2'b10;
          end else begin
            PE_wrapper_287__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_287__state == 2'b11) begin
        if(PE_wrapper_287__ap_done) begin
          PE_wrapper_287__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_287__state == 2'b10) begin
        if(PE_wrapper_287__ap_done_global__q0) begin
          PE_wrapper_287__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_287__ap_start = (PE_wrapper_287__state == 2'b01);
  assign PE_wrapper_288__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_288__is_done__q0 = (PE_wrapper_288__state == 2'b10);
  assign PE_wrapper_288__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_288__state <= 2'b00;
    end else begin
      if(PE_wrapper_288__state == 2'b00) begin
        if(PE_wrapper_288__ap_start_global__q0) begin
          PE_wrapper_288__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_288__state == 2'b01) begin
        if(PE_wrapper_288__ap_ready) begin
          if(PE_wrapper_288__ap_done) begin
            PE_wrapper_288__state <= 2'b10;
          end else begin
            PE_wrapper_288__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_288__state == 2'b11) begin
        if(PE_wrapper_288__ap_done) begin
          PE_wrapper_288__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_288__state == 2'b10) begin
        if(PE_wrapper_288__ap_done_global__q0) begin
          PE_wrapper_288__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_288__ap_start = (PE_wrapper_288__state == 2'b01);
  assign PE_wrapper_289__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_289__is_done__q0 = (PE_wrapper_289__state == 2'b10);
  assign PE_wrapper_289__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_289__state <= 2'b00;
    end else begin
      if(PE_wrapper_289__state == 2'b00) begin
        if(PE_wrapper_289__ap_start_global__q0) begin
          PE_wrapper_289__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_289__state == 2'b01) begin
        if(PE_wrapper_289__ap_ready) begin
          if(PE_wrapper_289__ap_done) begin
            PE_wrapper_289__state <= 2'b10;
          end else begin
            PE_wrapper_289__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_289__state == 2'b11) begin
        if(PE_wrapper_289__ap_done) begin
          PE_wrapper_289__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_289__state == 2'b10) begin
        if(PE_wrapper_289__ap_done_global__q0) begin
          PE_wrapper_289__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_289__ap_start = (PE_wrapper_289__state == 2'b01);
  assign PE_wrapper_290__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_290__is_done__q0 = (PE_wrapper_290__state == 2'b10);
  assign PE_wrapper_290__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_290__state <= 2'b00;
    end else begin
      if(PE_wrapper_290__state == 2'b00) begin
        if(PE_wrapper_290__ap_start_global__q0) begin
          PE_wrapper_290__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_290__state == 2'b01) begin
        if(PE_wrapper_290__ap_ready) begin
          if(PE_wrapper_290__ap_done) begin
            PE_wrapper_290__state <= 2'b10;
          end else begin
            PE_wrapper_290__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_290__state == 2'b11) begin
        if(PE_wrapper_290__ap_done) begin
          PE_wrapper_290__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_290__state == 2'b10) begin
        if(PE_wrapper_290__ap_done_global__q0) begin
          PE_wrapper_290__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_290__ap_start = (PE_wrapper_290__state == 2'b01);
  assign PE_wrapper_291__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_291__is_done__q0 = (PE_wrapper_291__state == 2'b10);
  assign PE_wrapper_291__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_291__state <= 2'b00;
    end else begin
      if(PE_wrapper_291__state == 2'b00) begin
        if(PE_wrapper_291__ap_start_global__q0) begin
          PE_wrapper_291__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_291__state == 2'b01) begin
        if(PE_wrapper_291__ap_ready) begin
          if(PE_wrapper_291__ap_done) begin
            PE_wrapper_291__state <= 2'b10;
          end else begin
            PE_wrapper_291__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_291__state == 2'b11) begin
        if(PE_wrapper_291__ap_done) begin
          PE_wrapper_291__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_291__state == 2'b10) begin
        if(PE_wrapper_291__ap_done_global__q0) begin
          PE_wrapper_291__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_291__ap_start = (PE_wrapper_291__state == 2'b01);
  assign PE_wrapper_292__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_292__is_done__q0 = (PE_wrapper_292__state == 2'b10);
  assign PE_wrapper_292__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_292__state <= 2'b00;
    end else begin
      if(PE_wrapper_292__state == 2'b00) begin
        if(PE_wrapper_292__ap_start_global__q0) begin
          PE_wrapper_292__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_292__state == 2'b01) begin
        if(PE_wrapper_292__ap_ready) begin
          if(PE_wrapper_292__ap_done) begin
            PE_wrapper_292__state <= 2'b10;
          end else begin
            PE_wrapper_292__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_292__state == 2'b11) begin
        if(PE_wrapper_292__ap_done) begin
          PE_wrapper_292__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_292__state == 2'b10) begin
        if(PE_wrapper_292__ap_done_global__q0) begin
          PE_wrapper_292__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_292__ap_start = (PE_wrapper_292__state == 2'b01);
  assign PE_wrapper_293__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_293__is_done__q0 = (PE_wrapper_293__state == 2'b10);
  assign PE_wrapper_293__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_293__state <= 2'b00;
    end else begin
      if(PE_wrapper_293__state == 2'b00) begin
        if(PE_wrapper_293__ap_start_global__q0) begin
          PE_wrapper_293__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_293__state == 2'b01) begin
        if(PE_wrapper_293__ap_ready) begin
          if(PE_wrapper_293__ap_done) begin
            PE_wrapper_293__state <= 2'b10;
          end else begin
            PE_wrapper_293__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_293__state == 2'b11) begin
        if(PE_wrapper_293__ap_done) begin
          PE_wrapper_293__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_293__state == 2'b10) begin
        if(PE_wrapper_293__ap_done_global__q0) begin
          PE_wrapper_293__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_293__ap_start = (PE_wrapper_293__state == 2'b01);
  assign PE_wrapper_294__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_294__is_done__q0 = (PE_wrapper_294__state == 2'b10);
  assign PE_wrapper_294__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_294__state <= 2'b00;
    end else begin
      if(PE_wrapper_294__state == 2'b00) begin
        if(PE_wrapper_294__ap_start_global__q0) begin
          PE_wrapper_294__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_294__state == 2'b01) begin
        if(PE_wrapper_294__ap_ready) begin
          if(PE_wrapper_294__ap_done) begin
            PE_wrapper_294__state <= 2'b10;
          end else begin
            PE_wrapper_294__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_294__state == 2'b11) begin
        if(PE_wrapper_294__ap_done) begin
          PE_wrapper_294__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_294__state == 2'b10) begin
        if(PE_wrapper_294__ap_done_global__q0) begin
          PE_wrapper_294__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_294__ap_start = (PE_wrapper_294__state == 2'b01);
  assign PE_wrapper_295__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_295__is_done__q0 = (PE_wrapper_295__state == 2'b10);
  assign PE_wrapper_295__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_295__state <= 2'b00;
    end else begin
      if(PE_wrapper_295__state == 2'b00) begin
        if(PE_wrapper_295__ap_start_global__q0) begin
          PE_wrapper_295__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_295__state == 2'b01) begin
        if(PE_wrapper_295__ap_ready) begin
          if(PE_wrapper_295__ap_done) begin
            PE_wrapper_295__state <= 2'b10;
          end else begin
            PE_wrapper_295__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_295__state == 2'b11) begin
        if(PE_wrapper_295__ap_done) begin
          PE_wrapper_295__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_295__state == 2'b10) begin
        if(PE_wrapper_295__ap_done_global__q0) begin
          PE_wrapper_295__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_295__ap_start = (PE_wrapper_295__state == 2'b01);
  assign PE_wrapper_296__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_296__is_done__q0 = (PE_wrapper_296__state == 2'b10);
  assign PE_wrapper_296__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_296__state <= 2'b00;
    end else begin
      if(PE_wrapper_296__state == 2'b00) begin
        if(PE_wrapper_296__ap_start_global__q0) begin
          PE_wrapper_296__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_296__state == 2'b01) begin
        if(PE_wrapper_296__ap_ready) begin
          if(PE_wrapper_296__ap_done) begin
            PE_wrapper_296__state <= 2'b10;
          end else begin
            PE_wrapper_296__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_296__state == 2'b11) begin
        if(PE_wrapper_296__ap_done) begin
          PE_wrapper_296__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_296__state == 2'b10) begin
        if(PE_wrapper_296__ap_done_global__q0) begin
          PE_wrapper_296__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_296__ap_start = (PE_wrapper_296__state == 2'b01);
  assign PE_wrapper_297__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_297__is_done__q0 = (PE_wrapper_297__state == 2'b10);
  assign PE_wrapper_297__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_297__state <= 2'b00;
    end else begin
      if(PE_wrapper_297__state == 2'b00) begin
        if(PE_wrapper_297__ap_start_global__q0) begin
          PE_wrapper_297__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_297__state == 2'b01) begin
        if(PE_wrapper_297__ap_ready) begin
          if(PE_wrapper_297__ap_done) begin
            PE_wrapper_297__state <= 2'b10;
          end else begin
            PE_wrapper_297__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_297__state == 2'b11) begin
        if(PE_wrapper_297__ap_done) begin
          PE_wrapper_297__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_297__state == 2'b10) begin
        if(PE_wrapper_297__ap_done_global__q0) begin
          PE_wrapper_297__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_297__ap_start = (PE_wrapper_297__state == 2'b01);
  assign PE_wrapper_298__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_298__is_done__q0 = (PE_wrapper_298__state == 2'b10);
  assign PE_wrapper_298__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_298__state <= 2'b00;
    end else begin
      if(PE_wrapper_298__state == 2'b00) begin
        if(PE_wrapper_298__ap_start_global__q0) begin
          PE_wrapper_298__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_298__state == 2'b01) begin
        if(PE_wrapper_298__ap_ready) begin
          if(PE_wrapper_298__ap_done) begin
            PE_wrapper_298__state <= 2'b10;
          end else begin
            PE_wrapper_298__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_298__state == 2'b11) begin
        if(PE_wrapper_298__ap_done) begin
          PE_wrapper_298__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_298__state == 2'b10) begin
        if(PE_wrapper_298__ap_done_global__q0) begin
          PE_wrapper_298__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_298__ap_start = (PE_wrapper_298__state == 2'b01);
  assign PE_wrapper_299__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_299__is_done__q0 = (PE_wrapper_299__state == 2'b10);
  assign PE_wrapper_299__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_299__state <= 2'b00;
    end else begin
      if(PE_wrapper_299__state == 2'b00) begin
        if(PE_wrapper_299__ap_start_global__q0) begin
          PE_wrapper_299__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_299__state == 2'b01) begin
        if(PE_wrapper_299__ap_ready) begin
          if(PE_wrapper_299__ap_done) begin
            PE_wrapper_299__state <= 2'b10;
          end else begin
            PE_wrapper_299__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_299__state == 2'b11) begin
        if(PE_wrapper_299__ap_done) begin
          PE_wrapper_299__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_299__state == 2'b10) begin
        if(PE_wrapper_299__ap_done_global__q0) begin
          PE_wrapper_299__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_299__ap_start = (PE_wrapper_299__state == 2'b01);
  assign PE_wrapper_300__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_300__is_done__q0 = (PE_wrapper_300__state == 2'b10);
  assign PE_wrapper_300__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_300__state <= 2'b00;
    end else begin
      if(PE_wrapper_300__state == 2'b00) begin
        if(PE_wrapper_300__ap_start_global__q0) begin
          PE_wrapper_300__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_300__state == 2'b01) begin
        if(PE_wrapper_300__ap_ready) begin
          if(PE_wrapper_300__ap_done) begin
            PE_wrapper_300__state <= 2'b10;
          end else begin
            PE_wrapper_300__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_300__state == 2'b11) begin
        if(PE_wrapper_300__ap_done) begin
          PE_wrapper_300__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_300__state == 2'b10) begin
        if(PE_wrapper_300__ap_done_global__q0) begin
          PE_wrapper_300__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_300__ap_start = (PE_wrapper_300__state == 2'b01);
  assign PE_wrapper_301__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_301__is_done__q0 = (PE_wrapper_301__state == 2'b10);
  assign PE_wrapper_301__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_301__state <= 2'b00;
    end else begin
      if(PE_wrapper_301__state == 2'b00) begin
        if(PE_wrapper_301__ap_start_global__q0) begin
          PE_wrapper_301__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_301__state == 2'b01) begin
        if(PE_wrapper_301__ap_ready) begin
          if(PE_wrapper_301__ap_done) begin
            PE_wrapper_301__state <= 2'b10;
          end else begin
            PE_wrapper_301__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_301__state == 2'b11) begin
        if(PE_wrapper_301__ap_done) begin
          PE_wrapper_301__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_301__state == 2'b10) begin
        if(PE_wrapper_301__ap_done_global__q0) begin
          PE_wrapper_301__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_301__ap_start = (PE_wrapper_301__state == 2'b01);
  assign PE_wrapper_302__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_302__is_done__q0 = (PE_wrapper_302__state == 2'b10);
  assign PE_wrapper_302__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_302__state <= 2'b00;
    end else begin
      if(PE_wrapper_302__state == 2'b00) begin
        if(PE_wrapper_302__ap_start_global__q0) begin
          PE_wrapper_302__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_302__state == 2'b01) begin
        if(PE_wrapper_302__ap_ready) begin
          if(PE_wrapper_302__ap_done) begin
            PE_wrapper_302__state <= 2'b10;
          end else begin
            PE_wrapper_302__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_302__state == 2'b11) begin
        if(PE_wrapper_302__ap_done) begin
          PE_wrapper_302__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_302__state == 2'b10) begin
        if(PE_wrapper_302__ap_done_global__q0) begin
          PE_wrapper_302__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_302__ap_start = (PE_wrapper_302__state == 2'b01);
  assign PE_wrapper_303__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_303__is_done__q0 = (PE_wrapper_303__state == 2'b10);
  assign PE_wrapper_303__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_303__state <= 2'b00;
    end else begin
      if(PE_wrapper_303__state == 2'b00) begin
        if(PE_wrapper_303__ap_start_global__q0) begin
          PE_wrapper_303__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_303__state == 2'b01) begin
        if(PE_wrapper_303__ap_ready) begin
          if(PE_wrapper_303__ap_done) begin
            PE_wrapper_303__state <= 2'b10;
          end else begin
            PE_wrapper_303__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_303__state == 2'b11) begin
        if(PE_wrapper_303__ap_done) begin
          PE_wrapper_303__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_303__state == 2'b10) begin
        if(PE_wrapper_303__ap_done_global__q0) begin
          PE_wrapper_303__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_303__ap_start = (PE_wrapper_303__state == 2'b01);
  assign PE_wrapper_304__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_304__is_done__q0 = (PE_wrapper_304__state == 2'b10);
  assign PE_wrapper_304__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_304__state <= 2'b00;
    end else begin
      if(PE_wrapper_304__state == 2'b00) begin
        if(PE_wrapper_304__ap_start_global__q0) begin
          PE_wrapper_304__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_304__state == 2'b01) begin
        if(PE_wrapper_304__ap_ready) begin
          if(PE_wrapper_304__ap_done) begin
            PE_wrapper_304__state <= 2'b10;
          end else begin
            PE_wrapper_304__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_304__state == 2'b11) begin
        if(PE_wrapper_304__ap_done) begin
          PE_wrapper_304__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_304__state == 2'b10) begin
        if(PE_wrapper_304__ap_done_global__q0) begin
          PE_wrapper_304__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_304__ap_start = (PE_wrapper_304__state == 2'b01);
  assign PE_wrapper_305__ap_start_global__q0 = ap_start__q0;
  assign PE_wrapper_305__is_done__q0 = (PE_wrapper_305__state == 2'b10);
  assign PE_wrapper_305__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PE_wrapper_305__state <= 2'b00;
    end else begin
      if(PE_wrapper_305__state == 2'b00) begin
        if(PE_wrapper_305__ap_start_global__q0) begin
          PE_wrapper_305__state <= 2'b01;
        end 
      end 
      if(PE_wrapper_305__state == 2'b01) begin
        if(PE_wrapper_305__ap_ready) begin
          if(PE_wrapper_305__ap_done) begin
            PE_wrapper_305__state <= 2'b10;
          end else begin
            PE_wrapper_305__state <= 2'b11;
          end
        end 
      end 
      if(PE_wrapper_305__state == 2'b11) begin
        if(PE_wrapper_305__ap_done) begin
          PE_wrapper_305__state <= 2'b10;
        end 
      end 
      if(PE_wrapper_305__state == 2'b10) begin
        if(PE_wrapper_305__ap_done_global__q0) begin
          PE_wrapper_305__state <= 2'b00;
        end 
      end 
    end
  end

  assign PE_wrapper_305__ap_start = (PE_wrapper_305__state == 2'b01);

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      tapa_state <= 2'b00;
    end else begin
      case(tapa_state)
        2'b00: begin
          if(ap_start__q0) begin
            tapa_state <= 2'b01;
          end 
        end
        2'b01: begin
          if(A_IO_L2_in_0__is_done__q0 && A_IO_L2_in_1__is_done__q0 && A_IO_L2_in_2__is_done__q0 && A_IO_L2_in_3__is_done__q0 && A_IO_L2_in_4__is_done__q0 && A_IO_L2_in_5__is_done__q0 && A_IO_L2_in_6__is_done__q0 && A_IO_L2_in_7__is_done__q0 && A_IO_L2_in_8__is_done__q0 && A_IO_L2_in_9__is_done__q0 && A_IO_L2_in_10__is_done__q0 && A_IO_L2_in_11__is_done__q0 && A_IO_L2_in_12__is_done__q0 && A_IO_L2_in_13__is_done__q0 && A_IO_L2_in_14__is_done__q0 && A_IO_L2_in_15__is_done__q0 && A_IO_L2_in_16__is_done__q0 && A_IO_L2_in_boundary_0__is_done__q0 && A_IO_L3_in_0__is_done__q0 && A_IO_L3_in_serialize_0__is_done__q0 && A_PE_dummy_in_0__is_done__q0 && A_PE_dummy_in_1__is_done__q0 && A_PE_dummy_in_2__is_done__q0 && A_PE_dummy_in_3__is_done__q0 && A_PE_dummy_in_4__is_done__q0 && A_PE_dummy_in_5__is_done__q0 && A_PE_dummy_in_6__is_done__q0 && A_PE_dummy_in_7__is_done__q0 && A_PE_dummy_in_8__is_done__q0 && A_PE_dummy_in_9__is_done__q0 && A_PE_dummy_in_10__is_done__q0 && A_PE_dummy_in_11__is_done__q0 && A_PE_dummy_in_12__is_done__q0 && A_PE_dummy_in_13__is_done__q0 && A_PE_dummy_in_14__is_done__q0 && A_PE_dummy_in_15__is_done__q0 && A_PE_dummy_in_16__is_done__q0 && A_PE_dummy_in_17__is_done__q0 && B_IO_L2_in_0__is_done__q0 && B_IO_L2_in_1__is_done__q0 && B_IO_L2_in_2__is_done__q0 && B_IO_L2_in_3__is_done__q0 && B_IO_L2_in_4__is_done__q0 && B_IO_L2_in_5__is_done__q0 && B_IO_L2_in_6__is_done__q0 && B_IO_L2_in_7__is_done__q0 && B_IO_L2_in_8__is_done__q0 && B_IO_L2_in_9__is_done__q0 && B_IO_L2_in_10__is_done__q0 && B_IO_L2_in_11__is_done__q0 && B_IO_L2_in_12__is_done__q0 && B_IO_L2_in_13__is_done__q0 && B_IO_L2_in_14__is_done__q0 && B_IO_L2_in_15__is_done__q0 && B_IO_L2_in_boundary_0__is_done__q0 && B_IO_L3_in_0__is_done__q0 && B_IO_L3_in_serialize_0__is_done__q0 && B_PE_dummy_in_0__is_done__q0 && B_PE_dummy_in_1__is_done__q0 && B_PE_dummy_in_2__is_done__q0 && B_PE_dummy_in_3__is_done__q0 && B_PE_dummy_in_4__is_done__q0 && B_PE_dummy_in_5__is_done__q0 && B_PE_dummy_in_6__is_done__q0 && B_PE_dummy_in_7__is_done__q0 && B_PE_dummy_in_8__is_done__q0 && B_PE_dummy_in_9__is_done__q0 && B_PE_dummy_in_10__is_done__q0 && B_PE_dummy_in_11__is_done__q0 && B_PE_dummy_in_12__is_done__q0 && B_PE_dummy_in_13__is_done__q0 && B_PE_dummy_in_14__is_done__q0 && B_PE_dummy_in_15__is_done__q0 && B_PE_dummy_in_16__is_done__q0 && C_drain_IO_L1_out_boundary_wrapper_0__is_done__q0 && C_drain_IO_L1_out_boundary_wrapper_1__is_done__q0 && C_drain_IO_L1_out_boundary_wrapper_2__is_done__q0 && C_drain_IO_L1_out_boundary_wrapper_3__is_done__q0 && C_drain_IO_L1_out_boundary_wrapper_4__is_done__q0 && C_drain_IO_L1_out_boundary_wrapper_5__is_done__q0 && C_drain_IO_L1_out_boundary_wrapper_6__is_done__q0 && C_drain_IO_L1_out_boundary_wrapper_7__is_done__q0 && C_drain_IO_L1_out_boundary_wrapper_8__is_done__q0 && C_drain_IO_L1_out_boundary_wrapper_9__is_done__q0 && C_drain_IO_L1_out_boundary_wrapper_10__is_done__q0 && C_drain_IO_L1_out_boundary_wrapper_11__is_done__q0 && C_drain_IO_L1_out_boundary_wrapper_12__is_done__q0 && C_drain_IO_L1_out_boundary_wrapper_13__is_done__q0 && C_drain_IO_L1_out_boundary_wrapper_14__is_done__q0 && C_drain_IO_L1_out_boundary_wrapper_15__is_done__q0 && C_drain_IO_L1_out_boundary_wrapper_16__is_done__q0 && C_drain_IO_L1_out_wrapper_0__is_done__q0 && C_drain_IO_L1_out_wrapper_1__is_done__q0 && C_drain_IO_L1_out_wrapper_2__is_done__q0 && C_drain_IO_L1_out_wrapper_3__is_done__q0 && C_drain_IO_L1_out_wrapper_4__is_done__q0 && C_drain_IO_L1_out_wrapper_5__is_done__q0 && C_drain_IO_L1_out_wrapper_6__is_done__q0 && C_drain_IO_L1_out_wrapper_7__is_done__q0 && C_drain_IO_L1_out_wrapper_8__is_done__q0 && C_drain_IO_L1_out_wrapper_9__is_done__q0 && C_drain_IO_L1_out_wrapper_10__is_done__q0 && C_drain_IO_L1_out_wrapper_11__is_done__q0 && C_drain_IO_L1_out_wrapper_12__is_done__q0 && C_drain_IO_L1_out_wrapper_13__is_done__q0 && C_drain_IO_L1_out_wrapper_14__is_done__q0 && C_drain_IO_L1_out_wrapper_15__is_done__q0 && C_drain_IO_L1_out_wrapper_16__is_done__q0 && C_drain_IO_L1_out_wrapper_17__is_done__q0 && C_drain_IO_L1_out_wrapper_18__is_done__q0 && C_drain_IO_L1_out_wrapper_19__is_done__q0 && C_drain_IO_L1_out_wrapper_20__is_done__q0 && C_drain_IO_L1_out_wrapper_21__is_done__q0 && C_drain_IO_L1_out_wrapper_22__is_done__q0 && C_drain_IO_L1_out_wrapper_23__is_done__q0 && C_drain_IO_L1_out_wrapper_24__is_done__q0 && C_drain_IO_L1_out_wrapper_25__is_done__q0 && C_drain_IO_L1_out_wrapper_26__is_done__q0 && C_drain_IO_L1_out_wrapper_27__is_done__q0 && C_drain_IO_L1_out_wrapper_28__is_done__q0 && C_drain_IO_L1_out_wrapper_29__is_done__q0 && C_drain_IO_L1_out_wrapper_30__is_done__q0 && C_drain_IO_L1_out_wrapper_31__is_done__q0 && C_drain_IO_L1_out_wrapper_32__is_done__q0 && C_drain_IO_L1_out_wrapper_33__is_done__q0 && C_drain_IO_L1_out_wrapper_34__is_done__q0 && C_drain_IO_L1_out_wrapper_35__is_done__q0 && C_drain_IO_L1_out_wrapper_36__is_done__q0 && C_drain_IO_L1_out_wrapper_37__is_done__q0 && C_drain_IO_L1_out_wrapper_38__is_done__q0 && C_drain_IO_L1_out_wrapper_39__is_done__q0 && C_drain_IO_L1_out_wrapper_40__is_done__q0 && C_drain_IO_L1_out_wrapper_41__is_done__q0 && C_drain_IO_L1_out_wrapper_42__is_done__q0 && C_drain_IO_L1_out_wrapper_43__is_done__q0 && C_drain_IO_L1_out_wrapper_44__is_done__q0 && C_drain_IO_L1_out_wrapper_45__is_done__q0 && C_drain_IO_L1_out_wrapper_46__is_done__q0 && C_drain_IO_L1_out_wrapper_47__is_done__q0 && C_drain_IO_L1_out_wrapper_48__is_done__q0 && C_drain_IO_L1_out_wrapper_49__is_done__q0 && C_drain_IO_L1_out_wrapper_50__is_done__q0 && C_drain_IO_L1_out_wrapper_51__is_done__q0 && C_drain_IO_L1_out_wrapper_52__is_done__q0 && C_drain_IO_L1_out_wrapper_53__is_done__q0 && C_drain_IO_L1_out_wrapper_54__is_done__q0 && C_drain_IO_L1_out_wrapper_55__is_done__q0 && C_drain_IO_L1_out_wrapper_56__is_done__q0 && C_drain_IO_L1_out_wrapper_57__is_done__q0 && C_drain_IO_L1_out_wrapper_58__is_done__q0 && C_drain_IO_L1_out_wrapper_59__is_done__q0 && C_drain_IO_L1_out_wrapper_60__is_done__q0 && C_drain_IO_L1_out_wrapper_61__is_done__q0 && C_drain_IO_L1_out_wrapper_62__is_done__q0 && C_drain_IO_L1_out_wrapper_63__is_done__q0 && C_drain_IO_L1_out_wrapper_64__is_done__q0 && C_drain_IO_L1_out_wrapper_65__is_done__q0 && C_drain_IO_L1_out_wrapper_66__is_done__q0 && C_drain_IO_L1_out_wrapper_67__is_done__q0 && C_drain_IO_L1_out_wrapper_68__is_done__q0 && C_drain_IO_L1_out_wrapper_69__is_done__q0 && C_drain_IO_L1_out_wrapper_70__is_done__q0 && C_drain_IO_L1_out_wrapper_71__is_done__q0 && C_drain_IO_L1_out_wrapper_72__is_done__q0 && C_drain_IO_L1_out_wrapper_73__is_done__q0 && C_drain_IO_L1_out_wrapper_74__is_done__q0 && C_drain_IO_L1_out_wrapper_75__is_done__q0 && C_drain_IO_L1_out_wrapper_76__is_done__q0 && C_drain_IO_L1_out_wrapper_77__is_done__q0 && C_drain_IO_L1_out_wrapper_78__is_done__q0 && C_drain_IO_L1_out_wrapper_79__is_done__q0 && C_drain_IO_L1_out_wrapper_80__is_done__q0 && C_drain_IO_L1_out_wrapper_81__is_done__q0 && C_drain_IO_L1_out_wrapper_82__is_done__q0 && C_drain_IO_L1_out_wrapper_83__is_done__q0 && C_drain_IO_L1_out_wrapper_84__is_done__q0 && C_drain_IO_L1_out_wrapper_85__is_done__q0 && C_drain_IO_L1_out_wrapper_86__is_done__q0 && C_drain_IO_L1_out_wrapper_87__is_done__q0 && C_drain_IO_L1_out_wrapper_88__is_done__q0 && C_drain_IO_L1_out_wrapper_89__is_done__q0 && C_drain_IO_L1_out_wrapper_90__is_done__q0 && C_drain_IO_L1_out_wrapper_91__is_done__q0 && C_drain_IO_L1_out_wrapper_92__is_done__q0 && C_drain_IO_L1_out_wrapper_93__is_done__q0 && C_drain_IO_L1_out_wrapper_94__is_done__q0 && C_drain_IO_L1_out_wrapper_95__is_done__q0 && C_drain_IO_L1_out_wrapper_96__is_done__q0 && C_drain_IO_L1_out_wrapper_97__is_done__q0 && C_drain_IO_L1_out_wrapper_98__is_done__q0 && C_drain_IO_L1_out_wrapper_99__is_done__q0 && C_drain_IO_L1_out_wrapper_100__is_done__q0 && C_drain_IO_L1_out_wrapper_101__is_done__q0 && C_drain_IO_L1_out_wrapper_102__is_done__q0 && C_drain_IO_L1_out_wrapper_103__is_done__q0 && C_drain_IO_L1_out_wrapper_104__is_done__q0 && C_drain_IO_L1_out_wrapper_105__is_done__q0 && C_drain_IO_L1_out_wrapper_106__is_done__q0 && C_drain_IO_L1_out_wrapper_107__is_done__q0 && C_drain_IO_L1_out_wrapper_108__is_done__q0 && C_drain_IO_L1_out_wrapper_109__is_done__q0 && C_drain_IO_L1_out_wrapper_110__is_done__q0 && C_drain_IO_L1_out_wrapper_111__is_done__q0 && C_drain_IO_L1_out_wrapper_112__is_done__q0 && C_drain_IO_L1_out_wrapper_113__is_done__q0 && C_drain_IO_L1_out_wrapper_114__is_done__q0 && C_drain_IO_L1_out_wrapper_115__is_done__q0 && C_drain_IO_L1_out_wrapper_116__is_done__q0 && C_drain_IO_L1_out_wrapper_117__is_done__q0 && C_drain_IO_L1_out_wrapper_118__is_done__q0 && C_drain_IO_L1_out_wrapper_119__is_done__q0 && C_drain_IO_L1_out_wrapper_120__is_done__q0 && C_drain_IO_L1_out_wrapper_121__is_done__q0 && C_drain_IO_L1_out_wrapper_122__is_done__q0 && C_drain_IO_L1_out_wrapper_123__is_done__q0 && C_drain_IO_L1_out_wrapper_124__is_done__q0 && C_drain_IO_L1_out_wrapper_125__is_done__q0 && C_drain_IO_L1_out_wrapper_126__is_done__q0 && C_drain_IO_L1_out_wrapper_127__is_done__q0 && C_drain_IO_L1_out_wrapper_128__is_done__q0 && C_drain_IO_L1_out_wrapper_129__is_done__q0 && C_drain_IO_L1_out_wrapper_130__is_done__q0 && C_drain_IO_L1_out_wrapper_131__is_done__q0 && C_drain_IO_L1_out_wrapper_132__is_done__q0 && C_drain_IO_L1_out_wrapper_133__is_done__q0 && C_drain_IO_L1_out_wrapper_134__is_done__q0 && C_drain_IO_L1_out_wrapper_135__is_done__q0 && C_drain_IO_L1_out_wrapper_136__is_done__q0 && C_drain_IO_L1_out_wrapper_137__is_done__q0 && C_drain_IO_L1_out_wrapper_138__is_done__q0 && C_drain_IO_L1_out_wrapper_139__is_done__q0 && C_drain_IO_L1_out_wrapper_140__is_done__q0 && C_drain_IO_L1_out_wrapper_141__is_done__q0 && C_drain_IO_L1_out_wrapper_142__is_done__q0 && C_drain_IO_L1_out_wrapper_143__is_done__q0 && C_drain_IO_L1_out_wrapper_144__is_done__q0 && C_drain_IO_L1_out_wrapper_145__is_done__q0 && C_drain_IO_L1_out_wrapper_146__is_done__q0 && C_drain_IO_L1_out_wrapper_147__is_done__q0 && C_drain_IO_L1_out_wrapper_148__is_done__q0 && C_drain_IO_L1_out_wrapper_149__is_done__q0 && C_drain_IO_L1_out_wrapper_150__is_done__q0 && C_drain_IO_L1_out_wrapper_151__is_done__q0 && C_drain_IO_L1_out_wrapper_152__is_done__q0 && C_drain_IO_L1_out_wrapper_153__is_done__q0 && C_drain_IO_L1_out_wrapper_154__is_done__q0 && C_drain_IO_L1_out_wrapper_155__is_done__q0 && C_drain_IO_L1_out_wrapper_156__is_done__q0 && C_drain_IO_L1_out_wrapper_157__is_done__q0 && C_drain_IO_L1_out_wrapper_158__is_done__q0 && C_drain_IO_L1_out_wrapper_159__is_done__q0 && C_drain_IO_L1_out_wrapper_160__is_done__q0 && C_drain_IO_L1_out_wrapper_161__is_done__q0 && C_drain_IO_L1_out_wrapper_162__is_done__q0 && C_drain_IO_L1_out_wrapper_163__is_done__q0 && C_drain_IO_L1_out_wrapper_164__is_done__q0 && C_drain_IO_L1_out_wrapper_165__is_done__q0 && C_drain_IO_L1_out_wrapper_166__is_done__q0 && C_drain_IO_L1_out_wrapper_167__is_done__q0 && C_drain_IO_L1_out_wrapper_168__is_done__q0 && C_drain_IO_L1_out_wrapper_169__is_done__q0 && C_drain_IO_L1_out_wrapper_170__is_done__q0 && C_drain_IO_L1_out_wrapper_171__is_done__q0 && C_drain_IO_L1_out_wrapper_172__is_done__q0 && C_drain_IO_L1_out_wrapper_173__is_done__q0 && C_drain_IO_L1_out_wrapper_174__is_done__q0 && C_drain_IO_L1_out_wrapper_175__is_done__q0 && C_drain_IO_L1_out_wrapper_176__is_done__q0 && C_drain_IO_L1_out_wrapper_177__is_done__q0 && C_drain_IO_L1_out_wrapper_178__is_done__q0 && C_drain_IO_L1_out_wrapper_179__is_done__q0 && C_drain_IO_L1_out_wrapper_180__is_done__q0 && C_drain_IO_L1_out_wrapper_181__is_done__q0 && C_drain_IO_L1_out_wrapper_182__is_done__q0 && C_drain_IO_L1_out_wrapper_183__is_done__q0 && C_drain_IO_L1_out_wrapper_184__is_done__q0 && C_drain_IO_L1_out_wrapper_185__is_done__q0 && C_drain_IO_L1_out_wrapper_186__is_done__q0 && C_drain_IO_L1_out_wrapper_187__is_done__q0 && C_drain_IO_L1_out_wrapper_188__is_done__q0 && C_drain_IO_L1_out_wrapper_189__is_done__q0 && C_drain_IO_L1_out_wrapper_190__is_done__q0 && C_drain_IO_L1_out_wrapper_191__is_done__q0 && C_drain_IO_L1_out_wrapper_192__is_done__q0 && C_drain_IO_L1_out_wrapper_193__is_done__q0 && C_drain_IO_L1_out_wrapper_194__is_done__q0 && C_drain_IO_L1_out_wrapper_195__is_done__q0 && C_drain_IO_L1_out_wrapper_196__is_done__q0 && C_drain_IO_L1_out_wrapper_197__is_done__q0 && C_drain_IO_L1_out_wrapper_198__is_done__q0 && C_drain_IO_L1_out_wrapper_199__is_done__q0 && C_drain_IO_L1_out_wrapper_200__is_done__q0 && C_drain_IO_L1_out_wrapper_201__is_done__q0 && C_drain_IO_L1_out_wrapper_202__is_done__q0 && C_drain_IO_L1_out_wrapper_203__is_done__q0 && C_drain_IO_L1_out_wrapper_204__is_done__q0 && C_drain_IO_L1_out_wrapper_205__is_done__q0 && C_drain_IO_L1_out_wrapper_206__is_done__q0 && C_drain_IO_L1_out_wrapper_207__is_done__q0 && C_drain_IO_L1_out_wrapper_208__is_done__q0 && C_drain_IO_L1_out_wrapper_209__is_done__q0 && C_drain_IO_L1_out_wrapper_210__is_done__q0 && C_drain_IO_L1_out_wrapper_211__is_done__q0 && C_drain_IO_L1_out_wrapper_212__is_done__q0 && C_drain_IO_L1_out_wrapper_213__is_done__q0 && C_drain_IO_L1_out_wrapper_214__is_done__q0 && C_drain_IO_L1_out_wrapper_215__is_done__q0 && C_drain_IO_L1_out_wrapper_216__is_done__q0 && C_drain_IO_L1_out_wrapper_217__is_done__q0 && C_drain_IO_L1_out_wrapper_218__is_done__q0 && C_drain_IO_L1_out_wrapper_219__is_done__q0 && C_drain_IO_L1_out_wrapper_220__is_done__q0 && C_drain_IO_L1_out_wrapper_221__is_done__q0 && C_drain_IO_L1_out_wrapper_222__is_done__q0 && C_drain_IO_L1_out_wrapper_223__is_done__q0 && C_drain_IO_L1_out_wrapper_224__is_done__q0 && C_drain_IO_L1_out_wrapper_225__is_done__q0 && C_drain_IO_L1_out_wrapper_226__is_done__q0 && C_drain_IO_L1_out_wrapper_227__is_done__q0 && C_drain_IO_L1_out_wrapper_228__is_done__q0 && C_drain_IO_L1_out_wrapper_229__is_done__q0 && C_drain_IO_L1_out_wrapper_230__is_done__q0 && C_drain_IO_L1_out_wrapper_231__is_done__q0 && C_drain_IO_L1_out_wrapper_232__is_done__q0 && C_drain_IO_L1_out_wrapper_233__is_done__q0 && C_drain_IO_L1_out_wrapper_234__is_done__q0 && C_drain_IO_L1_out_wrapper_235__is_done__q0 && C_drain_IO_L1_out_wrapper_236__is_done__q0 && C_drain_IO_L1_out_wrapper_237__is_done__q0 && C_drain_IO_L1_out_wrapper_238__is_done__q0 && C_drain_IO_L1_out_wrapper_239__is_done__q0 && C_drain_IO_L1_out_wrapper_240__is_done__q0 && C_drain_IO_L1_out_wrapper_241__is_done__q0 && C_drain_IO_L1_out_wrapper_242__is_done__q0 && C_drain_IO_L1_out_wrapper_243__is_done__q0 && C_drain_IO_L1_out_wrapper_244__is_done__q0 && C_drain_IO_L1_out_wrapper_245__is_done__q0 && C_drain_IO_L1_out_wrapper_246__is_done__q0 && C_drain_IO_L1_out_wrapper_247__is_done__q0 && C_drain_IO_L1_out_wrapper_248__is_done__q0 && C_drain_IO_L1_out_wrapper_249__is_done__q0 && C_drain_IO_L1_out_wrapper_250__is_done__q0 && C_drain_IO_L1_out_wrapper_251__is_done__q0 && C_drain_IO_L1_out_wrapper_252__is_done__q0 && C_drain_IO_L1_out_wrapper_253__is_done__q0 && C_drain_IO_L1_out_wrapper_254__is_done__q0 && C_drain_IO_L1_out_wrapper_255__is_done__q0 && C_drain_IO_L1_out_wrapper_256__is_done__q0 && C_drain_IO_L1_out_wrapper_257__is_done__q0 && C_drain_IO_L1_out_wrapper_258__is_done__q0 && C_drain_IO_L1_out_wrapper_259__is_done__q0 && C_drain_IO_L1_out_wrapper_260__is_done__q0 && C_drain_IO_L1_out_wrapper_261__is_done__q0 && C_drain_IO_L1_out_wrapper_262__is_done__q0 && C_drain_IO_L1_out_wrapper_263__is_done__q0 && C_drain_IO_L1_out_wrapper_264__is_done__q0 && C_drain_IO_L1_out_wrapper_265__is_done__q0 && C_drain_IO_L1_out_wrapper_266__is_done__q0 && C_drain_IO_L1_out_wrapper_267__is_done__q0 && C_drain_IO_L1_out_wrapper_268__is_done__q0 && C_drain_IO_L1_out_wrapper_269__is_done__q0 && C_drain_IO_L1_out_wrapper_270__is_done__q0 && C_drain_IO_L1_out_wrapper_271__is_done__q0 && C_drain_IO_L1_out_wrapper_272__is_done__q0 && C_drain_IO_L1_out_wrapper_273__is_done__q0 && C_drain_IO_L1_out_wrapper_274__is_done__q0 && C_drain_IO_L1_out_wrapper_275__is_done__q0 && C_drain_IO_L1_out_wrapper_276__is_done__q0 && C_drain_IO_L1_out_wrapper_277__is_done__q0 && C_drain_IO_L1_out_wrapper_278__is_done__q0 && C_drain_IO_L1_out_wrapper_279__is_done__q0 && C_drain_IO_L1_out_wrapper_280__is_done__q0 && C_drain_IO_L1_out_wrapper_281__is_done__q0 && C_drain_IO_L1_out_wrapper_282__is_done__q0 && C_drain_IO_L1_out_wrapper_283__is_done__q0 && C_drain_IO_L1_out_wrapper_284__is_done__q0 && C_drain_IO_L1_out_wrapper_285__is_done__q0 && C_drain_IO_L1_out_wrapper_286__is_done__q0 && C_drain_IO_L1_out_wrapper_287__is_done__q0 && C_drain_IO_L1_out_wrapper_288__is_done__q0 && C_drain_IO_L2_out_0__is_done__q0 && C_drain_IO_L2_out_1__is_done__q0 && C_drain_IO_L2_out_2__is_done__q0 && C_drain_IO_L2_out_3__is_done__q0 && C_drain_IO_L2_out_4__is_done__q0 && C_drain_IO_L2_out_5__is_done__q0 && C_drain_IO_L2_out_6__is_done__q0 && C_drain_IO_L2_out_7__is_done__q0 && C_drain_IO_L2_out_8__is_done__q0 && C_drain_IO_L2_out_9__is_done__q0 && C_drain_IO_L2_out_10__is_done__q0 && C_drain_IO_L2_out_11__is_done__q0 && C_drain_IO_L2_out_12__is_done__q0 && C_drain_IO_L2_out_13__is_done__q0 && C_drain_IO_L2_out_14__is_done__q0 && C_drain_IO_L2_out_15__is_done__q0 && C_drain_IO_L2_out_boundary_0__is_done__q0 && C_drain_IO_L3_out_0__is_done__q0 && C_drain_IO_L3_out_serialize_0__is_done__q0 && PE_wrapper_0__is_done__q0 && PE_wrapper_1__is_done__q0 && PE_wrapper_2__is_done__q0 && PE_wrapper_3__is_done__q0 && PE_wrapper_4__is_done__q0 && PE_wrapper_5__is_done__q0 && PE_wrapper_6__is_done__q0 && PE_wrapper_7__is_done__q0 && PE_wrapper_8__is_done__q0 && PE_wrapper_9__is_done__q0 && PE_wrapper_10__is_done__q0 && PE_wrapper_11__is_done__q0 && PE_wrapper_12__is_done__q0 && PE_wrapper_13__is_done__q0 && PE_wrapper_14__is_done__q0 && PE_wrapper_15__is_done__q0 && PE_wrapper_16__is_done__q0 && PE_wrapper_17__is_done__q0 && PE_wrapper_18__is_done__q0 && PE_wrapper_19__is_done__q0 && PE_wrapper_20__is_done__q0 && PE_wrapper_21__is_done__q0 && PE_wrapper_22__is_done__q0 && PE_wrapper_23__is_done__q0 && PE_wrapper_24__is_done__q0 && PE_wrapper_25__is_done__q0 && PE_wrapper_26__is_done__q0 && PE_wrapper_27__is_done__q0 && PE_wrapper_28__is_done__q0 && PE_wrapper_29__is_done__q0 && PE_wrapper_30__is_done__q0 && PE_wrapper_31__is_done__q0 && PE_wrapper_32__is_done__q0 && PE_wrapper_33__is_done__q0 && PE_wrapper_34__is_done__q0 && PE_wrapper_35__is_done__q0 && PE_wrapper_36__is_done__q0 && PE_wrapper_37__is_done__q0 && PE_wrapper_38__is_done__q0 && PE_wrapper_39__is_done__q0 && PE_wrapper_40__is_done__q0 && PE_wrapper_41__is_done__q0 && PE_wrapper_42__is_done__q0 && PE_wrapper_43__is_done__q0 && PE_wrapper_44__is_done__q0 && PE_wrapper_45__is_done__q0 && PE_wrapper_46__is_done__q0 && PE_wrapper_47__is_done__q0 && PE_wrapper_48__is_done__q0 && PE_wrapper_49__is_done__q0 && PE_wrapper_50__is_done__q0 && PE_wrapper_51__is_done__q0 && PE_wrapper_52__is_done__q0 && PE_wrapper_53__is_done__q0 && PE_wrapper_54__is_done__q0 && PE_wrapper_55__is_done__q0 && PE_wrapper_56__is_done__q0 && PE_wrapper_57__is_done__q0 && PE_wrapper_58__is_done__q0 && PE_wrapper_59__is_done__q0 && PE_wrapper_60__is_done__q0 && PE_wrapper_61__is_done__q0 && PE_wrapper_62__is_done__q0 && PE_wrapper_63__is_done__q0 && PE_wrapper_64__is_done__q0 && PE_wrapper_65__is_done__q0 && PE_wrapper_66__is_done__q0 && PE_wrapper_67__is_done__q0 && PE_wrapper_68__is_done__q0 && PE_wrapper_69__is_done__q0 && PE_wrapper_70__is_done__q0 && PE_wrapper_71__is_done__q0 && PE_wrapper_72__is_done__q0 && PE_wrapper_73__is_done__q0 && PE_wrapper_74__is_done__q0 && PE_wrapper_75__is_done__q0 && PE_wrapper_76__is_done__q0 && PE_wrapper_77__is_done__q0 && PE_wrapper_78__is_done__q0 && PE_wrapper_79__is_done__q0 && PE_wrapper_80__is_done__q0 && PE_wrapper_81__is_done__q0 && PE_wrapper_82__is_done__q0 && PE_wrapper_83__is_done__q0 && PE_wrapper_84__is_done__q0 && PE_wrapper_85__is_done__q0 && PE_wrapper_86__is_done__q0 && PE_wrapper_87__is_done__q0 && PE_wrapper_88__is_done__q0 && PE_wrapper_89__is_done__q0 && PE_wrapper_90__is_done__q0 && PE_wrapper_91__is_done__q0 && PE_wrapper_92__is_done__q0 && PE_wrapper_93__is_done__q0 && PE_wrapper_94__is_done__q0 && PE_wrapper_95__is_done__q0 && PE_wrapper_96__is_done__q0 && PE_wrapper_97__is_done__q0 && PE_wrapper_98__is_done__q0 && PE_wrapper_99__is_done__q0 && PE_wrapper_100__is_done__q0 && PE_wrapper_101__is_done__q0 && PE_wrapper_102__is_done__q0 && PE_wrapper_103__is_done__q0 && PE_wrapper_104__is_done__q0 && PE_wrapper_105__is_done__q0 && PE_wrapper_106__is_done__q0 && PE_wrapper_107__is_done__q0 && PE_wrapper_108__is_done__q0 && PE_wrapper_109__is_done__q0 && PE_wrapper_110__is_done__q0 && PE_wrapper_111__is_done__q0 && PE_wrapper_112__is_done__q0 && PE_wrapper_113__is_done__q0 && PE_wrapper_114__is_done__q0 && PE_wrapper_115__is_done__q0 && PE_wrapper_116__is_done__q0 && PE_wrapper_117__is_done__q0 && PE_wrapper_118__is_done__q0 && PE_wrapper_119__is_done__q0 && PE_wrapper_120__is_done__q0 && PE_wrapper_121__is_done__q0 && PE_wrapper_122__is_done__q0 && PE_wrapper_123__is_done__q0 && PE_wrapper_124__is_done__q0 && PE_wrapper_125__is_done__q0 && PE_wrapper_126__is_done__q0 && PE_wrapper_127__is_done__q0 && PE_wrapper_128__is_done__q0 && PE_wrapper_129__is_done__q0 && PE_wrapper_130__is_done__q0 && PE_wrapper_131__is_done__q0 && PE_wrapper_132__is_done__q0 && PE_wrapper_133__is_done__q0 && PE_wrapper_134__is_done__q0 && PE_wrapper_135__is_done__q0 && PE_wrapper_136__is_done__q0 && PE_wrapper_137__is_done__q0 && PE_wrapper_138__is_done__q0 && PE_wrapper_139__is_done__q0 && PE_wrapper_140__is_done__q0 && PE_wrapper_141__is_done__q0 && PE_wrapper_142__is_done__q0 && PE_wrapper_143__is_done__q0 && PE_wrapper_144__is_done__q0 && PE_wrapper_145__is_done__q0 && PE_wrapper_146__is_done__q0 && PE_wrapper_147__is_done__q0 && PE_wrapper_148__is_done__q0 && PE_wrapper_149__is_done__q0 && PE_wrapper_150__is_done__q0 && PE_wrapper_151__is_done__q0 && PE_wrapper_152__is_done__q0 && PE_wrapper_153__is_done__q0 && PE_wrapper_154__is_done__q0 && PE_wrapper_155__is_done__q0 && PE_wrapper_156__is_done__q0 && PE_wrapper_157__is_done__q0 && PE_wrapper_158__is_done__q0 && PE_wrapper_159__is_done__q0 && PE_wrapper_160__is_done__q0 && PE_wrapper_161__is_done__q0 && PE_wrapper_162__is_done__q0 && PE_wrapper_163__is_done__q0 && PE_wrapper_164__is_done__q0 && PE_wrapper_165__is_done__q0 && PE_wrapper_166__is_done__q0 && PE_wrapper_167__is_done__q0 && PE_wrapper_168__is_done__q0 && PE_wrapper_169__is_done__q0 && PE_wrapper_170__is_done__q0 && PE_wrapper_171__is_done__q0 && PE_wrapper_172__is_done__q0 && PE_wrapper_173__is_done__q0 && PE_wrapper_174__is_done__q0 && PE_wrapper_175__is_done__q0 && PE_wrapper_176__is_done__q0 && PE_wrapper_177__is_done__q0 && PE_wrapper_178__is_done__q0 && PE_wrapper_179__is_done__q0 && PE_wrapper_180__is_done__q0 && PE_wrapper_181__is_done__q0 && PE_wrapper_182__is_done__q0 && PE_wrapper_183__is_done__q0 && PE_wrapper_184__is_done__q0 && PE_wrapper_185__is_done__q0 && PE_wrapper_186__is_done__q0 && PE_wrapper_187__is_done__q0 && PE_wrapper_188__is_done__q0 && PE_wrapper_189__is_done__q0 && PE_wrapper_190__is_done__q0 && PE_wrapper_191__is_done__q0 && PE_wrapper_192__is_done__q0 && PE_wrapper_193__is_done__q0 && PE_wrapper_194__is_done__q0 && PE_wrapper_195__is_done__q0 && PE_wrapper_196__is_done__q0 && PE_wrapper_197__is_done__q0 && PE_wrapper_198__is_done__q0 && PE_wrapper_199__is_done__q0 && PE_wrapper_200__is_done__q0 && PE_wrapper_201__is_done__q0 && PE_wrapper_202__is_done__q0 && PE_wrapper_203__is_done__q0 && PE_wrapper_204__is_done__q0 && PE_wrapper_205__is_done__q0 && PE_wrapper_206__is_done__q0 && PE_wrapper_207__is_done__q0 && PE_wrapper_208__is_done__q0 && PE_wrapper_209__is_done__q0 && PE_wrapper_210__is_done__q0 && PE_wrapper_211__is_done__q0 && PE_wrapper_212__is_done__q0 && PE_wrapper_213__is_done__q0 && PE_wrapper_214__is_done__q0 && PE_wrapper_215__is_done__q0 && PE_wrapper_216__is_done__q0 && PE_wrapper_217__is_done__q0 && PE_wrapper_218__is_done__q0 && PE_wrapper_219__is_done__q0 && PE_wrapper_220__is_done__q0 && PE_wrapper_221__is_done__q0 && PE_wrapper_222__is_done__q0 && PE_wrapper_223__is_done__q0 && PE_wrapper_224__is_done__q0 && PE_wrapper_225__is_done__q0 && PE_wrapper_226__is_done__q0 && PE_wrapper_227__is_done__q0 && PE_wrapper_228__is_done__q0 && PE_wrapper_229__is_done__q0 && PE_wrapper_230__is_done__q0 && PE_wrapper_231__is_done__q0 && PE_wrapper_232__is_done__q0 && PE_wrapper_233__is_done__q0 && PE_wrapper_234__is_done__q0 && PE_wrapper_235__is_done__q0 && PE_wrapper_236__is_done__q0 && PE_wrapper_237__is_done__q0 && PE_wrapper_238__is_done__q0 && PE_wrapper_239__is_done__q0 && PE_wrapper_240__is_done__q0 && PE_wrapper_241__is_done__q0 && PE_wrapper_242__is_done__q0 && PE_wrapper_243__is_done__q0 && PE_wrapper_244__is_done__q0 && PE_wrapper_245__is_done__q0 && PE_wrapper_246__is_done__q0 && PE_wrapper_247__is_done__q0 && PE_wrapper_248__is_done__q0 && PE_wrapper_249__is_done__q0 && PE_wrapper_250__is_done__q0 && PE_wrapper_251__is_done__q0 && PE_wrapper_252__is_done__q0 && PE_wrapper_253__is_done__q0 && PE_wrapper_254__is_done__q0 && PE_wrapper_255__is_done__q0 && PE_wrapper_256__is_done__q0 && PE_wrapper_257__is_done__q0 && PE_wrapper_258__is_done__q0 && PE_wrapper_259__is_done__q0 && PE_wrapper_260__is_done__q0 && PE_wrapper_261__is_done__q0 && PE_wrapper_262__is_done__q0 && PE_wrapper_263__is_done__q0 && PE_wrapper_264__is_done__q0 && PE_wrapper_265__is_done__q0 && PE_wrapper_266__is_done__q0 && PE_wrapper_267__is_done__q0 && PE_wrapper_268__is_done__q0 && PE_wrapper_269__is_done__q0 && PE_wrapper_270__is_done__q0 && PE_wrapper_271__is_done__q0 && PE_wrapper_272__is_done__q0 && PE_wrapper_273__is_done__q0 && PE_wrapper_274__is_done__q0 && PE_wrapper_275__is_done__q0 && PE_wrapper_276__is_done__q0 && PE_wrapper_277__is_done__q0 && PE_wrapper_278__is_done__q0 && PE_wrapper_279__is_done__q0 && PE_wrapper_280__is_done__q0 && PE_wrapper_281__is_done__q0 && PE_wrapper_282__is_done__q0 && PE_wrapper_283__is_done__q0 && PE_wrapper_284__is_done__q0 && PE_wrapper_285__is_done__q0 && PE_wrapper_286__is_done__q0 && PE_wrapper_287__is_done__q0 && PE_wrapper_288__is_done__q0 && PE_wrapper_289__is_done__q0 && PE_wrapper_290__is_done__q0 && PE_wrapper_291__is_done__q0 && PE_wrapper_292__is_done__q0 && PE_wrapper_293__is_done__q0 && PE_wrapper_294__is_done__q0 && PE_wrapper_295__is_done__q0 && PE_wrapper_296__is_done__q0 && PE_wrapper_297__is_done__q0 && PE_wrapper_298__is_done__q0 && PE_wrapper_299__is_done__q0 && PE_wrapper_300__is_done__q0 && PE_wrapper_301__is_done__q0 && PE_wrapper_302__is_done__q0 && PE_wrapper_303__is_done__q0 && PE_wrapper_304__is_done__q0 && PE_wrapper_305__is_done__q0) begin
            tapa_state <= 2'b10;
          end 
        end
        2'b10: begin
          tapa_state <= 2'b00;
          countdown <= 1'd0;
        end
        2'b11: begin
          if(countdown == 1'd0) begin
            tapa_state <= 2'b00;
          end else begin
            countdown <= (countdown - 1'd1);
          end
        end
      endcase
    end
  end

  assign ap_idle = (tapa_state == 2'b00);
  assign ap_done = ap_done__q0;
  assign ap_ready = ap_done__q0;
  assign ap_start__q0 = ap_start;
  assign ap_done__q0 = (tapa_state == 2'b10);

endmodule

