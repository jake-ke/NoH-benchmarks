

module Knn_fsm
(
  ap_clk,
  ap_rst_n,
  ap_start,
  ap_ready,
  ap_done,
  ap_idle,
  L3_out_dist,
  L3_out_id,
  in_0,
  in_1,
  in_10,
  in_11,
  in_12,
  in_13,
  in_14,
  in_15,
  in_16,
  in_17,
  in_18,
  in_19,
  in_2,
  in_20,
  in_21,
  in_22,
  in_23,
  in_24,
  in_25,
  in_26,
  in_3,
  in_4,
  in_5,
  in_6,
  in_7,
  in_8,
  in_9,
  krnl_globalSort_L1_L2_0__ap_start,
  krnl_globalSort_L1_L2_0__ap_ready,
  krnl_globalSort_L1_L2_0__ap_done,
  krnl_globalSort_L1_L2_0__ap_idle,
  krnl_globalSort_L1_L2_1__ap_start,
  krnl_globalSort_L1_L2_1__ap_ready,
  krnl_globalSort_L1_L2_1__ap_done,
  krnl_globalSort_L1_L2_1__ap_idle,
  krnl_globalSort_L1_L2_2__ap_start,
  krnl_globalSort_L1_L2_2__ap_ready,
  krnl_globalSort_L1_L2_2__ap_done,
  krnl_globalSort_L1_L2_2__ap_idle,
  krnl_globalSort_L1_L2_3__ap_start,
  krnl_globalSort_L1_L2_3__ap_ready,
  krnl_globalSort_L1_L2_3__ap_done,
  krnl_globalSort_L1_L2_3__ap_idle,
  krnl_globalSort_L1_L2_4__ap_start,
  krnl_globalSort_L1_L2_4__ap_ready,
  krnl_globalSort_L1_L2_4__ap_done,
  krnl_globalSort_L1_L2_4__ap_idle,
  krnl_globalSort_L1_L2_5__ap_start,
  krnl_globalSort_L1_L2_5__ap_ready,
  krnl_globalSort_L1_L2_5__ap_done,
  krnl_globalSort_L1_L2_5__ap_idle,
  krnl_globalSort_L1_L2_6__ap_start,
  krnl_globalSort_L1_L2_6__ap_ready,
  krnl_globalSort_L1_L2_6__ap_done,
  krnl_globalSort_L1_L2_6__ap_idle,
  krnl_globalSort_L1_L2_7__ap_start,
  krnl_globalSort_L1_L2_7__ap_ready,
  krnl_globalSort_L1_L2_7__ap_done,
  krnl_globalSort_L1_L2_7__ap_idle,
  krnl_globalSort_L1_L2_8__ap_start,
  krnl_globalSort_L1_L2_8__ap_ready,
  krnl_globalSort_L1_L2_8__ap_done,
  krnl_globalSort_L1_L2_8__ap_idle,
  krnl_globalSort_L1_L2_9__ap_start,
  krnl_globalSort_L1_L2_9__ap_ready,
  krnl_globalSort_L1_L2_9__ap_done,
  krnl_globalSort_L1_L2_9__ap_idle,
  krnl_globalSort_L1_L2_10__ap_start,
  krnl_globalSort_L1_L2_10__ap_ready,
  krnl_globalSort_L1_L2_10__ap_done,
  krnl_globalSort_L1_L2_10__ap_idle,
  krnl_globalSort_L1_L2_11__ap_start,
  krnl_globalSort_L1_L2_11__ap_ready,
  krnl_globalSort_L1_L2_11__ap_done,
  krnl_globalSort_L1_L2_11__ap_idle,
  krnl_globalSort_L1_L2_12__ap_start,
  krnl_globalSort_L1_L2_12__ap_ready,
  krnl_globalSort_L1_L2_12__ap_done,
  krnl_globalSort_L1_L2_12__ap_idle,
  krnl_output_dist_id_0___L3_out_dist__q0,
  krnl_output_dist_id_0___L3_out_id__q0,
  krnl_output_dist_id_0__ap_start,
  krnl_output_dist_id_0__ap_ready,
  krnl_output_dist_id_0__ap_done,
  krnl_output_dist_id_0__ap_idle,
  krnl_partialKnn_wrapper_0_0___in_0__q0,
  krnl_partialKnn_wrapper_0_0__ap_start,
  krnl_partialKnn_wrapper_0_0__ap_ready,
  krnl_partialKnn_wrapper_0_0__ap_done,
  krnl_partialKnn_wrapper_0_0__ap_idle,
  krnl_partialKnn_wrapper_1_0___in_1__q0,
  krnl_partialKnn_wrapper_1_0__ap_start,
  krnl_partialKnn_wrapper_1_0__ap_ready,
  krnl_partialKnn_wrapper_1_0__ap_done,
  krnl_partialKnn_wrapper_1_0__ap_idle,
  krnl_partialKnn_wrapper_10_0___in_10__q0,
  krnl_partialKnn_wrapper_10_0__ap_start,
  krnl_partialKnn_wrapper_10_0__ap_ready,
  krnl_partialKnn_wrapper_10_0__ap_done,
  krnl_partialKnn_wrapper_10_0__ap_idle,
  krnl_partialKnn_wrapper_11_0___in_11__q0,
  krnl_partialKnn_wrapper_11_0__ap_start,
  krnl_partialKnn_wrapper_11_0__ap_ready,
  krnl_partialKnn_wrapper_11_0__ap_done,
  krnl_partialKnn_wrapper_11_0__ap_idle,
  krnl_partialKnn_wrapper_12_0___in_12__q0,
  krnl_partialKnn_wrapper_12_0__ap_start,
  krnl_partialKnn_wrapper_12_0__ap_ready,
  krnl_partialKnn_wrapper_12_0__ap_done,
  krnl_partialKnn_wrapper_12_0__ap_idle,
  krnl_partialKnn_wrapper_13_0___in_13__q0,
  krnl_partialKnn_wrapper_13_0__ap_start,
  krnl_partialKnn_wrapper_13_0__ap_ready,
  krnl_partialKnn_wrapper_13_0__ap_done,
  krnl_partialKnn_wrapper_13_0__ap_idle,
  krnl_partialKnn_wrapper_14_0___in_14__q0,
  krnl_partialKnn_wrapper_14_0__ap_start,
  krnl_partialKnn_wrapper_14_0__ap_ready,
  krnl_partialKnn_wrapper_14_0__ap_done,
  krnl_partialKnn_wrapper_14_0__ap_idle,
  krnl_partialKnn_wrapper_15_0___in_15__q0,
  krnl_partialKnn_wrapper_15_0__ap_start,
  krnl_partialKnn_wrapper_15_0__ap_ready,
  krnl_partialKnn_wrapper_15_0__ap_done,
  krnl_partialKnn_wrapper_15_0__ap_idle,
  krnl_partialKnn_wrapper_16_0___in_16__q0,
  krnl_partialKnn_wrapper_16_0__ap_start,
  krnl_partialKnn_wrapper_16_0__ap_ready,
  krnl_partialKnn_wrapper_16_0__ap_done,
  krnl_partialKnn_wrapper_16_0__ap_idle,
  krnl_partialKnn_wrapper_17_0___in_17__q0,
  krnl_partialKnn_wrapper_17_0__ap_start,
  krnl_partialKnn_wrapper_17_0__ap_ready,
  krnl_partialKnn_wrapper_17_0__ap_done,
  krnl_partialKnn_wrapper_17_0__ap_idle,
  krnl_partialKnn_wrapper_18_0___in_18__q0,
  krnl_partialKnn_wrapper_18_0__ap_start,
  krnl_partialKnn_wrapper_18_0__ap_ready,
  krnl_partialKnn_wrapper_18_0__ap_done,
  krnl_partialKnn_wrapper_18_0__ap_idle,
  krnl_partialKnn_wrapper_19_0___in_19__q0,
  krnl_partialKnn_wrapper_19_0__ap_start,
  krnl_partialKnn_wrapper_19_0__ap_ready,
  krnl_partialKnn_wrapper_19_0__ap_done,
  krnl_partialKnn_wrapper_19_0__ap_idle,
  krnl_partialKnn_wrapper_2_0___in_2__q0,
  krnl_partialKnn_wrapper_2_0__ap_start,
  krnl_partialKnn_wrapper_2_0__ap_ready,
  krnl_partialKnn_wrapper_2_0__ap_done,
  krnl_partialKnn_wrapper_2_0__ap_idle,
  krnl_partialKnn_wrapper_20_0___in_20__q0,
  krnl_partialKnn_wrapper_20_0__ap_start,
  krnl_partialKnn_wrapper_20_0__ap_ready,
  krnl_partialKnn_wrapper_20_0__ap_done,
  krnl_partialKnn_wrapper_20_0__ap_idle,
  krnl_partialKnn_wrapper_21_0___in_21__q0,
  krnl_partialKnn_wrapper_21_0__ap_start,
  krnl_partialKnn_wrapper_21_0__ap_ready,
  krnl_partialKnn_wrapper_21_0__ap_done,
  krnl_partialKnn_wrapper_21_0__ap_idle,
  krnl_partialKnn_wrapper_22_0___in_22__q0,
  krnl_partialKnn_wrapper_22_0__ap_start,
  krnl_partialKnn_wrapper_22_0__ap_ready,
  krnl_partialKnn_wrapper_22_0__ap_done,
  krnl_partialKnn_wrapper_22_0__ap_idle,
  krnl_partialKnn_wrapper_23_0___in_23__q0,
  krnl_partialKnn_wrapper_23_0__ap_start,
  krnl_partialKnn_wrapper_23_0__ap_ready,
  krnl_partialKnn_wrapper_23_0__ap_done,
  krnl_partialKnn_wrapper_23_0__ap_idle,
  krnl_partialKnn_wrapper_24_0___in_24__q0,
  krnl_partialKnn_wrapper_24_0__ap_start,
  krnl_partialKnn_wrapper_24_0__ap_ready,
  krnl_partialKnn_wrapper_24_0__ap_done,
  krnl_partialKnn_wrapper_24_0__ap_idle,
  krnl_partialKnn_wrapper_25_0___in_25__q0,
  krnl_partialKnn_wrapper_25_0__ap_start,
  krnl_partialKnn_wrapper_25_0__ap_ready,
  krnl_partialKnn_wrapper_25_0__ap_done,
  krnl_partialKnn_wrapper_25_0__ap_idle,
  krnl_partialKnn_wrapper_26_0___in_26__q0,
  krnl_partialKnn_wrapper_26_0__ap_start,
  krnl_partialKnn_wrapper_26_0__ap_ready,
  krnl_partialKnn_wrapper_26_0__ap_done,
  krnl_partialKnn_wrapper_26_0__ap_idle,
  krnl_partialKnn_wrapper_3_0___in_3__q0,
  krnl_partialKnn_wrapper_3_0__ap_start,
  krnl_partialKnn_wrapper_3_0__ap_ready,
  krnl_partialKnn_wrapper_3_0__ap_done,
  krnl_partialKnn_wrapper_3_0__ap_idle,
  krnl_partialKnn_wrapper_4_0___in_4__q0,
  krnl_partialKnn_wrapper_4_0__ap_start,
  krnl_partialKnn_wrapper_4_0__ap_ready,
  krnl_partialKnn_wrapper_4_0__ap_done,
  krnl_partialKnn_wrapper_4_0__ap_idle,
  krnl_partialKnn_wrapper_5_0___in_5__q0,
  krnl_partialKnn_wrapper_5_0__ap_start,
  krnl_partialKnn_wrapper_5_0__ap_ready,
  krnl_partialKnn_wrapper_5_0__ap_done,
  krnl_partialKnn_wrapper_5_0__ap_idle,
  krnl_partialKnn_wrapper_6_0___in_6__q0,
  krnl_partialKnn_wrapper_6_0__ap_start,
  krnl_partialKnn_wrapper_6_0__ap_ready,
  krnl_partialKnn_wrapper_6_0__ap_done,
  krnl_partialKnn_wrapper_6_0__ap_idle,
  krnl_partialKnn_wrapper_7_0___in_7__q0,
  krnl_partialKnn_wrapper_7_0__ap_start,
  krnl_partialKnn_wrapper_7_0__ap_ready,
  krnl_partialKnn_wrapper_7_0__ap_done,
  krnl_partialKnn_wrapper_7_0__ap_idle,
  krnl_partialKnn_wrapper_8_0___in_8__q0,
  krnl_partialKnn_wrapper_8_0__ap_start,
  krnl_partialKnn_wrapper_8_0__ap_ready,
  krnl_partialKnn_wrapper_8_0__ap_done,
  krnl_partialKnn_wrapper_8_0__ap_idle,
  krnl_partialKnn_wrapper_9_0___in_9__q0,
  krnl_partialKnn_wrapper_9_0__ap_start,
  krnl_partialKnn_wrapper_9_0__ap_ready,
  krnl_partialKnn_wrapper_9_0__ap_done,
  krnl_partialKnn_wrapper_9_0__ap_idle
);

  // pragma RS clk port=ap_clk
  // pragma RS rst port=ap_rst_n active=low
  // pragma RS ap-ctrl ap_start=ap_start ap_done=ap_done ap_idle=ap_idle ap_ready=ap_ready scalar=(in_0|in_1|in_2|in_3|in_4|in_5|in_6|in_7|in_8|in_9|in_10|in_11|in_12|in_13|in_14|in_15|in_16|in_17|in_18|in_19|in_20|in_21|in_22|in_23|in_24|in_25|in_26|L3_out_dist|L3_out_id)
  // pragma RS ap-ctrl ap_start=krnl_globalSort_L1_L2_0__ap_start ap_done=krnl_globalSort_L1_L2_0__ap_done ap_idle=krnl_globalSort_L1_L2_0__ap_idle ap_ready=krnl_globalSort_L1_L2_0__ap_ready
  // pragma RS ap-ctrl ap_start=krnl_globalSort_L1_L2_1__ap_start ap_done=krnl_globalSort_L1_L2_1__ap_done ap_idle=krnl_globalSort_L1_L2_1__ap_idle ap_ready=krnl_globalSort_L1_L2_1__ap_ready
  // pragma RS ap-ctrl ap_start=krnl_globalSort_L1_L2_2__ap_start ap_done=krnl_globalSort_L1_L2_2__ap_done ap_idle=krnl_globalSort_L1_L2_2__ap_idle ap_ready=krnl_globalSort_L1_L2_2__ap_ready
  // pragma RS ap-ctrl ap_start=krnl_globalSort_L1_L2_3__ap_start ap_done=krnl_globalSort_L1_L2_3__ap_done ap_idle=krnl_globalSort_L1_L2_3__ap_idle ap_ready=krnl_globalSort_L1_L2_3__ap_ready
  // pragma RS ap-ctrl ap_start=krnl_globalSort_L1_L2_4__ap_start ap_done=krnl_globalSort_L1_L2_4__ap_done ap_idle=krnl_globalSort_L1_L2_4__ap_idle ap_ready=krnl_globalSort_L1_L2_4__ap_ready
  // pragma RS ap-ctrl ap_start=krnl_globalSort_L1_L2_5__ap_start ap_done=krnl_globalSort_L1_L2_5__ap_done ap_idle=krnl_globalSort_L1_L2_5__ap_idle ap_ready=krnl_globalSort_L1_L2_5__ap_ready
  // pragma RS ap-ctrl ap_start=krnl_globalSort_L1_L2_6__ap_start ap_done=krnl_globalSort_L1_L2_6__ap_done ap_idle=krnl_globalSort_L1_L2_6__ap_idle ap_ready=krnl_globalSort_L1_L2_6__ap_ready
  // pragma RS ap-ctrl ap_start=krnl_globalSort_L1_L2_7__ap_start ap_done=krnl_globalSort_L1_L2_7__ap_done ap_idle=krnl_globalSort_L1_L2_7__ap_idle ap_ready=krnl_globalSort_L1_L2_7__ap_ready
  // pragma RS ap-ctrl ap_start=krnl_globalSort_L1_L2_8__ap_start ap_done=krnl_globalSort_L1_L2_8__ap_done ap_idle=krnl_globalSort_L1_L2_8__ap_idle ap_ready=krnl_globalSort_L1_L2_8__ap_ready
  // pragma RS ap-ctrl ap_start=krnl_globalSort_L1_L2_9__ap_start ap_done=krnl_globalSort_L1_L2_9__ap_done ap_idle=krnl_globalSort_L1_L2_9__ap_idle ap_ready=krnl_globalSort_L1_L2_9__ap_ready
  // pragma RS ap-ctrl ap_start=krnl_globalSort_L1_L2_10__ap_start ap_done=krnl_globalSort_L1_L2_10__ap_done ap_idle=krnl_globalSort_L1_L2_10__ap_idle ap_ready=krnl_globalSort_L1_L2_10__ap_ready
  // pragma RS ap-ctrl ap_start=krnl_globalSort_L1_L2_11__ap_start ap_done=krnl_globalSort_L1_L2_11__ap_done ap_idle=krnl_globalSort_L1_L2_11__ap_idle ap_ready=krnl_globalSort_L1_L2_11__ap_ready
  // pragma RS ap-ctrl ap_start=krnl_globalSort_L1_L2_12__ap_start ap_done=krnl_globalSort_L1_L2_12__ap_done ap_idle=krnl_globalSort_L1_L2_12__ap_idle ap_ready=krnl_globalSort_L1_L2_12__ap_ready
  // pragma RS ap-ctrl ap_start=krnl_output_dist_id_0__ap_start ap_done=krnl_output_dist_id_0__ap_done ap_idle=krnl_output_dist_id_0__ap_idle ap_ready=krnl_output_dist_id_0__ap_ready scalar=krnl_output_dist_id_0___.*
  // pragma RS ap-ctrl ap_start=krnl_partialKnn_wrapper_0_0__ap_start ap_done=krnl_partialKnn_wrapper_0_0__ap_done ap_idle=krnl_partialKnn_wrapper_0_0__ap_idle ap_ready=krnl_partialKnn_wrapper_0_0__ap_ready scalar=krnl_partialKnn_wrapper_0_0___.*
  // pragma RS ap-ctrl ap_start=krnl_partialKnn_wrapper_1_0__ap_start ap_done=krnl_partialKnn_wrapper_1_0__ap_done ap_idle=krnl_partialKnn_wrapper_1_0__ap_idle ap_ready=krnl_partialKnn_wrapper_1_0__ap_ready scalar=krnl_partialKnn_wrapper_1_0___.*
  // pragma RS ap-ctrl ap_start=krnl_partialKnn_wrapper_10_0__ap_start ap_done=krnl_partialKnn_wrapper_10_0__ap_done ap_idle=krnl_partialKnn_wrapper_10_0__ap_idle ap_ready=krnl_partialKnn_wrapper_10_0__ap_ready scalar=krnl_partialKnn_wrapper_10_0___.*
  // pragma RS ap-ctrl ap_start=krnl_partialKnn_wrapper_11_0__ap_start ap_done=krnl_partialKnn_wrapper_11_0__ap_done ap_idle=krnl_partialKnn_wrapper_11_0__ap_idle ap_ready=krnl_partialKnn_wrapper_11_0__ap_ready scalar=krnl_partialKnn_wrapper_11_0___.*
  // pragma RS ap-ctrl ap_start=krnl_partialKnn_wrapper_12_0__ap_start ap_done=krnl_partialKnn_wrapper_12_0__ap_done ap_idle=krnl_partialKnn_wrapper_12_0__ap_idle ap_ready=krnl_partialKnn_wrapper_12_0__ap_ready scalar=krnl_partialKnn_wrapper_12_0___.*
  // pragma RS ap-ctrl ap_start=krnl_partialKnn_wrapper_13_0__ap_start ap_done=krnl_partialKnn_wrapper_13_0__ap_done ap_idle=krnl_partialKnn_wrapper_13_0__ap_idle ap_ready=krnl_partialKnn_wrapper_13_0__ap_ready scalar=krnl_partialKnn_wrapper_13_0___.*
  // pragma RS ap-ctrl ap_start=krnl_partialKnn_wrapper_14_0__ap_start ap_done=krnl_partialKnn_wrapper_14_0__ap_done ap_idle=krnl_partialKnn_wrapper_14_0__ap_idle ap_ready=krnl_partialKnn_wrapper_14_0__ap_ready scalar=krnl_partialKnn_wrapper_14_0___.*
  // pragma RS ap-ctrl ap_start=krnl_partialKnn_wrapper_15_0__ap_start ap_done=krnl_partialKnn_wrapper_15_0__ap_done ap_idle=krnl_partialKnn_wrapper_15_0__ap_idle ap_ready=krnl_partialKnn_wrapper_15_0__ap_ready scalar=krnl_partialKnn_wrapper_15_0___.*
  // pragma RS ap-ctrl ap_start=krnl_partialKnn_wrapper_16_0__ap_start ap_done=krnl_partialKnn_wrapper_16_0__ap_done ap_idle=krnl_partialKnn_wrapper_16_0__ap_idle ap_ready=krnl_partialKnn_wrapper_16_0__ap_ready scalar=krnl_partialKnn_wrapper_16_0___.*
  // pragma RS ap-ctrl ap_start=krnl_partialKnn_wrapper_17_0__ap_start ap_done=krnl_partialKnn_wrapper_17_0__ap_done ap_idle=krnl_partialKnn_wrapper_17_0__ap_idle ap_ready=krnl_partialKnn_wrapper_17_0__ap_ready scalar=krnl_partialKnn_wrapper_17_0___.*
  // pragma RS ap-ctrl ap_start=krnl_partialKnn_wrapper_18_0__ap_start ap_done=krnl_partialKnn_wrapper_18_0__ap_done ap_idle=krnl_partialKnn_wrapper_18_0__ap_idle ap_ready=krnl_partialKnn_wrapper_18_0__ap_ready scalar=krnl_partialKnn_wrapper_18_0___.*
  // pragma RS ap-ctrl ap_start=krnl_partialKnn_wrapper_19_0__ap_start ap_done=krnl_partialKnn_wrapper_19_0__ap_done ap_idle=krnl_partialKnn_wrapper_19_0__ap_idle ap_ready=krnl_partialKnn_wrapper_19_0__ap_ready scalar=krnl_partialKnn_wrapper_19_0___.*
  // pragma RS ap-ctrl ap_start=krnl_partialKnn_wrapper_2_0__ap_start ap_done=krnl_partialKnn_wrapper_2_0__ap_done ap_idle=krnl_partialKnn_wrapper_2_0__ap_idle ap_ready=krnl_partialKnn_wrapper_2_0__ap_ready scalar=krnl_partialKnn_wrapper_2_0___.*
  // pragma RS ap-ctrl ap_start=krnl_partialKnn_wrapper_20_0__ap_start ap_done=krnl_partialKnn_wrapper_20_0__ap_done ap_idle=krnl_partialKnn_wrapper_20_0__ap_idle ap_ready=krnl_partialKnn_wrapper_20_0__ap_ready scalar=krnl_partialKnn_wrapper_20_0___.*
  // pragma RS ap-ctrl ap_start=krnl_partialKnn_wrapper_21_0__ap_start ap_done=krnl_partialKnn_wrapper_21_0__ap_done ap_idle=krnl_partialKnn_wrapper_21_0__ap_idle ap_ready=krnl_partialKnn_wrapper_21_0__ap_ready scalar=krnl_partialKnn_wrapper_21_0___.*
  // pragma RS ap-ctrl ap_start=krnl_partialKnn_wrapper_22_0__ap_start ap_done=krnl_partialKnn_wrapper_22_0__ap_done ap_idle=krnl_partialKnn_wrapper_22_0__ap_idle ap_ready=krnl_partialKnn_wrapper_22_0__ap_ready scalar=krnl_partialKnn_wrapper_22_0___.*
  // pragma RS ap-ctrl ap_start=krnl_partialKnn_wrapper_23_0__ap_start ap_done=krnl_partialKnn_wrapper_23_0__ap_done ap_idle=krnl_partialKnn_wrapper_23_0__ap_idle ap_ready=krnl_partialKnn_wrapper_23_0__ap_ready scalar=krnl_partialKnn_wrapper_23_0___.*
  // pragma RS ap-ctrl ap_start=krnl_partialKnn_wrapper_24_0__ap_start ap_done=krnl_partialKnn_wrapper_24_0__ap_done ap_idle=krnl_partialKnn_wrapper_24_0__ap_idle ap_ready=krnl_partialKnn_wrapper_24_0__ap_ready scalar=krnl_partialKnn_wrapper_24_0___.*
  // pragma RS ap-ctrl ap_start=krnl_partialKnn_wrapper_25_0__ap_start ap_done=krnl_partialKnn_wrapper_25_0__ap_done ap_idle=krnl_partialKnn_wrapper_25_0__ap_idle ap_ready=krnl_partialKnn_wrapper_25_0__ap_ready scalar=krnl_partialKnn_wrapper_25_0___.*
  // pragma RS ap-ctrl ap_start=krnl_partialKnn_wrapper_26_0__ap_start ap_done=krnl_partialKnn_wrapper_26_0__ap_done ap_idle=krnl_partialKnn_wrapper_26_0__ap_idle ap_ready=krnl_partialKnn_wrapper_26_0__ap_ready scalar=krnl_partialKnn_wrapper_26_0___.*
  // pragma RS ap-ctrl ap_start=krnl_partialKnn_wrapper_3_0__ap_start ap_done=krnl_partialKnn_wrapper_3_0__ap_done ap_idle=krnl_partialKnn_wrapper_3_0__ap_idle ap_ready=krnl_partialKnn_wrapper_3_0__ap_ready scalar=krnl_partialKnn_wrapper_3_0___.*
  // pragma RS ap-ctrl ap_start=krnl_partialKnn_wrapper_4_0__ap_start ap_done=krnl_partialKnn_wrapper_4_0__ap_done ap_idle=krnl_partialKnn_wrapper_4_0__ap_idle ap_ready=krnl_partialKnn_wrapper_4_0__ap_ready scalar=krnl_partialKnn_wrapper_4_0___.*
  // pragma RS ap-ctrl ap_start=krnl_partialKnn_wrapper_5_0__ap_start ap_done=krnl_partialKnn_wrapper_5_0__ap_done ap_idle=krnl_partialKnn_wrapper_5_0__ap_idle ap_ready=krnl_partialKnn_wrapper_5_0__ap_ready scalar=krnl_partialKnn_wrapper_5_0___.*
  // pragma RS ap-ctrl ap_start=krnl_partialKnn_wrapper_6_0__ap_start ap_done=krnl_partialKnn_wrapper_6_0__ap_done ap_idle=krnl_partialKnn_wrapper_6_0__ap_idle ap_ready=krnl_partialKnn_wrapper_6_0__ap_ready scalar=krnl_partialKnn_wrapper_6_0___.*
  // pragma RS ap-ctrl ap_start=krnl_partialKnn_wrapper_7_0__ap_start ap_done=krnl_partialKnn_wrapper_7_0__ap_done ap_idle=krnl_partialKnn_wrapper_7_0__ap_idle ap_ready=krnl_partialKnn_wrapper_7_0__ap_ready scalar=krnl_partialKnn_wrapper_7_0___.*
  // pragma RS ap-ctrl ap_start=krnl_partialKnn_wrapper_8_0__ap_start ap_done=krnl_partialKnn_wrapper_8_0__ap_done ap_idle=krnl_partialKnn_wrapper_8_0__ap_idle ap_ready=krnl_partialKnn_wrapper_8_0__ap_ready scalar=krnl_partialKnn_wrapper_8_0___.*
  // pragma RS ap-ctrl ap_start=krnl_partialKnn_wrapper_9_0__ap_start ap_done=krnl_partialKnn_wrapper_9_0__ap_done ap_idle=krnl_partialKnn_wrapper_9_0__ap_idle ap_ready=krnl_partialKnn_wrapper_9_0__ap_ready scalar=krnl_partialKnn_wrapper_9_0___.*

  input ap_clk;
  input ap_rst_n;
  input ap_start;
  output ap_ready;
  output ap_done;
  output ap_idle;
  input [63:0] L3_out_dist;
  input [63:0] L3_out_id;
  input [63:0] in_0;
  input [63:0] in_1;
  input [63:0] in_10;
  input [63:0] in_11;
  input [63:0] in_12;
  input [63:0] in_13;
  input [63:0] in_14;
  input [63:0] in_15;
  input [63:0] in_16;
  input [63:0] in_17;
  input [63:0] in_18;
  input [63:0] in_19;
  input [63:0] in_2;
  input [63:0] in_20;
  input [63:0] in_21;
  input [63:0] in_22;
  input [63:0] in_23;
  input [63:0] in_24;
  input [63:0] in_25;
  input [63:0] in_26;
  input [63:0] in_3;
  input [63:0] in_4;
  input [63:0] in_5;
  input [63:0] in_6;
  input [63:0] in_7;
  input [63:0] in_8;
  input [63:0] in_9;
  output krnl_globalSort_L1_L2_0__ap_start;
  input krnl_globalSort_L1_L2_0__ap_ready;
  input krnl_globalSort_L1_L2_0__ap_done;
  input krnl_globalSort_L1_L2_0__ap_idle;
  output krnl_globalSort_L1_L2_1__ap_start;
  input krnl_globalSort_L1_L2_1__ap_ready;
  input krnl_globalSort_L1_L2_1__ap_done;
  input krnl_globalSort_L1_L2_1__ap_idle;
  output krnl_globalSort_L1_L2_2__ap_start;
  input krnl_globalSort_L1_L2_2__ap_ready;
  input krnl_globalSort_L1_L2_2__ap_done;
  input krnl_globalSort_L1_L2_2__ap_idle;
  output krnl_globalSort_L1_L2_3__ap_start;
  input krnl_globalSort_L1_L2_3__ap_ready;
  input krnl_globalSort_L1_L2_3__ap_done;
  input krnl_globalSort_L1_L2_3__ap_idle;
  output krnl_globalSort_L1_L2_4__ap_start;
  input krnl_globalSort_L1_L2_4__ap_ready;
  input krnl_globalSort_L1_L2_4__ap_done;
  input krnl_globalSort_L1_L2_4__ap_idle;
  output krnl_globalSort_L1_L2_5__ap_start;
  input krnl_globalSort_L1_L2_5__ap_ready;
  input krnl_globalSort_L1_L2_5__ap_done;
  input krnl_globalSort_L1_L2_5__ap_idle;
  output krnl_globalSort_L1_L2_6__ap_start;
  input krnl_globalSort_L1_L2_6__ap_ready;
  input krnl_globalSort_L1_L2_6__ap_done;
  input krnl_globalSort_L1_L2_6__ap_idle;
  output krnl_globalSort_L1_L2_7__ap_start;
  input krnl_globalSort_L1_L2_7__ap_ready;
  input krnl_globalSort_L1_L2_7__ap_done;
  input krnl_globalSort_L1_L2_7__ap_idle;
  output krnl_globalSort_L1_L2_8__ap_start;
  input krnl_globalSort_L1_L2_8__ap_ready;
  input krnl_globalSort_L1_L2_8__ap_done;
  input krnl_globalSort_L1_L2_8__ap_idle;
  output krnl_globalSort_L1_L2_9__ap_start;
  input krnl_globalSort_L1_L2_9__ap_ready;
  input krnl_globalSort_L1_L2_9__ap_done;
  input krnl_globalSort_L1_L2_9__ap_idle;
  output krnl_globalSort_L1_L2_10__ap_start;
  input krnl_globalSort_L1_L2_10__ap_ready;
  input krnl_globalSort_L1_L2_10__ap_done;
  input krnl_globalSort_L1_L2_10__ap_idle;
  output krnl_globalSort_L1_L2_11__ap_start;
  input krnl_globalSort_L1_L2_11__ap_ready;
  input krnl_globalSort_L1_L2_11__ap_done;
  input krnl_globalSort_L1_L2_11__ap_idle;
  output krnl_globalSort_L1_L2_12__ap_start;
  input krnl_globalSort_L1_L2_12__ap_ready;
  input krnl_globalSort_L1_L2_12__ap_done;
  input krnl_globalSort_L1_L2_12__ap_idle;
  output [63:0] krnl_output_dist_id_0___L3_out_dist__q0;
  output [63:0] krnl_output_dist_id_0___L3_out_id__q0;
  output krnl_output_dist_id_0__ap_start;
  input krnl_output_dist_id_0__ap_ready;
  input krnl_output_dist_id_0__ap_done;
  input krnl_output_dist_id_0__ap_idle;
  output [63:0] krnl_partialKnn_wrapper_0_0___in_0__q0;
  output krnl_partialKnn_wrapper_0_0__ap_start;
  input krnl_partialKnn_wrapper_0_0__ap_ready;
  input krnl_partialKnn_wrapper_0_0__ap_done;
  input krnl_partialKnn_wrapper_0_0__ap_idle;
  output [63:0] krnl_partialKnn_wrapper_1_0___in_1__q0;
  output krnl_partialKnn_wrapper_1_0__ap_start;
  input krnl_partialKnn_wrapper_1_0__ap_ready;
  input krnl_partialKnn_wrapper_1_0__ap_done;
  input krnl_partialKnn_wrapper_1_0__ap_idle;
  output [63:0] krnl_partialKnn_wrapper_10_0___in_10__q0;
  output krnl_partialKnn_wrapper_10_0__ap_start;
  input krnl_partialKnn_wrapper_10_0__ap_ready;
  input krnl_partialKnn_wrapper_10_0__ap_done;
  input krnl_partialKnn_wrapper_10_0__ap_idle;
  output [63:0] krnl_partialKnn_wrapper_11_0___in_11__q0;
  output krnl_partialKnn_wrapper_11_0__ap_start;
  input krnl_partialKnn_wrapper_11_0__ap_ready;
  input krnl_partialKnn_wrapper_11_0__ap_done;
  input krnl_partialKnn_wrapper_11_0__ap_idle;
  output [63:0] krnl_partialKnn_wrapper_12_0___in_12__q0;
  output krnl_partialKnn_wrapper_12_0__ap_start;
  input krnl_partialKnn_wrapper_12_0__ap_ready;
  input krnl_partialKnn_wrapper_12_0__ap_done;
  input krnl_partialKnn_wrapper_12_0__ap_idle;
  output [63:0] krnl_partialKnn_wrapper_13_0___in_13__q0;
  output krnl_partialKnn_wrapper_13_0__ap_start;
  input krnl_partialKnn_wrapper_13_0__ap_ready;
  input krnl_partialKnn_wrapper_13_0__ap_done;
  input krnl_partialKnn_wrapper_13_0__ap_idle;
  output [63:0] krnl_partialKnn_wrapper_14_0___in_14__q0;
  output krnl_partialKnn_wrapper_14_0__ap_start;
  input krnl_partialKnn_wrapper_14_0__ap_ready;
  input krnl_partialKnn_wrapper_14_0__ap_done;
  input krnl_partialKnn_wrapper_14_0__ap_idle;
  output [63:0] krnl_partialKnn_wrapper_15_0___in_15__q0;
  output krnl_partialKnn_wrapper_15_0__ap_start;
  input krnl_partialKnn_wrapper_15_0__ap_ready;
  input krnl_partialKnn_wrapper_15_0__ap_done;
  input krnl_partialKnn_wrapper_15_0__ap_idle;
  output [63:0] krnl_partialKnn_wrapper_16_0___in_16__q0;
  output krnl_partialKnn_wrapper_16_0__ap_start;
  input krnl_partialKnn_wrapper_16_0__ap_ready;
  input krnl_partialKnn_wrapper_16_0__ap_done;
  input krnl_partialKnn_wrapper_16_0__ap_idle;
  output [63:0] krnl_partialKnn_wrapper_17_0___in_17__q0;
  output krnl_partialKnn_wrapper_17_0__ap_start;
  input krnl_partialKnn_wrapper_17_0__ap_ready;
  input krnl_partialKnn_wrapper_17_0__ap_done;
  input krnl_partialKnn_wrapper_17_0__ap_idle;
  output [63:0] krnl_partialKnn_wrapper_18_0___in_18__q0;
  output krnl_partialKnn_wrapper_18_0__ap_start;
  input krnl_partialKnn_wrapper_18_0__ap_ready;
  input krnl_partialKnn_wrapper_18_0__ap_done;
  input krnl_partialKnn_wrapper_18_0__ap_idle;
  output [63:0] krnl_partialKnn_wrapper_19_0___in_19__q0;
  output krnl_partialKnn_wrapper_19_0__ap_start;
  input krnl_partialKnn_wrapper_19_0__ap_ready;
  input krnl_partialKnn_wrapper_19_0__ap_done;
  input krnl_partialKnn_wrapper_19_0__ap_idle;
  output [63:0] krnl_partialKnn_wrapper_2_0___in_2__q0;
  output krnl_partialKnn_wrapper_2_0__ap_start;
  input krnl_partialKnn_wrapper_2_0__ap_ready;
  input krnl_partialKnn_wrapper_2_0__ap_done;
  input krnl_partialKnn_wrapper_2_0__ap_idle;
  output [63:0] krnl_partialKnn_wrapper_20_0___in_20__q0;
  output krnl_partialKnn_wrapper_20_0__ap_start;
  input krnl_partialKnn_wrapper_20_0__ap_ready;
  input krnl_partialKnn_wrapper_20_0__ap_done;
  input krnl_partialKnn_wrapper_20_0__ap_idle;
  output [63:0] krnl_partialKnn_wrapper_21_0___in_21__q0;
  output krnl_partialKnn_wrapper_21_0__ap_start;
  input krnl_partialKnn_wrapper_21_0__ap_ready;
  input krnl_partialKnn_wrapper_21_0__ap_done;
  input krnl_partialKnn_wrapper_21_0__ap_idle;
  output [63:0] krnl_partialKnn_wrapper_22_0___in_22__q0;
  output krnl_partialKnn_wrapper_22_0__ap_start;
  input krnl_partialKnn_wrapper_22_0__ap_ready;
  input krnl_partialKnn_wrapper_22_0__ap_done;
  input krnl_partialKnn_wrapper_22_0__ap_idle;
  output [63:0] krnl_partialKnn_wrapper_23_0___in_23__q0;
  output krnl_partialKnn_wrapper_23_0__ap_start;
  input krnl_partialKnn_wrapper_23_0__ap_ready;
  input krnl_partialKnn_wrapper_23_0__ap_done;
  input krnl_partialKnn_wrapper_23_0__ap_idle;
  output [63:0] krnl_partialKnn_wrapper_24_0___in_24__q0;
  output krnl_partialKnn_wrapper_24_0__ap_start;
  input krnl_partialKnn_wrapper_24_0__ap_ready;
  input krnl_partialKnn_wrapper_24_0__ap_done;
  input krnl_partialKnn_wrapper_24_0__ap_idle;
  output [63:0] krnl_partialKnn_wrapper_25_0___in_25__q0;
  output krnl_partialKnn_wrapper_25_0__ap_start;
  input krnl_partialKnn_wrapper_25_0__ap_ready;
  input krnl_partialKnn_wrapper_25_0__ap_done;
  input krnl_partialKnn_wrapper_25_0__ap_idle;
  output [63:0] krnl_partialKnn_wrapper_26_0___in_26__q0;
  output krnl_partialKnn_wrapper_26_0__ap_start;
  input krnl_partialKnn_wrapper_26_0__ap_ready;
  input krnl_partialKnn_wrapper_26_0__ap_done;
  input krnl_partialKnn_wrapper_26_0__ap_idle;
  output [63:0] krnl_partialKnn_wrapper_3_0___in_3__q0;
  output krnl_partialKnn_wrapper_3_0__ap_start;
  input krnl_partialKnn_wrapper_3_0__ap_ready;
  input krnl_partialKnn_wrapper_3_0__ap_done;
  input krnl_partialKnn_wrapper_3_0__ap_idle;
  output [63:0] krnl_partialKnn_wrapper_4_0___in_4__q0;
  output krnl_partialKnn_wrapper_4_0__ap_start;
  input krnl_partialKnn_wrapper_4_0__ap_ready;
  input krnl_partialKnn_wrapper_4_0__ap_done;
  input krnl_partialKnn_wrapper_4_0__ap_idle;
  output [63:0] krnl_partialKnn_wrapper_5_0___in_5__q0;
  output krnl_partialKnn_wrapper_5_0__ap_start;
  input krnl_partialKnn_wrapper_5_0__ap_ready;
  input krnl_partialKnn_wrapper_5_0__ap_done;
  input krnl_partialKnn_wrapper_5_0__ap_idle;
  output [63:0] krnl_partialKnn_wrapper_6_0___in_6__q0;
  output krnl_partialKnn_wrapper_6_0__ap_start;
  input krnl_partialKnn_wrapper_6_0__ap_ready;
  input krnl_partialKnn_wrapper_6_0__ap_done;
  input krnl_partialKnn_wrapper_6_0__ap_idle;
  output [63:0] krnl_partialKnn_wrapper_7_0___in_7__q0;
  output krnl_partialKnn_wrapper_7_0__ap_start;
  input krnl_partialKnn_wrapper_7_0__ap_ready;
  input krnl_partialKnn_wrapper_7_0__ap_done;
  input krnl_partialKnn_wrapper_7_0__ap_idle;
  output [63:0] krnl_partialKnn_wrapper_8_0___in_8__q0;
  output krnl_partialKnn_wrapper_8_0__ap_start;
  input krnl_partialKnn_wrapper_8_0__ap_ready;
  input krnl_partialKnn_wrapper_8_0__ap_done;
  input krnl_partialKnn_wrapper_8_0__ap_idle;
  output [63:0] krnl_partialKnn_wrapper_9_0___in_9__q0;
  output krnl_partialKnn_wrapper_9_0__ap_start;
  input krnl_partialKnn_wrapper_9_0__ap_ready;
  input krnl_partialKnn_wrapper_9_0__ap_done;
  input krnl_partialKnn_wrapper_9_0__ap_idle;
  wire krnl_globalSort_L1_L2_0__ap_start_global__q0;
  wire krnl_globalSort_L1_L2_0__is_done__q0;
  wire krnl_globalSort_L1_L2_0__ap_done_global__q0;
  wire krnl_globalSort_L1_L2_0__ap_start;
  wire krnl_globalSort_L1_L2_0__ap_ready;
  wire krnl_globalSort_L1_L2_0__ap_done;
  wire krnl_globalSort_L1_L2_0__ap_idle;
  reg [1:0] krnl_globalSort_L1_L2_0__state;
  wire krnl_globalSort_L1_L2_1__ap_start_global__q0;
  wire krnl_globalSort_L1_L2_1__is_done__q0;
  wire krnl_globalSort_L1_L2_1__ap_done_global__q0;
  wire krnl_globalSort_L1_L2_1__ap_start;
  wire krnl_globalSort_L1_L2_1__ap_ready;
  wire krnl_globalSort_L1_L2_1__ap_done;
  wire krnl_globalSort_L1_L2_1__ap_idle;
  reg [1:0] krnl_globalSort_L1_L2_1__state;
  wire krnl_globalSort_L1_L2_2__ap_start_global__q0;
  wire krnl_globalSort_L1_L2_2__is_done__q0;
  wire krnl_globalSort_L1_L2_2__ap_done_global__q0;
  wire krnl_globalSort_L1_L2_2__ap_start;
  wire krnl_globalSort_L1_L2_2__ap_ready;
  wire krnl_globalSort_L1_L2_2__ap_done;
  wire krnl_globalSort_L1_L2_2__ap_idle;
  reg [1:0] krnl_globalSort_L1_L2_2__state;
  wire krnl_globalSort_L1_L2_3__ap_start_global__q0;
  wire krnl_globalSort_L1_L2_3__is_done__q0;
  wire krnl_globalSort_L1_L2_3__ap_done_global__q0;
  wire krnl_globalSort_L1_L2_3__ap_start;
  wire krnl_globalSort_L1_L2_3__ap_ready;
  wire krnl_globalSort_L1_L2_3__ap_done;
  wire krnl_globalSort_L1_L2_3__ap_idle;
  reg [1:0] krnl_globalSort_L1_L2_3__state;
  wire krnl_globalSort_L1_L2_4__ap_start_global__q0;
  wire krnl_globalSort_L1_L2_4__is_done__q0;
  wire krnl_globalSort_L1_L2_4__ap_done_global__q0;
  wire krnl_globalSort_L1_L2_4__ap_start;
  wire krnl_globalSort_L1_L2_4__ap_ready;
  wire krnl_globalSort_L1_L2_4__ap_done;
  wire krnl_globalSort_L1_L2_4__ap_idle;
  reg [1:0] krnl_globalSort_L1_L2_4__state;
  wire krnl_globalSort_L1_L2_5__ap_start_global__q0;
  wire krnl_globalSort_L1_L2_5__is_done__q0;
  wire krnl_globalSort_L1_L2_5__ap_done_global__q0;
  wire krnl_globalSort_L1_L2_5__ap_start;
  wire krnl_globalSort_L1_L2_5__ap_ready;
  wire krnl_globalSort_L1_L2_5__ap_done;
  wire krnl_globalSort_L1_L2_5__ap_idle;
  reg [1:0] krnl_globalSort_L1_L2_5__state;
  wire krnl_globalSort_L1_L2_6__ap_start_global__q0;
  wire krnl_globalSort_L1_L2_6__is_done__q0;
  wire krnl_globalSort_L1_L2_6__ap_done_global__q0;
  wire krnl_globalSort_L1_L2_6__ap_start;
  wire krnl_globalSort_L1_L2_6__ap_ready;
  wire krnl_globalSort_L1_L2_6__ap_done;
  wire krnl_globalSort_L1_L2_6__ap_idle;
  reg [1:0] krnl_globalSort_L1_L2_6__state;
  wire krnl_globalSort_L1_L2_7__ap_start_global__q0;
  wire krnl_globalSort_L1_L2_7__is_done__q0;
  wire krnl_globalSort_L1_L2_7__ap_done_global__q0;
  wire krnl_globalSort_L1_L2_7__ap_start;
  wire krnl_globalSort_L1_L2_7__ap_ready;
  wire krnl_globalSort_L1_L2_7__ap_done;
  wire krnl_globalSort_L1_L2_7__ap_idle;
  reg [1:0] krnl_globalSort_L1_L2_7__state;
  wire krnl_globalSort_L1_L2_8__ap_start_global__q0;
  wire krnl_globalSort_L1_L2_8__is_done__q0;
  wire krnl_globalSort_L1_L2_8__ap_done_global__q0;
  wire krnl_globalSort_L1_L2_8__ap_start;
  wire krnl_globalSort_L1_L2_8__ap_ready;
  wire krnl_globalSort_L1_L2_8__ap_done;
  wire krnl_globalSort_L1_L2_8__ap_idle;
  reg [1:0] krnl_globalSort_L1_L2_8__state;
  wire krnl_globalSort_L1_L2_9__ap_start_global__q0;
  wire krnl_globalSort_L1_L2_9__is_done__q0;
  wire krnl_globalSort_L1_L2_9__ap_done_global__q0;
  wire krnl_globalSort_L1_L2_9__ap_start;
  wire krnl_globalSort_L1_L2_9__ap_ready;
  wire krnl_globalSort_L1_L2_9__ap_done;
  wire krnl_globalSort_L1_L2_9__ap_idle;
  reg [1:0] krnl_globalSort_L1_L2_9__state;
  wire krnl_globalSort_L1_L2_10__ap_start_global__q0;
  wire krnl_globalSort_L1_L2_10__is_done__q0;
  wire krnl_globalSort_L1_L2_10__ap_done_global__q0;
  wire krnl_globalSort_L1_L2_10__ap_start;
  wire krnl_globalSort_L1_L2_10__ap_ready;
  wire krnl_globalSort_L1_L2_10__ap_done;
  wire krnl_globalSort_L1_L2_10__ap_idle;
  reg [1:0] krnl_globalSort_L1_L2_10__state;
  wire krnl_globalSort_L1_L2_11__ap_start_global__q0;
  wire krnl_globalSort_L1_L2_11__is_done__q0;
  wire krnl_globalSort_L1_L2_11__ap_done_global__q0;
  wire krnl_globalSort_L1_L2_11__ap_start;
  wire krnl_globalSort_L1_L2_11__ap_ready;
  wire krnl_globalSort_L1_L2_11__ap_done;
  wire krnl_globalSort_L1_L2_11__ap_idle;
  reg [1:0] krnl_globalSort_L1_L2_11__state;
  wire krnl_globalSort_L1_L2_12__ap_start_global__q0;
  wire krnl_globalSort_L1_L2_12__is_done__q0;
  wire krnl_globalSort_L1_L2_12__ap_done_global__q0;
  wire krnl_globalSort_L1_L2_12__ap_start;
  wire krnl_globalSort_L1_L2_12__ap_ready;
  wire krnl_globalSort_L1_L2_12__ap_done;
  wire krnl_globalSort_L1_L2_12__ap_idle;
  reg [1:0] krnl_globalSort_L1_L2_12__state;
  wire [63:0] krnl_output_dist_id_0___L3_out_dist__q0;
  wire [63:0] krnl_output_dist_id_0___L3_out_id__q0;
  wire krnl_output_dist_id_0__ap_start_global__q0;
  wire krnl_output_dist_id_0__is_done__q0;
  wire krnl_output_dist_id_0__ap_done_global__q0;
  wire krnl_output_dist_id_0__ap_start;
  wire krnl_output_dist_id_0__ap_ready;
  wire krnl_output_dist_id_0__ap_done;
  wire krnl_output_dist_id_0__ap_idle;
  reg [1:0] krnl_output_dist_id_0__state;
  wire [63:0] krnl_partialKnn_wrapper_0_0___in_0__q0;
  wire krnl_partialKnn_wrapper_0_0__ap_start_global__q0;
  wire krnl_partialKnn_wrapper_0_0__is_done__q0;
  wire krnl_partialKnn_wrapper_0_0__ap_done_global__q0;
  wire krnl_partialKnn_wrapper_0_0__ap_start;
  wire krnl_partialKnn_wrapper_0_0__ap_ready;
  wire krnl_partialKnn_wrapper_0_0__ap_done;
  wire krnl_partialKnn_wrapper_0_0__ap_idle;
  reg [1:0] krnl_partialKnn_wrapper_0_0__state;
  wire [63:0] krnl_partialKnn_wrapper_1_0___in_1__q0;
  wire krnl_partialKnn_wrapper_1_0__ap_start_global__q0;
  wire krnl_partialKnn_wrapper_1_0__is_done__q0;
  wire krnl_partialKnn_wrapper_1_0__ap_done_global__q0;
  wire krnl_partialKnn_wrapper_1_0__ap_start;
  wire krnl_partialKnn_wrapper_1_0__ap_ready;
  wire krnl_partialKnn_wrapper_1_0__ap_done;
  wire krnl_partialKnn_wrapper_1_0__ap_idle;
  reg [1:0] krnl_partialKnn_wrapper_1_0__state;
  wire [63:0] krnl_partialKnn_wrapper_10_0___in_10__q0;
  wire krnl_partialKnn_wrapper_10_0__ap_start_global__q0;
  wire krnl_partialKnn_wrapper_10_0__is_done__q0;
  wire krnl_partialKnn_wrapper_10_0__ap_done_global__q0;
  wire krnl_partialKnn_wrapper_10_0__ap_start;
  wire krnl_partialKnn_wrapper_10_0__ap_ready;
  wire krnl_partialKnn_wrapper_10_0__ap_done;
  wire krnl_partialKnn_wrapper_10_0__ap_idle;
  reg [1:0] krnl_partialKnn_wrapper_10_0__state;
  wire [63:0] krnl_partialKnn_wrapper_11_0___in_11__q0;
  wire krnl_partialKnn_wrapper_11_0__ap_start_global__q0;
  wire krnl_partialKnn_wrapper_11_0__is_done__q0;
  wire krnl_partialKnn_wrapper_11_0__ap_done_global__q0;
  wire krnl_partialKnn_wrapper_11_0__ap_start;
  wire krnl_partialKnn_wrapper_11_0__ap_ready;
  wire krnl_partialKnn_wrapper_11_0__ap_done;
  wire krnl_partialKnn_wrapper_11_0__ap_idle;
  reg [1:0] krnl_partialKnn_wrapper_11_0__state;
  wire [63:0] krnl_partialKnn_wrapper_12_0___in_12__q0;
  wire krnl_partialKnn_wrapper_12_0__ap_start_global__q0;
  wire krnl_partialKnn_wrapper_12_0__is_done__q0;
  wire krnl_partialKnn_wrapper_12_0__ap_done_global__q0;
  wire krnl_partialKnn_wrapper_12_0__ap_start;
  wire krnl_partialKnn_wrapper_12_0__ap_ready;
  wire krnl_partialKnn_wrapper_12_0__ap_done;
  wire krnl_partialKnn_wrapper_12_0__ap_idle;
  reg [1:0] krnl_partialKnn_wrapper_12_0__state;
  wire [63:0] krnl_partialKnn_wrapper_13_0___in_13__q0;
  wire krnl_partialKnn_wrapper_13_0__ap_start_global__q0;
  wire krnl_partialKnn_wrapper_13_0__is_done__q0;
  wire krnl_partialKnn_wrapper_13_0__ap_done_global__q0;
  wire krnl_partialKnn_wrapper_13_0__ap_start;
  wire krnl_partialKnn_wrapper_13_0__ap_ready;
  wire krnl_partialKnn_wrapper_13_0__ap_done;
  wire krnl_partialKnn_wrapper_13_0__ap_idle;
  reg [1:0] krnl_partialKnn_wrapper_13_0__state;
  wire [63:0] krnl_partialKnn_wrapper_14_0___in_14__q0;
  wire krnl_partialKnn_wrapper_14_0__ap_start_global__q0;
  wire krnl_partialKnn_wrapper_14_0__is_done__q0;
  wire krnl_partialKnn_wrapper_14_0__ap_done_global__q0;
  wire krnl_partialKnn_wrapper_14_0__ap_start;
  wire krnl_partialKnn_wrapper_14_0__ap_ready;
  wire krnl_partialKnn_wrapper_14_0__ap_done;
  wire krnl_partialKnn_wrapper_14_0__ap_idle;
  reg [1:0] krnl_partialKnn_wrapper_14_0__state;
  wire [63:0] krnl_partialKnn_wrapper_15_0___in_15__q0;
  wire krnl_partialKnn_wrapper_15_0__ap_start_global__q0;
  wire krnl_partialKnn_wrapper_15_0__is_done__q0;
  wire krnl_partialKnn_wrapper_15_0__ap_done_global__q0;
  wire krnl_partialKnn_wrapper_15_0__ap_start;
  wire krnl_partialKnn_wrapper_15_0__ap_ready;
  wire krnl_partialKnn_wrapper_15_0__ap_done;
  wire krnl_partialKnn_wrapper_15_0__ap_idle;
  reg [1:0] krnl_partialKnn_wrapper_15_0__state;
  wire [63:0] krnl_partialKnn_wrapper_16_0___in_16__q0;
  wire krnl_partialKnn_wrapper_16_0__ap_start_global__q0;
  wire krnl_partialKnn_wrapper_16_0__is_done__q0;
  wire krnl_partialKnn_wrapper_16_0__ap_done_global__q0;
  wire krnl_partialKnn_wrapper_16_0__ap_start;
  wire krnl_partialKnn_wrapper_16_0__ap_ready;
  wire krnl_partialKnn_wrapper_16_0__ap_done;
  wire krnl_partialKnn_wrapper_16_0__ap_idle;
  reg [1:0] krnl_partialKnn_wrapper_16_0__state;
  wire [63:0] krnl_partialKnn_wrapper_17_0___in_17__q0;
  wire krnl_partialKnn_wrapper_17_0__ap_start_global__q0;
  wire krnl_partialKnn_wrapper_17_0__is_done__q0;
  wire krnl_partialKnn_wrapper_17_0__ap_done_global__q0;
  wire krnl_partialKnn_wrapper_17_0__ap_start;
  wire krnl_partialKnn_wrapper_17_0__ap_ready;
  wire krnl_partialKnn_wrapper_17_0__ap_done;
  wire krnl_partialKnn_wrapper_17_0__ap_idle;
  reg [1:0] krnl_partialKnn_wrapper_17_0__state;
  wire [63:0] krnl_partialKnn_wrapper_18_0___in_18__q0;
  wire krnl_partialKnn_wrapper_18_0__ap_start_global__q0;
  wire krnl_partialKnn_wrapper_18_0__is_done__q0;
  wire krnl_partialKnn_wrapper_18_0__ap_done_global__q0;
  wire krnl_partialKnn_wrapper_18_0__ap_start;
  wire krnl_partialKnn_wrapper_18_0__ap_ready;
  wire krnl_partialKnn_wrapper_18_0__ap_done;
  wire krnl_partialKnn_wrapper_18_0__ap_idle;
  reg [1:0] krnl_partialKnn_wrapper_18_0__state;
  wire [63:0] krnl_partialKnn_wrapper_19_0___in_19__q0;
  wire krnl_partialKnn_wrapper_19_0__ap_start_global__q0;
  wire krnl_partialKnn_wrapper_19_0__is_done__q0;
  wire krnl_partialKnn_wrapper_19_0__ap_done_global__q0;
  wire krnl_partialKnn_wrapper_19_0__ap_start;
  wire krnl_partialKnn_wrapper_19_0__ap_ready;
  wire krnl_partialKnn_wrapper_19_0__ap_done;
  wire krnl_partialKnn_wrapper_19_0__ap_idle;
  reg [1:0] krnl_partialKnn_wrapper_19_0__state;
  wire [63:0] krnl_partialKnn_wrapper_2_0___in_2__q0;
  wire krnl_partialKnn_wrapper_2_0__ap_start_global__q0;
  wire krnl_partialKnn_wrapper_2_0__is_done__q0;
  wire krnl_partialKnn_wrapper_2_0__ap_done_global__q0;
  wire krnl_partialKnn_wrapper_2_0__ap_start;
  wire krnl_partialKnn_wrapper_2_0__ap_ready;
  wire krnl_partialKnn_wrapper_2_0__ap_done;
  wire krnl_partialKnn_wrapper_2_0__ap_idle;
  reg [1:0] krnl_partialKnn_wrapper_2_0__state;
  wire [63:0] krnl_partialKnn_wrapper_20_0___in_20__q0;
  wire krnl_partialKnn_wrapper_20_0__ap_start_global__q0;
  wire krnl_partialKnn_wrapper_20_0__is_done__q0;
  wire krnl_partialKnn_wrapper_20_0__ap_done_global__q0;
  wire krnl_partialKnn_wrapper_20_0__ap_start;
  wire krnl_partialKnn_wrapper_20_0__ap_ready;
  wire krnl_partialKnn_wrapper_20_0__ap_done;
  wire krnl_partialKnn_wrapper_20_0__ap_idle;
  reg [1:0] krnl_partialKnn_wrapper_20_0__state;
  wire [63:0] krnl_partialKnn_wrapper_21_0___in_21__q0;
  wire krnl_partialKnn_wrapper_21_0__ap_start_global__q0;
  wire krnl_partialKnn_wrapper_21_0__is_done__q0;
  wire krnl_partialKnn_wrapper_21_0__ap_done_global__q0;
  wire krnl_partialKnn_wrapper_21_0__ap_start;
  wire krnl_partialKnn_wrapper_21_0__ap_ready;
  wire krnl_partialKnn_wrapper_21_0__ap_done;
  wire krnl_partialKnn_wrapper_21_0__ap_idle;
  reg [1:0] krnl_partialKnn_wrapper_21_0__state;
  wire [63:0] krnl_partialKnn_wrapper_22_0___in_22__q0;
  wire krnl_partialKnn_wrapper_22_0__ap_start_global__q0;
  wire krnl_partialKnn_wrapper_22_0__is_done__q0;
  wire krnl_partialKnn_wrapper_22_0__ap_done_global__q0;
  wire krnl_partialKnn_wrapper_22_0__ap_start;
  wire krnl_partialKnn_wrapper_22_0__ap_ready;
  wire krnl_partialKnn_wrapper_22_0__ap_done;
  wire krnl_partialKnn_wrapper_22_0__ap_idle;
  reg [1:0] krnl_partialKnn_wrapper_22_0__state;
  wire [63:0] krnl_partialKnn_wrapper_23_0___in_23__q0;
  wire krnl_partialKnn_wrapper_23_0__ap_start_global__q0;
  wire krnl_partialKnn_wrapper_23_0__is_done__q0;
  wire krnl_partialKnn_wrapper_23_0__ap_done_global__q0;
  wire krnl_partialKnn_wrapper_23_0__ap_start;
  wire krnl_partialKnn_wrapper_23_0__ap_ready;
  wire krnl_partialKnn_wrapper_23_0__ap_done;
  wire krnl_partialKnn_wrapper_23_0__ap_idle;
  reg [1:0] krnl_partialKnn_wrapper_23_0__state;
  wire [63:0] krnl_partialKnn_wrapper_24_0___in_24__q0;
  wire krnl_partialKnn_wrapper_24_0__ap_start_global__q0;
  wire krnl_partialKnn_wrapper_24_0__is_done__q0;
  wire krnl_partialKnn_wrapper_24_0__ap_done_global__q0;
  wire krnl_partialKnn_wrapper_24_0__ap_start;
  wire krnl_partialKnn_wrapper_24_0__ap_ready;
  wire krnl_partialKnn_wrapper_24_0__ap_done;
  wire krnl_partialKnn_wrapper_24_0__ap_idle;
  reg [1:0] krnl_partialKnn_wrapper_24_0__state;
  wire [63:0] krnl_partialKnn_wrapper_25_0___in_25__q0;
  wire krnl_partialKnn_wrapper_25_0__ap_start_global__q0;
  wire krnl_partialKnn_wrapper_25_0__is_done__q0;
  wire krnl_partialKnn_wrapper_25_0__ap_done_global__q0;
  wire krnl_partialKnn_wrapper_25_0__ap_start;
  wire krnl_partialKnn_wrapper_25_0__ap_ready;
  wire krnl_partialKnn_wrapper_25_0__ap_done;
  wire krnl_partialKnn_wrapper_25_0__ap_idle;
  reg [1:0] krnl_partialKnn_wrapper_25_0__state;
  wire [63:0] krnl_partialKnn_wrapper_26_0___in_26__q0;
  wire krnl_partialKnn_wrapper_26_0__ap_start_global__q0;
  wire krnl_partialKnn_wrapper_26_0__is_done__q0;
  wire krnl_partialKnn_wrapper_26_0__ap_done_global__q0;
  wire krnl_partialKnn_wrapper_26_0__ap_start;
  wire krnl_partialKnn_wrapper_26_0__ap_ready;
  wire krnl_partialKnn_wrapper_26_0__ap_done;
  wire krnl_partialKnn_wrapper_26_0__ap_idle;
  reg [1:0] krnl_partialKnn_wrapper_26_0__state;
  wire [63:0] krnl_partialKnn_wrapper_3_0___in_3__q0;
  wire krnl_partialKnn_wrapper_3_0__ap_start_global__q0;
  wire krnl_partialKnn_wrapper_3_0__is_done__q0;
  wire krnl_partialKnn_wrapper_3_0__ap_done_global__q0;
  wire krnl_partialKnn_wrapper_3_0__ap_start;
  wire krnl_partialKnn_wrapper_3_0__ap_ready;
  wire krnl_partialKnn_wrapper_3_0__ap_done;
  wire krnl_partialKnn_wrapper_3_0__ap_idle;
  reg [1:0] krnl_partialKnn_wrapper_3_0__state;
  wire [63:0] krnl_partialKnn_wrapper_4_0___in_4__q0;
  wire krnl_partialKnn_wrapper_4_0__ap_start_global__q0;
  wire krnl_partialKnn_wrapper_4_0__is_done__q0;
  wire krnl_partialKnn_wrapper_4_0__ap_done_global__q0;
  wire krnl_partialKnn_wrapper_4_0__ap_start;
  wire krnl_partialKnn_wrapper_4_0__ap_ready;
  wire krnl_partialKnn_wrapper_4_0__ap_done;
  wire krnl_partialKnn_wrapper_4_0__ap_idle;
  reg [1:0] krnl_partialKnn_wrapper_4_0__state;
  wire [63:0] krnl_partialKnn_wrapper_5_0___in_5__q0;
  wire krnl_partialKnn_wrapper_5_0__ap_start_global__q0;
  wire krnl_partialKnn_wrapper_5_0__is_done__q0;
  wire krnl_partialKnn_wrapper_5_0__ap_done_global__q0;
  wire krnl_partialKnn_wrapper_5_0__ap_start;
  wire krnl_partialKnn_wrapper_5_0__ap_ready;
  wire krnl_partialKnn_wrapper_5_0__ap_done;
  wire krnl_partialKnn_wrapper_5_0__ap_idle;
  reg [1:0] krnl_partialKnn_wrapper_5_0__state;
  wire [63:0] krnl_partialKnn_wrapper_6_0___in_6__q0;
  wire krnl_partialKnn_wrapper_6_0__ap_start_global__q0;
  wire krnl_partialKnn_wrapper_6_0__is_done__q0;
  wire krnl_partialKnn_wrapper_6_0__ap_done_global__q0;
  wire krnl_partialKnn_wrapper_6_0__ap_start;
  wire krnl_partialKnn_wrapper_6_0__ap_ready;
  wire krnl_partialKnn_wrapper_6_0__ap_done;
  wire krnl_partialKnn_wrapper_6_0__ap_idle;
  reg [1:0] krnl_partialKnn_wrapper_6_0__state;
  wire [63:0] krnl_partialKnn_wrapper_7_0___in_7__q0;
  wire krnl_partialKnn_wrapper_7_0__ap_start_global__q0;
  wire krnl_partialKnn_wrapper_7_0__is_done__q0;
  wire krnl_partialKnn_wrapper_7_0__ap_done_global__q0;
  wire krnl_partialKnn_wrapper_7_0__ap_start;
  wire krnl_partialKnn_wrapper_7_0__ap_ready;
  wire krnl_partialKnn_wrapper_7_0__ap_done;
  wire krnl_partialKnn_wrapper_7_0__ap_idle;
  reg [1:0] krnl_partialKnn_wrapper_7_0__state;
  wire [63:0] krnl_partialKnn_wrapper_8_0___in_8__q0;
  wire krnl_partialKnn_wrapper_8_0__ap_start_global__q0;
  wire krnl_partialKnn_wrapper_8_0__is_done__q0;
  wire krnl_partialKnn_wrapper_8_0__ap_done_global__q0;
  wire krnl_partialKnn_wrapper_8_0__ap_start;
  wire krnl_partialKnn_wrapper_8_0__ap_ready;
  wire krnl_partialKnn_wrapper_8_0__ap_done;
  wire krnl_partialKnn_wrapper_8_0__ap_idle;
  reg [1:0] krnl_partialKnn_wrapper_8_0__state;
  wire [63:0] krnl_partialKnn_wrapper_9_0___in_9__q0;
  wire krnl_partialKnn_wrapper_9_0__ap_start_global__q0;
  wire krnl_partialKnn_wrapper_9_0__is_done__q0;
  wire krnl_partialKnn_wrapper_9_0__ap_done_global__q0;
  wire krnl_partialKnn_wrapper_9_0__ap_start;
  wire krnl_partialKnn_wrapper_9_0__ap_ready;
  wire krnl_partialKnn_wrapper_9_0__ap_done;
  wire krnl_partialKnn_wrapper_9_0__ap_idle;
  reg [1:0] krnl_partialKnn_wrapper_9_0__state;
  reg [1:0] tapa_state;
  reg [0:0] countdown;
  wire ap_start__q0;
  wire ap_done__q0;
  assign krnl_globalSort_L1_L2_0__ap_start_global__q0 = ap_start__q0;
  assign krnl_globalSort_L1_L2_0__is_done__q0 = (krnl_globalSort_L1_L2_0__state == 2'b10);
  assign krnl_globalSort_L1_L2_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      krnl_globalSort_L1_L2_0__state <= 2'b00;
    end else begin
      if(krnl_globalSort_L1_L2_0__state == 2'b00) begin
        if(krnl_globalSort_L1_L2_0__ap_start_global__q0) begin
          krnl_globalSort_L1_L2_0__state <= 2'b01;
        end 
      end 
      if(krnl_globalSort_L1_L2_0__state == 2'b01) begin
        if(krnl_globalSort_L1_L2_0__ap_ready) begin
          if(krnl_globalSort_L1_L2_0__ap_done) begin
            krnl_globalSort_L1_L2_0__state <= 2'b10;
          end else begin
            krnl_globalSort_L1_L2_0__state <= 2'b11;
          end
        end 
      end 
      if(krnl_globalSort_L1_L2_0__state == 2'b11) begin
        if(krnl_globalSort_L1_L2_0__ap_done) begin
          krnl_globalSort_L1_L2_0__state <= 2'b10;
        end 
      end 
      if(krnl_globalSort_L1_L2_0__state == 2'b10) begin
        if(krnl_globalSort_L1_L2_0__ap_done_global__q0) begin
          krnl_globalSort_L1_L2_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign krnl_globalSort_L1_L2_0__ap_start = (krnl_globalSort_L1_L2_0__state == 2'b01);
  assign krnl_globalSort_L1_L2_1__ap_start_global__q0 = ap_start__q0;
  assign krnl_globalSort_L1_L2_1__is_done__q0 = (krnl_globalSort_L1_L2_1__state == 2'b10);
  assign krnl_globalSort_L1_L2_1__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      krnl_globalSort_L1_L2_1__state <= 2'b00;
    end else begin
      if(krnl_globalSort_L1_L2_1__state == 2'b00) begin
        if(krnl_globalSort_L1_L2_1__ap_start_global__q0) begin
          krnl_globalSort_L1_L2_1__state <= 2'b01;
        end 
      end 
      if(krnl_globalSort_L1_L2_1__state == 2'b01) begin
        if(krnl_globalSort_L1_L2_1__ap_ready) begin
          if(krnl_globalSort_L1_L2_1__ap_done) begin
            krnl_globalSort_L1_L2_1__state <= 2'b10;
          end else begin
            krnl_globalSort_L1_L2_1__state <= 2'b11;
          end
        end 
      end 
      if(krnl_globalSort_L1_L2_1__state == 2'b11) begin
        if(krnl_globalSort_L1_L2_1__ap_done) begin
          krnl_globalSort_L1_L2_1__state <= 2'b10;
        end 
      end 
      if(krnl_globalSort_L1_L2_1__state == 2'b10) begin
        if(krnl_globalSort_L1_L2_1__ap_done_global__q0) begin
          krnl_globalSort_L1_L2_1__state <= 2'b00;
        end 
      end 
    end
  end

  assign krnl_globalSort_L1_L2_1__ap_start = (krnl_globalSort_L1_L2_1__state == 2'b01);
  assign krnl_globalSort_L1_L2_2__ap_start_global__q0 = ap_start__q0;
  assign krnl_globalSort_L1_L2_2__is_done__q0 = (krnl_globalSort_L1_L2_2__state == 2'b10);
  assign krnl_globalSort_L1_L2_2__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      krnl_globalSort_L1_L2_2__state <= 2'b00;
    end else begin
      if(krnl_globalSort_L1_L2_2__state == 2'b00) begin
        if(krnl_globalSort_L1_L2_2__ap_start_global__q0) begin
          krnl_globalSort_L1_L2_2__state <= 2'b01;
        end 
      end 
      if(krnl_globalSort_L1_L2_2__state == 2'b01) begin
        if(krnl_globalSort_L1_L2_2__ap_ready) begin
          if(krnl_globalSort_L1_L2_2__ap_done) begin
            krnl_globalSort_L1_L2_2__state <= 2'b10;
          end else begin
            krnl_globalSort_L1_L2_2__state <= 2'b11;
          end
        end 
      end 
      if(krnl_globalSort_L1_L2_2__state == 2'b11) begin
        if(krnl_globalSort_L1_L2_2__ap_done) begin
          krnl_globalSort_L1_L2_2__state <= 2'b10;
        end 
      end 
      if(krnl_globalSort_L1_L2_2__state == 2'b10) begin
        if(krnl_globalSort_L1_L2_2__ap_done_global__q0) begin
          krnl_globalSort_L1_L2_2__state <= 2'b00;
        end 
      end 
    end
  end

  assign krnl_globalSort_L1_L2_2__ap_start = (krnl_globalSort_L1_L2_2__state == 2'b01);
  assign krnl_globalSort_L1_L2_3__ap_start_global__q0 = ap_start__q0;
  assign krnl_globalSort_L1_L2_3__is_done__q0 = (krnl_globalSort_L1_L2_3__state == 2'b10);
  assign krnl_globalSort_L1_L2_3__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      krnl_globalSort_L1_L2_3__state <= 2'b00;
    end else begin
      if(krnl_globalSort_L1_L2_3__state == 2'b00) begin
        if(krnl_globalSort_L1_L2_3__ap_start_global__q0) begin
          krnl_globalSort_L1_L2_3__state <= 2'b01;
        end 
      end 
      if(krnl_globalSort_L1_L2_3__state == 2'b01) begin
        if(krnl_globalSort_L1_L2_3__ap_ready) begin
          if(krnl_globalSort_L1_L2_3__ap_done) begin
            krnl_globalSort_L1_L2_3__state <= 2'b10;
          end else begin
            krnl_globalSort_L1_L2_3__state <= 2'b11;
          end
        end 
      end 
      if(krnl_globalSort_L1_L2_3__state == 2'b11) begin
        if(krnl_globalSort_L1_L2_3__ap_done) begin
          krnl_globalSort_L1_L2_3__state <= 2'b10;
        end 
      end 
      if(krnl_globalSort_L1_L2_3__state == 2'b10) begin
        if(krnl_globalSort_L1_L2_3__ap_done_global__q0) begin
          krnl_globalSort_L1_L2_3__state <= 2'b00;
        end 
      end 
    end
  end

  assign krnl_globalSort_L1_L2_3__ap_start = (krnl_globalSort_L1_L2_3__state == 2'b01);
  assign krnl_globalSort_L1_L2_4__ap_start_global__q0 = ap_start__q0;
  assign krnl_globalSort_L1_L2_4__is_done__q0 = (krnl_globalSort_L1_L2_4__state == 2'b10);
  assign krnl_globalSort_L1_L2_4__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      krnl_globalSort_L1_L2_4__state <= 2'b00;
    end else begin
      if(krnl_globalSort_L1_L2_4__state == 2'b00) begin
        if(krnl_globalSort_L1_L2_4__ap_start_global__q0) begin
          krnl_globalSort_L1_L2_4__state <= 2'b01;
        end 
      end 
      if(krnl_globalSort_L1_L2_4__state == 2'b01) begin
        if(krnl_globalSort_L1_L2_4__ap_ready) begin
          if(krnl_globalSort_L1_L2_4__ap_done) begin
            krnl_globalSort_L1_L2_4__state <= 2'b10;
          end else begin
            krnl_globalSort_L1_L2_4__state <= 2'b11;
          end
        end 
      end 
      if(krnl_globalSort_L1_L2_4__state == 2'b11) begin
        if(krnl_globalSort_L1_L2_4__ap_done) begin
          krnl_globalSort_L1_L2_4__state <= 2'b10;
        end 
      end 
      if(krnl_globalSort_L1_L2_4__state == 2'b10) begin
        if(krnl_globalSort_L1_L2_4__ap_done_global__q0) begin
          krnl_globalSort_L1_L2_4__state <= 2'b00;
        end 
      end 
    end
  end

  assign krnl_globalSort_L1_L2_4__ap_start = (krnl_globalSort_L1_L2_4__state == 2'b01);
  assign krnl_globalSort_L1_L2_5__ap_start_global__q0 = ap_start__q0;
  assign krnl_globalSort_L1_L2_5__is_done__q0 = (krnl_globalSort_L1_L2_5__state == 2'b10);
  assign krnl_globalSort_L1_L2_5__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      krnl_globalSort_L1_L2_5__state <= 2'b00;
    end else begin
      if(krnl_globalSort_L1_L2_5__state == 2'b00) begin
        if(krnl_globalSort_L1_L2_5__ap_start_global__q0) begin
          krnl_globalSort_L1_L2_5__state <= 2'b01;
        end 
      end 
      if(krnl_globalSort_L1_L2_5__state == 2'b01) begin
        if(krnl_globalSort_L1_L2_5__ap_ready) begin
          if(krnl_globalSort_L1_L2_5__ap_done) begin
            krnl_globalSort_L1_L2_5__state <= 2'b10;
          end else begin
            krnl_globalSort_L1_L2_5__state <= 2'b11;
          end
        end 
      end 
      if(krnl_globalSort_L1_L2_5__state == 2'b11) begin
        if(krnl_globalSort_L1_L2_5__ap_done) begin
          krnl_globalSort_L1_L2_5__state <= 2'b10;
        end 
      end 
      if(krnl_globalSort_L1_L2_5__state == 2'b10) begin
        if(krnl_globalSort_L1_L2_5__ap_done_global__q0) begin
          krnl_globalSort_L1_L2_5__state <= 2'b00;
        end 
      end 
    end
  end

  assign krnl_globalSort_L1_L2_5__ap_start = (krnl_globalSort_L1_L2_5__state == 2'b01);
  assign krnl_globalSort_L1_L2_6__ap_start_global__q0 = ap_start__q0;
  assign krnl_globalSort_L1_L2_6__is_done__q0 = (krnl_globalSort_L1_L2_6__state == 2'b10);
  assign krnl_globalSort_L1_L2_6__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      krnl_globalSort_L1_L2_6__state <= 2'b00;
    end else begin
      if(krnl_globalSort_L1_L2_6__state == 2'b00) begin
        if(krnl_globalSort_L1_L2_6__ap_start_global__q0) begin
          krnl_globalSort_L1_L2_6__state <= 2'b01;
        end 
      end 
      if(krnl_globalSort_L1_L2_6__state == 2'b01) begin
        if(krnl_globalSort_L1_L2_6__ap_ready) begin
          if(krnl_globalSort_L1_L2_6__ap_done) begin
            krnl_globalSort_L1_L2_6__state <= 2'b10;
          end else begin
            krnl_globalSort_L1_L2_6__state <= 2'b11;
          end
        end 
      end 
      if(krnl_globalSort_L1_L2_6__state == 2'b11) begin
        if(krnl_globalSort_L1_L2_6__ap_done) begin
          krnl_globalSort_L1_L2_6__state <= 2'b10;
        end 
      end 
      if(krnl_globalSort_L1_L2_6__state == 2'b10) begin
        if(krnl_globalSort_L1_L2_6__ap_done_global__q0) begin
          krnl_globalSort_L1_L2_6__state <= 2'b00;
        end 
      end 
    end
  end

  assign krnl_globalSort_L1_L2_6__ap_start = (krnl_globalSort_L1_L2_6__state == 2'b01);
  assign krnl_globalSort_L1_L2_7__ap_start_global__q0 = ap_start__q0;
  assign krnl_globalSort_L1_L2_7__is_done__q0 = (krnl_globalSort_L1_L2_7__state == 2'b10);
  assign krnl_globalSort_L1_L2_7__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      krnl_globalSort_L1_L2_7__state <= 2'b00;
    end else begin
      if(krnl_globalSort_L1_L2_7__state == 2'b00) begin
        if(krnl_globalSort_L1_L2_7__ap_start_global__q0) begin
          krnl_globalSort_L1_L2_7__state <= 2'b01;
        end 
      end 
      if(krnl_globalSort_L1_L2_7__state == 2'b01) begin
        if(krnl_globalSort_L1_L2_7__ap_ready) begin
          if(krnl_globalSort_L1_L2_7__ap_done) begin
            krnl_globalSort_L1_L2_7__state <= 2'b10;
          end else begin
            krnl_globalSort_L1_L2_7__state <= 2'b11;
          end
        end 
      end 
      if(krnl_globalSort_L1_L2_7__state == 2'b11) begin
        if(krnl_globalSort_L1_L2_7__ap_done) begin
          krnl_globalSort_L1_L2_7__state <= 2'b10;
        end 
      end 
      if(krnl_globalSort_L1_L2_7__state == 2'b10) begin
        if(krnl_globalSort_L1_L2_7__ap_done_global__q0) begin
          krnl_globalSort_L1_L2_7__state <= 2'b00;
        end 
      end 
    end
  end

  assign krnl_globalSort_L1_L2_7__ap_start = (krnl_globalSort_L1_L2_7__state == 2'b01);
  assign krnl_globalSort_L1_L2_8__ap_start_global__q0 = ap_start__q0;
  assign krnl_globalSort_L1_L2_8__is_done__q0 = (krnl_globalSort_L1_L2_8__state == 2'b10);
  assign krnl_globalSort_L1_L2_8__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      krnl_globalSort_L1_L2_8__state <= 2'b00;
    end else begin
      if(krnl_globalSort_L1_L2_8__state == 2'b00) begin
        if(krnl_globalSort_L1_L2_8__ap_start_global__q0) begin
          krnl_globalSort_L1_L2_8__state <= 2'b01;
        end 
      end 
      if(krnl_globalSort_L1_L2_8__state == 2'b01) begin
        if(krnl_globalSort_L1_L2_8__ap_ready) begin
          if(krnl_globalSort_L1_L2_8__ap_done) begin
            krnl_globalSort_L1_L2_8__state <= 2'b10;
          end else begin
            krnl_globalSort_L1_L2_8__state <= 2'b11;
          end
        end 
      end 
      if(krnl_globalSort_L1_L2_8__state == 2'b11) begin
        if(krnl_globalSort_L1_L2_8__ap_done) begin
          krnl_globalSort_L1_L2_8__state <= 2'b10;
        end 
      end 
      if(krnl_globalSort_L1_L2_8__state == 2'b10) begin
        if(krnl_globalSort_L1_L2_8__ap_done_global__q0) begin
          krnl_globalSort_L1_L2_8__state <= 2'b00;
        end 
      end 
    end
  end

  assign krnl_globalSort_L1_L2_8__ap_start = (krnl_globalSort_L1_L2_8__state == 2'b01);
  assign krnl_globalSort_L1_L2_9__ap_start_global__q0 = ap_start__q0;
  assign krnl_globalSort_L1_L2_9__is_done__q0 = (krnl_globalSort_L1_L2_9__state == 2'b10);
  assign krnl_globalSort_L1_L2_9__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      krnl_globalSort_L1_L2_9__state <= 2'b00;
    end else begin
      if(krnl_globalSort_L1_L2_9__state == 2'b00) begin
        if(krnl_globalSort_L1_L2_9__ap_start_global__q0) begin
          krnl_globalSort_L1_L2_9__state <= 2'b01;
        end 
      end 
      if(krnl_globalSort_L1_L2_9__state == 2'b01) begin
        if(krnl_globalSort_L1_L2_9__ap_ready) begin
          if(krnl_globalSort_L1_L2_9__ap_done) begin
            krnl_globalSort_L1_L2_9__state <= 2'b10;
          end else begin
            krnl_globalSort_L1_L2_9__state <= 2'b11;
          end
        end 
      end 
      if(krnl_globalSort_L1_L2_9__state == 2'b11) begin
        if(krnl_globalSort_L1_L2_9__ap_done) begin
          krnl_globalSort_L1_L2_9__state <= 2'b10;
        end 
      end 
      if(krnl_globalSort_L1_L2_9__state == 2'b10) begin
        if(krnl_globalSort_L1_L2_9__ap_done_global__q0) begin
          krnl_globalSort_L1_L2_9__state <= 2'b00;
        end 
      end 
    end
  end

  assign krnl_globalSort_L1_L2_9__ap_start = (krnl_globalSort_L1_L2_9__state == 2'b01);
  assign krnl_globalSort_L1_L2_10__ap_start_global__q0 = ap_start__q0;
  assign krnl_globalSort_L1_L2_10__is_done__q0 = (krnl_globalSort_L1_L2_10__state == 2'b10);
  assign krnl_globalSort_L1_L2_10__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      krnl_globalSort_L1_L2_10__state <= 2'b00;
    end else begin
      if(krnl_globalSort_L1_L2_10__state == 2'b00) begin
        if(krnl_globalSort_L1_L2_10__ap_start_global__q0) begin
          krnl_globalSort_L1_L2_10__state <= 2'b01;
        end 
      end 
      if(krnl_globalSort_L1_L2_10__state == 2'b01) begin
        if(krnl_globalSort_L1_L2_10__ap_ready) begin
          if(krnl_globalSort_L1_L2_10__ap_done) begin
            krnl_globalSort_L1_L2_10__state <= 2'b10;
          end else begin
            krnl_globalSort_L1_L2_10__state <= 2'b11;
          end
        end 
      end 
      if(krnl_globalSort_L1_L2_10__state == 2'b11) begin
        if(krnl_globalSort_L1_L2_10__ap_done) begin
          krnl_globalSort_L1_L2_10__state <= 2'b10;
        end 
      end 
      if(krnl_globalSort_L1_L2_10__state == 2'b10) begin
        if(krnl_globalSort_L1_L2_10__ap_done_global__q0) begin
          krnl_globalSort_L1_L2_10__state <= 2'b00;
        end 
      end 
    end
  end

  assign krnl_globalSort_L1_L2_10__ap_start = (krnl_globalSort_L1_L2_10__state == 2'b01);
  assign krnl_globalSort_L1_L2_11__ap_start_global__q0 = ap_start__q0;
  assign krnl_globalSort_L1_L2_11__is_done__q0 = (krnl_globalSort_L1_L2_11__state == 2'b10);
  assign krnl_globalSort_L1_L2_11__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      krnl_globalSort_L1_L2_11__state <= 2'b00;
    end else begin
      if(krnl_globalSort_L1_L2_11__state == 2'b00) begin
        if(krnl_globalSort_L1_L2_11__ap_start_global__q0) begin
          krnl_globalSort_L1_L2_11__state <= 2'b01;
        end 
      end 
      if(krnl_globalSort_L1_L2_11__state == 2'b01) begin
        if(krnl_globalSort_L1_L2_11__ap_ready) begin
          if(krnl_globalSort_L1_L2_11__ap_done) begin
            krnl_globalSort_L1_L2_11__state <= 2'b10;
          end else begin
            krnl_globalSort_L1_L2_11__state <= 2'b11;
          end
        end 
      end 
      if(krnl_globalSort_L1_L2_11__state == 2'b11) begin
        if(krnl_globalSort_L1_L2_11__ap_done) begin
          krnl_globalSort_L1_L2_11__state <= 2'b10;
        end 
      end 
      if(krnl_globalSort_L1_L2_11__state == 2'b10) begin
        if(krnl_globalSort_L1_L2_11__ap_done_global__q0) begin
          krnl_globalSort_L1_L2_11__state <= 2'b00;
        end 
      end 
    end
  end

  assign krnl_globalSort_L1_L2_11__ap_start = (krnl_globalSort_L1_L2_11__state == 2'b01);
  assign krnl_globalSort_L1_L2_12__ap_start_global__q0 = ap_start__q0;
  assign krnl_globalSort_L1_L2_12__is_done__q0 = (krnl_globalSort_L1_L2_12__state == 2'b10);
  assign krnl_globalSort_L1_L2_12__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      krnl_globalSort_L1_L2_12__state <= 2'b00;
    end else begin
      if(krnl_globalSort_L1_L2_12__state == 2'b00) begin
        if(krnl_globalSort_L1_L2_12__ap_start_global__q0) begin
          krnl_globalSort_L1_L2_12__state <= 2'b01;
        end 
      end 
      if(krnl_globalSort_L1_L2_12__state == 2'b01) begin
        if(krnl_globalSort_L1_L2_12__ap_ready) begin
          if(krnl_globalSort_L1_L2_12__ap_done) begin
            krnl_globalSort_L1_L2_12__state <= 2'b10;
          end else begin
            krnl_globalSort_L1_L2_12__state <= 2'b11;
          end
        end 
      end 
      if(krnl_globalSort_L1_L2_12__state == 2'b11) begin
        if(krnl_globalSort_L1_L2_12__ap_done) begin
          krnl_globalSort_L1_L2_12__state <= 2'b10;
        end 
      end 
      if(krnl_globalSort_L1_L2_12__state == 2'b10) begin
        if(krnl_globalSort_L1_L2_12__ap_done_global__q0) begin
          krnl_globalSort_L1_L2_12__state <= 2'b00;
        end 
      end 
    end
  end

  assign krnl_globalSort_L1_L2_12__ap_start = (krnl_globalSort_L1_L2_12__state == 2'b01);
  assign krnl_output_dist_id_0___L3_out_dist__q0 = L3_out_dist;
  assign krnl_output_dist_id_0___L3_out_id__q0 = L3_out_id;
  assign krnl_output_dist_id_0__ap_start_global__q0 = ap_start__q0;
  assign krnl_output_dist_id_0__is_done__q0 = (krnl_output_dist_id_0__state == 2'b10);
  assign krnl_output_dist_id_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      krnl_output_dist_id_0__state <= 2'b00;
    end else begin
      if(krnl_output_dist_id_0__state == 2'b00) begin
        if(krnl_output_dist_id_0__ap_start_global__q0) begin
          krnl_output_dist_id_0__state <= 2'b01;
        end 
      end 
      if(krnl_output_dist_id_0__state == 2'b01) begin
        if(krnl_output_dist_id_0__ap_ready) begin
          if(krnl_output_dist_id_0__ap_done) begin
            krnl_output_dist_id_0__state <= 2'b10;
          end else begin
            krnl_output_dist_id_0__state <= 2'b11;
          end
        end 
      end 
      if(krnl_output_dist_id_0__state == 2'b11) begin
        if(krnl_output_dist_id_0__ap_done) begin
          krnl_output_dist_id_0__state <= 2'b10;
        end 
      end 
      if(krnl_output_dist_id_0__state == 2'b10) begin
        if(krnl_output_dist_id_0__ap_done_global__q0) begin
          krnl_output_dist_id_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign krnl_output_dist_id_0__ap_start = (krnl_output_dist_id_0__state == 2'b01);
  assign krnl_partialKnn_wrapper_0_0___in_0__q0 = in_0;
  assign krnl_partialKnn_wrapper_0_0__ap_start_global__q0 = ap_start__q0;
  assign krnl_partialKnn_wrapper_0_0__is_done__q0 = (krnl_partialKnn_wrapper_0_0__state == 2'b10);
  assign krnl_partialKnn_wrapper_0_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      krnl_partialKnn_wrapper_0_0__state <= 2'b00;
    end else begin
      if(krnl_partialKnn_wrapper_0_0__state == 2'b00) begin
        if(krnl_partialKnn_wrapper_0_0__ap_start_global__q0) begin
          krnl_partialKnn_wrapper_0_0__state <= 2'b01;
        end 
      end 
      if(krnl_partialKnn_wrapper_0_0__state == 2'b01) begin
        if(krnl_partialKnn_wrapper_0_0__ap_ready) begin
          if(krnl_partialKnn_wrapper_0_0__ap_done) begin
            krnl_partialKnn_wrapper_0_0__state <= 2'b10;
          end else begin
            krnl_partialKnn_wrapper_0_0__state <= 2'b11;
          end
        end 
      end 
      if(krnl_partialKnn_wrapper_0_0__state == 2'b11) begin
        if(krnl_partialKnn_wrapper_0_0__ap_done) begin
          krnl_partialKnn_wrapper_0_0__state <= 2'b10;
        end 
      end 
      if(krnl_partialKnn_wrapper_0_0__state == 2'b10) begin
        if(krnl_partialKnn_wrapper_0_0__ap_done_global__q0) begin
          krnl_partialKnn_wrapper_0_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign krnl_partialKnn_wrapper_0_0__ap_start = (krnl_partialKnn_wrapper_0_0__state == 2'b01);
  assign krnl_partialKnn_wrapper_1_0___in_1__q0 = in_1;
  assign krnl_partialKnn_wrapper_1_0__ap_start_global__q0 = ap_start__q0;
  assign krnl_partialKnn_wrapper_1_0__is_done__q0 = (krnl_partialKnn_wrapper_1_0__state == 2'b10);
  assign krnl_partialKnn_wrapper_1_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      krnl_partialKnn_wrapper_1_0__state <= 2'b00;
    end else begin
      if(krnl_partialKnn_wrapper_1_0__state == 2'b00) begin
        if(krnl_partialKnn_wrapper_1_0__ap_start_global__q0) begin
          krnl_partialKnn_wrapper_1_0__state <= 2'b01;
        end 
      end 
      if(krnl_partialKnn_wrapper_1_0__state == 2'b01) begin
        if(krnl_partialKnn_wrapper_1_0__ap_ready) begin
          if(krnl_partialKnn_wrapper_1_0__ap_done) begin
            krnl_partialKnn_wrapper_1_0__state <= 2'b10;
          end else begin
            krnl_partialKnn_wrapper_1_0__state <= 2'b11;
          end
        end 
      end 
      if(krnl_partialKnn_wrapper_1_0__state == 2'b11) begin
        if(krnl_partialKnn_wrapper_1_0__ap_done) begin
          krnl_partialKnn_wrapper_1_0__state <= 2'b10;
        end 
      end 
      if(krnl_partialKnn_wrapper_1_0__state == 2'b10) begin
        if(krnl_partialKnn_wrapper_1_0__ap_done_global__q0) begin
          krnl_partialKnn_wrapper_1_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign krnl_partialKnn_wrapper_1_0__ap_start = (krnl_partialKnn_wrapper_1_0__state == 2'b01);
  assign krnl_partialKnn_wrapper_10_0___in_10__q0 = in_10;
  assign krnl_partialKnn_wrapper_10_0__ap_start_global__q0 = ap_start__q0;
  assign krnl_partialKnn_wrapper_10_0__is_done__q0 = (krnl_partialKnn_wrapper_10_0__state == 2'b10);
  assign krnl_partialKnn_wrapper_10_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      krnl_partialKnn_wrapper_10_0__state <= 2'b00;
    end else begin
      if(krnl_partialKnn_wrapper_10_0__state == 2'b00) begin
        if(krnl_partialKnn_wrapper_10_0__ap_start_global__q0) begin
          krnl_partialKnn_wrapper_10_0__state <= 2'b01;
        end 
      end 
      if(krnl_partialKnn_wrapper_10_0__state == 2'b01) begin
        if(krnl_partialKnn_wrapper_10_0__ap_ready) begin
          if(krnl_partialKnn_wrapper_10_0__ap_done) begin
            krnl_partialKnn_wrapper_10_0__state <= 2'b10;
          end else begin
            krnl_partialKnn_wrapper_10_0__state <= 2'b11;
          end
        end 
      end 
      if(krnl_partialKnn_wrapper_10_0__state == 2'b11) begin
        if(krnl_partialKnn_wrapper_10_0__ap_done) begin
          krnl_partialKnn_wrapper_10_0__state <= 2'b10;
        end 
      end 
      if(krnl_partialKnn_wrapper_10_0__state == 2'b10) begin
        if(krnl_partialKnn_wrapper_10_0__ap_done_global__q0) begin
          krnl_partialKnn_wrapper_10_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign krnl_partialKnn_wrapper_10_0__ap_start = (krnl_partialKnn_wrapper_10_0__state == 2'b01);
  assign krnl_partialKnn_wrapper_11_0___in_11__q0 = in_11;
  assign krnl_partialKnn_wrapper_11_0__ap_start_global__q0 = ap_start__q0;
  assign krnl_partialKnn_wrapper_11_0__is_done__q0 = (krnl_partialKnn_wrapper_11_0__state == 2'b10);
  assign krnl_partialKnn_wrapper_11_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      krnl_partialKnn_wrapper_11_0__state <= 2'b00;
    end else begin
      if(krnl_partialKnn_wrapper_11_0__state == 2'b00) begin
        if(krnl_partialKnn_wrapper_11_0__ap_start_global__q0) begin
          krnl_partialKnn_wrapper_11_0__state <= 2'b01;
        end 
      end 
      if(krnl_partialKnn_wrapper_11_0__state == 2'b01) begin
        if(krnl_partialKnn_wrapper_11_0__ap_ready) begin
          if(krnl_partialKnn_wrapper_11_0__ap_done) begin
            krnl_partialKnn_wrapper_11_0__state <= 2'b10;
          end else begin
            krnl_partialKnn_wrapper_11_0__state <= 2'b11;
          end
        end 
      end 
      if(krnl_partialKnn_wrapper_11_0__state == 2'b11) begin
        if(krnl_partialKnn_wrapper_11_0__ap_done) begin
          krnl_partialKnn_wrapper_11_0__state <= 2'b10;
        end 
      end 
      if(krnl_partialKnn_wrapper_11_0__state == 2'b10) begin
        if(krnl_partialKnn_wrapper_11_0__ap_done_global__q0) begin
          krnl_partialKnn_wrapper_11_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign krnl_partialKnn_wrapper_11_0__ap_start = (krnl_partialKnn_wrapper_11_0__state == 2'b01);
  assign krnl_partialKnn_wrapper_12_0___in_12__q0 = in_12;
  assign krnl_partialKnn_wrapper_12_0__ap_start_global__q0 = ap_start__q0;
  assign krnl_partialKnn_wrapper_12_0__is_done__q0 = (krnl_partialKnn_wrapper_12_0__state == 2'b10);
  assign krnl_partialKnn_wrapper_12_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      krnl_partialKnn_wrapper_12_0__state <= 2'b00;
    end else begin
      if(krnl_partialKnn_wrapper_12_0__state == 2'b00) begin
        if(krnl_partialKnn_wrapper_12_0__ap_start_global__q0) begin
          krnl_partialKnn_wrapper_12_0__state <= 2'b01;
        end 
      end 
      if(krnl_partialKnn_wrapper_12_0__state == 2'b01) begin
        if(krnl_partialKnn_wrapper_12_0__ap_ready) begin
          if(krnl_partialKnn_wrapper_12_0__ap_done) begin
            krnl_partialKnn_wrapper_12_0__state <= 2'b10;
          end else begin
            krnl_partialKnn_wrapper_12_0__state <= 2'b11;
          end
        end 
      end 
      if(krnl_partialKnn_wrapper_12_0__state == 2'b11) begin
        if(krnl_partialKnn_wrapper_12_0__ap_done) begin
          krnl_partialKnn_wrapper_12_0__state <= 2'b10;
        end 
      end 
      if(krnl_partialKnn_wrapper_12_0__state == 2'b10) begin
        if(krnl_partialKnn_wrapper_12_0__ap_done_global__q0) begin
          krnl_partialKnn_wrapper_12_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign krnl_partialKnn_wrapper_12_0__ap_start = (krnl_partialKnn_wrapper_12_0__state == 2'b01);
  assign krnl_partialKnn_wrapper_13_0___in_13__q0 = in_13;
  assign krnl_partialKnn_wrapper_13_0__ap_start_global__q0 = ap_start__q0;
  assign krnl_partialKnn_wrapper_13_0__is_done__q0 = (krnl_partialKnn_wrapper_13_0__state == 2'b10);
  assign krnl_partialKnn_wrapper_13_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      krnl_partialKnn_wrapper_13_0__state <= 2'b00;
    end else begin
      if(krnl_partialKnn_wrapper_13_0__state == 2'b00) begin
        if(krnl_partialKnn_wrapper_13_0__ap_start_global__q0) begin
          krnl_partialKnn_wrapper_13_0__state <= 2'b01;
        end 
      end 
      if(krnl_partialKnn_wrapper_13_0__state == 2'b01) begin
        if(krnl_partialKnn_wrapper_13_0__ap_ready) begin
          if(krnl_partialKnn_wrapper_13_0__ap_done) begin
            krnl_partialKnn_wrapper_13_0__state <= 2'b10;
          end else begin
            krnl_partialKnn_wrapper_13_0__state <= 2'b11;
          end
        end 
      end 
      if(krnl_partialKnn_wrapper_13_0__state == 2'b11) begin
        if(krnl_partialKnn_wrapper_13_0__ap_done) begin
          krnl_partialKnn_wrapper_13_0__state <= 2'b10;
        end 
      end 
      if(krnl_partialKnn_wrapper_13_0__state == 2'b10) begin
        if(krnl_partialKnn_wrapper_13_0__ap_done_global__q0) begin
          krnl_partialKnn_wrapper_13_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign krnl_partialKnn_wrapper_13_0__ap_start = (krnl_partialKnn_wrapper_13_0__state == 2'b01);
  assign krnl_partialKnn_wrapper_14_0___in_14__q0 = in_14;
  assign krnl_partialKnn_wrapper_14_0__ap_start_global__q0 = ap_start__q0;
  assign krnl_partialKnn_wrapper_14_0__is_done__q0 = (krnl_partialKnn_wrapper_14_0__state == 2'b10);
  assign krnl_partialKnn_wrapper_14_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      krnl_partialKnn_wrapper_14_0__state <= 2'b00;
    end else begin
      if(krnl_partialKnn_wrapper_14_0__state == 2'b00) begin
        if(krnl_partialKnn_wrapper_14_0__ap_start_global__q0) begin
          krnl_partialKnn_wrapper_14_0__state <= 2'b01;
        end 
      end 
      if(krnl_partialKnn_wrapper_14_0__state == 2'b01) begin
        if(krnl_partialKnn_wrapper_14_0__ap_ready) begin
          if(krnl_partialKnn_wrapper_14_0__ap_done) begin
            krnl_partialKnn_wrapper_14_0__state <= 2'b10;
          end else begin
            krnl_partialKnn_wrapper_14_0__state <= 2'b11;
          end
        end 
      end 
      if(krnl_partialKnn_wrapper_14_0__state == 2'b11) begin
        if(krnl_partialKnn_wrapper_14_0__ap_done) begin
          krnl_partialKnn_wrapper_14_0__state <= 2'b10;
        end 
      end 
      if(krnl_partialKnn_wrapper_14_0__state == 2'b10) begin
        if(krnl_partialKnn_wrapper_14_0__ap_done_global__q0) begin
          krnl_partialKnn_wrapper_14_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign krnl_partialKnn_wrapper_14_0__ap_start = (krnl_partialKnn_wrapper_14_0__state == 2'b01);
  assign krnl_partialKnn_wrapper_15_0___in_15__q0 = in_15;
  assign krnl_partialKnn_wrapper_15_0__ap_start_global__q0 = ap_start__q0;
  assign krnl_partialKnn_wrapper_15_0__is_done__q0 = (krnl_partialKnn_wrapper_15_0__state == 2'b10);
  assign krnl_partialKnn_wrapper_15_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      krnl_partialKnn_wrapper_15_0__state <= 2'b00;
    end else begin
      if(krnl_partialKnn_wrapper_15_0__state == 2'b00) begin
        if(krnl_partialKnn_wrapper_15_0__ap_start_global__q0) begin
          krnl_partialKnn_wrapper_15_0__state <= 2'b01;
        end 
      end 
      if(krnl_partialKnn_wrapper_15_0__state == 2'b01) begin
        if(krnl_partialKnn_wrapper_15_0__ap_ready) begin
          if(krnl_partialKnn_wrapper_15_0__ap_done) begin
            krnl_partialKnn_wrapper_15_0__state <= 2'b10;
          end else begin
            krnl_partialKnn_wrapper_15_0__state <= 2'b11;
          end
        end 
      end 
      if(krnl_partialKnn_wrapper_15_0__state == 2'b11) begin
        if(krnl_partialKnn_wrapper_15_0__ap_done) begin
          krnl_partialKnn_wrapper_15_0__state <= 2'b10;
        end 
      end 
      if(krnl_partialKnn_wrapper_15_0__state == 2'b10) begin
        if(krnl_partialKnn_wrapper_15_0__ap_done_global__q0) begin
          krnl_partialKnn_wrapper_15_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign krnl_partialKnn_wrapper_15_0__ap_start = (krnl_partialKnn_wrapper_15_0__state == 2'b01);
  assign krnl_partialKnn_wrapper_16_0___in_16__q0 = in_16;
  assign krnl_partialKnn_wrapper_16_0__ap_start_global__q0 = ap_start__q0;
  assign krnl_partialKnn_wrapper_16_0__is_done__q0 = (krnl_partialKnn_wrapper_16_0__state == 2'b10);
  assign krnl_partialKnn_wrapper_16_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      krnl_partialKnn_wrapper_16_0__state <= 2'b00;
    end else begin
      if(krnl_partialKnn_wrapper_16_0__state == 2'b00) begin
        if(krnl_partialKnn_wrapper_16_0__ap_start_global__q0) begin
          krnl_partialKnn_wrapper_16_0__state <= 2'b01;
        end 
      end 
      if(krnl_partialKnn_wrapper_16_0__state == 2'b01) begin
        if(krnl_partialKnn_wrapper_16_0__ap_ready) begin
          if(krnl_partialKnn_wrapper_16_0__ap_done) begin
            krnl_partialKnn_wrapper_16_0__state <= 2'b10;
          end else begin
            krnl_partialKnn_wrapper_16_0__state <= 2'b11;
          end
        end 
      end 
      if(krnl_partialKnn_wrapper_16_0__state == 2'b11) begin
        if(krnl_partialKnn_wrapper_16_0__ap_done) begin
          krnl_partialKnn_wrapper_16_0__state <= 2'b10;
        end 
      end 
      if(krnl_partialKnn_wrapper_16_0__state == 2'b10) begin
        if(krnl_partialKnn_wrapper_16_0__ap_done_global__q0) begin
          krnl_partialKnn_wrapper_16_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign krnl_partialKnn_wrapper_16_0__ap_start = (krnl_partialKnn_wrapper_16_0__state == 2'b01);
  assign krnl_partialKnn_wrapper_17_0___in_17__q0 = in_17;
  assign krnl_partialKnn_wrapper_17_0__ap_start_global__q0 = ap_start__q0;
  assign krnl_partialKnn_wrapper_17_0__is_done__q0 = (krnl_partialKnn_wrapper_17_0__state == 2'b10);
  assign krnl_partialKnn_wrapper_17_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      krnl_partialKnn_wrapper_17_0__state <= 2'b00;
    end else begin
      if(krnl_partialKnn_wrapper_17_0__state == 2'b00) begin
        if(krnl_partialKnn_wrapper_17_0__ap_start_global__q0) begin
          krnl_partialKnn_wrapper_17_0__state <= 2'b01;
        end 
      end 
      if(krnl_partialKnn_wrapper_17_0__state == 2'b01) begin
        if(krnl_partialKnn_wrapper_17_0__ap_ready) begin
          if(krnl_partialKnn_wrapper_17_0__ap_done) begin
            krnl_partialKnn_wrapper_17_0__state <= 2'b10;
          end else begin
            krnl_partialKnn_wrapper_17_0__state <= 2'b11;
          end
        end 
      end 
      if(krnl_partialKnn_wrapper_17_0__state == 2'b11) begin
        if(krnl_partialKnn_wrapper_17_0__ap_done) begin
          krnl_partialKnn_wrapper_17_0__state <= 2'b10;
        end 
      end 
      if(krnl_partialKnn_wrapper_17_0__state == 2'b10) begin
        if(krnl_partialKnn_wrapper_17_0__ap_done_global__q0) begin
          krnl_partialKnn_wrapper_17_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign krnl_partialKnn_wrapper_17_0__ap_start = (krnl_partialKnn_wrapper_17_0__state == 2'b01);
  assign krnl_partialKnn_wrapper_18_0___in_18__q0 = in_18;
  assign krnl_partialKnn_wrapper_18_0__ap_start_global__q0 = ap_start__q0;
  assign krnl_partialKnn_wrapper_18_0__is_done__q0 = (krnl_partialKnn_wrapper_18_0__state == 2'b10);
  assign krnl_partialKnn_wrapper_18_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      krnl_partialKnn_wrapper_18_0__state <= 2'b00;
    end else begin
      if(krnl_partialKnn_wrapper_18_0__state == 2'b00) begin
        if(krnl_partialKnn_wrapper_18_0__ap_start_global__q0) begin
          krnl_partialKnn_wrapper_18_0__state <= 2'b01;
        end 
      end 
      if(krnl_partialKnn_wrapper_18_0__state == 2'b01) begin
        if(krnl_partialKnn_wrapper_18_0__ap_ready) begin
          if(krnl_partialKnn_wrapper_18_0__ap_done) begin
            krnl_partialKnn_wrapper_18_0__state <= 2'b10;
          end else begin
            krnl_partialKnn_wrapper_18_0__state <= 2'b11;
          end
        end 
      end 
      if(krnl_partialKnn_wrapper_18_0__state == 2'b11) begin
        if(krnl_partialKnn_wrapper_18_0__ap_done) begin
          krnl_partialKnn_wrapper_18_0__state <= 2'b10;
        end 
      end 
      if(krnl_partialKnn_wrapper_18_0__state == 2'b10) begin
        if(krnl_partialKnn_wrapper_18_0__ap_done_global__q0) begin
          krnl_partialKnn_wrapper_18_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign krnl_partialKnn_wrapper_18_0__ap_start = (krnl_partialKnn_wrapper_18_0__state == 2'b01);
  assign krnl_partialKnn_wrapper_19_0___in_19__q0 = in_19;
  assign krnl_partialKnn_wrapper_19_0__ap_start_global__q0 = ap_start__q0;
  assign krnl_partialKnn_wrapper_19_0__is_done__q0 = (krnl_partialKnn_wrapper_19_0__state == 2'b10);
  assign krnl_partialKnn_wrapper_19_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      krnl_partialKnn_wrapper_19_0__state <= 2'b00;
    end else begin
      if(krnl_partialKnn_wrapper_19_0__state == 2'b00) begin
        if(krnl_partialKnn_wrapper_19_0__ap_start_global__q0) begin
          krnl_partialKnn_wrapper_19_0__state <= 2'b01;
        end 
      end 
      if(krnl_partialKnn_wrapper_19_0__state == 2'b01) begin
        if(krnl_partialKnn_wrapper_19_0__ap_ready) begin
          if(krnl_partialKnn_wrapper_19_0__ap_done) begin
            krnl_partialKnn_wrapper_19_0__state <= 2'b10;
          end else begin
            krnl_partialKnn_wrapper_19_0__state <= 2'b11;
          end
        end 
      end 
      if(krnl_partialKnn_wrapper_19_0__state == 2'b11) begin
        if(krnl_partialKnn_wrapper_19_0__ap_done) begin
          krnl_partialKnn_wrapper_19_0__state <= 2'b10;
        end 
      end 
      if(krnl_partialKnn_wrapper_19_0__state == 2'b10) begin
        if(krnl_partialKnn_wrapper_19_0__ap_done_global__q0) begin
          krnl_partialKnn_wrapper_19_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign krnl_partialKnn_wrapper_19_0__ap_start = (krnl_partialKnn_wrapper_19_0__state == 2'b01);
  assign krnl_partialKnn_wrapper_2_0___in_2__q0 = in_2;
  assign krnl_partialKnn_wrapper_2_0__ap_start_global__q0 = ap_start__q0;
  assign krnl_partialKnn_wrapper_2_0__is_done__q0 = (krnl_partialKnn_wrapper_2_0__state == 2'b10);
  assign krnl_partialKnn_wrapper_2_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      krnl_partialKnn_wrapper_2_0__state <= 2'b00;
    end else begin
      if(krnl_partialKnn_wrapper_2_0__state == 2'b00) begin
        if(krnl_partialKnn_wrapper_2_0__ap_start_global__q0) begin
          krnl_partialKnn_wrapper_2_0__state <= 2'b01;
        end 
      end 
      if(krnl_partialKnn_wrapper_2_0__state == 2'b01) begin
        if(krnl_partialKnn_wrapper_2_0__ap_ready) begin
          if(krnl_partialKnn_wrapper_2_0__ap_done) begin
            krnl_partialKnn_wrapper_2_0__state <= 2'b10;
          end else begin
            krnl_partialKnn_wrapper_2_0__state <= 2'b11;
          end
        end 
      end 
      if(krnl_partialKnn_wrapper_2_0__state == 2'b11) begin
        if(krnl_partialKnn_wrapper_2_0__ap_done) begin
          krnl_partialKnn_wrapper_2_0__state <= 2'b10;
        end 
      end 
      if(krnl_partialKnn_wrapper_2_0__state == 2'b10) begin
        if(krnl_partialKnn_wrapper_2_0__ap_done_global__q0) begin
          krnl_partialKnn_wrapper_2_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign krnl_partialKnn_wrapper_2_0__ap_start = (krnl_partialKnn_wrapper_2_0__state == 2'b01);
  assign krnl_partialKnn_wrapper_20_0___in_20__q0 = in_20;
  assign krnl_partialKnn_wrapper_20_0__ap_start_global__q0 = ap_start__q0;
  assign krnl_partialKnn_wrapper_20_0__is_done__q0 = (krnl_partialKnn_wrapper_20_0__state == 2'b10);
  assign krnl_partialKnn_wrapper_20_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      krnl_partialKnn_wrapper_20_0__state <= 2'b00;
    end else begin
      if(krnl_partialKnn_wrapper_20_0__state == 2'b00) begin
        if(krnl_partialKnn_wrapper_20_0__ap_start_global__q0) begin
          krnl_partialKnn_wrapper_20_0__state <= 2'b01;
        end 
      end 
      if(krnl_partialKnn_wrapper_20_0__state == 2'b01) begin
        if(krnl_partialKnn_wrapper_20_0__ap_ready) begin
          if(krnl_partialKnn_wrapper_20_0__ap_done) begin
            krnl_partialKnn_wrapper_20_0__state <= 2'b10;
          end else begin
            krnl_partialKnn_wrapper_20_0__state <= 2'b11;
          end
        end 
      end 
      if(krnl_partialKnn_wrapper_20_0__state == 2'b11) begin
        if(krnl_partialKnn_wrapper_20_0__ap_done) begin
          krnl_partialKnn_wrapper_20_0__state <= 2'b10;
        end 
      end 
      if(krnl_partialKnn_wrapper_20_0__state == 2'b10) begin
        if(krnl_partialKnn_wrapper_20_0__ap_done_global__q0) begin
          krnl_partialKnn_wrapper_20_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign krnl_partialKnn_wrapper_20_0__ap_start = (krnl_partialKnn_wrapper_20_0__state == 2'b01);
  assign krnl_partialKnn_wrapper_21_0___in_21__q0 = in_21;
  assign krnl_partialKnn_wrapper_21_0__ap_start_global__q0 = ap_start__q0;
  assign krnl_partialKnn_wrapper_21_0__is_done__q0 = (krnl_partialKnn_wrapper_21_0__state == 2'b10);
  assign krnl_partialKnn_wrapper_21_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      krnl_partialKnn_wrapper_21_0__state <= 2'b00;
    end else begin
      if(krnl_partialKnn_wrapper_21_0__state == 2'b00) begin
        if(krnl_partialKnn_wrapper_21_0__ap_start_global__q0) begin
          krnl_partialKnn_wrapper_21_0__state <= 2'b01;
        end 
      end 
      if(krnl_partialKnn_wrapper_21_0__state == 2'b01) begin
        if(krnl_partialKnn_wrapper_21_0__ap_ready) begin
          if(krnl_partialKnn_wrapper_21_0__ap_done) begin
            krnl_partialKnn_wrapper_21_0__state <= 2'b10;
          end else begin
            krnl_partialKnn_wrapper_21_0__state <= 2'b11;
          end
        end 
      end 
      if(krnl_partialKnn_wrapper_21_0__state == 2'b11) begin
        if(krnl_partialKnn_wrapper_21_0__ap_done) begin
          krnl_partialKnn_wrapper_21_0__state <= 2'b10;
        end 
      end 
      if(krnl_partialKnn_wrapper_21_0__state == 2'b10) begin
        if(krnl_partialKnn_wrapper_21_0__ap_done_global__q0) begin
          krnl_partialKnn_wrapper_21_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign krnl_partialKnn_wrapper_21_0__ap_start = (krnl_partialKnn_wrapper_21_0__state == 2'b01);
  assign krnl_partialKnn_wrapper_22_0___in_22__q0 = in_22;
  assign krnl_partialKnn_wrapper_22_0__ap_start_global__q0 = ap_start__q0;
  assign krnl_partialKnn_wrapper_22_0__is_done__q0 = (krnl_partialKnn_wrapper_22_0__state == 2'b10);
  assign krnl_partialKnn_wrapper_22_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      krnl_partialKnn_wrapper_22_0__state <= 2'b00;
    end else begin
      if(krnl_partialKnn_wrapper_22_0__state == 2'b00) begin
        if(krnl_partialKnn_wrapper_22_0__ap_start_global__q0) begin
          krnl_partialKnn_wrapper_22_0__state <= 2'b01;
        end 
      end 
      if(krnl_partialKnn_wrapper_22_0__state == 2'b01) begin
        if(krnl_partialKnn_wrapper_22_0__ap_ready) begin
          if(krnl_partialKnn_wrapper_22_0__ap_done) begin
            krnl_partialKnn_wrapper_22_0__state <= 2'b10;
          end else begin
            krnl_partialKnn_wrapper_22_0__state <= 2'b11;
          end
        end 
      end 
      if(krnl_partialKnn_wrapper_22_0__state == 2'b11) begin
        if(krnl_partialKnn_wrapper_22_0__ap_done) begin
          krnl_partialKnn_wrapper_22_0__state <= 2'b10;
        end 
      end 
      if(krnl_partialKnn_wrapper_22_0__state == 2'b10) begin
        if(krnl_partialKnn_wrapper_22_0__ap_done_global__q0) begin
          krnl_partialKnn_wrapper_22_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign krnl_partialKnn_wrapper_22_0__ap_start = (krnl_partialKnn_wrapper_22_0__state == 2'b01);
  assign krnl_partialKnn_wrapper_23_0___in_23__q0 = in_23;
  assign krnl_partialKnn_wrapper_23_0__ap_start_global__q0 = ap_start__q0;
  assign krnl_partialKnn_wrapper_23_0__is_done__q0 = (krnl_partialKnn_wrapper_23_0__state == 2'b10);
  assign krnl_partialKnn_wrapper_23_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      krnl_partialKnn_wrapper_23_0__state <= 2'b00;
    end else begin
      if(krnl_partialKnn_wrapper_23_0__state == 2'b00) begin
        if(krnl_partialKnn_wrapper_23_0__ap_start_global__q0) begin
          krnl_partialKnn_wrapper_23_0__state <= 2'b01;
        end 
      end 
      if(krnl_partialKnn_wrapper_23_0__state == 2'b01) begin
        if(krnl_partialKnn_wrapper_23_0__ap_ready) begin
          if(krnl_partialKnn_wrapper_23_0__ap_done) begin
            krnl_partialKnn_wrapper_23_0__state <= 2'b10;
          end else begin
            krnl_partialKnn_wrapper_23_0__state <= 2'b11;
          end
        end 
      end 
      if(krnl_partialKnn_wrapper_23_0__state == 2'b11) begin
        if(krnl_partialKnn_wrapper_23_0__ap_done) begin
          krnl_partialKnn_wrapper_23_0__state <= 2'b10;
        end 
      end 
      if(krnl_partialKnn_wrapper_23_0__state == 2'b10) begin
        if(krnl_partialKnn_wrapper_23_0__ap_done_global__q0) begin
          krnl_partialKnn_wrapper_23_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign krnl_partialKnn_wrapper_23_0__ap_start = (krnl_partialKnn_wrapper_23_0__state == 2'b01);
  assign krnl_partialKnn_wrapper_24_0___in_24__q0 = in_24;
  assign krnl_partialKnn_wrapper_24_0__ap_start_global__q0 = ap_start__q0;
  assign krnl_partialKnn_wrapper_24_0__is_done__q0 = (krnl_partialKnn_wrapper_24_0__state == 2'b10);
  assign krnl_partialKnn_wrapper_24_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      krnl_partialKnn_wrapper_24_0__state <= 2'b00;
    end else begin
      if(krnl_partialKnn_wrapper_24_0__state == 2'b00) begin
        if(krnl_partialKnn_wrapper_24_0__ap_start_global__q0) begin
          krnl_partialKnn_wrapper_24_0__state <= 2'b01;
        end 
      end 
      if(krnl_partialKnn_wrapper_24_0__state == 2'b01) begin
        if(krnl_partialKnn_wrapper_24_0__ap_ready) begin
          if(krnl_partialKnn_wrapper_24_0__ap_done) begin
            krnl_partialKnn_wrapper_24_0__state <= 2'b10;
          end else begin
            krnl_partialKnn_wrapper_24_0__state <= 2'b11;
          end
        end 
      end 
      if(krnl_partialKnn_wrapper_24_0__state == 2'b11) begin
        if(krnl_partialKnn_wrapper_24_0__ap_done) begin
          krnl_partialKnn_wrapper_24_0__state <= 2'b10;
        end 
      end 
      if(krnl_partialKnn_wrapper_24_0__state == 2'b10) begin
        if(krnl_partialKnn_wrapper_24_0__ap_done_global__q0) begin
          krnl_partialKnn_wrapper_24_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign krnl_partialKnn_wrapper_24_0__ap_start = (krnl_partialKnn_wrapper_24_0__state == 2'b01);
  assign krnl_partialKnn_wrapper_25_0___in_25__q0 = in_25;
  assign krnl_partialKnn_wrapper_25_0__ap_start_global__q0 = ap_start__q0;
  assign krnl_partialKnn_wrapper_25_0__is_done__q0 = (krnl_partialKnn_wrapper_25_0__state == 2'b10);
  assign krnl_partialKnn_wrapper_25_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      krnl_partialKnn_wrapper_25_0__state <= 2'b00;
    end else begin
      if(krnl_partialKnn_wrapper_25_0__state == 2'b00) begin
        if(krnl_partialKnn_wrapper_25_0__ap_start_global__q0) begin
          krnl_partialKnn_wrapper_25_0__state <= 2'b01;
        end 
      end 
      if(krnl_partialKnn_wrapper_25_0__state == 2'b01) begin
        if(krnl_partialKnn_wrapper_25_0__ap_ready) begin
          if(krnl_partialKnn_wrapper_25_0__ap_done) begin
            krnl_partialKnn_wrapper_25_0__state <= 2'b10;
          end else begin
            krnl_partialKnn_wrapper_25_0__state <= 2'b11;
          end
        end 
      end 
      if(krnl_partialKnn_wrapper_25_0__state == 2'b11) begin
        if(krnl_partialKnn_wrapper_25_0__ap_done) begin
          krnl_partialKnn_wrapper_25_0__state <= 2'b10;
        end 
      end 
      if(krnl_partialKnn_wrapper_25_0__state == 2'b10) begin
        if(krnl_partialKnn_wrapper_25_0__ap_done_global__q0) begin
          krnl_partialKnn_wrapper_25_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign krnl_partialKnn_wrapper_25_0__ap_start = (krnl_partialKnn_wrapper_25_0__state == 2'b01);
  assign krnl_partialKnn_wrapper_26_0___in_26__q0 = in_26;
  assign krnl_partialKnn_wrapper_26_0__ap_start_global__q0 = ap_start__q0;
  assign krnl_partialKnn_wrapper_26_0__is_done__q0 = (krnl_partialKnn_wrapper_26_0__state == 2'b10);
  assign krnl_partialKnn_wrapper_26_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      krnl_partialKnn_wrapper_26_0__state <= 2'b00;
    end else begin
      if(krnl_partialKnn_wrapper_26_0__state == 2'b00) begin
        if(krnl_partialKnn_wrapper_26_0__ap_start_global__q0) begin
          krnl_partialKnn_wrapper_26_0__state <= 2'b01;
        end 
      end 
      if(krnl_partialKnn_wrapper_26_0__state == 2'b01) begin
        if(krnl_partialKnn_wrapper_26_0__ap_ready) begin
          if(krnl_partialKnn_wrapper_26_0__ap_done) begin
            krnl_partialKnn_wrapper_26_0__state <= 2'b10;
          end else begin
            krnl_partialKnn_wrapper_26_0__state <= 2'b11;
          end
        end 
      end 
      if(krnl_partialKnn_wrapper_26_0__state == 2'b11) begin
        if(krnl_partialKnn_wrapper_26_0__ap_done) begin
          krnl_partialKnn_wrapper_26_0__state <= 2'b10;
        end 
      end 
      if(krnl_partialKnn_wrapper_26_0__state == 2'b10) begin
        if(krnl_partialKnn_wrapper_26_0__ap_done_global__q0) begin
          krnl_partialKnn_wrapper_26_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign krnl_partialKnn_wrapper_26_0__ap_start = (krnl_partialKnn_wrapper_26_0__state == 2'b01);
  assign krnl_partialKnn_wrapper_3_0___in_3__q0 = in_3;
  assign krnl_partialKnn_wrapper_3_0__ap_start_global__q0 = ap_start__q0;
  assign krnl_partialKnn_wrapper_3_0__is_done__q0 = (krnl_partialKnn_wrapper_3_0__state == 2'b10);
  assign krnl_partialKnn_wrapper_3_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      krnl_partialKnn_wrapper_3_0__state <= 2'b00;
    end else begin
      if(krnl_partialKnn_wrapper_3_0__state == 2'b00) begin
        if(krnl_partialKnn_wrapper_3_0__ap_start_global__q0) begin
          krnl_partialKnn_wrapper_3_0__state <= 2'b01;
        end 
      end 
      if(krnl_partialKnn_wrapper_3_0__state == 2'b01) begin
        if(krnl_partialKnn_wrapper_3_0__ap_ready) begin
          if(krnl_partialKnn_wrapper_3_0__ap_done) begin
            krnl_partialKnn_wrapper_3_0__state <= 2'b10;
          end else begin
            krnl_partialKnn_wrapper_3_0__state <= 2'b11;
          end
        end 
      end 
      if(krnl_partialKnn_wrapper_3_0__state == 2'b11) begin
        if(krnl_partialKnn_wrapper_3_0__ap_done) begin
          krnl_partialKnn_wrapper_3_0__state <= 2'b10;
        end 
      end 
      if(krnl_partialKnn_wrapper_3_0__state == 2'b10) begin
        if(krnl_partialKnn_wrapper_3_0__ap_done_global__q0) begin
          krnl_partialKnn_wrapper_3_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign krnl_partialKnn_wrapper_3_0__ap_start = (krnl_partialKnn_wrapper_3_0__state == 2'b01);
  assign krnl_partialKnn_wrapper_4_0___in_4__q0 = in_4;
  assign krnl_partialKnn_wrapper_4_0__ap_start_global__q0 = ap_start__q0;
  assign krnl_partialKnn_wrapper_4_0__is_done__q0 = (krnl_partialKnn_wrapper_4_0__state == 2'b10);
  assign krnl_partialKnn_wrapper_4_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      krnl_partialKnn_wrapper_4_0__state <= 2'b00;
    end else begin
      if(krnl_partialKnn_wrapper_4_0__state == 2'b00) begin
        if(krnl_partialKnn_wrapper_4_0__ap_start_global__q0) begin
          krnl_partialKnn_wrapper_4_0__state <= 2'b01;
        end 
      end 
      if(krnl_partialKnn_wrapper_4_0__state == 2'b01) begin
        if(krnl_partialKnn_wrapper_4_0__ap_ready) begin
          if(krnl_partialKnn_wrapper_4_0__ap_done) begin
            krnl_partialKnn_wrapper_4_0__state <= 2'b10;
          end else begin
            krnl_partialKnn_wrapper_4_0__state <= 2'b11;
          end
        end 
      end 
      if(krnl_partialKnn_wrapper_4_0__state == 2'b11) begin
        if(krnl_partialKnn_wrapper_4_0__ap_done) begin
          krnl_partialKnn_wrapper_4_0__state <= 2'b10;
        end 
      end 
      if(krnl_partialKnn_wrapper_4_0__state == 2'b10) begin
        if(krnl_partialKnn_wrapper_4_0__ap_done_global__q0) begin
          krnl_partialKnn_wrapper_4_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign krnl_partialKnn_wrapper_4_0__ap_start = (krnl_partialKnn_wrapper_4_0__state == 2'b01);
  assign krnl_partialKnn_wrapper_5_0___in_5__q0 = in_5;
  assign krnl_partialKnn_wrapper_5_0__ap_start_global__q0 = ap_start__q0;
  assign krnl_partialKnn_wrapper_5_0__is_done__q0 = (krnl_partialKnn_wrapper_5_0__state == 2'b10);
  assign krnl_partialKnn_wrapper_5_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      krnl_partialKnn_wrapper_5_0__state <= 2'b00;
    end else begin
      if(krnl_partialKnn_wrapper_5_0__state == 2'b00) begin
        if(krnl_partialKnn_wrapper_5_0__ap_start_global__q0) begin
          krnl_partialKnn_wrapper_5_0__state <= 2'b01;
        end 
      end 
      if(krnl_partialKnn_wrapper_5_0__state == 2'b01) begin
        if(krnl_partialKnn_wrapper_5_0__ap_ready) begin
          if(krnl_partialKnn_wrapper_5_0__ap_done) begin
            krnl_partialKnn_wrapper_5_0__state <= 2'b10;
          end else begin
            krnl_partialKnn_wrapper_5_0__state <= 2'b11;
          end
        end 
      end 
      if(krnl_partialKnn_wrapper_5_0__state == 2'b11) begin
        if(krnl_partialKnn_wrapper_5_0__ap_done) begin
          krnl_partialKnn_wrapper_5_0__state <= 2'b10;
        end 
      end 
      if(krnl_partialKnn_wrapper_5_0__state == 2'b10) begin
        if(krnl_partialKnn_wrapper_5_0__ap_done_global__q0) begin
          krnl_partialKnn_wrapper_5_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign krnl_partialKnn_wrapper_5_0__ap_start = (krnl_partialKnn_wrapper_5_0__state == 2'b01);
  assign krnl_partialKnn_wrapper_6_0___in_6__q0 = in_6;
  assign krnl_partialKnn_wrapper_6_0__ap_start_global__q0 = ap_start__q0;
  assign krnl_partialKnn_wrapper_6_0__is_done__q0 = (krnl_partialKnn_wrapper_6_0__state == 2'b10);
  assign krnl_partialKnn_wrapper_6_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      krnl_partialKnn_wrapper_6_0__state <= 2'b00;
    end else begin
      if(krnl_partialKnn_wrapper_6_0__state == 2'b00) begin
        if(krnl_partialKnn_wrapper_6_0__ap_start_global__q0) begin
          krnl_partialKnn_wrapper_6_0__state <= 2'b01;
        end 
      end 
      if(krnl_partialKnn_wrapper_6_0__state == 2'b01) begin
        if(krnl_partialKnn_wrapper_6_0__ap_ready) begin
          if(krnl_partialKnn_wrapper_6_0__ap_done) begin
            krnl_partialKnn_wrapper_6_0__state <= 2'b10;
          end else begin
            krnl_partialKnn_wrapper_6_0__state <= 2'b11;
          end
        end 
      end 
      if(krnl_partialKnn_wrapper_6_0__state == 2'b11) begin
        if(krnl_partialKnn_wrapper_6_0__ap_done) begin
          krnl_partialKnn_wrapper_6_0__state <= 2'b10;
        end 
      end 
      if(krnl_partialKnn_wrapper_6_0__state == 2'b10) begin
        if(krnl_partialKnn_wrapper_6_0__ap_done_global__q0) begin
          krnl_partialKnn_wrapper_6_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign krnl_partialKnn_wrapper_6_0__ap_start = (krnl_partialKnn_wrapper_6_0__state == 2'b01);
  assign krnl_partialKnn_wrapper_7_0___in_7__q0 = in_7;
  assign krnl_partialKnn_wrapper_7_0__ap_start_global__q0 = ap_start__q0;
  assign krnl_partialKnn_wrapper_7_0__is_done__q0 = (krnl_partialKnn_wrapper_7_0__state == 2'b10);
  assign krnl_partialKnn_wrapper_7_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      krnl_partialKnn_wrapper_7_0__state <= 2'b00;
    end else begin
      if(krnl_partialKnn_wrapper_7_0__state == 2'b00) begin
        if(krnl_partialKnn_wrapper_7_0__ap_start_global__q0) begin
          krnl_partialKnn_wrapper_7_0__state <= 2'b01;
        end 
      end 
      if(krnl_partialKnn_wrapper_7_0__state == 2'b01) begin
        if(krnl_partialKnn_wrapper_7_0__ap_ready) begin
          if(krnl_partialKnn_wrapper_7_0__ap_done) begin
            krnl_partialKnn_wrapper_7_0__state <= 2'b10;
          end else begin
            krnl_partialKnn_wrapper_7_0__state <= 2'b11;
          end
        end 
      end 
      if(krnl_partialKnn_wrapper_7_0__state == 2'b11) begin
        if(krnl_partialKnn_wrapper_7_0__ap_done) begin
          krnl_partialKnn_wrapper_7_0__state <= 2'b10;
        end 
      end 
      if(krnl_partialKnn_wrapper_7_0__state == 2'b10) begin
        if(krnl_partialKnn_wrapper_7_0__ap_done_global__q0) begin
          krnl_partialKnn_wrapper_7_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign krnl_partialKnn_wrapper_7_0__ap_start = (krnl_partialKnn_wrapper_7_0__state == 2'b01);
  assign krnl_partialKnn_wrapper_8_0___in_8__q0 = in_8;
  assign krnl_partialKnn_wrapper_8_0__ap_start_global__q0 = ap_start__q0;
  assign krnl_partialKnn_wrapper_8_0__is_done__q0 = (krnl_partialKnn_wrapper_8_0__state == 2'b10);
  assign krnl_partialKnn_wrapper_8_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      krnl_partialKnn_wrapper_8_0__state <= 2'b00;
    end else begin
      if(krnl_partialKnn_wrapper_8_0__state == 2'b00) begin
        if(krnl_partialKnn_wrapper_8_0__ap_start_global__q0) begin
          krnl_partialKnn_wrapper_8_0__state <= 2'b01;
        end 
      end 
      if(krnl_partialKnn_wrapper_8_0__state == 2'b01) begin
        if(krnl_partialKnn_wrapper_8_0__ap_ready) begin
          if(krnl_partialKnn_wrapper_8_0__ap_done) begin
            krnl_partialKnn_wrapper_8_0__state <= 2'b10;
          end else begin
            krnl_partialKnn_wrapper_8_0__state <= 2'b11;
          end
        end 
      end 
      if(krnl_partialKnn_wrapper_8_0__state == 2'b11) begin
        if(krnl_partialKnn_wrapper_8_0__ap_done) begin
          krnl_partialKnn_wrapper_8_0__state <= 2'b10;
        end 
      end 
      if(krnl_partialKnn_wrapper_8_0__state == 2'b10) begin
        if(krnl_partialKnn_wrapper_8_0__ap_done_global__q0) begin
          krnl_partialKnn_wrapper_8_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign krnl_partialKnn_wrapper_8_0__ap_start = (krnl_partialKnn_wrapper_8_0__state == 2'b01);
  assign krnl_partialKnn_wrapper_9_0___in_9__q0 = in_9;
  assign krnl_partialKnn_wrapper_9_0__ap_start_global__q0 = ap_start__q0;
  assign krnl_partialKnn_wrapper_9_0__is_done__q0 = (krnl_partialKnn_wrapper_9_0__state == 2'b10);
  assign krnl_partialKnn_wrapper_9_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      krnl_partialKnn_wrapper_9_0__state <= 2'b00;
    end else begin
      if(krnl_partialKnn_wrapper_9_0__state == 2'b00) begin
        if(krnl_partialKnn_wrapper_9_0__ap_start_global__q0) begin
          krnl_partialKnn_wrapper_9_0__state <= 2'b01;
        end 
      end 
      if(krnl_partialKnn_wrapper_9_0__state == 2'b01) begin
        if(krnl_partialKnn_wrapper_9_0__ap_ready) begin
          if(krnl_partialKnn_wrapper_9_0__ap_done) begin
            krnl_partialKnn_wrapper_9_0__state <= 2'b10;
          end else begin
            krnl_partialKnn_wrapper_9_0__state <= 2'b11;
          end
        end 
      end 
      if(krnl_partialKnn_wrapper_9_0__state == 2'b11) begin
        if(krnl_partialKnn_wrapper_9_0__ap_done) begin
          krnl_partialKnn_wrapper_9_0__state <= 2'b10;
        end 
      end 
      if(krnl_partialKnn_wrapper_9_0__state == 2'b10) begin
        if(krnl_partialKnn_wrapper_9_0__ap_done_global__q0) begin
          krnl_partialKnn_wrapper_9_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign krnl_partialKnn_wrapper_9_0__ap_start = (krnl_partialKnn_wrapper_9_0__state == 2'b01);

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      tapa_state <= 2'b00;
    end else begin
      case(tapa_state)
        2'b00: begin
          if(ap_start__q0) begin
            tapa_state <= 2'b01;
          end 
        end
        2'b01: begin
          if(krnl_globalSort_L1_L2_0__is_done__q0 && krnl_globalSort_L1_L2_1__is_done__q0 && krnl_globalSort_L1_L2_2__is_done__q0 && krnl_globalSort_L1_L2_3__is_done__q0 && krnl_globalSort_L1_L2_4__is_done__q0 && krnl_globalSort_L1_L2_5__is_done__q0 && krnl_globalSort_L1_L2_6__is_done__q0 && krnl_globalSort_L1_L2_7__is_done__q0 && krnl_globalSort_L1_L2_8__is_done__q0 && krnl_globalSort_L1_L2_9__is_done__q0 && krnl_globalSort_L1_L2_10__is_done__q0 && krnl_globalSort_L1_L2_11__is_done__q0 && krnl_globalSort_L1_L2_12__is_done__q0 && krnl_output_dist_id_0__is_done__q0 && krnl_partialKnn_wrapper_0_0__is_done__q0 && krnl_partialKnn_wrapper_1_0__is_done__q0 && krnl_partialKnn_wrapper_10_0__is_done__q0 && krnl_partialKnn_wrapper_11_0__is_done__q0 && krnl_partialKnn_wrapper_12_0__is_done__q0 && krnl_partialKnn_wrapper_13_0__is_done__q0 && krnl_partialKnn_wrapper_14_0__is_done__q0 && krnl_partialKnn_wrapper_15_0__is_done__q0 && krnl_partialKnn_wrapper_16_0__is_done__q0 && krnl_partialKnn_wrapper_17_0__is_done__q0 && krnl_partialKnn_wrapper_18_0__is_done__q0 && krnl_partialKnn_wrapper_19_0__is_done__q0 && krnl_partialKnn_wrapper_2_0__is_done__q0 && krnl_partialKnn_wrapper_20_0__is_done__q0 && krnl_partialKnn_wrapper_21_0__is_done__q0 && krnl_partialKnn_wrapper_22_0__is_done__q0 && krnl_partialKnn_wrapper_23_0__is_done__q0 && krnl_partialKnn_wrapper_24_0__is_done__q0 && krnl_partialKnn_wrapper_25_0__is_done__q0 && krnl_partialKnn_wrapper_26_0__is_done__q0 && krnl_partialKnn_wrapper_3_0__is_done__q0 && krnl_partialKnn_wrapper_4_0__is_done__q0 && krnl_partialKnn_wrapper_5_0__is_done__q0 && krnl_partialKnn_wrapper_6_0__is_done__q0 && krnl_partialKnn_wrapper_7_0__is_done__q0 && krnl_partialKnn_wrapper_8_0__is_done__q0 && krnl_partialKnn_wrapper_9_0__is_done__q0) begin
            tapa_state <= 2'b10;
          end 
        end
        2'b10: begin
          tapa_state <= 2'b00;
          countdown <= 1'd0;
        end
        2'b11: begin
          if(countdown == 1'd0) begin
            tapa_state <= 2'b00;
          end else begin
            countdown <= (countdown - 1'd1);
          end
        end
      endcase
    end
  end

  assign ap_idle = (tapa_state == 2'b00);
  assign ap_done = ap_done__q0;
  assign ap_ready = ap_done__q0;
  assign ap_start__q0 = ap_start;
  assign ap_done__q0 = (tapa_state == 2'b10);

endmodule

