`timescale 1 ns / 1 ps 

(* CORE_GENERATION_INFO = "jacobi3d_kernel_jacobi3d_kernel,hls_ip_2023_2_2,{HLS_INPUT_TYPE=cxx,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=0,HLS_INPUT_PART=xcvp1802-lsvc4072-2MP-e-S,HLS_INPUT_CLOCK=3.330000,HLS_INPUT_ARCH=others,HLS_SYN_CLOCK=1.000000,HLS_SYN_LAT=0,HLS_SYN_TPT=none,HLS_SYN_MEM=0,HLS_SYN_DSP=0,HLS_SYN_FF=246,HLS_SYN_LUT=424,HLS_VERSION=2023_2_2}" *)


module jacobi3d_kernel
(
  s_axi_control_AWVALID,
  s_axi_control_AWREADY,
  s_axi_control_AWADDR,
  s_axi_control_WVALID,
  s_axi_control_WREADY,
  s_axi_control_WDATA,
  s_axi_control_WSTRB,
  s_axi_control_ARVALID,
  s_axi_control_ARREADY,
  s_axi_control_ARADDR,
  s_axi_control_RVALID,
  s_axi_control_RREADY,
  s_axi_control_RDATA,
  s_axi_control_RRESP,
  s_axi_control_BVALID,
  s_axi_control_BREADY,
  s_axi_control_BRESP,
  ap_clk,
  ap_rst_n,
  interrupt,
  m_axi_bank_0_t1_ARADDR,
  m_axi_bank_0_t1_ARBURST,
  m_axi_bank_0_t1_ARCACHE,
  m_axi_bank_0_t1_ARID,
  m_axi_bank_0_t1_ARLEN,
  m_axi_bank_0_t1_ARLOCK,
  m_axi_bank_0_t1_ARPROT,
  m_axi_bank_0_t1_ARQOS,
  m_axi_bank_0_t1_ARREADY,
  m_axi_bank_0_t1_ARSIZE,
  m_axi_bank_0_t1_ARVALID,
  m_axi_bank_0_t1_AWADDR,
  m_axi_bank_0_t1_AWBURST,
  m_axi_bank_0_t1_AWCACHE,
  m_axi_bank_0_t1_AWID,
  m_axi_bank_0_t1_AWLEN,
  m_axi_bank_0_t1_AWLOCK,
  m_axi_bank_0_t1_AWPROT,
  m_axi_bank_0_t1_AWQOS,
  m_axi_bank_0_t1_AWREADY,
  m_axi_bank_0_t1_AWSIZE,
  m_axi_bank_0_t1_AWVALID,
  m_axi_bank_0_t1_BID,
  m_axi_bank_0_t1_BREADY,
  m_axi_bank_0_t1_BRESP,
  m_axi_bank_0_t1_BVALID,
  m_axi_bank_0_t1_RDATA,
  m_axi_bank_0_t1_RID,
  m_axi_bank_0_t1_RLAST,
  m_axi_bank_0_t1_RREADY,
  m_axi_bank_0_t1_RRESP,
  m_axi_bank_0_t1_RVALID,
  m_axi_bank_0_t1_WDATA,
  m_axi_bank_0_t1_WLAST,
  m_axi_bank_0_t1_WREADY,
  m_axi_bank_0_t1_WSTRB,
  m_axi_bank_0_t1_WVALID,
  m_axi_bank_1_t0_ARADDR,
  m_axi_bank_1_t0_ARBURST,
  m_axi_bank_1_t0_ARCACHE,
  m_axi_bank_1_t0_ARID,
  m_axi_bank_1_t0_ARLEN,
  m_axi_bank_1_t0_ARLOCK,
  m_axi_bank_1_t0_ARPROT,
  m_axi_bank_1_t0_ARQOS,
  m_axi_bank_1_t0_ARREADY,
  m_axi_bank_1_t0_ARSIZE,
  m_axi_bank_1_t0_ARVALID,
  m_axi_bank_1_t0_AWADDR,
  m_axi_bank_1_t0_AWBURST,
  m_axi_bank_1_t0_AWCACHE,
  m_axi_bank_1_t0_AWID,
  m_axi_bank_1_t0_AWLEN,
  m_axi_bank_1_t0_AWLOCK,
  m_axi_bank_1_t0_AWPROT,
  m_axi_bank_1_t0_AWQOS,
  m_axi_bank_1_t0_AWREADY,
  m_axi_bank_1_t0_AWSIZE,
  m_axi_bank_1_t0_AWVALID,
  m_axi_bank_1_t0_BID,
  m_axi_bank_1_t0_BREADY,
  m_axi_bank_1_t0_BRESP,
  m_axi_bank_1_t0_BVALID,
  m_axi_bank_1_t0_RDATA,
  m_axi_bank_1_t0_RID,
  m_axi_bank_1_t0_RLAST,
  m_axi_bank_1_t0_RREADY,
  m_axi_bank_1_t0_RRESP,
  m_axi_bank_1_t0_RVALID,
  m_axi_bank_1_t0_WDATA,
  m_axi_bank_1_t0_WLAST,
  m_axi_bank_1_t0_WREADY,
  m_axi_bank_1_t0_WSTRB,
  m_axi_bank_1_t0_WVALID
);

  parameter C_S_AXI_CONTROL_DATA_WIDTH = 32;
  parameter C_S_AXI_CONTROL_ADDR_WIDTH = 6;
  parameter C_S_AXI_DATA_WIDTH = 32;
  parameter C_S_AXI_CONTROL_WSTRB_WIDTH = 32 / 8;
  parameter C_S_AXI_WSTRB_WIDTH = 32 / 8;
  (* RS_HS = "s_axi_control_AW.valid" *)input s_axi_control_AWVALID;
  (* RS_HS = "s_axi_control_AW.ready" *)output s_axi_control_AWREADY;
  (* RS_HS = "s_axi_control_AW.data" *)input [C_S_AXI_CONTROL_ADDR_WIDTH-1:0] s_axi_control_AWADDR;
  (* RS_HS = "s_axi_control_W.valid" *)input s_axi_control_WVALID;
  (* RS_HS = "s_axi_control_W.ready" *)output s_axi_control_WREADY;
  (* RS_HS = "s_axi_control_W.data" *)input [C_S_AXI_CONTROL_DATA_WIDTH-1:0] s_axi_control_WDATA;
  (* RS_HS = "s_axi_control_W.data" *)input [C_S_AXI_CONTROL_WSTRB_WIDTH-1:0] s_axi_control_WSTRB;
  (* RS_HS = "s_axi_control_AR.valid" *)input s_axi_control_ARVALID;
  (* RS_HS = "s_axi_control_AR.ready" *)output s_axi_control_ARREADY;
  (* RS_HS = "s_axi_control_AR.data" *)input [C_S_AXI_CONTROL_ADDR_WIDTH-1:0] s_axi_control_ARADDR;
  (* RS_HS = "s_axi_control_R.valid" *)output s_axi_control_RVALID;
  (* RS_HS = "s_axi_control_R.ready" *)input s_axi_control_RREADY;
  (* RS_HS = "s_axi_control_R.data" *)output [C_S_AXI_CONTROL_DATA_WIDTH-1:0] s_axi_control_RDATA;
  (* RS_HS = "s_axi_control_R.data" *)output [1:0] s_axi_control_RRESP;
  (* RS_HS = "s_axi_control_B.valid" *)output s_axi_control_BVALID;
  (* RS_HS = "s_axi_control_B.ready" *)input s_axi_control_BREADY;
  (* RS_HS = "s_axi_control_B.data" *)output [1:0] s_axi_control_BRESP;
  (* RS_CLK *)input ap_clk;
  (* RS_RST = "ff" *)input ap_rst_n;
  (* RS_FF = "interrupt" *)output interrupt;
  (* RS_HS = "m_axi_bank_0_t1_AR.data" *)output [63:0] m_axi_bank_0_t1_ARADDR;
  (* RS_HS = "m_axi_bank_0_t1_AR.data" *)output [1:0] m_axi_bank_0_t1_ARBURST;
  (* RS_HS = "m_axi_bank_0_t1_AR.data" *)output [3:0] m_axi_bank_0_t1_ARCACHE;
  (* RS_HS = "m_axi_bank_0_t1_AR.data" *)output [0:0] m_axi_bank_0_t1_ARID;
  (* RS_HS = "m_axi_bank_0_t1_AR.data" *)output [7:0] m_axi_bank_0_t1_ARLEN;
  (* RS_HS = "m_axi_bank_0_t1_AR.data" *)output m_axi_bank_0_t1_ARLOCK;
  (* RS_HS = "m_axi_bank_0_t1_AR.data" *)output [2:0] m_axi_bank_0_t1_ARPROT;
  (* RS_HS = "m_axi_bank_0_t1_AR.data" *)output [3:0] m_axi_bank_0_t1_ARQOS;
  (* RS_HS = "m_axi_bank_0_t1_AR.ready" *)input m_axi_bank_0_t1_ARREADY;
  (* RS_HS = "m_axi_bank_0_t1_AR.data" *)output [2:0] m_axi_bank_0_t1_ARSIZE;
  (* RS_HS = "m_axi_bank_0_t1_AR.valid" *)output m_axi_bank_0_t1_ARVALID;
  (* RS_HS = "m_axi_bank_0_t1_AW.data" *)output [63:0] m_axi_bank_0_t1_AWADDR;
  (* RS_HS = "m_axi_bank_0_t1_AW.data" *)output [1:0] m_axi_bank_0_t1_AWBURST;
  (* RS_HS = "m_axi_bank_0_t1_AW.data" *)output [3:0] m_axi_bank_0_t1_AWCACHE;
  (* RS_HS = "m_axi_bank_0_t1_AW.data" *)output [0:0] m_axi_bank_0_t1_AWID;
  (* RS_HS = "m_axi_bank_0_t1_AW.data" *)output [7:0] m_axi_bank_0_t1_AWLEN;
  (* RS_HS = "m_axi_bank_0_t1_AW.data" *)output m_axi_bank_0_t1_AWLOCK;
  (* RS_HS = "m_axi_bank_0_t1_AW.data" *)output [2:0] m_axi_bank_0_t1_AWPROT;
  (* RS_HS = "m_axi_bank_0_t1_AW.data" *)output [3:0] m_axi_bank_0_t1_AWQOS;
  (* RS_HS = "m_axi_bank_0_t1_AW.ready" *)input m_axi_bank_0_t1_AWREADY;
  (* RS_HS = "m_axi_bank_0_t1_AW.data" *)output [2:0] m_axi_bank_0_t1_AWSIZE;
  (* RS_HS = "m_axi_bank_0_t1_AW.valid" *)output m_axi_bank_0_t1_AWVALID;
  (* RS_HS = "m_axi_bank_0_t1_B.data" *)input [0:0] m_axi_bank_0_t1_BID;
  (* RS_HS = "m_axi_bank_0_t1_B.ready" *)output m_axi_bank_0_t1_BREADY;
  (* RS_HS = "m_axi_bank_0_t1_B.data" *)input [1:0] m_axi_bank_0_t1_BRESP;
  (* RS_HS = "m_axi_bank_0_t1_B.valid" *)input m_axi_bank_0_t1_BVALID;
  (* RS_HS = "m_axi_bank_0_t1_R.data" *)input [511:0] m_axi_bank_0_t1_RDATA;
  (* RS_HS = "m_axi_bank_0_t1_R.data" *)input [0:0] m_axi_bank_0_t1_RID;
  (* RS_HS = "m_axi_bank_0_t1_R.data" *)input m_axi_bank_0_t1_RLAST;
  (* RS_HS = "m_axi_bank_0_t1_R.ready" *)output m_axi_bank_0_t1_RREADY;
  (* RS_HS = "m_axi_bank_0_t1_R.data" *)input [1:0] m_axi_bank_0_t1_RRESP;
  (* RS_HS = "m_axi_bank_0_t1_R.valid" *)input m_axi_bank_0_t1_RVALID;
  (* RS_HS = "m_axi_bank_0_t1_W.data" *)output [511:0] m_axi_bank_0_t1_WDATA;
  (* RS_HS = "m_axi_bank_0_t1_W.data" *)output m_axi_bank_0_t1_WLAST;
  (* RS_HS = "m_axi_bank_0_t1_W.ready" *)input m_axi_bank_0_t1_WREADY;
  (* RS_HS = "m_axi_bank_0_t1_W.data" *)output [63:0] m_axi_bank_0_t1_WSTRB;
  (* RS_HS = "m_axi_bank_0_t1_W.valid" *)output m_axi_bank_0_t1_WVALID;
  (* RS_HS = "m_axi_bank_1_t0_AR.data" *)output [63:0] m_axi_bank_1_t0_ARADDR;
  (* RS_HS = "m_axi_bank_1_t0_AR.data" *)output [1:0] m_axi_bank_1_t0_ARBURST;
  (* RS_HS = "m_axi_bank_1_t0_AR.data" *)output [3:0] m_axi_bank_1_t0_ARCACHE;
  (* RS_HS = "m_axi_bank_1_t0_AR.data" *)output [0:0] m_axi_bank_1_t0_ARID;
  (* RS_HS = "m_axi_bank_1_t0_AR.data" *)output [7:0] m_axi_bank_1_t0_ARLEN;
  (* RS_HS = "m_axi_bank_1_t0_AR.data" *)output m_axi_bank_1_t0_ARLOCK;
  (* RS_HS = "m_axi_bank_1_t0_AR.data" *)output [2:0] m_axi_bank_1_t0_ARPROT;
  (* RS_HS = "m_axi_bank_1_t0_AR.data" *)output [3:0] m_axi_bank_1_t0_ARQOS;
  (* RS_HS = "m_axi_bank_1_t0_AR.ready" *)input m_axi_bank_1_t0_ARREADY;
  (* RS_HS = "m_axi_bank_1_t0_AR.data" *)output [2:0] m_axi_bank_1_t0_ARSIZE;
  (* RS_HS = "m_axi_bank_1_t0_AR.valid" *)output m_axi_bank_1_t0_ARVALID;
  (* RS_HS = "m_axi_bank_1_t0_AW.data" *)output [63:0] m_axi_bank_1_t0_AWADDR;
  (* RS_HS = "m_axi_bank_1_t0_AW.data" *)output [1:0] m_axi_bank_1_t0_AWBURST;
  (* RS_HS = "m_axi_bank_1_t0_AW.data" *)output [3:0] m_axi_bank_1_t0_AWCACHE;
  (* RS_HS = "m_axi_bank_1_t0_AW.data" *)output [0:0] m_axi_bank_1_t0_AWID;
  (* RS_HS = "m_axi_bank_1_t0_AW.data" *)output [7:0] m_axi_bank_1_t0_AWLEN;
  (* RS_HS = "m_axi_bank_1_t0_AW.data" *)output m_axi_bank_1_t0_AWLOCK;
  (* RS_HS = "m_axi_bank_1_t0_AW.data" *)output [2:0] m_axi_bank_1_t0_AWPROT;
  (* RS_HS = "m_axi_bank_1_t0_AW.data" *)output [3:0] m_axi_bank_1_t0_AWQOS;
  (* RS_HS = "m_axi_bank_1_t0_AW.ready" *)input m_axi_bank_1_t0_AWREADY;
  (* RS_HS = "m_axi_bank_1_t0_AW.data" *)output [2:0] m_axi_bank_1_t0_AWSIZE;
  (* RS_HS = "m_axi_bank_1_t0_AW.valid" *)output m_axi_bank_1_t0_AWVALID;
  (* RS_HS = "m_axi_bank_1_t0_B.data" *)input [0:0] m_axi_bank_1_t0_BID;
  (* RS_HS = "m_axi_bank_1_t0_B.ready" *)output m_axi_bank_1_t0_BREADY;
  (* RS_HS = "m_axi_bank_1_t0_B.data" *)input [1:0] m_axi_bank_1_t0_BRESP;
  (* RS_HS = "m_axi_bank_1_t0_B.valid" *)input m_axi_bank_1_t0_BVALID;
  (* RS_HS = "m_axi_bank_1_t0_R.data" *)input [511:0] m_axi_bank_1_t0_RDATA;
  (* RS_HS = "m_axi_bank_1_t0_R.data" *)input [0:0] m_axi_bank_1_t0_RID;
  (* RS_HS = "m_axi_bank_1_t0_R.data" *)input m_axi_bank_1_t0_RLAST;
  (* RS_HS = "m_axi_bank_1_t0_R.ready" *)output m_axi_bank_1_t0_RREADY;
  (* RS_HS = "m_axi_bank_1_t0_R.data" *)input [1:0] m_axi_bank_1_t0_RRESP;
  (* RS_HS = "m_axi_bank_1_t0_R.valid" *)input m_axi_bank_1_t0_RVALID;
  (* RS_HS = "m_axi_bank_1_t0_W.data" *)output [511:0] m_axi_bank_1_t0_WDATA;
  (* RS_HS = "m_axi_bank_1_t0_W.data" *)output m_axi_bank_1_t0_WLAST;
  (* RS_HS = "m_axi_bank_1_t0_W.ready" *)input m_axi_bank_1_t0_WREADY;
  (* RS_HS = "m_axi_bank_1_t0_W.data" *)output [63:0] m_axi_bank_1_t0_WSTRB;
  (* RS_HS = "m_axi_bank_1_t0_W.valid" *)output m_axi_bank_1_t0_WVALID;
  wire ap_start;
  wire [63:0] bank_1_t0;
  wire [63:0] bank_0_t1;
  wire [63:0] coalesced_data_num;
  wire [512:0] bank_0_t1_buf__dout;
  wire bank_0_t1_buf__empty_n;
  wire bank_0_t1_buf__read;
  wire [512:0] bank_0_t1_buf__din;
  wire bank_0_t1_buf__full_n;
  wire bank_0_t1_buf__write;
  wire [512:0] bank_1_t0_buf__dout;
  wire bank_1_t0_buf__empty_n;
  wire bank_1_t0_buf__read;
  wire [512:0] bank_1_t0_buf__din;
  wire bank_1_t0_buf__full_n;
  wire bank_1_t0_buf__write;
  wire [512:0] from_t0_to_t0_bank_1__dout;
  wire from_t0_to_t0_bank_1__empty_n;
  wire from_t0_to_t0_bank_1__read;
  wire [512:0] from_t0_to_t0_bank_1__din;
  wire from_t0_to_t0_bank_1__full_n;
  wire from_t0_to_t0_bank_1__write;
  wire [512:0] from_t1_bank_0_to_t1_iter1__dout;
  wire from_t1_bank_0_to_t1_iter1__empty_n;
  wire from_t1_bank_0_to_t1_iter1__read;
  wire [512:0] from_t1_bank_0_to_t1_iter1__din;
  wire from_t1_bank_0_to_t1_iter1__full_n;
  wire from_t1_bank_0_to_t1_iter1__write;
  wire [512:0] from_t1_iter100_to_t1_iter101__dout;
  wire from_t1_iter100_to_t1_iter101__empty_n;
  wire from_t1_iter100_to_t1_iter101__read;
  wire [512:0] from_t1_iter100_to_t1_iter101__din;
  wire from_t1_iter100_to_t1_iter101__full_n;
  wire from_t1_iter100_to_t1_iter101__write;
  wire [512:0] from_t1_iter101_to_t1_iter102__dout;
  wire from_t1_iter101_to_t1_iter102__empty_n;
  wire from_t1_iter101_to_t1_iter102__read;
  wire [512:0] from_t1_iter101_to_t1_iter102__din;
  wire from_t1_iter101_to_t1_iter102__full_n;
  wire from_t1_iter101_to_t1_iter102__write;
  wire [512:0] from_t1_iter102_to_t1_iter103__dout;
  wire from_t1_iter102_to_t1_iter103__empty_n;
  wire from_t1_iter102_to_t1_iter103__read;
  wire [512:0] from_t1_iter102_to_t1_iter103__din;
  wire from_t1_iter102_to_t1_iter103__full_n;
  wire from_t1_iter102_to_t1_iter103__write;
  wire [512:0] from_t1_iter103_to_t1_iter104__dout;
  wire from_t1_iter103_to_t1_iter104__empty_n;
  wire from_t1_iter103_to_t1_iter104__read;
  wire [512:0] from_t1_iter103_to_t1_iter104__din;
  wire from_t1_iter103_to_t1_iter104__full_n;
  wire from_t1_iter103_to_t1_iter104__write;
  wire [512:0] from_t1_iter104_to_t1_iter105__dout;
  wire from_t1_iter104_to_t1_iter105__empty_n;
  wire from_t1_iter104_to_t1_iter105__read;
  wire [512:0] from_t1_iter104_to_t1_iter105__din;
  wire from_t1_iter104_to_t1_iter105__full_n;
  wire from_t1_iter104_to_t1_iter105__write;
  wire [512:0] from_t1_iter105_to_t1_iter106__dout;
  wire from_t1_iter105_to_t1_iter106__empty_n;
  wire from_t1_iter105_to_t1_iter106__read;
  wire [512:0] from_t1_iter105_to_t1_iter106__din;
  wire from_t1_iter105_to_t1_iter106__full_n;
  wire from_t1_iter105_to_t1_iter106__write;
  wire [512:0] from_t1_iter106_to_t1_iter107__dout;
  wire from_t1_iter106_to_t1_iter107__empty_n;
  wire from_t1_iter106_to_t1_iter107__read;
  wire [512:0] from_t1_iter106_to_t1_iter107__din;
  wire from_t1_iter106_to_t1_iter107__full_n;
  wire from_t1_iter106_to_t1_iter107__write;
  wire [512:0] from_t1_iter107_to_t1_iter108__dout;
  wire from_t1_iter107_to_t1_iter108__empty_n;
  wire from_t1_iter107_to_t1_iter108__read;
  wire [512:0] from_t1_iter107_to_t1_iter108__din;
  wire from_t1_iter107_to_t1_iter108__full_n;
  wire from_t1_iter107_to_t1_iter108__write;
  wire [512:0] from_t1_iter108_to_t0__dout;
  wire from_t1_iter108_to_t0__empty_n;
  wire from_t1_iter108_to_t0__read;
  wire [512:0] from_t1_iter108_to_t0__din;
  wire from_t1_iter108_to_t0__full_n;
  wire from_t1_iter108_to_t0__write;
  wire [512:0] from_t1_iter10_to_t1_iter11__dout;
  wire from_t1_iter10_to_t1_iter11__empty_n;
  wire from_t1_iter10_to_t1_iter11__read;
  wire [512:0] from_t1_iter10_to_t1_iter11__din;
  wire from_t1_iter10_to_t1_iter11__full_n;
  wire from_t1_iter10_to_t1_iter11__write;
  wire [512:0] from_t1_iter11_to_t1_iter12__dout;
  wire from_t1_iter11_to_t1_iter12__empty_n;
  wire from_t1_iter11_to_t1_iter12__read;
  wire [512:0] from_t1_iter11_to_t1_iter12__din;
  wire from_t1_iter11_to_t1_iter12__full_n;
  wire from_t1_iter11_to_t1_iter12__write;
  wire [512:0] from_t1_iter12_to_t1_iter13__dout;
  wire from_t1_iter12_to_t1_iter13__empty_n;
  wire from_t1_iter12_to_t1_iter13__read;
  wire [512:0] from_t1_iter12_to_t1_iter13__din;
  wire from_t1_iter12_to_t1_iter13__full_n;
  wire from_t1_iter12_to_t1_iter13__write;
  wire [512:0] from_t1_iter13_to_t1_iter14__dout;
  wire from_t1_iter13_to_t1_iter14__empty_n;
  wire from_t1_iter13_to_t1_iter14__read;
  wire [512:0] from_t1_iter13_to_t1_iter14__din;
  wire from_t1_iter13_to_t1_iter14__full_n;
  wire from_t1_iter13_to_t1_iter14__write;
  wire [512:0] from_t1_iter14_to_t1_iter15__dout;
  wire from_t1_iter14_to_t1_iter15__empty_n;
  wire from_t1_iter14_to_t1_iter15__read;
  wire [512:0] from_t1_iter14_to_t1_iter15__din;
  wire from_t1_iter14_to_t1_iter15__full_n;
  wire from_t1_iter14_to_t1_iter15__write;
  wire [512:0] from_t1_iter15_to_t1_iter16__dout;
  wire from_t1_iter15_to_t1_iter16__empty_n;
  wire from_t1_iter15_to_t1_iter16__read;
  wire [512:0] from_t1_iter15_to_t1_iter16__din;
  wire from_t1_iter15_to_t1_iter16__full_n;
  wire from_t1_iter15_to_t1_iter16__write;
  wire [512:0] from_t1_iter16_to_t1_iter17__dout;
  wire from_t1_iter16_to_t1_iter17__empty_n;
  wire from_t1_iter16_to_t1_iter17__read;
  wire [512:0] from_t1_iter16_to_t1_iter17__din;
  wire from_t1_iter16_to_t1_iter17__full_n;
  wire from_t1_iter16_to_t1_iter17__write;
  wire [512:0] from_t1_iter17_to_t1_iter18__dout;
  wire from_t1_iter17_to_t1_iter18__empty_n;
  wire from_t1_iter17_to_t1_iter18__read;
  wire [512:0] from_t1_iter17_to_t1_iter18__din;
  wire from_t1_iter17_to_t1_iter18__full_n;
  wire from_t1_iter17_to_t1_iter18__write;
  wire [512:0] from_t1_iter18_to_t1_iter19__dout;
  wire from_t1_iter18_to_t1_iter19__empty_n;
  wire from_t1_iter18_to_t1_iter19__read;
  wire [512:0] from_t1_iter18_to_t1_iter19__din;
  wire from_t1_iter18_to_t1_iter19__full_n;
  wire from_t1_iter18_to_t1_iter19__write;
  wire [512:0] from_t1_iter19_to_t1_iter20__dout;
  wire from_t1_iter19_to_t1_iter20__empty_n;
  wire from_t1_iter19_to_t1_iter20__read;
  wire [512:0] from_t1_iter19_to_t1_iter20__din;
  wire from_t1_iter19_to_t1_iter20__full_n;
  wire from_t1_iter19_to_t1_iter20__write;
  wire [512:0] from_t1_iter1_to_t1_iter2__dout;
  wire from_t1_iter1_to_t1_iter2__empty_n;
  wire from_t1_iter1_to_t1_iter2__read;
  wire [512:0] from_t1_iter1_to_t1_iter2__din;
  wire from_t1_iter1_to_t1_iter2__full_n;
  wire from_t1_iter1_to_t1_iter2__write;
  wire [512:0] from_t1_iter20_to_t1_iter21__dout;
  wire from_t1_iter20_to_t1_iter21__empty_n;
  wire from_t1_iter20_to_t1_iter21__read;
  wire [512:0] from_t1_iter20_to_t1_iter21__din;
  wire from_t1_iter20_to_t1_iter21__full_n;
  wire from_t1_iter20_to_t1_iter21__write;
  wire [512:0] from_t1_iter21_to_t1_iter22__dout;
  wire from_t1_iter21_to_t1_iter22__empty_n;
  wire from_t1_iter21_to_t1_iter22__read;
  wire [512:0] from_t1_iter21_to_t1_iter22__din;
  wire from_t1_iter21_to_t1_iter22__full_n;
  wire from_t1_iter21_to_t1_iter22__write;
  wire [512:0] from_t1_iter22_to_t1_iter23__dout;
  wire from_t1_iter22_to_t1_iter23__empty_n;
  wire from_t1_iter22_to_t1_iter23__read;
  wire [512:0] from_t1_iter22_to_t1_iter23__din;
  wire from_t1_iter22_to_t1_iter23__full_n;
  wire from_t1_iter22_to_t1_iter23__write;
  wire [512:0] from_t1_iter23_to_t1_iter24__dout;
  wire from_t1_iter23_to_t1_iter24__empty_n;
  wire from_t1_iter23_to_t1_iter24__read;
  wire [512:0] from_t1_iter23_to_t1_iter24__din;
  wire from_t1_iter23_to_t1_iter24__full_n;
  wire from_t1_iter23_to_t1_iter24__write;
  wire [512:0] from_t1_iter24_to_t1_iter25__dout;
  wire from_t1_iter24_to_t1_iter25__empty_n;
  wire from_t1_iter24_to_t1_iter25__read;
  wire [512:0] from_t1_iter24_to_t1_iter25__din;
  wire from_t1_iter24_to_t1_iter25__full_n;
  wire from_t1_iter24_to_t1_iter25__write;
  wire [512:0] from_t1_iter25_to_t1_iter26__dout;
  wire from_t1_iter25_to_t1_iter26__empty_n;
  wire from_t1_iter25_to_t1_iter26__read;
  wire [512:0] from_t1_iter25_to_t1_iter26__din;
  wire from_t1_iter25_to_t1_iter26__full_n;
  wire from_t1_iter25_to_t1_iter26__write;
  wire [512:0] from_t1_iter26_to_t1_iter27__dout;
  wire from_t1_iter26_to_t1_iter27__empty_n;
  wire from_t1_iter26_to_t1_iter27__read;
  wire [512:0] from_t1_iter26_to_t1_iter27__din;
  wire from_t1_iter26_to_t1_iter27__full_n;
  wire from_t1_iter26_to_t1_iter27__write;
  wire [512:0] from_t1_iter27_to_t1_iter28__dout;
  wire from_t1_iter27_to_t1_iter28__empty_n;
  wire from_t1_iter27_to_t1_iter28__read;
  wire [512:0] from_t1_iter27_to_t1_iter28__din;
  wire from_t1_iter27_to_t1_iter28__full_n;
  wire from_t1_iter27_to_t1_iter28__write;
  wire [512:0] from_t1_iter28_to_t1_iter29__dout;
  wire from_t1_iter28_to_t1_iter29__empty_n;
  wire from_t1_iter28_to_t1_iter29__read;
  wire [512:0] from_t1_iter28_to_t1_iter29__din;
  wire from_t1_iter28_to_t1_iter29__full_n;
  wire from_t1_iter28_to_t1_iter29__write;
  wire [512:0] from_t1_iter29_to_t1_iter30__dout;
  wire from_t1_iter29_to_t1_iter30__empty_n;
  wire from_t1_iter29_to_t1_iter30__read;
  wire [512:0] from_t1_iter29_to_t1_iter30__din;
  wire from_t1_iter29_to_t1_iter30__full_n;
  wire from_t1_iter29_to_t1_iter30__write;
  wire [512:0] from_t1_iter2_to_t1_iter3__dout;
  wire from_t1_iter2_to_t1_iter3__empty_n;
  wire from_t1_iter2_to_t1_iter3__read;
  wire [512:0] from_t1_iter2_to_t1_iter3__din;
  wire from_t1_iter2_to_t1_iter3__full_n;
  wire from_t1_iter2_to_t1_iter3__write;
  wire [512:0] from_t1_iter30_to_t1_iter31__dout;
  wire from_t1_iter30_to_t1_iter31__empty_n;
  wire from_t1_iter30_to_t1_iter31__read;
  wire [512:0] from_t1_iter30_to_t1_iter31__din;
  wire from_t1_iter30_to_t1_iter31__full_n;
  wire from_t1_iter30_to_t1_iter31__write;
  wire [512:0] from_t1_iter31_to_t1_iter32__dout;
  wire from_t1_iter31_to_t1_iter32__empty_n;
  wire from_t1_iter31_to_t1_iter32__read;
  wire [512:0] from_t1_iter31_to_t1_iter32__din;
  wire from_t1_iter31_to_t1_iter32__full_n;
  wire from_t1_iter31_to_t1_iter32__write;
  wire [512:0] from_t1_iter32_to_t1_iter33__dout;
  wire from_t1_iter32_to_t1_iter33__empty_n;
  wire from_t1_iter32_to_t1_iter33__read;
  wire [512:0] from_t1_iter32_to_t1_iter33__din;
  wire from_t1_iter32_to_t1_iter33__full_n;
  wire from_t1_iter32_to_t1_iter33__write;
  wire [512:0] from_t1_iter33_to_t1_iter34__dout;
  wire from_t1_iter33_to_t1_iter34__empty_n;
  wire from_t1_iter33_to_t1_iter34__read;
  wire [512:0] from_t1_iter33_to_t1_iter34__din;
  wire from_t1_iter33_to_t1_iter34__full_n;
  wire from_t1_iter33_to_t1_iter34__write;
  wire [512:0] from_t1_iter34_to_t1_iter35__dout;
  wire from_t1_iter34_to_t1_iter35__empty_n;
  wire from_t1_iter34_to_t1_iter35__read;
  wire [512:0] from_t1_iter34_to_t1_iter35__din;
  wire from_t1_iter34_to_t1_iter35__full_n;
  wire from_t1_iter34_to_t1_iter35__write;
  wire [512:0] from_t1_iter35_to_t1_iter36__dout;
  wire from_t1_iter35_to_t1_iter36__empty_n;
  wire from_t1_iter35_to_t1_iter36__read;
  wire [512:0] from_t1_iter35_to_t1_iter36__din;
  wire from_t1_iter35_to_t1_iter36__full_n;
  wire from_t1_iter35_to_t1_iter36__write;
  wire [512:0] from_t1_iter36_to_t1_iter37__dout;
  wire from_t1_iter36_to_t1_iter37__empty_n;
  wire from_t1_iter36_to_t1_iter37__read;
  wire [512:0] from_t1_iter36_to_t1_iter37__din;
  wire from_t1_iter36_to_t1_iter37__full_n;
  wire from_t1_iter36_to_t1_iter37__write;
  wire [512:0] from_t1_iter37_to_t1_iter38__dout;
  wire from_t1_iter37_to_t1_iter38__empty_n;
  wire from_t1_iter37_to_t1_iter38__read;
  wire [512:0] from_t1_iter37_to_t1_iter38__din;
  wire from_t1_iter37_to_t1_iter38__full_n;
  wire from_t1_iter37_to_t1_iter38__write;
  wire [512:0] from_t1_iter38_to_t1_iter39__dout;
  wire from_t1_iter38_to_t1_iter39__empty_n;
  wire from_t1_iter38_to_t1_iter39__read;
  wire [512:0] from_t1_iter38_to_t1_iter39__din;
  wire from_t1_iter38_to_t1_iter39__full_n;
  wire from_t1_iter38_to_t1_iter39__write;
  wire [512:0] from_t1_iter39_to_t1_iter40__dout;
  wire from_t1_iter39_to_t1_iter40__empty_n;
  wire from_t1_iter39_to_t1_iter40__read;
  wire [512:0] from_t1_iter39_to_t1_iter40__din;
  wire from_t1_iter39_to_t1_iter40__full_n;
  wire from_t1_iter39_to_t1_iter40__write;
  wire [512:0] from_t1_iter3_to_t1_iter4__dout;
  wire from_t1_iter3_to_t1_iter4__empty_n;
  wire from_t1_iter3_to_t1_iter4__read;
  wire [512:0] from_t1_iter3_to_t1_iter4__din;
  wire from_t1_iter3_to_t1_iter4__full_n;
  wire from_t1_iter3_to_t1_iter4__write;
  wire [512:0] from_t1_iter40_to_t1_iter41__dout;
  wire from_t1_iter40_to_t1_iter41__empty_n;
  wire from_t1_iter40_to_t1_iter41__read;
  wire [512:0] from_t1_iter40_to_t1_iter41__din;
  wire from_t1_iter40_to_t1_iter41__full_n;
  wire from_t1_iter40_to_t1_iter41__write;
  wire [512:0] from_t1_iter41_to_t1_iter42__dout;
  wire from_t1_iter41_to_t1_iter42__empty_n;
  wire from_t1_iter41_to_t1_iter42__read;
  wire [512:0] from_t1_iter41_to_t1_iter42__din;
  wire from_t1_iter41_to_t1_iter42__full_n;
  wire from_t1_iter41_to_t1_iter42__write;
  wire [512:0] from_t1_iter42_to_t1_iter43__dout;
  wire from_t1_iter42_to_t1_iter43__empty_n;
  wire from_t1_iter42_to_t1_iter43__read;
  wire [512:0] from_t1_iter42_to_t1_iter43__din;
  wire from_t1_iter42_to_t1_iter43__full_n;
  wire from_t1_iter42_to_t1_iter43__write;
  wire [512:0] from_t1_iter43_to_t1_iter44__dout;
  wire from_t1_iter43_to_t1_iter44__empty_n;
  wire from_t1_iter43_to_t1_iter44__read;
  wire [512:0] from_t1_iter43_to_t1_iter44__din;
  wire from_t1_iter43_to_t1_iter44__full_n;
  wire from_t1_iter43_to_t1_iter44__write;
  wire [512:0] from_t1_iter44_to_t1_iter45__dout;
  wire from_t1_iter44_to_t1_iter45__empty_n;
  wire from_t1_iter44_to_t1_iter45__read;
  wire [512:0] from_t1_iter44_to_t1_iter45__din;
  wire from_t1_iter44_to_t1_iter45__full_n;
  wire from_t1_iter44_to_t1_iter45__write;
  wire [512:0] from_t1_iter45_to_t1_iter46__dout;
  wire from_t1_iter45_to_t1_iter46__empty_n;
  wire from_t1_iter45_to_t1_iter46__read;
  wire [512:0] from_t1_iter45_to_t1_iter46__din;
  wire from_t1_iter45_to_t1_iter46__full_n;
  wire from_t1_iter45_to_t1_iter46__write;
  wire [512:0] from_t1_iter46_to_t1_iter47__dout;
  wire from_t1_iter46_to_t1_iter47__empty_n;
  wire from_t1_iter46_to_t1_iter47__read;
  wire [512:0] from_t1_iter46_to_t1_iter47__din;
  wire from_t1_iter46_to_t1_iter47__full_n;
  wire from_t1_iter46_to_t1_iter47__write;
  wire [512:0] from_t1_iter47_to_t1_iter48__dout;
  wire from_t1_iter47_to_t1_iter48__empty_n;
  wire from_t1_iter47_to_t1_iter48__read;
  wire [512:0] from_t1_iter47_to_t1_iter48__din;
  wire from_t1_iter47_to_t1_iter48__full_n;
  wire from_t1_iter47_to_t1_iter48__write;
  wire [512:0] from_t1_iter48_to_t1_iter49__dout;
  wire from_t1_iter48_to_t1_iter49__empty_n;
  wire from_t1_iter48_to_t1_iter49__read;
  wire [512:0] from_t1_iter48_to_t1_iter49__din;
  wire from_t1_iter48_to_t1_iter49__full_n;
  wire from_t1_iter48_to_t1_iter49__write;
  wire [512:0] from_t1_iter49_to_t1_iter50__dout;
  wire from_t1_iter49_to_t1_iter50__empty_n;
  wire from_t1_iter49_to_t1_iter50__read;
  wire [512:0] from_t1_iter49_to_t1_iter50__din;
  wire from_t1_iter49_to_t1_iter50__full_n;
  wire from_t1_iter49_to_t1_iter50__write;
  wire [512:0] from_t1_iter4_to_t1_iter5__dout;
  wire from_t1_iter4_to_t1_iter5__empty_n;
  wire from_t1_iter4_to_t1_iter5__read;
  wire [512:0] from_t1_iter4_to_t1_iter5__din;
  wire from_t1_iter4_to_t1_iter5__full_n;
  wire from_t1_iter4_to_t1_iter5__write;
  wire [512:0] from_t1_iter50_to_t1_iter51__dout;
  wire from_t1_iter50_to_t1_iter51__empty_n;
  wire from_t1_iter50_to_t1_iter51__read;
  wire [512:0] from_t1_iter50_to_t1_iter51__din;
  wire from_t1_iter50_to_t1_iter51__full_n;
  wire from_t1_iter50_to_t1_iter51__write;
  wire [512:0] from_t1_iter51_to_t1_iter52__dout;
  wire from_t1_iter51_to_t1_iter52__empty_n;
  wire from_t1_iter51_to_t1_iter52__read;
  wire [512:0] from_t1_iter51_to_t1_iter52__din;
  wire from_t1_iter51_to_t1_iter52__full_n;
  wire from_t1_iter51_to_t1_iter52__write;
  wire [512:0] from_t1_iter52_to_t1_iter53__dout;
  wire from_t1_iter52_to_t1_iter53__empty_n;
  wire from_t1_iter52_to_t1_iter53__read;
  wire [512:0] from_t1_iter52_to_t1_iter53__din;
  wire from_t1_iter52_to_t1_iter53__full_n;
  wire from_t1_iter52_to_t1_iter53__write;
  wire [512:0] from_t1_iter53_to_t1_iter54__dout;
  wire from_t1_iter53_to_t1_iter54__empty_n;
  wire from_t1_iter53_to_t1_iter54__read;
  wire [512:0] from_t1_iter53_to_t1_iter54__din;
  wire from_t1_iter53_to_t1_iter54__full_n;
  wire from_t1_iter53_to_t1_iter54__write;
  wire [512:0] from_t1_iter54_to_t1_iter55__dout;
  wire from_t1_iter54_to_t1_iter55__empty_n;
  wire from_t1_iter54_to_t1_iter55__read;
  wire [512:0] from_t1_iter54_to_t1_iter55__din;
  wire from_t1_iter54_to_t1_iter55__full_n;
  wire from_t1_iter54_to_t1_iter55__write;
  wire [512:0] from_t1_iter55_to_t1_iter56__dout;
  wire from_t1_iter55_to_t1_iter56__empty_n;
  wire from_t1_iter55_to_t1_iter56__read;
  wire [512:0] from_t1_iter55_to_t1_iter56__din;
  wire from_t1_iter55_to_t1_iter56__full_n;
  wire from_t1_iter55_to_t1_iter56__write;
  wire [512:0] from_t1_iter56_to_t1_iter57__dout;
  wire from_t1_iter56_to_t1_iter57__empty_n;
  wire from_t1_iter56_to_t1_iter57__read;
  wire [512:0] from_t1_iter56_to_t1_iter57__din;
  wire from_t1_iter56_to_t1_iter57__full_n;
  wire from_t1_iter56_to_t1_iter57__write;
  wire [512:0] from_t1_iter57_to_t1_iter58__dout;
  wire from_t1_iter57_to_t1_iter58__empty_n;
  wire from_t1_iter57_to_t1_iter58__read;
  wire [512:0] from_t1_iter57_to_t1_iter58__din;
  wire from_t1_iter57_to_t1_iter58__full_n;
  wire from_t1_iter57_to_t1_iter58__write;
  wire [512:0] from_t1_iter58_to_t1_iter59__dout;
  wire from_t1_iter58_to_t1_iter59__empty_n;
  wire from_t1_iter58_to_t1_iter59__read;
  wire [512:0] from_t1_iter58_to_t1_iter59__din;
  wire from_t1_iter58_to_t1_iter59__full_n;
  wire from_t1_iter58_to_t1_iter59__write;
  wire [512:0] from_t1_iter59_to_t1_iter60__dout;
  wire from_t1_iter59_to_t1_iter60__empty_n;
  wire from_t1_iter59_to_t1_iter60__read;
  wire [512:0] from_t1_iter59_to_t1_iter60__din;
  wire from_t1_iter59_to_t1_iter60__full_n;
  wire from_t1_iter59_to_t1_iter60__write;
  wire [512:0] from_t1_iter5_to_t1_iter6__dout;
  wire from_t1_iter5_to_t1_iter6__empty_n;
  wire from_t1_iter5_to_t1_iter6__read;
  wire [512:0] from_t1_iter5_to_t1_iter6__din;
  wire from_t1_iter5_to_t1_iter6__full_n;
  wire from_t1_iter5_to_t1_iter6__write;
  wire [512:0] from_t1_iter60_to_t1_iter61__dout;
  wire from_t1_iter60_to_t1_iter61__empty_n;
  wire from_t1_iter60_to_t1_iter61__read;
  wire [512:0] from_t1_iter60_to_t1_iter61__din;
  wire from_t1_iter60_to_t1_iter61__full_n;
  wire from_t1_iter60_to_t1_iter61__write;
  wire [512:0] from_t1_iter61_to_t1_iter62__dout;
  wire from_t1_iter61_to_t1_iter62__empty_n;
  wire from_t1_iter61_to_t1_iter62__read;
  wire [512:0] from_t1_iter61_to_t1_iter62__din;
  wire from_t1_iter61_to_t1_iter62__full_n;
  wire from_t1_iter61_to_t1_iter62__write;
  wire [512:0] from_t1_iter62_to_t1_iter63__dout;
  wire from_t1_iter62_to_t1_iter63__empty_n;
  wire from_t1_iter62_to_t1_iter63__read;
  wire [512:0] from_t1_iter62_to_t1_iter63__din;
  wire from_t1_iter62_to_t1_iter63__full_n;
  wire from_t1_iter62_to_t1_iter63__write;
  wire [512:0] from_t1_iter63_to_t1_iter64__dout;
  wire from_t1_iter63_to_t1_iter64__empty_n;
  wire from_t1_iter63_to_t1_iter64__read;
  wire [512:0] from_t1_iter63_to_t1_iter64__din;
  wire from_t1_iter63_to_t1_iter64__full_n;
  wire from_t1_iter63_to_t1_iter64__write;
  wire [512:0] from_t1_iter64_to_t1_iter65__dout;
  wire from_t1_iter64_to_t1_iter65__empty_n;
  wire from_t1_iter64_to_t1_iter65__read;
  wire [512:0] from_t1_iter64_to_t1_iter65__din;
  wire from_t1_iter64_to_t1_iter65__full_n;
  wire from_t1_iter64_to_t1_iter65__write;
  wire [512:0] from_t1_iter65_to_t1_iter66__dout;
  wire from_t1_iter65_to_t1_iter66__empty_n;
  wire from_t1_iter65_to_t1_iter66__read;
  wire [512:0] from_t1_iter65_to_t1_iter66__din;
  wire from_t1_iter65_to_t1_iter66__full_n;
  wire from_t1_iter65_to_t1_iter66__write;
  wire [512:0] from_t1_iter66_to_t1_iter67__dout;
  wire from_t1_iter66_to_t1_iter67__empty_n;
  wire from_t1_iter66_to_t1_iter67__read;
  wire [512:0] from_t1_iter66_to_t1_iter67__din;
  wire from_t1_iter66_to_t1_iter67__full_n;
  wire from_t1_iter66_to_t1_iter67__write;
  wire [512:0] from_t1_iter67_to_t1_iter68__dout;
  wire from_t1_iter67_to_t1_iter68__empty_n;
  wire from_t1_iter67_to_t1_iter68__read;
  wire [512:0] from_t1_iter67_to_t1_iter68__din;
  wire from_t1_iter67_to_t1_iter68__full_n;
  wire from_t1_iter67_to_t1_iter68__write;
  wire [512:0] from_t1_iter68_to_t1_iter69__dout;
  wire from_t1_iter68_to_t1_iter69__empty_n;
  wire from_t1_iter68_to_t1_iter69__read;
  wire [512:0] from_t1_iter68_to_t1_iter69__din;
  wire from_t1_iter68_to_t1_iter69__full_n;
  wire from_t1_iter68_to_t1_iter69__write;
  wire [512:0] from_t1_iter69_to_t1_iter70__dout;
  wire from_t1_iter69_to_t1_iter70__empty_n;
  wire from_t1_iter69_to_t1_iter70__read;
  wire [512:0] from_t1_iter69_to_t1_iter70__din;
  wire from_t1_iter69_to_t1_iter70__full_n;
  wire from_t1_iter69_to_t1_iter70__write;
  wire [512:0] from_t1_iter6_to_t1_iter7__dout;
  wire from_t1_iter6_to_t1_iter7__empty_n;
  wire from_t1_iter6_to_t1_iter7__read;
  wire [512:0] from_t1_iter6_to_t1_iter7__din;
  wire from_t1_iter6_to_t1_iter7__full_n;
  wire from_t1_iter6_to_t1_iter7__write;
  wire [512:0] from_t1_iter70_to_t1_iter71__dout;
  wire from_t1_iter70_to_t1_iter71__empty_n;
  wire from_t1_iter70_to_t1_iter71__read;
  wire [512:0] from_t1_iter70_to_t1_iter71__din;
  wire from_t1_iter70_to_t1_iter71__full_n;
  wire from_t1_iter70_to_t1_iter71__write;
  wire [512:0] from_t1_iter71_to_t1_iter72__dout;
  wire from_t1_iter71_to_t1_iter72__empty_n;
  wire from_t1_iter71_to_t1_iter72__read;
  wire [512:0] from_t1_iter71_to_t1_iter72__din;
  wire from_t1_iter71_to_t1_iter72__full_n;
  wire from_t1_iter71_to_t1_iter72__write;
  wire [512:0] from_t1_iter72_to_t1_iter73__dout;
  wire from_t1_iter72_to_t1_iter73__empty_n;
  wire from_t1_iter72_to_t1_iter73__read;
  wire [512:0] from_t1_iter72_to_t1_iter73__din;
  wire from_t1_iter72_to_t1_iter73__full_n;
  wire from_t1_iter72_to_t1_iter73__write;
  wire [512:0] from_t1_iter73_to_t1_iter74__dout;
  wire from_t1_iter73_to_t1_iter74__empty_n;
  wire from_t1_iter73_to_t1_iter74__read;
  wire [512:0] from_t1_iter73_to_t1_iter74__din;
  wire from_t1_iter73_to_t1_iter74__full_n;
  wire from_t1_iter73_to_t1_iter74__write;
  wire [512:0] from_t1_iter74_to_t1_iter75__dout;
  wire from_t1_iter74_to_t1_iter75__empty_n;
  wire from_t1_iter74_to_t1_iter75__read;
  wire [512:0] from_t1_iter74_to_t1_iter75__din;
  wire from_t1_iter74_to_t1_iter75__full_n;
  wire from_t1_iter74_to_t1_iter75__write;
  wire [512:0] from_t1_iter75_to_t1_iter76__dout;
  wire from_t1_iter75_to_t1_iter76__empty_n;
  wire from_t1_iter75_to_t1_iter76__read;
  wire [512:0] from_t1_iter75_to_t1_iter76__din;
  wire from_t1_iter75_to_t1_iter76__full_n;
  wire from_t1_iter75_to_t1_iter76__write;
  wire [512:0] from_t1_iter76_to_t1_iter77__dout;
  wire from_t1_iter76_to_t1_iter77__empty_n;
  wire from_t1_iter76_to_t1_iter77__read;
  wire [512:0] from_t1_iter76_to_t1_iter77__din;
  wire from_t1_iter76_to_t1_iter77__full_n;
  wire from_t1_iter76_to_t1_iter77__write;
  wire [512:0] from_t1_iter77_to_t1_iter78__dout;
  wire from_t1_iter77_to_t1_iter78__empty_n;
  wire from_t1_iter77_to_t1_iter78__read;
  wire [512:0] from_t1_iter77_to_t1_iter78__din;
  wire from_t1_iter77_to_t1_iter78__full_n;
  wire from_t1_iter77_to_t1_iter78__write;
  wire [512:0] from_t1_iter78_to_t1_iter79__dout;
  wire from_t1_iter78_to_t1_iter79__empty_n;
  wire from_t1_iter78_to_t1_iter79__read;
  wire [512:0] from_t1_iter78_to_t1_iter79__din;
  wire from_t1_iter78_to_t1_iter79__full_n;
  wire from_t1_iter78_to_t1_iter79__write;
  wire [512:0] from_t1_iter79_to_t1_iter80__dout;
  wire from_t1_iter79_to_t1_iter80__empty_n;
  wire from_t1_iter79_to_t1_iter80__read;
  wire [512:0] from_t1_iter79_to_t1_iter80__din;
  wire from_t1_iter79_to_t1_iter80__full_n;
  wire from_t1_iter79_to_t1_iter80__write;
  wire [512:0] from_t1_iter7_to_t1_iter8__dout;
  wire from_t1_iter7_to_t1_iter8__empty_n;
  wire from_t1_iter7_to_t1_iter8__read;
  wire [512:0] from_t1_iter7_to_t1_iter8__din;
  wire from_t1_iter7_to_t1_iter8__full_n;
  wire from_t1_iter7_to_t1_iter8__write;
  wire [512:0] from_t1_iter80_to_t1_iter81__dout;
  wire from_t1_iter80_to_t1_iter81__empty_n;
  wire from_t1_iter80_to_t1_iter81__read;
  wire [512:0] from_t1_iter80_to_t1_iter81__din;
  wire from_t1_iter80_to_t1_iter81__full_n;
  wire from_t1_iter80_to_t1_iter81__write;
  wire [512:0] from_t1_iter81_to_t1_iter82__dout;
  wire from_t1_iter81_to_t1_iter82__empty_n;
  wire from_t1_iter81_to_t1_iter82__read;
  wire [512:0] from_t1_iter81_to_t1_iter82__din;
  wire from_t1_iter81_to_t1_iter82__full_n;
  wire from_t1_iter81_to_t1_iter82__write;
  wire [512:0] from_t1_iter82_to_t1_iter83__dout;
  wire from_t1_iter82_to_t1_iter83__empty_n;
  wire from_t1_iter82_to_t1_iter83__read;
  wire [512:0] from_t1_iter82_to_t1_iter83__din;
  wire from_t1_iter82_to_t1_iter83__full_n;
  wire from_t1_iter82_to_t1_iter83__write;
  wire [512:0] from_t1_iter83_to_t1_iter84__dout;
  wire from_t1_iter83_to_t1_iter84__empty_n;
  wire from_t1_iter83_to_t1_iter84__read;
  wire [512:0] from_t1_iter83_to_t1_iter84__din;
  wire from_t1_iter83_to_t1_iter84__full_n;
  wire from_t1_iter83_to_t1_iter84__write;
  wire [512:0] from_t1_iter84_to_t1_iter85__dout;
  wire from_t1_iter84_to_t1_iter85__empty_n;
  wire from_t1_iter84_to_t1_iter85__read;
  wire [512:0] from_t1_iter84_to_t1_iter85__din;
  wire from_t1_iter84_to_t1_iter85__full_n;
  wire from_t1_iter84_to_t1_iter85__write;
  wire [512:0] from_t1_iter85_to_t1_iter86__dout;
  wire from_t1_iter85_to_t1_iter86__empty_n;
  wire from_t1_iter85_to_t1_iter86__read;
  wire [512:0] from_t1_iter85_to_t1_iter86__din;
  wire from_t1_iter85_to_t1_iter86__full_n;
  wire from_t1_iter85_to_t1_iter86__write;
  wire [512:0] from_t1_iter86_to_t1_iter87__dout;
  wire from_t1_iter86_to_t1_iter87__empty_n;
  wire from_t1_iter86_to_t1_iter87__read;
  wire [512:0] from_t1_iter86_to_t1_iter87__din;
  wire from_t1_iter86_to_t1_iter87__full_n;
  wire from_t1_iter86_to_t1_iter87__write;
  wire [512:0] from_t1_iter87_to_t1_iter88__dout;
  wire from_t1_iter87_to_t1_iter88__empty_n;
  wire from_t1_iter87_to_t1_iter88__read;
  wire [512:0] from_t1_iter87_to_t1_iter88__din;
  wire from_t1_iter87_to_t1_iter88__full_n;
  wire from_t1_iter87_to_t1_iter88__write;
  wire [512:0] from_t1_iter88_to_t1_iter89__dout;
  wire from_t1_iter88_to_t1_iter89__empty_n;
  wire from_t1_iter88_to_t1_iter89__read;
  wire [512:0] from_t1_iter88_to_t1_iter89__din;
  wire from_t1_iter88_to_t1_iter89__full_n;
  wire from_t1_iter88_to_t1_iter89__write;
  wire [512:0] from_t1_iter89_to_t1_iter90__dout;
  wire from_t1_iter89_to_t1_iter90__empty_n;
  wire from_t1_iter89_to_t1_iter90__read;
  wire [512:0] from_t1_iter89_to_t1_iter90__din;
  wire from_t1_iter89_to_t1_iter90__full_n;
  wire from_t1_iter89_to_t1_iter90__write;
  wire [512:0] from_t1_iter8_to_t1_iter9__dout;
  wire from_t1_iter8_to_t1_iter9__empty_n;
  wire from_t1_iter8_to_t1_iter9__read;
  wire [512:0] from_t1_iter8_to_t1_iter9__din;
  wire from_t1_iter8_to_t1_iter9__full_n;
  wire from_t1_iter8_to_t1_iter9__write;
  wire [512:0] from_t1_iter90_to_t1_iter91__dout;
  wire from_t1_iter90_to_t1_iter91__empty_n;
  wire from_t1_iter90_to_t1_iter91__read;
  wire [512:0] from_t1_iter90_to_t1_iter91__din;
  wire from_t1_iter90_to_t1_iter91__full_n;
  wire from_t1_iter90_to_t1_iter91__write;
  wire [512:0] from_t1_iter91_to_t1_iter92__dout;
  wire from_t1_iter91_to_t1_iter92__empty_n;
  wire from_t1_iter91_to_t1_iter92__read;
  wire [512:0] from_t1_iter91_to_t1_iter92__din;
  wire from_t1_iter91_to_t1_iter92__full_n;
  wire from_t1_iter91_to_t1_iter92__write;
  wire [512:0] from_t1_iter92_to_t1_iter93__dout;
  wire from_t1_iter92_to_t1_iter93__empty_n;
  wire from_t1_iter92_to_t1_iter93__read;
  wire [512:0] from_t1_iter92_to_t1_iter93__din;
  wire from_t1_iter92_to_t1_iter93__full_n;
  wire from_t1_iter92_to_t1_iter93__write;
  wire [512:0] from_t1_iter93_to_t1_iter94__dout;
  wire from_t1_iter93_to_t1_iter94__empty_n;
  wire from_t1_iter93_to_t1_iter94__read;
  wire [512:0] from_t1_iter93_to_t1_iter94__din;
  wire from_t1_iter93_to_t1_iter94__full_n;
  wire from_t1_iter93_to_t1_iter94__write;
  wire [512:0] from_t1_iter94_to_t1_iter95__dout;
  wire from_t1_iter94_to_t1_iter95__empty_n;
  wire from_t1_iter94_to_t1_iter95__read;
  wire [512:0] from_t1_iter94_to_t1_iter95__din;
  wire from_t1_iter94_to_t1_iter95__full_n;
  wire from_t1_iter94_to_t1_iter95__write;
  wire [512:0] from_t1_iter95_to_t1_iter96__dout;
  wire from_t1_iter95_to_t1_iter96__empty_n;
  wire from_t1_iter95_to_t1_iter96__read;
  wire [512:0] from_t1_iter95_to_t1_iter96__din;
  wire from_t1_iter95_to_t1_iter96__full_n;
  wire from_t1_iter95_to_t1_iter96__write;
  wire [512:0] from_t1_iter96_to_t1_iter97__dout;
  wire from_t1_iter96_to_t1_iter97__empty_n;
  wire from_t1_iter96_to_t1_iter97__read;
  wire [512:0] from_t1_iter96_to_t1_iter97__din;
  wire from_t1_iter96_to_t1_iter97__full_n;
  wire from_t1_iter96_to_t1_iter97__write;
  wire [512:0] from_t1_iter97_to_t1_iter98__dout;
  wire from_t1_iter97_to_t1_iter98__empty_n;
  wire from_t1_iter97_to_t1_iter98__read;
  wire [512:0] from_t1_iter97_to_t1_iter98__din;
  wire from_t1_iter97_to_t1_iter98__full_n;
  wire from_t1_iter97_to_t1_iter98__write;
  wire [512:0] from_t1_iter98_to_t1_iter99__dout;
  wire from_t1_iter98_to_t1_iter99__empty_n;
  wire from_t1_iter98_to_t1_iter99__read;
  wire [512:0] from_t1_iter98_to_t1_iter99__din;
  wire from_t1_iter98_to_t1_iter99__full_n;
  wire from_t1_iter98_to_t1_iter99__write;
  wire [512:0] from_t1_iter99_to_t1_iter100__dout;
  wire from_t1_iter99_to_t1_iter100__empty_n;
  wire from_t1_iter99_to_t1_iter100__read;
  wire [512:0] from_t1_iter99_to_t1_iter100__din;
  wire from_t1_iter99_to_t1_iter100__full_n;
  wire from_t1_iter99_to_t1_iter100__write;
  wire [512:0] from_t1_iter9_to_t1_iter10__dout;
  wire from_t1_iter9_to_t1_iter10__empty_n;
  wire from_t1_iter9_to_t1_iter10__read;
  wire [512:0] from_t1_iter9_to_t1_iter10__din;
  wire from_t1_iter9_to_t1_iter10__full_n;
  wire from_t1_iter9_to_t1_iter10__write;
  wire [63:0] BurstRead_floatx16_0___bank_0_t1__q0;
  wire [63:0] bank_0_t1_read_addr__din;
  wire bank_0_t1_read_addr__full_n;
  wire bank_0_t1_read_addr__write;
  wire [511:0] bank_0_t1_read_data__dout;
  wire bank_0_t1_read_data__empty_n;
  wire bank_0_t1_read_data__read;
  wire [63:0] bank_0_t1_write_addr__din;
  wire bank_0_t1_write_addr__full_n;
  wire bank_0_t1_write_addr__write;
  wire [511:0] bank_0_t1_write_data__din;
  wire bank_0_t1_write_data__full_n;
  wire bank_0_t1_write_data__write;
  wire [7:0] bank_0_t1_write_resp__dout;
  wire bank_0_t1_write_resp__empty_n;
  wire bank_0_t1_write_resp__read;
  wire [63:0] BurstRead_floatx16_0___coalesced_data_num__q0;
  wire BurstRead_floatx16_0__ap_start;
  wire BurstRead_floatx16_0__ap_ready;
  wire BurstRead_floatx16_0__ap_done;
  wire BurstRead_floatx16_0__ap_idle;
  wire [63:0] BurstWrite_floatx16_0___bank_1_t0__q0;
  wire [63:0] bank_1_t0_read_addr__din;
  wire bank_1_t0_read_addr__full_n;
  wire bank_1_t0_read_addr__write;
  wire [511:0] bank_1_t0_read_data__dout;
  wire bank_1_t0_read_data__empty_n;
  wire bank_1_t0_read_data__read;
  wire [63:0] bank_1_t0_write_addr__din;
  wire bank_1_t0_write_addr__full_n;
  wire bank_1_t0_write_addr__write;
  wire [511:0] bank_1_t0_write_data__din;
  wire bank_1_t0_write_data__full_n;
  wire bank_1_t0_write_data__write;
  wire [7:0] bank_1_t0_write_resp__dout;
  wire bank_1_t0_write_resp__empty_n;
  wire bank_1_t0_write_resp__read;
  wire [63:0] BurstWrite_floatx16_0___coalesced_data_num__q0;
  wire BurstWrite_floatx16_0__ap_start;
  wire BurstWrite_floatx16_0__ap_ready;
  wire BurstWrite_floatx16_0__ap_done;
  wire BurstWrite_floatx16_0__ap_idle;
  wire Module0Func_0__ap_start;
  wire Module1Func_0__ap_start;
  wire Module2Func_0__ap_start;
  wire Module2Func_1__ap_start;
  wire Module2Func_2__ap_start;
  wire Module2Func_3__ap_start;
  wire Module2Func_4__ap_start;
  wire Module2Func_5__ap_start;
  wire Module2Func_6__ap_start;
  wire Module2Func_7__ap_start;
  wire Module2Func_8__ap_start;
  wire Module2Func_9__ap_start;
  wire Module2Func_10__ap_start;
  wire Module2Func_11__ap_start;
  wire Module2Func_12__ap_start;
  wire Module2Func_13__ap_start;
  wire Module2Func_14__ap_start;
  wire Module2Func_15__ap_start;
  wire Module2Func_16__ap_start;
  wire Module2Func_17__ap_start;
  wire Module2Func_18__ap_start;
  wire Module2Func_19__ap_start;
  wire Module2Func_20__ap_start;
  wire Module2Func_21__ap_start;
  wire Module2Func_22__ap_start;
  wire Module2Func_23__ap_start;
  wire Module2Func_24__ap_start;
  wire Module2Func_25__ap_start;
  wire Module2Func_26__ap_start;
  wire Module2Func_27__ap_start;
  wire Module2Func_28__ap_start;
  wire Module2Func_29__ap_start;
  wire Module2Func_30__ap_start;
  wire Module2Func_31__ap_start;
  wire Module2Func_32__ap_start;
  wire Module2Func_33__ap_start;
  wire Module2Func_34__ap_start;
  wire Module2Func_35__ap_start;
  wire Module2Func_36__ap_start;
  wire Module2Func_37__ap_start;
  wire Module2Func_38__ap_start;
  wire Module2Func_39__ap_start;
  wire Module2Func_40__ap_start;
  wire Module2Func_41__ap_start;
  wire Module2Func_42__ap_start;
  wire Module2Func_43__ap_start;
  wire Module2Func_44__ap_start;
  wire Module2Func_45__ap_start;
  wire Module2Func_46__ap_start;
  wire Module2Func_47__ap_start;
  wire Module2Func_48__ap_start;
  wire Module2Func_49__ap_start;
  wire Module2Func_50__ap_start;
  wire Module2Func_51__ap_start;
  wire Module2Func_52__ap_start;
  wire Module2Func_53__ap_start;
  wire Module2Func_54__ap_start;
  wire Module2Func_55__ap_start;
  wire Module2Func_56__ap_start;
  wire Module2Func_57__ap_start;
  wire Module2Func_58__ap_start;
  wire Module2Func_59__ap_start;
  wire Module2Func_60__ap_start;
  wire Module2Func_61__ap_start;
  wire Module2Func_62__ap_start;
  wire Module2Func_63__ap_start;
  wire Module2Func_64__ap_start;
  wire Module2Func_65__ap_start;
  wire Module2Func_66__ap_start;
  wire Module2Func_67__ap_start;
  wire Module2Func_68__ap_start;
  wire Module2Func_69__ap_start;
  wire Module2Func_70__ap_start;
  wire Module2Func_71__ap_start;
  wire Module2Func_72__ap_start;
  wire Module2Func_73__ap_start;
  wire Module2Func_74__ap_start;
  wire Module2Func_75__ap_start;
  wire Module2Func_76__ap_start;
  wire Module2Func_77__ap_start;
  wire Module2Func_78__ap_start;
  wire Module2Func_79__ap_start;
  wire Module2Func_80__ap_start;
  wire Module2Func_81__ap_start;
  wire Module2Func_82__ap_start;
  wire Module2Func_83__ap_start;
  wire Module2Func_84__ap_start;
  wire Module2Func_85__ap_start;
  wire Module2Func_86__ap_start;
  wire Module2Func_87__ap_start;
  wire Module2Func_88__ap_start;
  wire Module2Func_89__ap_start;
  wire Module2Func_90__ap_start;
  wire Module2Func_91__ap_start;
  wire Module2Func_92__ap_start;
  wire Module2Func_93__ap_start;
  wire Module2Func_94__ap_start;
  wire Module2Func_95__ap_start;
  wire Module2Func_96__ap_start;
  wire Module2Func_97__ap_start;
  wire Module2Func_98__ap_start;
  wire Module2Func_99__ap_start;
  wire Module2Func_100__ap_start;
  wire Module2Func_101__ap_start;
  wire Module2Func_102__ap_start;
  wire Module2Func_103__ap_start;
  wire Module2Func_104__ap_start;
  wire Module2Func_105__ap_start;
  wire Module2Func_106__ap_start;
  wire Module2Func_107__ap_start;
  wire Module3Func_0__ap_start;
  wire ap_rst_n_inv;
  wire ap_done;
  wire ap_idle;
  wire ap_ready;

  jacobi3d_kernel_control_s_axi
  #(
    .C_S_AXI_ADDR_WIDTH(C_S_AXI_CONTROL_ADDR_WIDTH),
    .C_S_AXI_DATA_WIDTH(C_S_AXI_CONTROL_DATA_WIDTH)
  )
  control_s_axi_U
  (
    .AWVALID(s_axi_control_AWVALID),
    .AWREADY(s_axi_control_AWREADY),
    .AWADDR(s_axi_control_AWADDR),
    .WVALID(s_axi_control_WVALID),
    .WREADY(s_axi_control_WREADY),
    .WDATA(s_axi_control_WDATA),
    .WSTRB(s_axi_control_WSTRB),
    .ARVALID(s_axi_control_ARVALID),
    .ARREADY(s_axi_control_ARREADY),
    .ARADDR(s_axi_control_ARADDR),
    .RVALID(s_axi_control_RVALID),
    .RREADY(s_axi_control_RREADY),
    .RDATA(s_axi_control_RDATA),
    .RRESP(s_axi_control_RRESP),
    .BVALID(s_axi_control_BVALID),
    .BREADY(s_axi_control_BREADY),
    .BRESP(s_axi_control_BRESP),
    .ACLK(ap_clk),
    .ARESET(ap_rst_n_inv),
    .ACLK_EN(1'b1),
    .bank_1_t0(bank_1_t0),
    .bank_0_t1(bank_0_t1),
    .coalesced_data_num(coalesced_data_num),
    .ap_start(ap_start),
    .interrupt(interrupt),
    .ap_ready(ap_ready),
    .ap_done(ap_done),
    .ap_idle(ap_idle)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(12),
    .DEPTH(4096)
  )
  bank_0_t1_buf
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(bank_0_t1_buf__dout),
    .if_empty_n(bank_0_t1_buf__empty_n),
    .if_read(bank_0_t1_buf__read),
    .if_read_ce(1'b1),
    .if_din(bank_0_t1_buf__din),
    .if_full_n(bank_0_t1_buf__full_n),
    .if_write(bank_0_t1_buf__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(12),
    .DEPTH(4096)
  )
  bank_1_t0_buf
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(bank_1_t0_buf__dout),
    .if_empty_n(bank_1_t0_buf__empty_n),
    .if_read(bank_1_t0_buf__read),
    .if_read_ce(1'b1),
    .if_din(bank_1_t0_buf__din),
    .if_full_n(bank_1_t0_buf__full_n),
    .if_write(bank_1_t0_buf__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t0_to_t0_bank_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t0_to_t0_bank_1__dout),
    .if_empty_n(from_t0_to_t0_bank_1__empty_n),
    .if_read(from_t0_to_t0_bank_1__read),
    .if_read_ce(1'b1),
    .if_din(from_t0_to_t0_bank_1__din),
    .if_full_n(from_t0_to_t0_bank_1__full_n),
    .if_write(from_t0_to_t0_bank_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_bank_0_to_t1_iter1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_bank_0_to_t1_iter1__dout),
    .if_empty_n(from_t1_bank_0_to_t1_iter1__empty_n),
    .if_read(from_t1_bank_0_to_t1_iter1__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_bank_0_to_t1_iter1__din),
    .if_full_n(from_t1_bank_0_to_t1_iter1__full_n),
    .if_write(from_t1_bank_0_to_t1_iter1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter100_to_t1_iter101
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter100_to_t1_iter101__dout),
    .if_empty_n(from_t1_iter100_to_t1_iter101__empty_n),
    .if_read(from_t1_iter100_to_t1_iter101__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter100_to_t1_iter101__din),
    .if_full_n(from_t1_iter100_to_t1_iter101__full_n),
    .if_write(from_t1_iter100_to_t1_iter101__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter101_to_t1_iter102
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter101_to_t1_iter102__dout),
    .if_empty_n(from_t1_iter101_to_t1_iter102__empty_n),
    .if_read(from_t1_iter101_to_t1_iter102__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter101_to_t1_iter102__din),
    .if_full_n(from_t1_iter101_to_t1_iter102__full_n),
    .if_write(from_t1_iter101_to_t1_iter102__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(136)
  )
  from_t1_iter102_to_t1_iter103
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter102_to_t1_iter103__dout),
    .if_empty_n(from_t1_iter102_to_t1_iter103__empty_n),
    .if_read(from_t1_iter102_to_t1_iter103__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter102_to_t1_iter103__din),
    .if_full_n(from_t1_iter102_to_t1_iter103__full_n),
    .if_write(from_t1_iter102_to_t1_iter103__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter103_to_t1_iter104
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter103_to_t1_iter104__dout),
    .if_empty_n(from_t1_iter103_to_t1_iter104__empty_n),
    .if_read(from_t1_iter103_to_t1_iter104__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter103_to_t1_iter104__din),
    .if_full_n(from_t1_iter103_to_t1_iter104__full_n),
    .if_write(from_t1_iter103_to_t1_iter104__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter104_to_t1_iter105
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter104_to_t1_iter105__dout),
    .if_empty_n(from_t1_iter104_to_t1_iter105__empty_n),
    .if_read(from_t1_iter104_to_t1_iter105__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter104_to_t1_iter105__din),
    .if_full_n(from_t1_iter104_to_t1_iter105__full_n),
    .if_write(from_t1_iter104_to_t1_iter105__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter105_to_t1_iter106
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter105_to_t1_iter106__dout),
    .if_empty_n(from_t1_iter105_to_t1_iter106__empty_n),
    .if_read(from_t1_iter105_to_t1_iter106__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter105_to_t1_iter106__din),
    .if_full_n(from_t1_iter105_to_t1_iter106__full_n),
    .if_write(from_t1_iter105_to_t1_iter106__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(140)
  )
  from_t1_iter106_to_t1_iter107
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter106_to_t1_iter107__dout),
    .if_empty_n(from_t1_iter106_to_t1_iter107__empty_n),
    .if_read(from_t1_iter106_to_t1_iter107__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter106_to_t1_iter107__din),
    .if_full_n(from_t1_iter106_to_t1_iter107__full_n),
    .if_write(from_t1_iter106_to_t1_iter107__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter107_to_t1_iter108
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter107_to_t1_iter108__dout),
    .if_empty_n(from_t1_iter107_to_t1_iter108__empty_n),
    .if_read(from_t1_iter107_to_t1_iter108__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter107_to_t1_iter108__din),
    .if_full_n(from_t1_iter107_to_t1_iter108__full_n),
    .if_write(from_t1_iter107_to_t1_iter108__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter108_to_t0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter108_to_t0__dout),
    .if_empty_n(from_t1_iter108_to_t0__empty_n),
    .if_read(from_t1_iter108_to_t0__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter108_to_t0__din),
    .if_full_n(from_t1_iter108_to_t0__full_n),
    .if_write(from_t1_iter108_to_t0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(130)
  )
  from_t1_iter10_to_t1_iter11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter10_to_t1_iter11__dout),
    .if_empty_n(from_t1_iter10_to_t1_iter11__empty_n),
    .if_read(from_t1_iter10_to_t1_iter11__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter10_to_t1_iter11__din),
    .if_full_n(from_t1_iter10_to_t1_iter11__full_n),
    .if_write(from_t1_iter10_to_t1_iter11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(132)
  )
  from_t1_iter11_to_t1_iter12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter11_to_t1_iter12__dout),
    .if_empty_n(from_t1_iter11_to_t1_iter12__empty_n),
    .if_read(from_t1_iter11_to_t1_iter12__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter11_to_t1_iter12__din),
    .if_full_n(from_t1_iter11_to_t1_iter12__full_n),
    .if_write(from_t1_iter11_to_t1_iter12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter12_to_t1_iter13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter12_to_t1_iter13__dout),
    .if_empty_n(from_t1_iter12_to_t1_iter13__empty_n),
    .if_read(from_t1_iter12_to_t1_iter13__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter12_to_t1_iter13__din),
    .if_full_n(from_t1_iter12_to_t1_iter13__full_n),
    .if_write(from_t1_iter12_to_t1_iter13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(140)
  )
  from_t1_iter13_to_t1_iter14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter13_to_t1_iter14__dout),
    .if_empty_n(from_t1_iter13_to_t1_iter14__empty_n),
    .if_read(from_t1_iter13_to_t1_iter14__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter13_to_t1_iter14__din),
    .if_full_n(from_t1_iter13_to_t1_iter14__full_n),
    .if_write(from_t1_iter13_to_t1_iter14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(130)
  )
  from_t1_iter14_to_t1_iter15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter14_to_t1_iter15__dout),
    .if_empty_n(from_t1_iter14_to_t1_iter15__empty_n),
    .if_read(from_t1_iter14_to_t1_iter15__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter14_to_t1_iter15__din),
    .if_full_n(from_t1_iter14_to_t1_iter15__full_n),
    .if_write(from_t1_iter14_to_t1_iter15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter15_to_t1_iter16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter15_to_t1_iter16__dout),
    .if_empty_n(from_t1_iter15_to_t1_iter16__empty_n),
    .if_read(from_t1_iter15_to_t1_iter16__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter15_to_t1_iter16__din),
    .if_full_n(from_t1_iter15_to_t1_iter16__full_n),
    .if_write(from_t1_iter15_to_t1_iter16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter16_to_t1_iter17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter16_to_t1_iter17__dout),
    .if_empty_n(from_t1_iter16_to_t1_iter17__empty_n),
    .if_read(from_t1_iter16_to_t1_iter17__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter16_to_t1_iter17__din),
    .if_full_n(from_t1_iter16_to_t1_iter17__full_n),
    .if_write(from_t1_iter16_to_t1_iter17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter17_to_t1_iter18
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter17_to_t1_iter18__dout),
    .if_empty_n(from_t1_iter17_to_t1_iter18__empty_n),
    .if_read(from_t1_iter17_to_t1_iter18__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter17_to_t1_iter18__din),
    .if_full_n(from_t1_iter17_to_t1_iter18__full_n),
    .if_write(from_t1_iter17_to_t1_iter18__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter18_to_t1_iter19
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter18_to_t1_iter19__dout),
    .if_empty_n(from_t1_iter18_to_t1_iter19__empty_n),
    .if_read(from_t1_iter18_to_t1_iter19__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter18_to_t1_iter19__din),
    .if_full_n(from_t1_iter18_to_t1_iter19__full_n),
    .if_write(from_t1_iter18_to_t1_iter19__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter19_to_t1_iter20
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter19_to_t1_iter20__dout),
    .if_empty_n(from_t1_iter19_to_t1_iter20__empty_n),
    .if_read(from_t1_iter19_to_t1_iter20__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter19_to_t1_iter20__din),
    .if_full_n(from_t1_iter19_to_t1_iter20__full_n),
    .if_write(from_t1_iter19_to_t1_iter20__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter1_to_t1_iter2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter1_to_t1_iter2__dout),
    .if_empty_n(from_t1_iter1_to_t1_iter2__empty_n),
    .if_read(from_t1_iter1_to_t1_iter2__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter1_to_t1_iter2__din),
    .if_full_n(from_t1_iter1_to_t1_iter2__full_n),
    .if_write(from_t1_iter1_to_t1_iter2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(130)
  )
  from_t1_iter20_to_t1_iter21
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter20_to_t1_iter21__dout),
    .if_empty_n(from_t1_iter20_to_t1_iter21__empty_n),
    .if_read(from_t1_iter20_to_t1_iter21__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter20_to_t1_iter21__din),
    .if_full_n(from_t1_iter20_to_t1_iter21__full_n),
    .if_write(from_t1_iter20_to_t1_iter21__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(132)
  )
  from_t1_iter21_to_t1_iter22
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter21_to_t1_iter22__dout),
    .if_empty_n(from_t1_iter21_to_t1_iter22__empty_n),
    .if_read(from_t1_iter21_to_t1_iter22__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter21_to_t1_iter22__din),
    .if_full_n(from_t1_iter21_to_t1_iter22__full_n),
    .if_write(from_t1_iter21_to_t1_iter22__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter22_to_t1_iter23
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter22_to_t1_iter23__dout),
    .if_empty_n(from_t1_iter22_to_t1_iter23__empty_n),
    .if_read(from_t1_iter22_to_t1_iter23__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter22_to_t1_iter23__din),
    .if_full_n(from_t1_iter22_to_t1_iter23__full_n),
    .if_write(from_t1_iter22_to_t1_iter23__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(130)
  )
  from_t1_iter23_to_t1_iter24
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter23_to_t1_iter24__dout),
    .if_empty_n(from_t1_iter23_to_t1_iter24__empty_n),
    .if_read(from_t1_iter23_to_t1_iter24__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter23_to_t1_iter24__din),
    .if_full_n(from_t1_iter23_to_t1_iter24__full_n),
    .if_write(from_t1_iter23_to_t1_iter24__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(130)
  )
  from_t1_iter24_to_t1_iter25
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter24_to_t1_iter25__dout),
    .if_empty_n(from_t1_iter24_to_t1_iter25__empty_n),
    .if_read(from_t1_iter24_to_t1_iter25__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter24_to_t1_iter25__din),
    .if_full_n(from_t1_iter24_to_t1_iter25__full_n),
    .if_write(from_t1_iter24_to_t1_iter25__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(130)
  )
  from_t1_iter25_to_t1_iter26
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter25_to_t1_iter26__dout),
    .if_empty_n(from_t1_iter25_to_t1_iter26__empty_n),
    .if_read(from_t1_iter25_to_t1_iter26__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter25_to_t1_iter26__din),
    .if_full_n(from_t1_iter25_to_t1_iter26__full_n),
    .if_write(from_t1_iter25_to_t1_iter26__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(134)
  )
  from_t1_iter26_to_t1_iter27
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter26_to_t1_iter27__dout),
    .if_empty_n(from_t1_iter26_to_t1_iter27__empty_n),
    .if_read(from_t1_iter26_to_t1_iter27__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter26_to_t1_iter27__din),
    .if_full_n(from_t1_iter26_to_t1_iter27__full_n),
    .if_write(from_t1_iter26_to_t1_iter27__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter27_to_t1_iter28
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter27_to_t1_iter28__dout),
    .if_empty_n(from_t1_iter27_to_t1_iter28__empty_n),
    .if_read(from_t1_iter27_to_t1_iter28__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter27_to_t1_iter28__din),
    .if_full_n(from_t1_iter27_to_t1_iter28__full_n),
    .if_write(from_t1_iter27_to_t1_iter28__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter28_to_t1_iter29
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter28_to_t1_iter29__dout),
    .if_empty_n(from_t1_iter28_to_t1_iter29__empty_n),
    .if_read(from_t1_iter28_to_t1_iter29__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter28_to_t1_iter29__din),
    .if_full_n(from_t1_iter28_to_t1_iter29__full_n),
    .if_write(from_t1_iter28_to_t1_iter29__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(130)
  )
  from_t1_iter29_to_t1_iter30
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter29_to_t1_iter30__dout),
    .if_empty_n(from_t1_iter29_to_t1_iter30__empty_n),
    .if_read(from_t1_iter29_to_t1_iter30__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter29_to_t1_iter30__din),
    .if_full_n(from_t1_iter29_to_t1_iter30__full_n),
    .if_write(from_t1_iter29_to_t1_iter30__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter2_to_t1_iter3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter2_to_t1_iter3__dout),
    .if_empty_n(from_t1_iter2_to_t1_iter3__empty_n),
    .if_read(from_t1_iter2_to_t1_iter3__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter2_to_t1_iter3__din),
    .if_full_n(from_t1_iter2_to_t1_iter3__full_n),
    .if_write(from_t1_iter2_to_t1_iter3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(130)
  )
  from_t1_iter30_to_t1_iter31
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter30_to_t1_iter31__dout),
    .if_empty_n(from_t1_iter30_to_t1_iter31__empty_n),
    .if_read(from_t1_iter30_to_t1_iter31__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter30_to_t1_iter31__din),
    .if_full_n(from_t1_iter30_to_t1_iter31__full_n),
    .if_write(from_t1_iter30_to_t1_iter31__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(130)
  )
  from_t1_iter31_to_t1_iter32
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter31_to_t1_iter32__dout),
    .if_empty_n(from_t1_iter31_to_t1_iter32__empty_n),
    .if_read(from_t1_iter31_to_t1_iter32__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter31_to_t1_iter32__din),
    .if_full_n(from_t1_iter31_to_t1_iter32__full_n),
    .if_write(from_t1_iter31_to_t1_iter32__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(130)
  )
  from_t1_iter32_to_t1_iter33
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter32_to_t1_iter33__dout),
    .if_empty_n(from_t1_iter32_to_t1_iter33__empty_n),
    .if_read(from_t1_iter32_to_t1_iter33__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter32_to_t1_iter33__din),
    .if_full_n(from_t1_iter32_to_t1_iter33__full_n),
    .if_write(from_t1_iter32_to_t1_iter33__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(130)
  )
  from_t1_iter33_to_t1_iter34
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter33_to_t1_iter34__dout),
    .if_empty_n(from_t1_iter33_to_t1_iter34__empty_n),
    .if_read(from_t1_iter33_to_t1_iter34__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter33_to_t1_iter34__din),
    .if_full_n(from_t1_iter33_to_t1_iter34__full_n),
    .if_write(from_t1_iter33_to_t1_iter34__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(130)
  )
  from_t1_iter34_to_t1_iter35
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter34_to_t1_iter35__dout),
    .if_empty_n(from_t1_iter34_to_t1_iter35__empty_n),
    .if_read(from_t1_iter34_to_t1_iter35__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter34_to_t1_iter35__din),
    .if_full_n(from_t1_iter34_to_t1_iter35__full_n),
    .if_write(from_t1_iter34_to_t1_iter35__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(130)
  )
  from_t1_iter35_to_t1_iter36
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter35_to_t1_iter36__dout),
    .if_empty_n(from_t1_iter35_to_t1_iter36__empty_n),
    .if_read(from_t1_iter35_to_t1_iter36__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter35_to_t1_iter36__din),
    .if_full_n(from_t1_iter35_to_t1_iter36__full_n),
    .if_write(from_t1_iter35_to_t1_iter36__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(130)
  )
  from_t1_iter36_to_t1_iter37
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter36_to_t1_iter37__dout),
    .if_empty_n(from_t1_iter36_to_t1_iter37__empty_n),
    .if_read(from_t1_iter36_to_t1_iter37__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter36_to_t1_iter37__din),
    .if_full_n(from_t1_iter36_to_t1_iter37__full_n),
    .if_write(from_t1_iter36_to_t1_iter37__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(130)
  )
  from_t1_iter37_to_t1_iter38
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter37_to_t1_iter38__dout),
    .if_empty_n(from_t1_iter37_to_t1_iter38__empty_n),
    .if_read(from_t1_iter37_to_t1_iter38__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter37_to_t1_iter38__din),
    .if_full_n(from_t1_iter37_to_t1_iter38__full_n),
    .if_write(from_t1_iter37_to_t1_iter38__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(130)
  )
  from_t1_iter38_to_t1_iter39
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter38_to_t1_iter39__dout),
    .if_empty_n(from_t1_iter38_to_t1_iter39__empty_n),
    .if_read(from_t1_iter38_to_t1_iter39__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter38_to_t1_iter39__din),
    .if_full_n(from_t1_iter38_to_t1_iter39__full_n),
    .if_write(from_t1_iter38_to_t1_iter39__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(130)
  )
  from_t1_iter39_to_t1_iter40
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter39_to_t1_iter40__dout),
    .if_empty_n(from_t1_iter39_to_t1_iter40__empty_n),
    .if_read(from_t1_iter39_to_t1_iter40__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter39_to_t1_iter40__din),
    .if_full_n(from_t1_iter39_to_t1_iter40__full_n),
    .if_write(from_t1_iter39_to_t1_iter40__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(130)
  )
  from_t1_iter3_to_t1_iter4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter3_to_t1_iter4__dout),
    .if_empty_n(from_t1_iter3_to_t1_iter4__empty_n),
    .if_read(from_t1_iter3_to_t1_iter4__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter3_to_t1_iter4__din),
    .if_full_n(from_t1_iter3_to_t1_iter4__full_n),
    .if_write(from_t1_iter3_to_t1_iter4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(130)
  )
  from_t1_iter40_to_t1_iter41
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter40_to_t1_iter41__dout),
    .if_empty_n(from_t1_iter40_to_t1_iter41__empty_n),
    .if_read(from_t1_iter40_to_t1_iter41__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter40_to_t1_iter41__din),
    .if_full_n(from_t1_iter40_to_t1_iter41__full_n),
    .if_write(from_t1_iter40_to_t1_iter41__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(132)
  )
  from_t1_iter41_to_t1_iter42
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter41_to_t1_iter42__dout),
    .if_empty_n(from_t1_iter41_to_t1_iter42__empty_n),
    .if_read(from_t1_iter41_to_t1_iter42__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter41_to_t1_iter42__din),
    .if_full_n(from_t1_iter41_to_t1_iter42__full_n),
    .if_write(from_t1_iter41_to_t1_iter42__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter42_to_t1_iter43
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter42_to_t1_iter43__dout),
    .if_empty_n(from_t1_iter42_to_t1_iter43__empty_n),
    .if_read(from_t1_iter42_to_t1_iter43__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter42_to_t1_iter43__din),
    .if_full_n(from_t1_iter42_to_t1_iter43__full_n),
    .if_write(from_t1_iter42_to_t1_iter43__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(134)
  )
  from_t1_iter43_to_t1_iter44
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter43_to_t1_iter44__dout),
    .if_empty_n(from_t1_iter43_to_t1_iter44__empty_n),
    .if_read(from_t1_iter43_to_t1_iter44__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter43_to_t1_iter44__din),
    .if_full_n(from_t1_iter43_to_t1_iter44__full_n),
    .if_write(from_t1_iter43_to_t1_iter44__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter44_to_t1_iter45
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter44_to_t1_iter45__dout),
    .if_empty_n(from_t1_iter44_to_t1_iter45__empty_n),
    .if_read(from_t1_iter44_to_t1_iter45__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter44_to_t1_iter45__din),
    .if_full_n(from_t1_iter44_to_t1_iter45__full_n),
    .if_write(from_t1_iter44_to_t1_iter45__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter45_to_t1_iter46
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter45_to_t1_iter46__dout),
    .if_empty_n(from_t1_iter45_to_t1_iter46__empty_n),
    .if_read(from_t1_iter45_to_t1_iter46__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter45_to_t1_iter46__din),
    .if_full_n(from_t1_iter45_to_t1_iter46__full_n),
    .if_write(from_t1_iter45_to_t1_iter46__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(130)
  )
  from_t1_iter46_to_t1_iter47
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter46_to_t1_iter47__dout),
    .if_empty_n(from_t1_iter46_to_t1_iter47__empty_n),
    .if_read(from_t1_iter46_to_t1_iter47__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter46_to_t1_iter47__din),
    .if_full_n(from_t1_iter46_to_t1_iter47__full_n),
    .if_write(from_t1_iter46_to_t1_iter47__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(132)
  )
  from_t1_iter47_to_t1_iter48
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter47_to_t1_iter48__dout),
    .if_empty_n(from_t1_iter47_to_t1_iter48__empty_n),
    .if_read(from_t1_iter47_to_t1_iter48__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter47_to_t1_iter48__din),
    .if_full_n(from_t1_iter47_to_t1_iter48__full_n),
    .if_write(from_t1_iter47_to_t1_iter48__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter48_to_t1_iter49
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter48_to_t1_iter49__dout),
    .if_empty_n(from_t1_iter48_to_t1_iter49__empty_n),
    .if_read(from_t1_iter48_to_t1_iter49__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter48_to_t1_iter49__din),
    .if_full_n(from_t1_iter48_to_t1_iter49__full_n),
    .if_write(from_t1_iter48_to_t1_iter49__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(130)
  )
  from_t1_iter49_to_t1_iter50
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter49_to_t1_iter50__dout),
    .if_empty_n(from_t1_iter49_to_t1_iter50__empty_n),
    .if_read(from_t1_iter49_to_t1_iter50__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter49_to_t1_iter50__din),
    .if_full_n(from_t1_iter49_to_t1_iter50__full_n),
    .if_write(from_t1_iter49_to_t1_iter50__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(130)
  )
  from_t1_iter4_to_t1_iter5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter4_to_t1_iter5__dout),
    .if_empty_n(from_t1_iter4_to_t1_iter5__empty_n),
    .if_read(from_t1_iter4_to_t1_iter5__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter4_to_t1_iter5__din),
    .if_full_n(from_t1_iter4_to_t1_iter5__full_n),
    .if_write(from_t1_iter4_to_t1_iter5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(134)
  )
  from_t1_iter50_to_t1_iter51
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter50_to_t1_iter51__dout),
    .if_empty_n(from_t1_iter50_to_t1_iter51__empty_n),
    .if_read(from_t1_iter50_to_t1_iter51__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter50_to_t1_iter51__din),
    .if_full_n(from_t1_iter50_to_t1_iter51__full_n),
    .if_write(from_t1_iter50_to_t1_iter51__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter51_to_t1_iter52
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter51_to_t1_iter52__dout),
    .if_empty_n(from_t1_iter51_to_t1_iter52__empty_n),
    .if_read(from_t1_iter51_to_t1_iter52__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter51_to_t1_iter52__din),
    .if_full_n(from_t1_iter51_to_t1_iter52__full_n),
    .if_write(from_t1_iter51_to_t1_iter52__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter52_to_t1_iter53
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter52_to_t1_iter53__dout),
    .if_empty_n(from_t1_iter52_to_t1_iter53__empty_n),
    .if_read(from_t1_iter52_to_t1_iter53__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter52_to_t1_iter53__din),
    .if_full_n(from_t1_iter52_to_t1_iter53__full_n),
    .if_write(from_t1_iter52_to_t1_iter53__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(130)
  )
  from_t1_iter53_to_t1_iter54
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter53_to_t1_iter54__dout),
    .if_empty_n(from_t1_iter53_to_t1_iter54__empty_n),
    .if_read(from_t1_iter53_to_t1_iter54__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter53_to_t1_iter54__din),
    .if_full_n(from_t1_iter53_to_t1_iter54__full_n),
    .if_write(from_t1_iter53_to_t1_iter54__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(130)
  )
  from_t1_iter54_to_t1_iter55
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter54_to_t1_iter55__dout),
    .if_empty_n(from_t1_iter54_to_t1_iter55__empty_n),
    .if_read(from_t1_iter54_to_t1_iter55__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter54_to_t1_iter55__din),
    .if_full_n(from_t1_iter54_to_t1_iter55__full_n),
    .if_write(from_t1_iter54_to_t1_iter55__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(130)
  )
  from_t1_iter55_to_t1_iter56
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter55_to_t1_iter56__dout),
    .if_empty_n(from_t1_iter55_to_t1_iter56__empty_n),
    .if_read(from_t1_iter55_to_t1_iter56__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter55_to_t1_iter56__din),
    .if_full_n(from_t1_iter55_to_t1_iter56__full_n),
    .if_write(from_t1_iter55_to_t1_iter56__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(130)
  )
  from_t1_iter56_to_t1_iter57
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter56_to_t1_iter57__dout),
    .if_empty_n(from_t1_iter56_to_t1_iter57__empty_n),
    .if_read(from_t1_iter56_to_t1_iter57__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter56_to_t1_iter57__din),
    .if_full_n(from_t1_iter56_to_t1_iter57__full_n),
    .if_write(from_t1_iter56_to_t1_iter57__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(130)
  )
  from_t1_iter57_to_t1_iter58
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter57_to_t1_iter58__dout),
    .if_empty_n(from_t1_iter57_to_t1_iter58__empty_n),
    .if_read(from_t1_iter57_to_t1_iter58__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter57_to_t1_iter58__din),
    .if_full_n(from_t1_iter57_to_t1_iter58__full_n),
    .if_write(from_t1_iter57_to_t1_iter58__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(130)
  )
  from_t1_iter58_to_t1_iter59
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter58_to_t1_iter59__dout),
    .if_empty_n(from_t1_iter58_to_t1_iter59__empty_n),
    .if_read(from_t1_iter58_to_t1_iter59__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter58_to_t1_iter59__din),
    .if_full_n(from_t1_iter58_to_t1_iter59__full_n),
    .if_write(from_t1_iter58_to_t1_iter59__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(130)
  )
  from_t1_iter59_to_t1_iter60
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter59_to_t1_iter60__dout),
    .if_empty_n(from_t1_iter59_to_t1_iter60__empty_n),
    .if_read(from_t1_iter59_to_t1_iter60__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter59_to_t1_iter60__din),
    .if_full_n(from_t1_iter59_to_t1_iter60__full_n),
    .if_write(from_t1_iter59_to_t1_iter60__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(130)
  )
  from_t1_iter5_to_t1_iter6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter5_to_t1_iter6__dout),
    .if_empty_n(from_t1_iter5_to_t1_iter6__empty_n),
    .if_read(from_t1_iter5_to_t1_iter6__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter5_to_t1_iter6__din),
    .if_full_n(from_t1_iter5_to_t1_iter6__full_n),
    .if_write(from_t1_iter5_to_t1_iter6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(130)
  )
  from_t1_iter60_to_t1_iter61
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter60_to_t1_iter61__dout),
    .if_empty_n(from_t1_iter60_to_t1_iter61__empty_n),
    .if_read(from_t1_iter60_to_t1_iter61__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter60_to_t1_iter61__din),
    .if_full_n(from_t1_iter60_to_t1_iter61__full_n),
    .if_write(from_t1_iter60_to_t1_iter61__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(136)
  )
  from_t1_iter61_to_t1_iter62
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter61_to_t1_iter62__dout),
    .if_empty_n(from_t1_iter61_to_t1_iter62__empty_n),
    .if_read(from_t1_iter61_to_t1_iter62__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter61_to_t1_iter62__din),
    .if_full_n(from_t1_iter61_to_t1_iter62__full_n),
    .if_write(from_t1_iter61_to_t1_iter62__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter62_to_t1_iter63
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter62_to_t1_iter63__dout),
    .if_empty_n(from_t1_iter62_to_t1_iter63__empty_n),
    .if_read(from_t1_iter62_to_t1_iter63__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter62_to_t1_iter63__din),
    .if_full_n(from_t1_iter62_to_t1_iter63__full_n),
    .if_write(from_t1_iter62_to_t1_iter63__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter63_to_t1_iter64
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter63_to_t1_iter64__dout),
    .if_empty_n(from_t1_iter63_to_t1_iter64__empty_n),
    .if_read(from_t1_iter63_to_t1_iter64__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter63_to_t1_iter64__din),
    .if_full_n(from_t1_iter63_to_t1_iter64__full_n),
    .if_write(from_t1_iter63_to_t1_iter64__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter64_to_t1_iter65
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter64_to_t1_iter65__dout),
    .if_empty_n(from_t1_iter64_to_t1_iter65__empty_n),
    .if_read(from_t1_iter64_to_t1_iter65__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter64_to_t1_iter65__din),
    .if_full_n(from_t1_iter64_to_t1_iter65__full_n),
    .if_write(from_t1_iter64_to_t1_iter65__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(130)
  )
  from_t1_iter65_to_t1_iter66
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter65_to_t1_iter66__dout),
    .if_empty_n(from_t1_iter65_to_t1_iter66__empty_n),
    .if_read(from_t1_iter65_to_t1_iter66__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter65_to_t1_iter66__din),
    .if_full_n(from_t1_iter65_to_t1_iter66__full_n),
    .if_write(from_t1_iter65_to_t1_iter66__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(130)
  )
  from_t1_iter66_to_t1_iter67
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter66_to_t1_iter67__dout),
    .if_empty_n(from_t1_iter66_to_t1_iter67__empty_n),
    .if_read(from_t1_iter66_to_t1_iter67__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter66_to_t1_iter67__din),
    .if_full_n(from_t1_iter66_to_t1_iter67__full_n),
    .if_write(from_t1_iter66_to_t1_iter67__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(130)
  )
  from_t1_iter67_to_t1_iter68
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter67_to_t1_iter68__dout),
    .if_empty_n(from_t1_iter67_to_t1_iter68__empty_n),
    .if_read(from_t1_iter67_to_t1_iter68__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter67_to_t1_iter68__din),
    .if_full_n(from_t1_iter67_to_t1_iter68__full_n),
    .if_write(from_t1_iter67_to_t1_iter68__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(130)
  )
  from_t1_iter68_to_t1_iter69
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter68_to_t1_iter69__dout),
    .if_empty_n(from_t1_iter68_to_t1_iter69__empty_n),
    .if_read(from_t1_iter68_to_t1_iter69__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter68_to_t1_iter69__din),
    .if_full_n(from_t1_iter68_to_t1_iter69__full_n),
    .if_write(from_t1_iter68_to_t1_iter69__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(134)
  )
  from_t1_iter69_to_t1_iter70
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter69_to_t1_iter70__dout),
    .if_empty_n(from_t1_iter69_to_t1_iter70__empty_n),
    .if_read(from_t1_iter69_to_t1_iter70__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter69_to_t1_iter70__din),
    .if_full_n(from_t1_iter69_to_t1_iter70__full_n),
    .if_write(from_t1_iter69_to_t1_iter70__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(134)
  )
  from_t1_iter6_to_t1_iter7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter6_to_t1_iter7__dout),
    .if_empty_n(from_t1_iter6_to_t1_iter7__empty_n),
    .if_read(from_t1_iter6_to_t1_iter7__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter6_to_t1_iter7__din),
    .if_full_n(from_t1_iter6_to_t1_iter7__full_n),
    .if_write(from_t1_iter6_to_t1_iter7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter70_to_t1_iter71
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter70_to_t1_iter71__dout),
    .if_empty_n(from_t1_iter70_to_t1_iter71__empty_n),
    .if_read(from_t1_iter70_to_t1_iter71__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter70_to_t1_iter71__din),
    .if_full_n(from_t1_iter70_to_t1_iter71__full_n),
    .if_write(from_t1_iter70_to_t1_iter71__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter71_to_t1_iter72
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter71_to_t1_iter72__dout),
    .if_empty_n(from_t1_iter71_to_t1_iter72__empty_n),
    .if_read(from_t1_iter71_to_t1_iter72__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter71_to_t1_iter72__din),
    .if_full_n(from_t1_iter71_to_t1_iter72__full_n),
    .if_write(from_t1_iter71_to_t1_iter72__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(132)
  )
  from_t1_iter72_to_t1_iter73
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter72_to_t1_iter73__dout),
    .if_empty_n(from_t1_iter72_to_t1_iter73__empty_n),
    .if_read(from_t1_iter72_to_t1_iter73__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter72_to_t1_iter73__din),
    .if_full_n(from_t1_iter72_to_t1_iter73__full_n),
    .if_write(from_t1_iter72_to_t1_iter73__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter73_to_t1_iter74
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter73_to_t1_iter74__dout),
    .if_empty_n(from_t1_iter73_to_t1_iter74__empty_n),
    .if_read(from_t1_iter73_to_t1_iter74__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter73_to_t1_iter74__din),
    .if_full_n(from_t1_iter73_to_t1_iter74__full_n),
    .if_write(from_t1_iter73_to_t1_iter74__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(134)
  )
  from_t1_iter74_to_t1_iter75
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter74_to_t1_iter75__dout),
    .if_empty_n(from_t1_iter74_to_t1_iter75__empty_n),
    .if_read(from_t1_iter74_to_t1_iter75__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter74_to_t1_iter75__din),
    .if_full_n(from_t1_iter74_to_t1_iter75__full_n),
    .if_write(from_t1_iter74_to_t1_iter75__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter75_to_t1_iter76
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter75_to_t1_iter76__dout),
    .if_empty_n(from_t1_iter75_to_t1_iter76__empty_n),
    .if_read(from_t1_iter75_to_t1_iter76__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter75_to_t1_iter76__din),
    .if_full_n(from_t1_iter75_to_t1_iter76__full_n),
    .if_write(from_t1_iter75_to_t1_iter76__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(132)
  )
  from_t1_iter76_to_t1_iter77
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter76_to_t1_iter77__dout),
    .if_empty_n(from_t1_iter76_to_t1_iter77__empty_n),
    .if_read(from_t1_iter76_to_t1_iter77__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter76_to_t1_iter77__din),
    .if_full_n(from_t1_iter76_to_t1_iter77__full_n),
    .if_write(from_t1_iter76_to_t1_iter77__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter77_to_t1_iter78
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter77_to_t1_iter78__dout),
    .if_empty_n(from_t1_iter77_to_t1_iter78__empty_n),
    .if_read(from_t1_iter77_to_t1_iter78__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter77_to_t1_iter78__din),
    .if_full_n(from_t1_iter77_to_t1_iter78__full_n),
    .if_write(from_t1_iter77_to_t1_iter78__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter78_to_t1_iter79
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter78_to_t1_iter79__dout),
    .if_empty_n(from_t1_iter78_to_t1_iter79__empty_n),
    .if_read(from_t1_iter78_to_t1_iter79__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter78_to_t1_iter79__din),
    .if_full_n(from_t1_iter78_to_t1_iter79__full_n),
    .if_write(from_t1_iter78_to_t1_iter79__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(130)
  )
  from_t1_iter79_to_t1_iter80
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter79_to_t1_iter80__dout),
    .if_empty_n(from_t1_iter79_to_t1_iter80__empty_n),
    .if_read(from_t1_iter79_to_t1_iter80__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter79_to_t1_iter80__din),
    .if_full_n(from_t1_iter79_to_t1_iter80__full_n),
    .if_write(from_t1_iter79_to_t1_iter80__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter7_to_t1_iter8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter7_to_t1_iter8__dout),
    .if_empty_n(from_t1_iter7_to_t1_iter8__empty_n),
    .if_read(from_t1_iter7_to_t1_iter8__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter7_to_t1_iter8__din),
    .if_full_n(from_t1_iter7_to_t1_iter8__full_n),
    .if_write(from_t1_iter7_to_t1_iter8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(132)
  )
  from_t1_iter80_to_t1_iter81
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter80_to_t1_iter81__dout),
    .if_empty_n(from_t1_iter80_to_t1_iter81__empty_n),
    .if_read(from_t1_iter80_to_t1_iter81__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter80_to_t1_iter81__din),
    .if_full_n(from_t1_iter80_to_t1_iter81__full_n),
    .if_write(from_t1_iter80_to_t1_iter81__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter81_to_t1_iter82
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter81_to_t1_iter82__dout),
    .if_empty_n(from_t1_iter81_to_t1_iter82__empty_n),
    .if_read(from_t1_iter81_to_t1_iter82__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter81_to_t1_iter82__din),
    .if_full_n(from_t1_iter81_to_t1_iter82__full_n),
    .if_write(from_t1_iter81_to_t1_iter82__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(130)
  )
  from_t1_iter82_to_t1_iter83
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter82_to_t1_iter83__dout),
    .if_empty_n(from_t1_iter82_to_t1_iter83__empty_n),
    .if_read(from_t1_iter82_to_t1_iter83__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter82_to_t1_iter83__din),
    .if_full_n(from_t1_iter82_to_t1_iter83__full_n),
    .if_write(from_t1_iter82_to_t1_iter83__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(130)
  )
  from_t1_iter83_to_t1_iter84
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter83_to_t1_iter84__dout),
    .if_empty_n(from_t1_iter83_to_t1_iter84__empty_n),
    .if_read(from_t1_iter83_to_t1_iter84__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter83_to_t1_iter84__din),
    .if_full_n(from_t1_iter83_to_t1_iter84__full_n),
    .if_write(from_t1_iter83_to_t1_iter84__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(136)
  )
  from_t1_iter84_to_t1_iter85
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter84_to_t1_iter85__dout),
    .if_empty_n(from_t1_iter84_to_t1_iter85__empty_n),
    .if_read(from_t1_iter84_to_t1_iter85__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter84_to_t1_iter85__din),
    .if_full_n(from_t1_iter84_to_t1_iter85__full_n),
    .if_write(from_t1_iter84_to_t1_iter85__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter85_to_t1_iter86
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter85_to_t1_iter86__dout),
    .if_empty_n(from_t1_iter85_to_t1_iter86__empty_n),
    .if_read(from_t1_iter85_to_t1_iter86__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter85_to_t1_iter86__din),
    .if_full_n(from_t1_iter85_to_t1_iter86__full_n),
    .if_write(from_t1_iter85_to_t1_iter86__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(136)
  )
  from_t1_iter86_to_t1_iter87
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter86_to_t1_iter87__dout),
    .if_empty_n(from_t1_iter86_to_t1_iter87__empty_n),
    .if_read(from_t1_iter86_to_t1_iter87__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter86_to_t1_iter87__din),
    .if_full_n(from_t1_iter86_to_t1_iter87__full_n),
    .if_write(from_t1_iter86_to_t1_iter87__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter87_to_t1_iter88
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter87_to_t1_iter88__dout),
    .if_empty_n(from_t1_iter87_to_t1_iter88__empty_n),
    .if_read(from_t1_iter87_to_t1_iter88__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter87_to_t1_iter88__din),
    .if_full_n(from_t1_iter87_to_t1_iter88__full_n),
    .if_write(from_t1_iter87_to_t1_iter88__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter88_to_t1_iter89
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter88_to_t1_iter89__dout),
    .if_empty_n(from_t1_iter88_to_t1_iter89__empty_n),
    .if_read(from_t1_iter88_to_t1_iter89__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter88_to_t1_iter89__din),
    .if_full_n(from_t1_iter88_to_t1_iter89__full_n),
    .if_write(from_t1_iter88_to_t1_iter89__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(134)
  )
  from_t1_iter89_to_t1_iter90
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter89_to_t1_iter90__dout),
    .if_empty_n(from_t1_iter89_to_t1_iter90__empty_n),
    .if_read(from_t1_iter89_to_t1_iter90__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter89_to_t1_iter90__din),
    .if_full_n(from_t1_iter89_to_t1_iter90__full_n),
    .if_write(from_t1_iter89_to_t1_iter90__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter8_to_t1_iter9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter8_to_t1_iter9__dout),
    .if_empty_n(from_t1_iter8_to_t1_iter9__empty_n),
    .if_read(from_t1_iter8_to_t1_iter9__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter8_to_t1_iter9__din),
    .if_full_n(from_t1_iter8_to_t1_iter9__full_n),
    .if_write(from_t1_iter8_to_t1_iter9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(130)
  )
  from_t1_iter90_to_t1_iter91
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter90_to_t1_iter91__dout),
    .if_empty_n(from_t1_iter90_to_t1_iter91__empty_n),
    .if_read(from_t1_iter90_to_t1_iter91__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter90_to_t1_iter91__din),
    .if_full_n(from_t1_iter90_to_t1_iter91__full_n),
    .if_write(from_t1_iter90_to_t1_iter91__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter91_to_t1_iter92
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter91_to_t1_iter92__dout),
    .if_empty_n(from_t1_iter91_to_t1_iter92__empty_n),
    .if_read(from_t1_iter91_to_t1_iter92__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter91_to_t1_iter92__din),
    .if_full_n(from_t1_iter91_to_t1_iter92__full_n),
    .if_write(from_t1_iter91_to_t1_iter92__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter92_to_t1_iter93
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter92_to_t1_iter93__dout),
    .if_empty_n(from_t1_iter92_to_t1_iter93__empty_n),
    .if_read(from_t1_iter92_to_t1_iter93__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter92_to_t1_iter93__din),
    .if_full_n(from_t1_iter92_to_t1_iter93__full_n),
    .if_write(from_t1_iter92_to_t1_iter93__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter93_to_t1_iter94
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter93_to_t1_iter94__dout),
    .if_empty_n(from_t1_iter93_to_t1_iter94__empty_n),
    .if_read(from_t1_iter93_to_t1_iter94__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter93_to_t1_iter94__din),
    .if_full_n(from_t1_iter93_to_t1_iter94__full_n),
    .if_write(from_t1_iter93_to_t1_iter94__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter94_to_t1_iter95
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter94_to_t1_iter95__dout),
    .if_empty_n(from_t1_iter94_to_t1_iter95__empty_n),
    .if_read(from_t1_iter94_to_t1_iter95__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter94_to_t1_iter95__din),
    .if_full_n(from_t1_iter94_to_t1_iter95__full_n),
    .if_write(from_t1_iter94_to_t1_iter95__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(136)
  )
  from_t1_iter95_to_t1_iter96
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter95_to_t1_iter96__dout),
    .if_empty_n(from_t1_iter95_to_t1_iter96__empty_n),
    .if_read(from_t1_iter95_to_t1_iter96__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter95_to_t1_iter96__din),
    .if_full_n(from_t1_iter95_to_t1_iter96__full_n),
    .if_write(from_t1_iter95_to_t1_iter96__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter96_to_t1_iter97
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter96_to_t1_iter97__dout),
    .if_empty_n(from_t1_iter96_to_t1_iter97__empty_n),
    .if_read(from_t1_iter96_to_t1_iter97__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter96_to_t1_iter97__din),
    .if_full_n(from_t1_iter96_to_t1_iter97__full_n),
    .if_write(from_t1_iter96_to_t1_iter97__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter97_to_t1_iter98
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter97_to_t1_iter98__dout),
    .if_empty_n(from_t1_iter97_to_t1_iter98__empty_n),
    .if_read(from_t1_iter97_to_t1_iter98__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter97_to_t1_iter98__din),
    .if_full_n(from_t1_iter97_to_t1_iter98__full_n),
    .if_write(from_t1_iter97_to_t1_iter98__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(132)
  )
  from_t1_iter98_to_t1_iter99
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter98_to_t1_iter99__dout),
    .if_empty_n(from_t1_iter98_to_t1_iter99__empty_n),
    .if_read(from_t1_iter98_to_t1_iter99__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter98_to_t1_iter99__din),
    .if_full_n(from_t1_iter98_to_t1_iter99__full_n),
    .if_write(from_t1_iter98_to_t1_iter99__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(7),
    .DEPTH(128)
  )
  from_t1_iter99_to_t1_iter100
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter99_to_t1_iter100__dout),
    .if_empty_n(from_t1_iter99_to_t1_iter100__empty_n),
    .if_read(from_t1_iter99_to_t1_iter100__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter99_to_t1_iter100__din),
    .if_full_n(from_t1_iter99_to_t1_iter100__full_n),
    .if_write(from_t1_iter99_to_t1_iter100__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(8),
    .DEPTH(130)
  )
  from_t1_iter9_to_t1_iter10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(from_t1_iter9_to_t1_iter10__dout),
    .if_empty_n(from_t1_iter9_to_t1_iter10__empty_n),
    .if_read(from_t1_iter9_to_t1_iter10__read),
    .if_read_ce(1'b1),
    .if_din(from_t1_iter9_to_t1_iter10__din),
    .if_full_n(from_t1_iter9_to_t1_iter10__full_n),
    .if_write(from_t1_iter9_to_t1_iter10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) BurstRead_floatx16
  BurstRead_floatx16_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(BurstRead_floatx16_0__ap_start),
    .ap_done(BurstRead_floatx16_0__ap_done),
    .ap_idle(BurstRead_floatx16_0__ap_idle),
    .ap_ready(BurstRead_floatx16_0__ap_ready),
    .src_read_addr_s_din(bank_0_t1_read_addr__din),
    .src_read_addr_s_full_n(bank_0_t1_read_addr__full_n),
    .src_read_addr_s_write(bank_0_t1_read_addr__write),
    .src_read_addr_offset(BurstRead_floatx16_0___bank_0_t1__q0),
    .src_read_data_s_dout({1'b0, bank_0_t1_read_data__dout}),
    .src_read_data_peek_dout({1'b0, bank_0_t1_read_data__dout}),
    .src_read_data_s_empty_n(bank_0_t1_read_data__empty_n),
    .src_read_data_peek_empty_n(bank_0_t1_read_data__empty_n),
    .src_read_data_s_read(bank_0_t1_read_data__read),
    .src_read_data_peek_read(),
    .src_write_addr_s_din(bank_0_t1_write_addr__din),
    .src_write_addr_s_full_n(bank_0_t1_write_addr__full_n),
    .src_write_addr_s_write(bank_0_t1_write_addr__write),
    .src_write_addr_offset(BurstRead_floatx16_0___bank_0_t1__q0),
    .src_write_data_din(bank_0_t1_write_data__din),
    .src_write_data_full_n(bank_0_t1_write_data__full_n),
    .src_write_data_write(bank_0_t1_write_data__write),
    .src_write_resp_s_dout({1'b0, bank_0_t1_write_resp__dout}),
    .src_write_resp_peek_dout({1'b0, bank_0_t1_write_resp__dout}),
    .src_write_resp_s_empty_n(bank_0_t1_write_resp__empty_n),
    .src_write_resp_peek_empty_n(bank_0_t1_write_resp__empty_n),
    .src_write_resp_s_read(bank_0_t1_write_resp__read),
    .src_write_resp_peek_read(),
    .dest_din(bank_0_t1_buf__din),
    .dest_full_n(bank_0_t1_buf__full_n),
    .dest_write(bank_0_t1_buf__write),
    .n(BurstRead_floatx16_0___coalesced_data_num__q0)
  );


  (* keep_hierarchy = "yes" *) BurstWrite_floatx16
  BurstWrite_floatx16_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(BurstWrite_floatx16_0__ap_start),
    .ap_done(BurstWrite_floatx16_0__ap_done),
    .ap_idle(BurstWrite_floatx16_0__ap_idle),
    .ap_ready(BurstWrite_floatx16_0__ap_ready),
    .dest_read_addr_s_din(bank_1_t0_read_addr__din),
    .dest_read_addr_s_full_n(bank_1_t0_read_addr__full_n),
    .dest_read_addr_s_write(bank_1_t0_read_addr__write),
    .dest_read_addr_offset(BurstWrite_floatx16_0___bank_1_t0__q0),
    .dest_read_data_s_dout({1'b0, bank_1_t0_read_data__dout}),
    .dest_read_data_peek_dout({1'b0, bank_1_t0_read_data__dout}),
    .dest_read_data_s_empty_n(bank_1_t0_read_data__empty_n),
    .dest_read_data_peek_empty_n(bank_1_t0_read_data__empty_n),
    .dest_read_data_s_read(bank_1_t0_read_data__read),
    .dest_read_data_peek_read(),
    .dest_write_addr_s_din(bank_1_t0_write_addr__din),
    .dest_write_addr_s_full_n(bank_1_t0_write_addr__full_n),
    .dest_write_addr_s_write(bank_1_t0_write_addr__write),
    .dest_write_addr_offset(BurstWrite_floatx16_0___bank_1_t0__q0),
    .dest_write_data_din(bank_1_t0_write_data__din),
    .dest_write_data_full_n(bank_1_t0_write_data__full_n),
    .dest_write_data_write(bank_1_t0_write_data__write),
    .dest_write_resp_s_dout({1'b0, bank_1_t0_write_resp__dout}),
    .dest_write_resp_peek_dout({1'b0, bank_1_t0_write_resp__dout}),
    .dest_write_resp_s_empty_n(bank_1_t0_write_resp__empty_n),
    .dest_write_resp_peek_empty_n(bank_1_t0_write_resp__empty_n),
    .dest_write_resp_s_read(bank_1_t0_write_resp__read),
    .dest_write_resp_peek_read(),
    .src_s_dout(bank_1_t0_buf__dout),
    .src_peek_dout(bank_1_t0_buf__dout),
    .src_s_empty_n(bank_1_t0_buf__empty_n),
    .src_peek_empty_n(bank_1_t0_buf__empty_n),
    .src_s_read(bank_1_t0_buf__read),
    .src_peek_read(),
    .n(BurstWrite_floatx16_0___coalesced_data_num__q0)
  );


  (* keep_hierarchy = "yes" *) Module0Func
  Module0Func_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module0Func_0__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .dram_t1_bank_0_fifo_s_dout(bank_0_t1_buf__dout),
    .dram_t1_bank_0_fifo_peek_dout(bank_0_t1_buf__dout),
    .dram_t1_bank_0_fifo_s_empty_n(bank_0_t1_buf__empty_n),
    .dram_t1_bank_0_fifo_peek_empty_n(bank_0_t1_buf__empty_n),
    .dram_t1_bank_0_fifo_s_read(bank_0_t1_buf__read),
    .dram_t1_bank_0_fifo_peek_read(),
    .fifo_st_0_din(from_t1_bank_0_to_t1_iter1__din),
    .fifo_st_0_full_n(from_t1_bank_0_to_t1_iter1__full_n),
    .fifo_st_0_write(from_t1_bank_0_to_t1_iter1__write)
  );


  (* keep_hierarchy = "yes" *) Module1Func
  Module1Func_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module1Func_0__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_bank_0_to_t1_iter1__dout),
    .fifo_ld_0_peek_dout(from_t1_bank_0_to_t1_iter1__dout),
    .fifo_ld_0_s_empty_n(from_t1_bank_0_to_t1_iter1__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_bank_0_to_t1_iter1__empty_n),
    .fifo_ld_0_s_read(from_t1_bank_0_to_t1_iter1__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter1_to_t1_iter2__din),
    .fifo_st_0_full_n(from_t1_iter1_to_t1_iter2__full_n),
    .fifo_st_0_write(from_t1_iter1_to_t1_iter2__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_0__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter1_to_t1_iter2__dout),
    .fifo_ld_0_peek_dout(from_t1_iter1_to_t1_iter2__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter1_to_t1_iter2__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter1_to_t1_iter2__empty_n),
    .fifo_ld_0_s_read(from_t1_iter1_to_t1_iter2__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter2_to_t1_iter3__din),
    .fifo_st_0_full_n(from_t1_iter2_to_t1_iter3__full_n),
    .fifo_st_0_write(from_t1_iter2_to_t1_iter3__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_1
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_1__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter2_to_t1_iter3__dout),
    .fifo_ld_0_peek_dout(from_t1_iter2_to_t1_iter3__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter2_to_t1_iter3__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter2_to_t1_iter3__empty_n),
    .fifo_ld_0_s_read(from_t1_iter2_to_t1_iter3__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter3_to_t1_iter4__din),
    .fifo_st_0_full_n(from_t1_iter3_to_t1_iter4__full_n),
    .fifo_st_0_write(from_t1_iter3_to_t1_iter4__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_2
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_2__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter3_to_t1_iter4__dout),
    .fifo_ld_0_peek_dout(from_t1_iter3_to_t1_iter4__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter3_to_t1_iter4__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter3_to_t1_iter4__empty_n),
    .fifo_ld_0_s_read(from_t1_iter3_to_t1_iter4__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter4_to_t1_iter5__din),
    .fifo_st_0_full_n(from_t1_iter4_to_t1_iter5__full_n),
    .fifo_st_0_write(from_t1_iter4_to_t1_iter5__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_3
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_3__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter4_to_t1_iter5__dout),
    .fifo_ld_0_peek_dout(from_t1_iter4_to_t1_iter5__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter4_to_t1_iter5__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter4_to_t1_iter5__empty_n),
    .fifo_ld_0_s_read(from_t1_iter4_to_t1_iter5__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter5_to_t1_iter6__din),
    .fifo_st_0_full_n(from_t1_iter5_to_t1_iter6__full_n),
    .fifo_st_0_write(from_t1_iter5_to_t1_iter6__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_4
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_4__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter5_to_t1_iter6__dout),
    .fifo_ld_0_peek_dout(from_t1_iter5_to_t1_iter6__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter5_to_t1_iter6__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter5_to_t1_iter6__empty_n),
    .fifo_ld_0_s_read(from_t1_iter5_to_t1_iter6__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter6_to_t1_iter7__din),
    .fifo_st_0_full_n(from_t1_iter6_to_t1_iter7__full_n),
    .fifo_st_0_write(from_t1_iter6_to_t1_iter7__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_5
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_5__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter6_to_t1_iter7__dout),
    .fifo_ld_0_peek_dout(from_t1_iter6_to_t1_iter7__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter6_to_t1_iter7__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter6_to_t1_iter7__empty_n),
    .fifo_ld_0_s_read(from_t1_iter6_to_t1_iter7__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter7_to_t1_iter8__din),
    .fifo_st_0_full_n(from_t1_iter7_to_t1_iter8__full_n),
    .fifo_st_0_write(from_t1_iter7_to_t1_iter8__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_6
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_6__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter7_to_t1_iter8__dout),
    .fifo_ld_0_peek_dout(from_t1_iter7_to_t1_iter8__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter7_to_t1_iter8__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter7_to_t1_iter8__empty_n),
    .fifo_ld_0_s_read(from_t1_iter7_to_t1_iter8__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter8_to_t1_iter9__din),
    .fifo_st_0_full_n(from_t1_iter8_to_t1_iter9__full_n),
    .fifo_st_0_write(from_t1_iter8_to_t1_iter9__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_7
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_7__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter8_to_t1_iter9__dout),
    .fifo_ld_0_peek_dout(from_t1_iter8_to_t1_iter9__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter8_to_t1_iter9__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter8_to_t1_iter9__empty_n),
    .fifo_ld_0_s_read(from_t1_iter8_to_t1_iter9__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter9_to_t1_iter10__din),
    .fifo_st_0_full_n(from_t1_iter9_to_t1_iter10__full_n),
    .fifo_st_0_write(from_t1_iter9_to_t1_iter10__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_8
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_8__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_st_0_din(from_t1_iter10_to_t1_iter11__din),
    .fifo_st_0_full_n(from_t1_iter10_to_t1_iter11__full_n),
    .fifo_st_0_write(from_t1_iter10_to_t1_iter11__write),
    .fifo_ld_0_s_dout(from_t1_iter9_to_t1_iter10__dout),
    .fifo_ld_0_peek_dout(from_t1_iter9_to_t1_iter10__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter9_to_t1_iter10__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter9_to_t1_iter10__empty_n),
    .fifo_ld_0_s_read(from_t1_iter9_to_t1_iter10__read),
    .fifo_ld_0_peek_read()
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_9
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_9__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter10_to_t1_iter11__dout),
    .fifo_ld_0_peek_dout(from_t1_iter10_to_t1_iter11__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter10_to_t1_iter11__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter10_to_t1_iter11__empty_n),
    .fifo_ld_0_s_read(from_t1_iter10_to_t1_iter11__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter11_to_t1_iter12__din),
    .fifo_st_0_full_n(from_t1_iter11_to_t1_iter12__full_n),
    .fifo_st_0_write(from_t1_iter11_to_t1_iter12__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_10
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_10__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter11_to_t1_iter12__dout),
    .fifo_ld_0_peek_dout(from_t1_iter11_to_t1_iter12__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter11_to_t1_iter12__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter11_to_t1_iter12__empty_n),
    .fifo_ld_0_s_read(from_t1_iter11_to_t1_iter12__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter12_to_t1_iter13__din),
    .fifo_st_0_full_n(from_t1_iter12_to_t1_iter13__full_n),
    .fifo_st_0_write(from_t1_iter12_to_t1_iter13__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_11
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_11__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter12_to_t1_iter13__dout),
    .fifo_ld_0_peek_dout(from_t1_iter12_to_t1_iter13__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter12_to_t1_iter13__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter12_to_t1_iter13__empty_n),
    .fifo_ld_0_s_read(from_t1_iter12_to_t1_iter13__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter13_to_t1_iter14__din),
    .fifo_st_0_full_n(from_t1_iter13_to_t1_iter14__full_n),
    .fifo_st_0_write(from_t1_iter13_to_t1_iter14__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_12
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_12__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter13_to_t1_iter14__dout),
    .fifo_ld_0_peek_dout(from_t1_iter13_to_t1_iter14__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter13_to_t1_iter14__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter13_to_t1_iter14__empty_n),
    .fifo_ld_0_s_read(from_t1_iter13_to_t1_iter14__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter14_to_t1_iter15__din),
    .fifo_st_0_full_n(from_t1_iter14_to_t1_iter15__full_n),
    .fifo_st_0_write(from_t1_iter14_to_t1_iter15__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_13
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_13__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter14_to_t1_iter15__dout),
    .fifo_ld_0_peek_dout(from_t1_iter14_to_t1_iter15__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter14_to_t1_iter15__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter14_to_t1_iter15__empty_n),
    .fifo_ld_0_s_read(from_t1_iter14_to_t1_iter15__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter15_to_t1_iter16__din),
    .fifo_st_0_full_n(from_t1_iter15_to_t1_iter16__full_n),
    .fifo_st_0_write(from_t1_iter15_to_t1_iter16__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_14
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_14__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter15_to_t1_iter16__dout),
    .fifo_ld_0_peek_dout(from_t1_iter15_to_t1_iter16__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter15_to_t1_iter16__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter15_to_t1_iter16__empty_n),
    .fifo_ld_0_s_read(from_t1_iter15_to_t1_iter16__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter16_to_t1_iter17__din),
    .fifo_st_0_full_n(from_t1_iter16_to_t1_iter17__full_n),
    .fifo_st_0_write(from_t1_iter16_to_t1_iter17__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_15
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_15__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter16_to_t1_iter17__dout),
    .fifo_ld_0_peek_dout(from_t1_iter16_to_t1_iter17__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter16_to_t1_iter17__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter16_to_t1_iter17__empty_n),
    .fifo_ld_0_s_read(from_t1_iter16_to_t1_iter17__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter17_to_t1_iter18__din),
    .fifo_st_0_full_n(from_t1_iter17_to_t1_iter18__full_n),
    .fifo_st_0_write(from_t1_iter17_to_t1_iter18__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_16
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_16__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter17_to_t1_iter18__dout),
    .fifo_ld_0_peek_dout(from_t1_iter17_to_t1_iter18__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter17_to_t1_iter18__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter17_to_t1_iter18__empty_n),
    .fifo_ld_0_s_read(from_t1_iter17_to_t1_iter18__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter18_to_t1_iter19__din),
    .fifo_st_0_full_n(from_t1_iter18_to_t1_iter19__full_n),
    .fifo_st_0_write(from_t1_iter18_to_t1_iter19__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_17
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_17__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter18_to_t1_iter19__dout),
    .fifo_ld_0_peek_dout(from_t1_iter18_to_t1_iter19__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter18_to_t1_iter19__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter18_to_t1_iter19__empty_n),
    .fifo_ld_0_s_read(from_t1_iter18_to_t1_iter19__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter19_to_t1_iter20__din),
    .fifo_st_0_full_n(from_t1_iter19_to_t1_iter20__full_n),
    .fifo_st_0_write(from_t1_iter19_to_t1_iter20__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_18
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_18__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter19_to_t1_iter20__dout),
    .fifo_ld_0_peek_dout(from_t1_iter19_to_t1_iter20__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter19_to_t1_iter20__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter19_to_t1_iter20__empty_n),
    .fifo_ld_0_s_read(from_t1_iter19_to_t1_iter20__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter20_to_t1_iter21__din),
    .fifo_st_0_full_n(from_t1_iter20_to_t1_iter21__full_n),
    .fifo_st_0_write(from_t1_iter20_to_t1_iter21__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_19
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_19__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter20_to_t1_iter21__dout),
    .fifo_ld_0_peek_dout(from_t1_iter20_to_t1_iter21__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter20_to_t1_iter21__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter20_to_t1_iter21__empty_n),
    .fifo_ld_0_s_read(from_t1_iter20_to_t1_iter21__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter21_to_t1_iter22__din),
    .fifo_st_0_full_n(from_t1_iter21_to_t1_iter22__full_n),
    .fifo_st_0_write(from_t1_iter21_to_t1_iter22__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_20
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_20__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter21_to_t1_iter22__dout),
    .fifo_ld_0_peek_dout(from_t1_iter21_to_t1_iter22__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter21_to_t1_iter22__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter21_to_t1_iter22__empty_n),
    .fifo_ld_0_s_read(from_t1_iter21_to_t1_iter22__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter22_to_t1_iter23__din),
    .fifo_st_0_full_n(from_t1_iter22_to_t1_iter23__full_n),
    .fifo_st_0_write(from_t1_iter22_to_t1_iter23__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_21
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_21__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter22_to_t1_iter23__dout),
    .fifo_ld_0_peek_dout(from_t1_iter22_to_t1_iter23__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter22_to_t1_iter23__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter22_to_t1_iter23__empty_n),
    .fifo_ld_0_s_read(from_t1_iter22_to_t1_iter23__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter23_to_t1_iter24__din),
    .fifo_st_0_full_n(from_t1_iter23_to_t1_iter24__full_n),
    .fifo_st_0_write(from_t1_iter23_to_t1_iter24__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_22
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_22__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter23_to_t1_iter24__dout),
    .fifo_ld_0_peek_dout(from_t1_iter23_to_t1_iter24__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter23_to_t1_iter24__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter23_to_t1_iter24__empty_n),
    .fifo_ld_0_s_read(from_t1_iter23_to_t1_iter24__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter24_to_t1_iter25__din),
    .fifo_st_0_full_n(from_t1_iter24_to_t1_iter25__full_n),
    .fifo_st_0_write(from_t1_iter24_to_t1_iter25__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_23
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_23__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter24_to_t1_iter25__dout),
    .fifo_ld_0_peek_dout(from_t1_iter24_to_t1_iter25__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter24_to_t1_iter25__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter24_to_t1_iter25__empty_n),
    .fifo_ld_0_s_read(from_t1_iter24_to_t1_iter25__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter25_to_t1_iter26__din),
    .fifo_st_0_full_n(from_t1_iter25_to_t1_iter26__full_n),
    .fifo_st_0_write(from_t1_iter25_to_t1_iter26__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_24
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_24__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter25_to_t1_iter26__dout),
    .fifo_ld_0_peek_dout(from_t1_iter25_to_t1_iter26__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter25_to_t1_iter26__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter25_to_t1_iter26__empty_n),
    .fifo_ld_0_s_read(from_t1_iter25_to_t1_iter26__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter26_to_t1_iter27__din),
    .fifo_st_0_full_n(from_t1_iter26_to_t1_iter27__full_n),
    .fifo_st_0_write(from_t1_iter26_to_t1_iter27__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_25
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_25__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter26_to_t1_iter27__dout),
    .fifo_ld_0_peek_dout(from_t1_iter26_to_t1_iter27__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter26_to_t1_iter27__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter26_to_t1_iter27__empty_n),
    .fifo_ld_0_s_read(from_t1_iter26_to_t1_iter27__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter27_to_t1_iter28__din),
    .fifo_st_0_full_n(from_t1_iter27_to_t1_iter28__full_n),
    .fifo_st_0_write(from_t1_iter27_to_t1_iter28__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_26
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_26__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter27_to_t1_iter28__dout),
    .fifo_ld_0_peek_dout(from_t1_iter27_to_t1_iter28__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter27_to_t1_iter28__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter27_to_t1_iter28__empty_n),
    .fifo_ld_0_s_read(from_t1_iter27_to_t1_iter28__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter28_to_t1_iter29__din),
    .fifo_st_0_full_n(from_t1_iter28_to_t1_iter29__full_n),
    .fifo_st_0_write(from_t1_iter28_to_t1_iter29__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_27
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_27__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter28_to_t1_iter29__dout),
    .fifo_ld_0_peek_dout(from_t1_iter28_to_t1_iter29__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter28_to_t1_iter29__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter28_to_t1_iter29__empty_n),
    .fifo_ld_0_s_read(from_t1_iter28_to_t1_iter29__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter29_to_t1_iter30__din),
    .fifo_st_0_full_n(from_t1_iter29_to_t1_iter30__full_n),
    .fifo_st_0_write(from_t1_iter29_to_t1_iter30__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_28
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_28__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter29_to_t1_iter30__dout),
    .fifo_ld_0_peek_dout(from_t1_iter29_to_t1_iter30__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter29_to_t1_iter30__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter29_to_t1_iter30__empty_n),
    .fifo_ld_0_s_read(from_t1_iter29_to_t1_iter30__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter30_to_t1_iter31__din),
    .fifo_st_0_full_n(from_t1_iter30_to_t1_iter31__full_n),
    .fifo_st_0_write(from_t1_iter30_to_t1_iter31__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_29
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_29__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter30_to_t1_iter31__dout),
    .fifo_ld_0_peek_dout(from_t1_iter30_to_t1_iter31__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter30_to_t1_iter31__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter30_to_t1_iter31__empty_n),
    .fifo_ld_0_s_read(from_t1_iter30_to_t1_iter31__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter31_to_t1_iter32__din),
    .fifo_st_0_full_n(from_t1_iter31_to_t1_iter32__full_n),
    .fifo_st_0_write(from_t1_iter31_to_t1_iter32__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_30
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_30__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter31_to_t1_iter32__dout),
    .fifo_ld_0_peek_dout(from_t1_iter31_to_t1_iter32__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter31_to_t1_iter32__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter31_to_t1_iter32__empty_n),
    .fifo_ld_0_s_read(from_t1_iter31_to_t1_iter32__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter32_to_t1_iter33__din),
    .fifo_st_0_full_n(from_t1_iter32_to_t1_iter33__full_n),
    .fifo_st_0_write(from_t1_iter32_to_t1_iter33__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_31
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_31__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter32_to_t1_iter33__dout),
    .fifo_ld_0_peek_dout(from_t1_iter32_to_t1_iter33__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter32_to_t1_iter33__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter32_to_t1_iter33__empty_n),
    .fifo_ld_0_s_read(from_t1_iter32_to_t1_iter33__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter33_to_t1_iter34__din),
    .fifo_st_0_full_n(from_t1_iter33_to_t1_iter34__full_n),
    .fifo_st_0_write(from_t1_iter33_to_t1_iter34__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_32
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_32__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter33_to_t1_iter34__dout),
    .fifo_ld_0_peek_dout(from_t1_iter33_to_t1_iter34__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter33_to_t1_iter34__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter33_to_t1_iter34__empty_n),
    .fifo_ld_0_s_read(from_t1_iter33_to_t1_iter34__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter34_to_t1_iter35__din),
    .fifo_st_0_full_n(from_t1_iter34_to_t1_iter35__full_n),
    .fifo_st_0_write(from_t1_iter34_to_t1_iter35__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_33
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_33__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter34_to_t1_iter35__dout),
    .fifo_ld_0_peek_dout(from_t1_iter34_to_t1_iter35__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter34_to_t1_iter35__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter34_to_t1_iter35__empty_n),
    .fifo_ld_0_s_read(from_t1_iter34_to_t1_iter35__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter35_to_t1_iter36__din),
    .fifo_st_0_full_n(from_t1_iter35_to_t1_iter36__full_n),
    .fifo_st_0_write(from_t1_iter35_to_t1_iter36__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_34
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_34__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter35_to_t1_iter36__dout),
    .fifo_ld_0_peek_dout(from_t1_iter35_to_t1_iter36__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter35_to_t1_iter36__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter35_to_t1_iter36__empty_n),
    .fifo_ld_0_s_read(from_t1_iter35_to_t1_iter36__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter36_to_t1_iter37__din),
    .fifo_st_0_full_n(from_t1_iter36_to_t1_iter37__full_n),
    .fifo_st_0_write(from_t1_iter36_to_t1_iter37__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_35
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_35__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter36_to_t1_iter37__dout),
    .fifo_ld_0_peek_dout(from_t1_iter36_to_t1_iter37__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter36_to_t1_iter37__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter36_to_t1_iter37__empty_n),
    .fifo_ld_0_s_read(from_t1_iter36_to_t1_iter37__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter37_to_t1_iter38__din),
    .fifo_st_0_full_n(from_t1_iter37_to_t1_iter38__full_n),
    .fifo_st_0_write(from_t1_iter37_to_t1_iter38__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_36
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_36__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter37_to_t1_iter38__dout),
    .fifo_ld_0_peek_dout(from_t1_iter37_to_t1_iter38__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter37_to_t1_iter38__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter37_to_t1_iter38__empty_n),
    .fifo_ld_0_s_read(from_t1_iter37_to_t1_iter38__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter38_to_t1_iter39__din),
    .fifo_st_0_full_n(from_t1_iter38_to_t1_iter39__full_n),
    .fifo_st_0_write(from_t1_iter38_to_t1_iter39__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_37
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_37__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter38_to_t1_iter39__dout),
    .fifo_ld_0_peek_dout(from_t1_iter38_to_t1_iter39__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter38_to_t1_iter39__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter38_to_t1_iter39__empty_n),
    .fifo_ld_0_s_read(from_t1_iter38_to_t1_iter39__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter39_to_t1_iter40__din),
    .fifo_st_0_full_n(from_t1_iter39_to_t1_iter40__full_n),
    .fifo_st_0_write(from_t1_iter39_to_t1_iter40__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_38
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_38__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter39_to_t1_iter40__dout),
    .fifo_ld_0_peek_dout(from_t1_iter39_to_t1_iter40__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter39_to_t1_iter40__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter39_to_t1_iter40__empty_n),
    .fifo_ld_0_s_read(from_t1_iter39_to_t1_iter40__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter40_to_t1_iter41__din),
    .fifo_st_0_full_n(from_t1_iter40_to_t1_iter41__full_n),
    .fifo_st_0_write(from_t1_iter40_to_t1_iter41__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_39
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_39__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter40_to_t1_iter41__dout),
    .fifo_ld_0_peek_dout(from_t1_iter40_to_t1_iter41__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter40_to_t1_iter41__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter40_to_t1_iter41__empty_n),
    .fifo_ld_0_s_read(from_t1_iter40_to_t1_iter41__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter41_to_t1_iter42__din),
    .fifo_st_0_full_n(from_t1_iter41_to_t1_iter42__full_n),
    .fifo_st_0_write(from_t1_iter41_to_t1_iter42__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_40
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_40__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter41_to_t1_iter42__dout),
    .fifo_ld_0_peek_dout(from_t1_iter41_to_t1_iter42__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter41_to_t1_iter42__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter41_to_t1_iter42__empty_n),
    .fifo_ld_0_s_read(from_t1_iter41_to_t1_iter42__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter42_to_t1_iter43__din),
    .fifo_st_0_full_n(from_t1_iter42_to_t1_iter43__full_n),
    .fifo_st_0_write(from_t1_iter42_to_t1_iter43__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_41
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_41__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter42_to_t1_iter43__dout),
    .fifo_ld_0_peek_dout(from_t1_iter42_to_t1_iter43__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter42_to_t1_iter43__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter42_to_t1_iter43__empty_n),
    .fifo_ld_0_s_read(from_t1_iter42_to_t1_iter43__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter43_to_t1_iter44__din),
    .fifo_st_0_full_n(from_t1_iter43_to_t1_iter44__full_n),
    .fifo_st_0_write(from_t1_iter43_to_t1_iter44__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_42
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_42__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter43_to_t1_iter44__dout),
    .fifo_ld_0_peek_dout(from_t1_iter43_to_t1_iter44__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter43_to_t1_iter44__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter43_to_t1_iter44__empty_n),
    .fifo_ld_0_s_read(from_t1_iter43_to_t1_iter44__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter44_to_t1_iter45__din),
    .fifo_st_0_full_n(from_t1_iter44_to_t1_iter45__full_n),
    .fifo_st_0_write(from_t1_iter44_to_t1_iter45__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_43
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_43__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter44_to_t1_iter45__dout),
    .fifo_ld_0_peek_dout(from_t1_iter44_to_t1_iter45__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter44_to_t1_iter45__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter44_to_t1_iter45__empty_n),
    .fifo_ld_0_s_read(from_t1_iter44_to_t1_iter45__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter45_to_t1_iter46__din),
    .fifo_st_0_full_n(from_t1_iter45_to_t1_iter46__full_n),
    .fifo_st_0_write(from_t1_iter45_to_t1_iter46__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_44
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_44__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter45_to_t1_iter46__dout),
    .fifo_ld_0_peek_dout(from_t1_iter45_to_t1_iter46__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter45_to_t1_iter46__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter45_to_t1_iter46__empty_n),
    .fifo_ld_0_s_read(from_t1_iter45_to_t1_iter46__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter46_to_t1_iter47__din),
    .fifo_st_0_full_n(from_t1_iter46_to_t1_iter47__full_n),
    .fifo_st_0_write(from_t1_iter46_to_t1_iter47__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_45
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_45__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter46_to_t1_iter47__dout),
    .fifo_ld_0_peek_dout(from_t1_iter46_to_t1_iter47__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter46_to_t1_iter47__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter46_to_t1_iter47__empty_n),
    .fifo_ld_0_s_read(from_t1_iter46_to_t1_iter47__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter47_to_t1_iter48__din),
    .fifo_st_0_full_n(from_t1_iter47_to_t1_iter48__full_n),
    .fifo_st_0_write(from_t1_iter47_to_t1_iter48__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_46
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_46__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter47_to_t1_iter48__dout),
    .fifo_ld_0_peek_dout(from_t1_iter47_to_t1_iter48__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter47_to_t1_iter48__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter47_to_t1_iter48__empty_n),
    .fifo_ld_0_s_read(from_t1_iter47_to_t1_iter48__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter48_to_t1_iter49__din),
    .fifo_st_0_full_n(from_t1_iter48_to_t1_iter49__full_n),
    .fifo_st_0_write(from_t1_iter48_to_t1_iter49__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_47
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_47__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter48_to_t1_iter49__dout),
    .fifo_ld_0_peek_dout(from_t1_iter48_to_t1_iter49__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter48_to_t1_iter49__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter48_to_t1_iter49__empty_n),
    .fifo_ld_0_s_read(from_t1_iter48_to_t1_iter49__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter49_to_t1_iter50__din),
    .fifo_st_0_full_n(from_t1_iter49_to_t1_iter50__full_n),
    .fifo_st_0_write(from_t1_iter49_to_t1_iter50__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_48
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_48__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter49_to_t1_iter50__dout),
    .fifo_ld_0_peek_dout(from_t1_iter49_to_t1_iter50__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter49_to_t1_iter50__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter49_to_t1_iter50__empty_n),
    .fifo_ld_0_s_read(from_t1_iter49_to_t1_iter50__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter50_to_t1_iter51__din),
    .fifo_st_0_full_n(from_t1_iter50_to_t1_iter51__full_n),
    .fifo_st_0_write(from_t1_iter50_to_t1_iter51__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_49
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_49__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter50_to_t1_iter51__dout),
    .fifo_ld_0_peek_dout(from_t1_iter50_to_t1_iter51__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter50_to_t1_iter51__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter50_to_t1_iter51__empty_n),
    .fifo_ld_0_s_read(from_t1_iter50_to_t1_iter51__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter51_to_t1_iter52__din),
    .fifo_st_0_full_n(from_t1_iter51_to_t1_iter52__full_n),
    .fifo_st_0_write(from_t1_iter51_to_t1_iter52__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_50
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_50__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter51_to_t1_iter52__dout),
    .fifo_ld_0_peek_dout(from_t1_iter51_to_t1_iter52__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter51_to_t1_iter52__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter51_to_t1_iter52__empty_n),
    .fifo_ld_0_s_read(from_t1_iter51_to_t1_iter52__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter52_to_t1_iter53__din),
    .fifo_st_0_full_n(from_t1_iter52_to_t1_iter53__full_n),
    .fifo_st_0_write(from_t1_iter52_to_t1_iter53__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_51
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_51__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter52_to_t1_iter53__dout),
    .fifo_ld_0_peek_dout(from_t1_iter52_to_t1_iter53__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter52_to_t1_iter53__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter52_to_t1_iter53__empty_n),
    .fifo_ld_0_s_read(from_t1_iter52_to_t1_iter53__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter53_to_t1_iter54__din),
    .fifo_st_0_full_n(from_t1_iter53_to_t1_iter54__full_n),
    .fifo_st_0_write(from_t1_iter53_to_t1_iter54__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_52
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_52__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter53_to_t1_iter54__dout),
    .fifo_ld_0_peek_dout(from_t1_iter53_to_t1_iter54__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter53_to_t1_iter54__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter53_to_t1_iter54__empty_n),
    .fifo_ld_0_s_read(from_t1_iter53_to_t1_iter54__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter54_to_t1_iter55__din),
    .fifo_st_0_full_n(from_t1_iter54_to_t1_iter55__full_n),
    .fifo_st_0_write(from_t1_iter54_to_t1_iter55__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_53
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_53__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter54_to_t1_iter55__dout),
    .fifo_ld_0_peek_dout(from_t1_iter54_to_t1_iter55__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter54_to_t1_iter55__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter54_to_t1_iter55__empty_n),
    .fifo_ld_0_s_read(from_t1_iter54_to_t1_iter55__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter55_to_t1_iter56__din),
    .fifo_st_0_full_n(from_t1_iter55_to_t1_iter56__full_n),
    .fifo_st_0_write(from_t1_iter55_to_t1_iter56__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_54
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_54__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter55_to_t1_iter56__dout),
    .fifo_ld_0_peek_dout(from_t1_iter55_to_t1_iter56__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter55_to_t1_iter56__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter55_to_t1_iter56__empty_n),
    .fifo_ld_0_s_read(from_t1_iter55_to_t1_iter56__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter56_to_t1_iter57__din),
    .fifo_st_0_full_n(from_t1_iter56_to_t1_iter57__full_n),
    .fifo_st_0_write(from_t1_iter56_to_t1_iter57__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_55
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_55__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter56_to_t1_iter57__dout),
    .fifo_ld_0_peek_dout(from_t1_iter56_to_t1_iter57__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter56_to_t1_iter57__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter56_to_t1_iter57__empty_n),
    .fifo_ld_0_s_read(from_t1_iter56_to_t1_iter57__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter57_to_t1_iter58__din),
    .fifo_st_0_full_n(from_t1_iter57_to_t1_iter58__full_n),
    .fifo_st_0_write(from_t1_iter57_to_t1_iter58__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_56
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_56__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter57_to_t1_iter58__dout),
    .fifo_ld_0_peek_dout(from_t1_iter57_to_t1_iter58__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter57_to_t1_iter58__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter57_to_t1_iter58__empty_n),
    .fifo_ld_0_s_read(from_t1_iter57_to_t1_iter58__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter58_to_t1_iter59__din),
    .fifo_st_0_full_n(from_t1_iter58_to_t1_iter59__full_n),
    .fifo_st_0_write(from_t1_iter58_to_t1_iter59__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_57
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_57__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter58_to_t1_iter59__dout),
    .fifo_ld_0_peek_dout(from_t1_iter58_to_t1_iter59__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter58_to_t1_iter59__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter58_to_t1_iter59__empty_n),
    .fifo_ld_0_s_read(from_t1_iter58_to_t1_iter59__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter59_to_t1_iter60__din),
    .fifo_st_0_full_n(from_t1_iter59_to_t1_iter60__full_n),
    .fifo_st_0_write(from_t1_iter59_to_t1_iter60__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_58
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_58__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter59_to_t1_iter60__dout),
    .fifo_ld_0_peek_dout(from_t1_iter59_to_t1_iter60__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter59_to_t1_iter60__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter59_to_t1_iter60__empty_n),
    .fifo_ld_0_s_read(from_t1_iter59_to_t1_iter60__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter60_to_t1_iter61__din),
    .fifo_st_0_full_n(from_t1_iter60_to_t1_iter61__full_n),
    .fifo_st_0_write(from_t1_iter60_to_t1_iter61__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_59
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_59__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter60_to_t1_iter61__dout),
    .fifo_ld_0_peek_dout(from_t1_iter60_to_t1_iter61__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter60_to_t1_iter61__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter60_to_t1_iter61__empty_n),
    .fifo_ld_0_s_read(from_t1_iter60_to_t1_iter61__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter61_to_t1_iter62__din),
    .fifo_st_0_full_n(from_t1_iter61_to_t1_iter62__full_n),
    .fifo_st_0_write(from_t1_iter61_to_t1_iter62__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_60
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_60__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter61_to_t1_iter62__dout),
    .fifo_ld_0_peek_dout(from_t1_iter61_to_t1_iter62__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter61_to_t1_iter62__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter61_to_t1_iter62__empty_n),
    .fifo_ld_0_s_read(from_t1_iter61_to_t1_iter62__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter62_to_t1_iter63__din),
    .fifo_st_0_full_n(from_t1_iter62_to_t1_iter63__full_n),
    .fifo_st_0_write(from_t1_iter62_to_t1_iter63__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_61
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_61__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter62_to_t1_iter63__dout),
    .fifo_ld_0_peek_dout(from_t1_iter62_to_t1_iter63__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter62_to_t1_iter63__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter62_to_t1_iter63__empty_n),
    .fifo_ld_0_s_read(from_t1_iter62_to_t1_iter63__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter63_to_t1_iter64__din),
    .fifo_st_0_full_n(from_t1_iter63_to_t1_iter64__full_n),
    .fifo_st_0_write(from_t1_iter63_to_t1_iter64__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_62
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_62__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter63_to_t1_iter64__dout),
    .fifo_ld_0_peek_dout(from_t1_iter63_to_t1_iter64__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter63_to_t1_iter64__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter63_to_t1_iter64__empty_n),
    .fifo_ld_0_s_read(from_t1_iter63_to_t1_iter64__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter64_to_t1_iter65__din),
    .fifo_st_0_full_n(from_t1_iter64_to_t1_iter65__full_n),
    .fifo_st_0_write(from_t1_iter64_to_t1_iter65__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_63
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_63__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter64_to_t1_iter65__dout),
    .fifo_ld_0_peek_dout(from_t1_iter64_to_t1_iter65__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter64_to_t1_iter65__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter64_to_t1_iter65__empty_n),
    .fifo_ld_0_s_read(from_t1_iter64_to_t1_iter65__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter65_to_t1_iter66__din),
    .fifo_st_0_full_n(from_t1_iter65_to_t1_iter66__full_n),
    .fifo_st_0_write(from_t1_iter65_to_t1_iter66__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_64
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_64__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter65_to_t1_iter66__dout),
    .fifo_ld_0_peek_dout(from_t1_iter65_to_t1_iter66__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter65_to_t1_iter66__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter65_to_t1_iter66__empty_n),
    .fifo_ld_0_s_read(from_t1_iter65_to_t1_iter66__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter66_to_t1_iter67__din),
    .fifo_st_0_full_n(from_t1_iter66_to_t1_iter67__full_n),
    .fifo_st_0_write(from_t1_iter66_to_t1_iter67__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_65
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_65__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter66_to_t1_iter67__dout),
    .fifo_ld_0_peek_dout(from_t1_iter66_to_t1_iter67__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter66_to_t1_iter67__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter66_to_t1_iter67__empty_n),
    .fifo_ld_0_s_read(from_t1_iter66_to_t1_iter67__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter67_to_t1_iter68__din),
    .fifo_st_0_full_n(from_t1_iter67_to_t1_iter68__full_n),
    .fifo_st_0_write(from_t1_iter67_to_t1_iter68__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_66
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_66__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter67_to_t1_iter68__dout),
    .fifo_ld_0_peek_dout(from_t1_iter67_to_t1_iter68__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter67_to_t1_iter68__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter67_to_t1_iter68__empty_n),
    .fifo_ld_0_s_read(from_t1_iter67_to_t1_iter68__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter68_to_t1_iter69__din),
    .fifo_st_0_full_n(from_t1_iter68_to_t1_iter69__full_n),
    .fifo_st_0_write(from_t1_iter68_to_t1_iter69__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_67
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_67__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter68_to_t1_iter69__dout),
    .fifo_ld_0_peek_dout(from_t1_iter68_to_t1_iter69__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter68_to_t1_iter69__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter68_to_t1_iter69__empty_n),
    .fifo_ld_0_s_read(from_t1_iter68_to_t1_iter69__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter69_to_t1_iter70__din),
    .fifo_st_0_full_n(from_t1_iter69_to_t1_iter70__full_n),
    .fifo_st_0_write(from_t1_iter69_to_t1_iter70__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_68
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_68__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter69_to_t1_iter70__dout),
    .fifo_ld_0_peek_dout(from_t1_iter69_to_t1_iter70__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter69_to_t1_iter70__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter69_to_t1_iter70__empty_n),
    .fifo_ld_0_s_read(from_t1_iter69_to_t1_iter70__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter70_to_t1_iter71__din),
    .fifo_st_0_full_n(from_t1_iter70_to_t1_iter71__full_n),
    .fifo_st_0_write(from_t1_iter70_to_t1_iter71__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_69
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_69__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter70_to_t1_iter71__dout),
    .fifo_ld_0_peek_dout(from_t1_iter70_to_t1_iter71__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter70_to_t1_iter71__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter70_to_t1_iter71__empty_n),
    .fifo_ld_0_s_read(from_t1_iter70_to_t1_iter71__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter71_to_t1_iter72__din),
    .fifo_st_0_full_n(from_t1_iter71_to_t1_iter72__full_n),
    .fifo_st_0_write(from_t1_iter71_to_t1_iter72__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_70
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_70__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter71_to_t1_iter72__dout),
    .fifo_ld_0_peek_dout(from_t1_iter71_to_t1_iter72__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter71_to_t1_iter72__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter71_to_t1_iter72__empty_n),
    .fifo_ld_0_s_read(from_t1_iter71_to_t1_iter72__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter72_to_t1_iter73__din),
    .fifo_st_0_full_n(from_t1_iter72_to_t1_iter73__full_n),
    .fifo_st_0_write(from_t1_iter72_to_t1_iter73__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_71
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_71__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter72_to_t1_iter73__dout),
    .fifo_ld_0_peek_dout(from_t1_iter72_to_t1_iter73__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter72_to_t1_iter73__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter72_to_t1_iter73__empty_n),
    .fifo_ld_0_s_read(from_t1_iter72_to_t1_iter73__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter73_to_t1_iter74__din),
    .fifo_st_0_full_n(from_t1_iter73_to_t1_iter74__full_n),
    .fifo_st_0_write(from_t1_iter73_to_t1_iter74__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_72
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_72__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter73_to_t1_iter74__dout),
    .fifo_ld_0_peek_dout(from_t1_iter73_to_t1_iter74__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter73_to_t1_iter74__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter73_to_t1_iter74__empty_n),
    .fifo_ld_0_s_read(from_t1_iter73_to_t1_iter74__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter74_to_t1_iter75__din),
    .fifo_st_0_full_n(from_t1_iter74_to_t1_iter75__full_n),
    .fifo_st_0_write(from_t1_iter74_to_t1_iter75__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_73
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_73__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter74_to_t1_iter75__dout),
    .fifo_ld_0_peek_dout(from_t1_iter74_to_t1_iter75__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter74_to_t1_iter75__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter74_to_t1_iter75__empty_n),
    .fifo_ld_0_s_read(from_t1_iter74_to_t1_iter75__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter75_to_t1_iter76__din),
    .fifo_st_0_full_n(from_t1_iter75_to_t1_iter76__full_n),
    .fifo_st_0_write(from_t1_iter75_to_t1_iter76__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_74
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_74__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter75_to_t1_iter76__dout),
    .fifo_ld_0_peek_dout(from_t1_iter75_to_t1_iter76__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter75_to_t1_iter76__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter75_to_t1_iter76__empty_n),
    .fifo_ld_0_s_read(from_t1_iter75_to_t1_iter76__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter76_to_t1_iter77__din),
    .fifo_st_0_full_n(from_t1_iter76_to_t1_iter77__full_n),
    .fifo_st_0_write(from_t1_iter76_to_t1_iter77__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_75
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_75__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter76_to_t1_iter77__dout),
    .fifo_ld_0_peek_dout(from_t1_iter76_to_t1_iter77__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter76_to_t1_iter77__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter76_to_t1_iter77__empty_n),
    .fifo_ld_0_s_read(from_t1_iter76_to_t1_iter77__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter77_to_t1_iter78__din),
    .fifo_st_0_full_n(from_t1_iter77_to_t1_iter78__full_n),
    .fifo_st_0_write(from_t1_iter77_to_t1_iter78__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_76
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_76__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter77_to_t1_iter78__dout),
    .fifo_ld_0_peek_dout(from_t1_iter77_to_t1_iter78__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter77_to_t1_iter78__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter77_to_t1_iter78__empty_n),
    .fifo_ld_0_s_read(from_t1_iter77_to_t1_iter78__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter78_to_t1_iter79__din),
    .fifo_st_0_full_n(from_t1_iter78_to_t1_iter79__full_n),
    .fifo_st_0_write(from_t1_iter78_to_t1_iter79__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_77
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_77__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter78_to_t1_iter79__dout),
    .fifo_ld_0_peek_dout(from_t1_iter78_to_t1_iter79__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter78_to_t1_iter79__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter78_to_t1_iter79__empty_n),
    .fifo_ld_0_s_read(from_t1_iter78_to_t1_iter79__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter79_to_t1_iter80__din),
    .fifo_st_0_full_n(from_t1_iter79_to_t1_iter80__full_n),
    .fifo_st_0_write(from_t1_iter79_to_t1_iter80__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_78
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_78__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter79_to_t1_iter80__dout),
    .fifo_ld_0_peek_dout(from_t1_iter79_to_t1_iter80__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter79_to_t1_iter80__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter79_to_t1_iter80__empty_n),
    .fifo_ld_0_s_read(from_t1_iter79_to_t1_iter80__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter80_to_t1_iter81__din),
    .fifo_st_0_full_n(from_t1_iter80_to_t1_iter81__full_n),
    .fifo_st_0_write(from_t1_iter80_to_t1_iter81__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_79
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_79__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter80_to_t1_iter81__dout),
    .fifo_ld_0_peek_dout(from_t1_iter80_to_t1_iter81__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter80_to_t1_iter81__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter80_to_t1_iter81__empty_n),
    .fifo_ld_0_s_read(from_t1_iter80_to_t1_iter81__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter81_to_t1_iter82__din),
    .fifo_st_0_full_n(from_t1_iter81_to_t1_iter82__full_n),
    .fifo_st_0_write(from_t1_iter81_to_t1_iter82__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_80
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_80__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter81_to_t1_iter82__dout),
    .fifo_ld_0_peek_dout(from_t1_iter81_to_t1_iter82__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter81_to_t1_iter82__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter81_to_t1_iter82__empty_n),
    .fifo_ld_0_s_read(from_t1_iter81_to_t1_iter82__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter82_to_t1_iter83__din),
    .fifo_st_0_full_n(from_t1_iter82_to_t1_iter83__full_n),
    .fifo_st_0_write(from_t1_iter82_to_t1_iter83__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_81
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_81__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter82_to_t1_iter83__dout),
    .fifo_ld_0_peek_dout(from_t1_iter82_to_t1_iter83__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter82_to_t1_iter83__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter82_to_t1_iter83__empty_n),
    .fifo_ld_0_s_read(from_t1_iter82_to_t1_iter83__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter83_to_t1_iter84__din),
    .fifo_st_0_full_n(from_t1_iter83_to_t1_iter84__full_n),
    .fifo_st_0_write(from_t1_iter83_to_t1_iter84__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_82
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_82__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter83_to_t1_iter84__dout),
    .fifo_ld_0_peek_dout(from_t1_iter83_to_t1_iter84__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter83_to_t1_iter84__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter83_to_t1_iter84__empty_n),
    .fifo_ld_0_s_read(from_t1_iter83_to_t1_iter84__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter84_to_t1_iter85__din),
    .fifo_st_0_full_n(from_t1_iter84_to_t1_iter85__full_n),
    .fifo_st_0_write(from_t1_iter84_to_t1_iter85__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_83
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_83__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter84_to_t1_iter85__dout),
    .fifo_ld_0_peek_dout(from_t1_iter84_to_t1_iter85__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter84_to_t1_iter85__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter84_to_t1_iter85__empty_n),
    .fifo_ld_0_s_read(from_t1_iter84_to_t1_iter85__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter85_to_t1_iter86__din),
    .fifo_st_0_full_n(from_t1_iter85_to_t1_iter86__full_n),
    .fifo_st_0_write(from_t1_iter85_to_t1_iter86__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_84
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_84__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter85_to_t1_iter86__dout),
    .fifo_ld_0_peek_dout(from_t1_iter85_to_t1_iter86__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter85_to_t1_iter86__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter85_to_t1_iter86__empty_n),
    .fifo_ld_0_s_read(from_t1_iter85_to_t1_iter86__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter86_to_t1_iter87__din),
    .fifo_st_0_full_n(from_t1_iter86_to_t1_iter87__full_n),
    .fifo_st_0_write(from_t1_iter86_to_t1_iter87__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_85
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_85__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter86_to_t1_iter87__dout),
    .fifo_ld_0_peek_dout(from_t1_iter86_to_t1_iter87__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter86_to_t1_iter87__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter86_to_t1_iter87__empty_n),
    .fifo_ld_0_s_read(from_t1_iter86_to_t1_iter87__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter87_to_t1_iter88__din),
    .fifo_st_0_full_n(from_t1_iter87_to_t1_iter88__full_n),
    .fifo_st_0_write(from_t1_iter87_to_t1_iter88__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_86
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_86__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter87_to_t1_iter88__dout),
    .fifo_ld_0_peek_dout(from_t1_iter87_to_t1_iter88__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter87_to_t1_iter88__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter87_to_t1_iter88__empty_n),
    .fifo_ld_0_s_read(from_t1_iter87_to_t1_iter88__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter88_to_t1_iter89__din),
    .fifo_st_0_full_n(from_t1_iter88_to_t1_iter89__full_n),
    .fifo_st_0_write(from_t1_iter88_to_t1_iter89__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_87
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_87__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter88_to_t1_iter89__dout),
    .fifo_ld_0_peek_dout(from_t1_iter88_to_t1_iter89__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter88_to_t1_iter89__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter88_to_t1_iter89__empty_n),
    .fifo_ld_0_s_read(from_t1_iter88_to_t1_iter89__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter89_to_t1_iter90__din),
    .fifo_st_0_full_n(from_t1_iter89_to_t1_iter90__full_n),
    .fifo_st_0_write(from_t1_iter89_to_t1_iter90__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_88
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_88__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter89_to_t1_iter90__dout),
    .fifo_ld_0_peek_dout(from_t1_iter89_to_t1_iter90__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter89_to_t1_iter90__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter89_to_t1_iter90__empty_n),
    .fifo_ld_0_s_read(from_t1_iter89_to_t1_iter90__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter90_to_t1_iter91__din),
    .fifo_st_0_full_n(from_t1_iter90_to_t1_iter91__full_n),
    .fifo_st_0_write(from_t1_iter90_to_t1_iter91__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_89
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_89__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter90_to_t1_iter91__dout),
    .fifo_ld_0_peek_dout(from_t1_iter90_to_t1_iter91__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter90_to_t1_iter91__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter90_to_t1_iter91__empty_n),
    .fifo_ld_0_s_read(from_t1_iter90_to_t1_iter91__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter91_to_t1_iter92__din),
    .fifo_st_0_full_n(from_t1_iter91_to_t1_iter92__full_n),
    .fifo_st_0_write(from_t1_iter91_to_t1_iter92__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_90
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_90__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter91_to_t1_iter92__dout),
    .fifo_ld_0_peek_dout(from_t1_iter91_to_t1_iter92__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter91_to_t1_iter92__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter91_to_t1_iter92__empty_n),
    .fifo_ld_0_s_read(from_t1_iter91_to_t1_iter92__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter92_to_t1_iter93__din),
    .fifo_st_0_full_n(from_t1_iter92_to_t1_iter93__full_n),
    .fifo_st_0_write(from_t1_iter92_to_t1_iter93__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_91
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_91__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter92_to_t1_iter93__dout),
    .fifo_ld_0_peek_dout(from_t1_iter92_to_t1_iter93__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter92_to_t1_iter93__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter92_to_t1_iter93__empty_n),
    .fifo_ld_0_s_read(from_t1_iter92_to_t1_iter93__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter93_to_t1_iter94__din),
    .fifo_st_0_full_n(from_t1_iter93_to_t1_iter94__full_n),
    .fifo_st_0_write(from_t1_iter93_to_t1_iter94__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_92
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_92__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter93_to_t1_iter94__dout),
    .fifo_ld_0_peek_dout(from_t1_iter93_to_t1_iter94__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter93_to_t1_iter94__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter93_to_t1_iter94__empty_n),
    .fifo_ld_0_s_read(from_t1_iter93_to_t1_iter94__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter94_to_t1_iter95__din),
    .fifo_st_0_full_n(from_t1_iter94_to_t1_iter95__full_n),
    .fifo_st_0_write(from_t1_iter94_to_t1_iter95__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_93
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_93__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter94_to_t1_iter95__dout),
    .fifo_ld_0_peek_dout(from_t1_iter94_to_t1_iter95__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter94_to_t1_iter95__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter94_to_t1_iter95__empty_n),
    .fifo_ld_0_s_read(from_t1_iter94_to_t1_iter95__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter95_to_t1_iter96__din),
    .fifo_st_0_full_n(from_t1_iter95_to_t1_iter96__full_n),
    .fifo_st_0_write(from_t1_iter95_to_t1_iter96__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_94
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_94__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter95_to_t1_iter96__dout),
    .fifo_ld_0_peek_dout(from_t1_iter95_to_t1_iter96__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter95_to_t1_iter96__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter95_to_t1_iter96__empty_n),
    .fifo_ld_0_s_read(from_t1_iter95_to_t1_iter96__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter96_to_t1_iter97__din),
    .fifo_st_0_full_n(from_t1_iter96_to_t1_iter97__full_n),
    .fifo_st_0_write(from_t1_iter96_to_t1_iter97__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_95
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_95__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter96_to_t1_iter97__dout),
    .fifo_ld_0_peek_dout(from_t1_iter96_to_t1_iter97__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter96_to_t1_iter97__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter96_to_t1_iter97__empty_n),
    .fifo_ld_0_s_read(from_t1_iter96_to_t1_iter97__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter97_to_t1_iter98__din),
    .fifo_st_0_full_n(from_t1_iter97_to_t1_iter98__full_n),
    .fifo_st_0_write(from_t1_iter97_to_t1_iter98__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_96
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_96__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter97_to_t1_iter98__dout),
    .fifo_ld_0_peek_dout(from_t1_iter97_to_t1_iter98__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter97_to_t1_iter98__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter97_to_t1_iter98__empty_n),
    .fifo_ld_0_s_read(from_t1_iter97_to_t1_iter98__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter98_to_t1_iter99__din),
    .fifo_st_0_full_n(from_t1_iter98_to_t1_iter99__full_n),
    .fifo_st_0_write(from_t1_iter98_to_t1_iter99__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_97
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_97__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter98_to_t1_iter99__dout),
    .fifo_ld_0_peek_dout(from_t1_iter98_to_t1_iter99__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter98_to_t1_iter99__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter98_to_t1_iter99__empty_n),
    .fifo_ld_0_s_read(from_t1_iter98_to_t1_iter99__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter99_to_t1_iter100__din),
    .fifo_st_0_full_n(from_t1_iter99_to_t1_iter100__full_n),
    .fifo_st_0_write(from_t1_iter99_to_t1_iter100__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_98
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_98__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_st_0_din(from_t1_iter100_to_t1_iter101__din),
    .fifo_st_0_full_n(from_t1_iter100_to_t1_iter101__full_n),
    .fifo_st_0_write(from_t1_iter100_to_t1_iter101__write),
    .fifo_ld_0_s_dout(from_t1_iter99_to_t1_iter100__dout),
    .fifo_ld_0_peek_dout(from_t1_iter99_to_t1_iter100__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter99_to_t1_iter100__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter99_to_t1_iter100__empty_n),
    .fifo_ld_0_s_read(from_t1_iter99_to_t1_iter100__read),
    .fifo_ld_0_peek_read()
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_99
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_99__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter100_to_t1_iter101__dout),
    .fifo_ld_0_peek_dout(from_t1_iter100_to_t1_iter101__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter100_to_t1_iter101__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter100_to_t1_iter101__empty_n),
    .fifo_ld_0_s_read(from_t1_iter100_to_t1_iter101__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter101_to_t1_iter102__din),
    .fifo_st_0_full_n(from_t1_iter101_to_t1_iter102__full_n),
    .fifo_st_0_write(from_t1_iter101_to_t1_iter102__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_100
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_100__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter101_to_t1_iter102__dout),
    .fifo_ld_0_peek_dout(from_t1_iter101_to_t1_iter102__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter101_to_t1_iter102__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter101_to_t1_iter102__empty_n),
    .fifo_ld_0_s_read(from_t1_iter101_to_t1_iter102__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter102_to_t1_iter103__din),
    .fifo_st_0_full_n(from_t1_iter102_to_t1_iter103__full_n),
    .fifo_st_0_write(from_t1_iter102_to_t1_iter103__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_101
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_101__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter102_to_t1_iter103__dout),
    .fifo_ld_0_peek_dout(from_t1_iter102_to_t1_iter103__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter102_to_t1_iter103__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter102_to_t1_iter103__empty_n),
    .fifo_ld_0_s_read(from_t1_iter102_to_t1_iter103__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter103_to_t1_iter104__din),
    .fifo_st_0_full_n(from_t1_iter103_to_t1_iter104__full_n),
    .fifo_st_0_write(from_t1_iter103_to_t1_iter104__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_102
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_102__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter103_to_t1_iter104__dout),
    .fifo_ld_0_peek_dout(from_t1_iter103_to_t1_iter104__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter103_to_t1_iter104__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter103_to_t1_iter104__empty_n),
    .fifo_ld_0_s_read(from_t1_iter103_to_t1_iter104__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter104_to_t1_iter105__din),
    .fifo_st_0_full_n(from_t1_iter104_to_t1_iter105__full_n),
    .fifo_st_0_write(from_t1_iter104_to_t1_iter105__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_103
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_103__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter104_to_t1_iter105__dout),
    .fifo_ld_0_peek_dout(from_t1_iter104_to_t1_iter105__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter104_to_t1_iter105__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter104_to_t1_iter105__empty_n),
    .fifo_ld_0_s_read(from_t1_iter104_to_t1_iter105__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter105_to_t1_iter106__din),
    .fifo_st_0_full_n(from_t1_iter105_to_t1_iter106__full_n),
    .fifo_st_0_write(from_t1_iter105_to_t1_iter106__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_104
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_104__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter105_to_t1_iter106__dout),
    .fifo_ld_0_peek_dout(from_t1_iter105_to_t1_iter106__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter105_to_t1_iter106__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter105_to_t1_iter106__empty_n),
    .fifo_ld_0_s_read(from_t1_iter105_to_t1_iter106__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter106_to_t1_iter107__din),
    .fifo_st_0_full_n(from_t1_iter106_to_t1_iter107__full_n),
    .fifo_st_0_write(from_t1_iter106_to_t1_iter107__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_105
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_105__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter106_to_t1_iter107__dout),
    .fifo_ld_0_peek_dout(from_t1_iter106_to_t1_iter107__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter106_to_t1_iter107__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter106_to_t1_iter107__empty_n),
    .fifo_ld_0_s_read(from_t1_iter106_to_t1_iter107__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter107_to_t1_iter108__din),
    .fifo_st_0_full_n(from_t1_iter107_to_t1_iter108__full_n),
    .fifo_st_0_write(from_t1_iter107_to_t1_iter108__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_106
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_106__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_ld_0_s_dout(from_t1_iter107_to_t1_iter108__dout),
    .fifo_ld_0_peek_dout(from_t1_iter107_to_t1_iter108__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter107_to_t1_iter108__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter107_to_t1_iter108__empty_n),
    .fifo_ld_0_s_read(from_t1_iter107_to_t1_iter108__read),
    .fifo_ld_0_peek_read(),
    .fifo_st_0_din(from_t1_iter108_to_t0__din),
    .fifo_st_0_full_n(from_t1_iter108_to_t0__full_n),
    .fifo_st_0_write(from_t1_iter108_to_t0__write)
  );


  (* keep_hierarchy = "yes" *) Module2Func
  Module2Func_107
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module2Func_107__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .fifo_st_0_din(from_t0_to_t0_bank_1__din),
    .fifo_st_0_full_n(from_t0_to_t0_bank_1__full_n),
    .fifo_st_0_write(from_t0_to_t0_bank_1__write),
    .fifo_ld_0_s_dout(from_t1_iter108_to_t0__dout),
    .fifo_ld_0_peek_dout(from_t1_iter108_to_t0__dout),
    .fifo_ld_0_s_empty_n(from_t1_iter108_to_t0__empty_n),
    .fifo_ld_0_peek_empty_n(from_t1_iter108_to_t0__empty_n),
    .fifo_ld_0_s_read(from_t1_iter108_to_t0__read),
    .fifo_ld_0_peek_read()
  );


  (* keep_hierarchy = "yes" *) Module3Func
  Module3Func_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(Module3Func_0__ap_start),
    .ap_done(),
    .ap_idle(),
    .ap_ready(),
    .dram_t0_bank_1_fifo_din(bank_1_t0_buf__din),
    .dram_t0_bank_1_fifo_full_n(bank_1_t0_buf__full_n),
    .dram_t0_bank_1_fifo_write(bank_1_t0_buf__write),
    .fifo_ld_0_s_dout(from_t0_to_t0_bank_1__dout),
    .fifo_ld_0_peek_dout(from_t0_to_t0_bank_1__dout),
    .fifo_ld_0_s_empty_n(from_t0_to_t0_bank_1__empty_n),
    .fifo_ld_0_peek_empty_n(from_t0_to_t0_bank_1__empty_n),
    .fifo_ld_0_s_read(from_t0_to_t0_bank_1__read),
    .fifo_ld_0_peek_read()
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  bank_0_t1__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_bank_0_t1_ARADDR),
    .m_axi_ARBURST(m_axi_bank_0_t1_ARBURST),
    .m_axi_ARCACHE(m_axi_bank_0_t1_ARCACHE),
    .m_axi_ARID(m_axi_bank_0_t1_ARID),
    .m_axi_ARLEN(m_axi_bank_0_t1_ARLEN),
    .m_axi_ARLOCK(m_axi_bank_0_t1_ARLOCK),
    .m_axi_ARPROT(m_axi_bank_0_t1_ARPROT),
    .m_axi_ARQOS(m_axi_bank_0_t1_ARQOS),
    .m_axi_ARREADY(m_axi_bank_0_t1_ARREADY),
    .m_axi_ARSIZE(m_axi_bank_0_t1_ARSIZE),
    .m_axi_ARVALID(m_axi_bank_0_t1_ARVALID),
    .m_axi_AWADDR(m_axi_bank_0_t1_AWADDR),
    .m_axi_AWBURST(m_axi_bank_0_t1_AWBURST),
    .m_axi_AWCACHE(m_axi_bank_0_t1_AWCACHE),
    .m_axi_AWID(m_axi_bank_0_t1_AWID),
    .m_axi_AWLEN(m_axi_bank_0_t1_AWLEN),
    .m_axi_AWLOCK(m_axi_bank_0_t1_AWLOCK),
    .m_axi_AWPROT(m_axi_bank_0_t1_AWPROT),
    .m_axi_AWQOS(m_axi_bank_0_t1_AWQOS),
    .m_axi_AWREADY(m_axi_bank_0_t1_AWREADY),
    .m_axi_AWSIZE(m_axi_bank_0_t1_AWSIZE),
    .m_axi_AWVALID(m_axi_bank_0_t1_AWVALID),
    .m_axi_BID(m_axi_bank_0_t1_BID),
    .m_axi_BREADY(m_axi_bank_0_t1_BREADY),
    .m_axi_BRESP(m_axi_bank_0_t1_BRESP),
    .m_axi_BVALID(m_axi_bank_0_t1_BVALID),
    .m_axi_RDATA(m_axi_bank_0_t1_RDATA),
    .m_axi_RID(m_axi_bank_0_t1_RID),
    .m_axi_RLAST(m_axi_bank_0_t1_RLAST),
    .m_axi_RREADY(m_axi_bank_0_t1_RREADY),
    .m_axi_RRESP(m_axi_bank_0_t1_RRESP),
    .m_axi_RVALID(m_axi_bank_0_t1_RVALID),
    .m_axi_WDATA(m_axi_bank_0_t1_WDATA),
    .m_axi_WLAST(m_axi_bank_0_t1_WLAST),
    .m_axi_WREADY(m_axi_bank_0_t1_WREADY),
    .m_axi_WSTRB(m_axi_bank_0_t1_WSTRB),
    .m_axi_WVALID(m_axi_bank_0_t1_WVALID),
    .read_addr_din(bank_0_t1_read_addr__din),
    .read_addr_full_n(bank_0_t1_read_addr__full_n),
    .read_addr_write(bank_0_t1_read_addr__write),
    .read_data_dout(bank_0_t1_read_data__dout),
    .read_data_empty_n(bank_0_t1_read_data__empty_n),
    .read_data_read(bank_0_t1_read_data__read),
    .write_addr_din(bank_0_t1_write_addr__din),
    .write_addr_full_n(bank_0_t1_write_addr__full_n),
    .write_addr_write(bank_0_t1_write_addr__write),
    .write_data_din(bank_0_t1_write_data__din),
    .write_data_full_n(bank_0_t1_write_data__full_n),
    .write_data_write(bank_0_t1_write_data__write),
    .write_resp_dout(bank_0_t1_write_resp__dout),
    .write_resp_empty_n(bank_0_t1_write_resp__empty_n),
    .write_resp_read(bank_0_t1_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(512),
    .DataWidthBytesLog(6),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(15)
  )
  bank_1_t0__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_bank_1_t0_ARADDR),
    .m_axi_ARBURST(m_axi_bank_1_t0_ARBURST),
    .m_axi_ARCACHE(m_axi_bank_1_t0_ARCACHE),
    .m_axi_ARID(m_axi_bank_1_t0_ARID),
    .m_axi_ARLEN(m_axi_bank_1_t0_ARLEN),
    .m_axi_ARLOCK(m_axi_bank_1_t0_ARLOCK),
    .m_axi_ARPROT(m_axi_bank_1_t0_ARPROT),
    .m_axi_ARQOS(m_axi_bank_1_t0_ARQOS),
    .m_axi_ARREADY(m_axi_bank_1_t0_ARREADY),
    .m_axi_ARSIZE(m_axi_bank_1_t0_ARSIZE),
    .m_axi_ARVALID(m_axi_bank_1_t0_ARVALID),
    .m_axi_AWADDR(m_axi_bank_1_t0_AWADDR),
    .m_axi_AWBURST(m_axi_bank_1_t0_AWBURST),
    .m_axi_AWCACHE(m_axi_bank_1_t0_AWCACHE),
    .m_axi_AWID(m_axi_bank_1_t0_AWID),
    .m_axi_AWLEN(m_axi_bank_1_t0_AWLEN),
    .m_axi_AWLOCK(m_axi_bank_1_t0_AWLOCK),
    .m_axi_AWPROT(m_axi_bank_1_t0_AWPROT),
    .m_axi_AWQOS(m_axi_bank_1_t0_AWQOS),
    .m_axi_AWREADY(m_axi_bank_1_t0_AWREADY),
    .m_axi_AWSIZE(m_axi_bank_1_t0_AWSIZE),
    .m_axi_AWVALID(m_axi_bank_1_t0_AWVALID),
    .m_axi_BID(m_axi_bank_1_t0_BID),
    .m_axi_BREADY(m_axi_bank_1_t0_BREADY),
    .m_axi_BRESP(m_axi_bank_1_t0_BRESP),
    .m_axi_BVALID(m_axi_bank_1_t0_BVALID),
    .m_axi_RDATA(m_axi_bank_1_t0_RDATA),
    .m_axi_RID(m_axi_bank_1_t0_RID),
    .m_axi_RLAST(m_axi_bank_1_t0_RLAST),
    .m_axi_RREADY(m_axi_bank_1_t0_RREADY),
    .m_axi_RRESP(m_axi_bank_1_t0_RRESP),
    .m_axi_RVALID(m_axi_bank_1_t0_RVALID),
    .m_axi_WDATA(m_axi_bank_1_t0_WDATA),
    .m_axi_WLAST(m_axi_bank_1_t0_WLAST),
    .m_axi_WREADY(m_axi_bank_1_t0_WREADY),
    .m_axi_WSTRB(m_axi_bank_1_t0_WSTRB),
    .m_axi_WVALID(m_axi_bank_1_t0_WVALID),
    .read_addr_din(bank_1_t0_read_addr__din),
    .read_addr_full_n(bank_1_t0_read_addr__full_n),
    .read_addr_write(bank_1_t0_read_addr__write),
    .read_data_dout(bank_1_t0_read_data__dout),
    .read_data_empty_n(bank_1_t0_read_data__empty_n),
    .read_data_read(bank_1_t0_read_data__read),
    .write_addr_din(bank_1_t0_write_addr__din),
    .write_addr_full_n(bank_1_t0_write_addr__full_n),
    .write_addr_write(bank_1_t0_write_addr__write),
    .write_data_din(bank_1_t0_write_data__din),
    .write_data_full_n(bank_1_t0_write_data__full_n),
    .write_data_write(bank_1_t0_write_data__write),
    .write_resp_dout(bank_1_t0_write_resp__dout),
    .write_resp_empty_n(bank_1_t0_write_resp__empty_n),
    .write_resp_read(bank_1_t0_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) jacobi3d_kernel_fsm
  __tapa_fsm_unit
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(ap_start),
    .ap_done(ap_done),
    .ap_idle(ap_idle),
    .ap_ready(ap_ready),
    .bank_0_t1(bank_0_t1),
    .coalesced_data_num(coalesced_data_num),
    .bank_1_t0(bank_1_t0),
    .BurstRead_floatx16_0___bank_0_t1__q0(BurstRead_floatx16_0___bank_0_t1__q0),
    .BurstRead_floatx16_0___coalesced_data_num__q0(BurstRead_floatx16_0___coalesced_data_num__q0),
    .BurstRead_floatx16_0__ap_start(BurstRead_floatx16_0__ap_start),
    .BurstRead_floatx16_0__ap_ready(BurstRead_floatx16_0__ap_ready),
    .BurstRead_floatx16_0__ap_done(BurstRead_floatx16_0__ap_done),
    .BurstRead_floatx16_0__ap_idle(BurstRead_floatx16_0__ap_idle),
    .BurstWrite_floatx16_0___bank_1_t0__q0(BurstWrite_floatx16_0___bank_1_t0__q0),
    .BurstWrite_floatx16_0___coalesced_data_num__q0(BurstWrite_floatx16_0___coalesced_data_num__q0),
    .BurstWrite_floatx16_0__ap_start(BurstWrite_floatx16_0__ap_start),
    .BurstWrite_floatx16_0__ap_ready(BurstWrite_floatx16_0__ap_ready),
    .BurstWrite_floatx16_0__ap_done(BurstWrite_floatx16_0__ap_done),
    .BurstWrite_floatx16_0__ap_idle(BurstWrite_floatx16_0__ap_idle),
    .Module0Func_0__ap_start(Module0Func_0__ap_start),
    .Module1Func_0__ap_start(Module1Func_0__ap_start),
    .Module2Func_0__ap_start(Module2Func_0__ap_start),
    .Module2Func_1__ap_start(Module2Func_1__ap_start),
    .Module2Func_2__ap_start(Module2Func_2__ap_start),
    .Module2Func_3__ap_start(Module2Func_3__ap_start),
    .Module2Func_4__ap_start(Module2Func_4__ap_start),
    .Module2Func_5__ap_start(Module2Func_5__ap_start),
    .Module2Func_6__ap_start(Module2Func_6__ap_start),
    .Module2Func_7__ap_start(Module2Func_7__ap_start),
    .Module2Func_8__ap_start(Module2Func_8__ap_start),
    .Module2Func_9__ap_start(Module2Func_9__ap_start),
    .Module2Func_10__ap_start(Module2Func_10__ap_start),
    .Module2Func_11__ap_start(Module2Func_11__ap_start),
    .Module2Func_12__ap_start(Module2Func_12__ap_start),
    .Module2Func_13__ap_start(Module2Func_13__ap_start),
    .Module2Func_14__ap_start(Module2Func_14__ap_start),
    .Module2Func_15__ap_start(Module2Func_15__ap_start),
    .Module2Func_16__ap_start(Module2Func_16__ap_start),
    .Module2Func_17__ap_start(Module2Func_17__ap_start),
    .Module2Func_18__ap_start(Module2Func_18__ap_start),
    .Module2Func_19__ap_start(Module2Func_19__ap_start),
    .Module2Func_20__ap_start(Module2Func_20__ap_start),
    .Module2Func_21__ap_start(Module2Func_21__ap_start),
    .Module2Func_22__ap_start(Module2Func_22__ap_start),
    .Module2Func_23__ap_start(Module2Func_23__ap_start),
    .Module2Func_24__ap_start(Module2Func_24__ap_start),
    .Module2Func_25__ap_start(Module2Func_25__ap_start),
    .Module2Func_26__ap_start(Module2Func_26__ap_start),
    .Module2Func_27__ap_start(Module2Func_27__ap_start),
    .Module2Func_28__ap_start(Module2Func_28__ap_start),
    .Module2Func_29__ap_start(Module2Func_29__ap_start),
    .Module2Func_30__ap_start(Module2Func_30__ap_start),
    .Module2Func_31__ap_start(Module2Func_31__ap_start),
    .Module2Func_32__ap_start(Module2Func_32__ap_start),
    .Module2Func_33__ap_start(Module2Func_33__ap_start),
    .Module2Func_34__ap_start(Module2Func_34__ap_start),
    .Module2Func_35__ap_start(Module2Func_35__ap_start),
    .Module2Func_36__ap_start(Module2Func_36__ap_start),
    .Module2Func_37__ap_start(Module2Func_37__ap_start),
    .Module2Func_38__ap_start(Module2Func_38__ap_start),
    .Module2Func_39__ap_start(Module2Func_39__ap_start),
    .Module2Func_40__ap_start(Module2Func_40__ap_start),
    .Module2Func_41__ap_start(Module2Func_41__ap_start),
    .Module2Func_42__ap_start(Module2Func_42__ap_start),
    .Module2Func_43__ap_start(Module2Func_43__ap_start),
    .Module2Func_44__ap_start(Module2Func_44__ap_start),
    .Module2Func_45__ap_start(Module2Func_45__ap_start),
    .Module2Func_46__ap_start(Module2Func_46__ap_start),
    .Module2Func_47__ap_start(Module2Func_47__ap_start),
    .Module2Func_48__ap_start(Module2Func_48__ap_start),
    .Module2Func_49__ap_start(Module2Func_49__ap_start),
    .Module2Func_50__ap_start(Module2Func_50__ap_start),
    .Module2Func_51__ap_start(Module2Func_51__ap_start),
    .Module2Func_52__ap_start(Module2Func_52__ap_start),
    .Module2Func_53__ap_start(Module2Func_53__ap_start),
    .Module2Func_54__ap_start(Module2Func_54__ap_start),
    .Module2Func_55__ap_start(Module2Func_55__ap_start),
    .Module2Func_56__ap_start(Module2Func_56__ap_start),
    .Module2Func_57__ap_start(Module2Func_57__ap_start),
    .Module2Func_58__ap_start(Module2Func_58__ap_start),
    .Module2Func_59__ap_start(Module2Func_59__ap_start),
    .Module2Func_60__ap_start(Module2Func_60__ap_start),
    .Module2Func_61__ap_start(Module2Func_61__ap_start),
    .Module2Func_62__ap_start(Module2Func_62__ap_start),
    .Module2Func_63__ap_start(Module2Func_63__ap_start),
    .Module2Func_64__ap_start(Module2Func_64__ap_start),
    .Module2Func_65__ap_start(Module2Func_65__ap_start),
    .Module2Func_66__ap_start(Module2Func_66__ap_start),
    .Module2Func_67__ap_start(Module2Func_67__ap_start),
    .Module2Func_68__ap_start(Module2Func_68__ap_start),
    .Module2Func_69__ap_start(Module2Func_69__ap_start),
    .Module2Func_70__ap_start(Module2Func_70__ap_start),
    .Module2Func_71__ap_start(Module2Func_71__ap_start),
    .Module2Func_72__ap_start(Module2Func_72__ap_start),
    .Module2Func_73__ap_start(Module2Func_73__ap_start),
    .Module2Func_74__ap_start(Module2Func_74__ap_start),
    .Module2Func_75__ap_start(Module2Func_75__ap_start),
    .Module2Func_76__ap_start(Module2Func_76__ap_start),
    .Module2Func_77__ap_start(Module2Func_77__ap_start),
    .Module2Func_78__ap_start(Module2Func_78__ap_start),
    .Module2Func_79__ap_start(Module2Func_79__ap_start),
    .Module2Func_80__ap_start(Module2Func_80__ap_start),
    .Module2Func_81__ap_start(Module2Func_81__ap_start),
    .Module2Func_82__ap_start(Module2Func_82__ap_start),
    .Module2Func_83__ap_start(Module2Func_83__ap_start),
    .Module2Func_84__ap_start(Module2Func_84__ap_start),
    .Module2Func_85__ap_start(Module2Func_85__ap_start),
    .Module2Func_86__ap_start(Module2Func_86__ap_start),
    .Module2Func_87__ap_start(Module2Func_87__ap_start),
    .Module2Func_88__ap_start(Module2Func_88__ap_start),
    .Module2Func_89__ap_start(Module2Func_89__ap_start),
    .Module2Func_90__ap_start(Module2Func_90__ap_start),
    .Module2Func_91__ap_start(Module2Func_91__ap_start),
    .Module2Func_92__ap_start(Module2Func_92__ap_start),
    .Module2Func_93__ap_start(Module2Func_93__ap_start),
    .Module2Func_94__ap_start(Module2Func_94__ap_start),
    .Module2Func_95__ap_start(Module2Func_95__ap_start),
    .Module2Func_96__ap_start(Module2Func_96__ap_start),
    .Module2Func_97__ap_start(Module2Func_97__ap_start),
    .Module2Func_98__ap_start(Module2Func_98__ap_start),
    .Module2Func_99__ap_start(Module2Func_99__ap_start),
    .Module2Func_100__ap_start(Module2Func_100__ap_start),
    .Module2Func_101__ap_start(Module2Func_101__ap_start),
    .Module2Func_102__ap_start(Module2Func_102__ap_start),
    .Module2Func_103__ap_start(Module2Func_103__ap_start),
    .Module2Func_104__ap_start(Module2Func_104__ap_start),
    .Module2Func_105__ap_start(Module2Func_105__ap_start),
    .Module2Func_106__ap_start(Module2Func_106__ap_start),
    .Module2Func_107__ap_start(Module2Func_107__ap_start),
    .Module3Func_0__ap_start(Module3Func_0__ap_start)
  );

  assign ap_rst_n_inv = (~ap_rst_n);

endmodule

