// This stub module is excluded from exporting