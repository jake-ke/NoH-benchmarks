`timescale 1 ns / 1 ps 

(* CORE_GENERATION_INFO = "kernel0_kernel0,hls_ip_2023_2_2,{HLS_INPUT_TYPE=cxx,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=0,HLS_INPUT_PART=xcvp1802-lsvc4072-2MP-e-S,HLS_INPUT_CLOCK=3.330000,HLS_INPUT_ARCH=others,HLS_SYN_CLOCK=1.000000,HLS_SYN_LAT=0,HLS_SYN_TPT=none,HLS_SYN_MEM=0,HLS_SYN_DSP=0,HLS_SYN_FF=246,HLS_SYN_LUT=424,HLS_VERSION=2023_2_2}" *)


module kernel0
(
  s_axi_control_AWVALID,
  s_axi_control_AWREADY,
  s_axi_control_AWADDR,
  s_axi_control_WVALID,
  s_axi_control_WREADY,
  s_axi_control_WDATA,
  s_axi_control_WSTRB,
  s_axi_control_ARVALID,
  s_axi_control_ARREADY,
  s_axi_control_ARADDR,
  s_axi_control_RVALID,
  s_axi_control_RREADY,
  s_axi_control_RDATA,
  s_axi_control_RRESP,
  s_axi_control_BVALID,
  s_axi_control_BREADY,
  s_axi_control_BRESP,
  ap_clk,
  ap_rst_n,
  interrupt,
  m_axi_A_ARADDR,
  m_axi_A_ARBURST,
  m_axi_A_ARCACHE,
  m_axi_A_ARID,
  m_axi_A_ARLEN,
  m_axi_A_ARLOCK,
  m_axi_A_ARPROT,
  m_axi_A_ARQOS,
  m_axi_A_ARREADY,
  m_axi_A_ARSIZE,
  m_axi_A_ARVALID,
  m_axi_A_AWADDR,
  m_axi_A_AWBURST,
  m_axi_A_AWCACHE,
  m_axi_A_AWID,
  m_axi_A_AWLEN,
  m_axi_A_AWLOCK,
  m_axi_A_AWPROT,
  m_axi_A_AWQOS,
  m_axi_A_AWREADY,
  m_axi_A_AWSIZE,
  m_axi_A_AWVALID,
  m_axi_A_BID,
  m_axi_A_BREADY,
  m_axi_A_BRESP,
  m_axi_A_BVALID,
  m_axi_A_RDATA,
  m_axi_A_RID,
  m_axi_A_RLAST,
  m_axi_A_RREADY,
  m_axi_A_RRESP,
  m_axi_A_RVALID,
  m_axi_A_WDATA,
  m_axi_A_WLAST,
  m_axi_A_WREADY,
  m_axi_A_WSTRB,
  m_axi_A_WVALID,
  m_axi_B_ARADDR,
  m_axi_B_ARBURST,
  m_axi_B_ARCACHE,
  m_axi_B_ARID,
  m_axi_B_ARLEN,
  m_axi_B_ARLOCK,
  m_axi_B_ARPROT,
  m_axi_B_ARQOS,
  m_axi_B_ARREADY,
  m_axi_B_ARSIZE,
  m_axi_B_ARVALID,
  m_axi_B_AWADDR,
  m_axi_B_AWBURST,
  m_axi_B_AWCACHE,
  m_axi_B_AWID,
  m_axi_B_AWLEN,
  m_axi_B_AWLOCK,
  m_axi_B_AWPROT,
  m_axi_B_AWQOS,
  m_axi_B_AWREADY,
  m_axi_B_AWSIZE,
  m_axi_B_AWVALID,
  m_axi_B_BID,
  m_axi_B_BREADY,
  m_axi_B_BRESP,
  m_axi_B_BVALID,
  m_axi_B_RDATA,
  m_axi_B_RID,
  m_axi_B_RLAST,
  m_axi_B_RREADY,
  m_axi_B_RRESP,
  m_axi_B_RVALID,
  m_axi_B_WDATA,
  m_axi_B_WLAST,
  m_axi_B_WREADY,
  m_axi_B_WSTRB,
  m_axi_B_WVALID,
  m_axi_C_ARADDR,
  m_axi_C_ARBURST,
  m_axi_C_ARCACHE,
  m_axi_C_ARID,
  m_axi_C_ARLEN,
  m_axi_C_ARLOCK,
  m_axi_C_ARPROT,
  m_axi_C_ARQOS,
  m_axi_C_ARREADY,
  m_axi_C_ARSIZE,
  m_axi_C_ARVALID,
  m_axi_C_AWADDR,
  m_axi_C_AWBURST,
  m_axi_C_AWCACHE,
  m_axi_C_AWID,
  m_axi_C_AWLEN,
  m_axi_C_AWLOCK,
  m_axi_C_AWPROT,
  m_axi_C_AWQOS,
  m_axi_C_AWREADY,
  m_axi_C_AWSIZE,
  m_axi_C_AWVALID,
  m_axi_C_BID,
  m_axi_C_BREADY,
  m_axi_C_BRESP,
  m_axi_C_BVALID,
  m_axi_C_RDATA,
  m_axi_C_RID,
  m_axi_C_RLAST,
  m_axi_C_RREADY,
  m_axi_C_RRESP,
  m_axi_C_RVALID,
  m_axi_C_WDATA,
  m_axi_C_WLAST,
  m_axi_C_WREADY,
  m_axi_C_WSTRB,
  m_axi_C_WVALID
);

  parameter C_S_AXI_CONTROL_DATA_WIDTH = 32;
  parameter C_S_AXI_CONTROL_ADDR_WIDTH = 6;
  parameter C_S_AXI_DATA_WIDTH = 32;
  parameter C_S_AXI_CONTROL_WSTRB_WIDTH = 32 / 8;
  parameter C_S_AXI_WSTRB_WIDTH = 32 / 8;
  (* RS_HS = "s_axi_control_AW.valid" *)input s_axi_control_AWVALID;
  (* RS_HS = "s_axi_control_AW.ready" *)output s_axi_control_AWREADY;
  (* RS_HS = "s_axi_control_AW.data" *)input [C_S_AXI_CONTROL_ADDR_WIDTH-1:0] s_axi_control_AWADDR;
  (* RS_HS = "s_axi_control_W.valid" *)input s_axi_control_WVALID;
  (* RS_HS = "s_axi_control_W.ready" *)output s_axi_control_WREADY;
  (* RS_HS = "s_axi_control_W.data" *)input [C_S_AXI_CONTROL_DATA_WIDTH-1:0] s_axi_control_WDATA;
  (* RS_HS = "s_axi_control_W.data" *)input [C_S_AXI_CONTROL_WSTRB_WIDTH-1:0] s_axi_control_WSTRB;
  (* RS_HS = "s_axi_control_AR.valid" *)input s_axi_control_ARVALID;
  (* RS_HS = "s_axi_control_AR.ready" *)output s_axi_control_ARREADY;
  (* RS_HS = "s_axi_control_AR.data" *)input [C_S_AXI_CONTROL_ADDR_WIDTH-1:0] s_axi_control_ARADDR;
  (* RS_HS = "s_axi_control_R.valid" *)output s_axi_control_RVALID;
  (* RS_HS = "s_axi_control_R.ready" *)input s_axi_control_RREADY;
  (* RS_HS = "s_axi_control_R.data" *)output [C_S_AXI_CONTROL_DATA_WIDTH-1:0] s_axi_control_RDATA;
  (* RS_HS = "s_axi_control_R.data" *)output [1:0] s_axi_control_RRESP;
  (* RS_HS = "s_axi_control_B.valid" *)output s_axi_control_BVALID;
  (* RS_HS = "s_axi_control_B.ready" *)input s_axi_control_BREADY;
  (* RS_HS = "s_axi_control_B.data" *)output [1:0] s_axi_control_BRESP;
  (* RS_CLK *)input ap_clk;
  (* RS_RST = "ff" *)input ap_rst_n;
  (* RS_FF = "interrupt" *)output interrupt;
  (* RS_HS = "m_axi_A_AR.data" *)output [63:0] m_axi_A_ARADDR;
  (* RS_HS = "m_axi_A_AR.data" *)output [1:0] m_axi_A_ARBURST;
  (* RS_HS = "m_axi_A_AR.data" *)output [3:0] m_axi_A_ARCACHE;
  (* RS_HS = "m_axi_A_AR.data" *)output [0:0] m_axi_A_ARID;
  (* RS_HS = "m_axi_A_AR.data" *)output [7:0] m_axi_A_ARLEN;
  (* RS_HS = "m_axi_A_AR.data" *)output m_axi_A_ARLOCK;
  (* RS_HS = "m_axi_A_AR.data" *)output [2:0] m_axi_A_ARPROT;
  (* RS_HS = "m_axi_A_AR.data" *)output [3:0] m_axi_A_ARQOS;
  (* RS_HS = "m_axi_A_AR.ready" *)input m_axi_A_ARREADY;
  (* RS_HS = "m_axi_A_AR.data" *)output [2:0] m_axi_A_ARSIZE;
  (* RS_HS = "m_axi_A_AR.valid" *)output m_axi_A_ARVALID;
  (* RS_HS = "m_axi_A_AW.data" *)output [63:0] m_axi_A_AWADDR;
  (* RS_HS = "m_axi_A_AW.data" *)output [1:0] m_axi_A_AWBURST;
  (* RS_HS = "m_axi_A_AW.data" *)output [3:0] m_axi_A_AWCACHE;
  (* RS_HS = "m_axi_A_AW.data" *)output [0:0] m_axi_A_AWID;
  (* RS_HS = "m_axi_A_AW.data" *)output [7:0] m_axi_A_AWLEN;
  (* RS_HS = "m_axi_A_AW.data" *)output m_axi_A_AWLOCK;
  (* RS_HS = "m_axi_A_AW.data" *)output [2:0] m_axi_A_AWPROT;
  (* RS_HS = "m_axi_A_AW.data" *)output [3:0] m_axi_A_AWQOS;
  (* RS_HS = "m_axi_A_AW.ready" *)input m_axi_A_AWREADY;
  (* RS_HS = "m_axi_A_AW.data" *)output [2:0] m_axi_A_AWSIZE;
  (* RS_HS = "m_axi_A_AW.valid" *)output m_axi_A_AWVALID;
  (* RS_HS = "m_axi_A_B.data" *)input [0:0] m_axi_A_BID;
  (* RS_HS = "m_axi_A_B.ready" *)output m_axi_A_BREADY;
  (* RS_HS = "m_axi_A_B.data" *)input [1:0] m_axi_A_BRESP;
  (* RS_HS = "m_axi_A_B.valid" *)input m_axi_A_BVALID;
  (* RS_HS = "m_axi_A_R.data" *)input [511:0] m_axi_A_RDATA;
  (* RS_HS = "m_axi_A_R.data" *)input [0:0] m_axi_A_RID;
  (* RS_HS = "m_axi_A_R.data" *)input m_axi_A_RLAST;
  (* RS_HS = "m_axi_A_R.ready" *)output m_axi_A_RREADY;
  (* RS_HS = "m_axi_A_R.data" *)input [1:0] m_axi_A_RRESP;
  (* RS_HS = "m_axi_A_R.valid" *)input m_axi_A_RVALID;
  (* RS_HS = "m_axi_A_W.data" *)output [511:0] m_axi_A_WDATA;
  (* RS_HS = "m_axi_A_W.data" *)output m_axi_A_WLAST;
  (* RS_HS = "m_axi_A_W.ready" *)input m_axi_A_WREADY;
  (* RS_HS = "m_axi_A_W.data" *)output [63:0] m_axi_A_WSTRB;
  (* RS_HS = "m_axi_A_W.valid" *)output m_axi_A_WVALID;
  (* RS_HS = "m_axi_B_AR.data" *)output [63:0] m_axi_B_ARADDR;
  (* RS_HS = "m_axi_B_AR.data" *)output [1:0] m_axi_B_ARBURST;
  (* RS_HS = "m_axi_B_AR.data" *)output [3:0] m_axi_B_ARCACHE;
  (* RS_HS = "m_axi_B_AR.data" *)output [0:0] m_axi_B_ARID;
  (* RS_HS = "m_axi_B_AR.data" *)output [7:0] m_axi_B_ARLEN;
  (* RS_HS = "m_axi_B_AR.data" *)output m_axi_B_ARLOCK;
  (* RS_HS = "m_axi_B_AR.data" *)output [2:0] m_axi_B_ARPROT;
  (* RS_HS = "m_axi_B_AR.data" *)output [3:0] m_axi_B_ARQOS;
  (* RS_HS = "m_axi_B_AR.ready" *)input m_axi_B_ARREADY;
  (* RS_HS = "m_axi_B_AR.data" *)output [2:0] m_axi_B_ARSIZE;
  (* RS_HS = "m_axi_B_AR.valid" *)output m_axi_B_ARVALID;
  (* RS_HS = "m_axi_B_AW.data" *)output [63:0] m_axi_B_AWADDR;
  (* RS_HS = "m_axi_B_AW.data" *)output [1:0] m_axi_B_AWBURST;
  (* RS_HS = "m_axi_B_AW.data" *)output [3:0] m_axi_B_AWCACHE;
  (* RS_HS = "m_axi_B_AW.data" *)output [0:0] m_axi_B_AWID;
  (* RS_HS = "m_axi_B_AW.data" *)output [7:0] m_axi_B_AWLEN;
  (* RS_HS = "m_axi_B_AW.data" *)output m_axi_B_AWLOCK;
  (* RS_HS = "m_axi_B_AW.data" *)output [2:0] m_axi_B_AWPROT;
  (* RS_HS = "m_axi_B_AW.data" *)output [3:0] m_axi_B_AWQOS;
  (* RS_HS = "m_axi_B_AW.ready" *)input m_axi_B_AWREADY;
  (* RS_HS = "m_axi_B_AW.data" *)output [2:0] m_axi_B_AWSIZE;
  (* RS_HS = "m_axi_B_AW.valid" *)output m_axi_B_AWVALID;
  (* RS_HS = "m_axi_B_B.data" *)input [0:0] m_axi_B_BID;
  (* RS_HS = "m_axi_B_B.ready" *)output m_axi_B_BREADY;
  (* RS_HS = "m_axi_B_B.data" *)input [1:0] m_axi_B_BRESP;
  (* RS_HS = "m_axi_B_B.valid" *)input m_axi_B_BVALID;
  (* RS_HS = "m_axi_B_R.data" *)input [511:0] m_axi_B_RDATA;
  (* RS_HS = "m_axi_B_R.data" *)input [0:0] m_axi_B_RID;
  (* RS_HS = "m_axi_B_R.data" *)input m_axi_B_RLAST;
  (* RS_HS = "m_axi_B_R.ready" *)output m_axi_B_RREADY;
  (* RS_HS = "m_axi_B_R.data" *)input [1:0] m_axi_B_RRESP;
  (* RS_HS = "m_axi_B_R.valid" *)input m_axi_B_RVALID;
  (* RS_HS = "m_axi_B_W.data" *)output [511:0] m_axi_B_WDATA;
  (* RS_HS = "m_axi_B_W.data" *)output m_axi_B_WLAST;
  (* RS_HS = "m_axi_B_W.ready" *)input m_axi_B_WREADY;
  (* RS_HS = "m_axi_B_W.data" *)output [63:0] m_axi_B_WSTRB;
  (* RS_HS = "m_axi_B_W.valid" *)output m_axi_B_WVALID;
  (* RS_HS = "m_axi_C_AR.data" *)output [63:0] m_axi_C_ARADDR;
  (* RS_HS = "m_axi_C_AR.data" *)output [1:0] m_axi_C_ARBURST;
  (* RS_HS = "m_axi_C_AR.data" *)output [3:0] m_axi_C_ARCACHE;
  (* RS_HS = "m_axi_C_AR.data" *)output [0:0] m_axi_C_ARID;
  (* RS_HS = "m_axi_C_AR.data" *)output [7:0] m_axi_C_ARLEN;
  (* RS_HS = "m_axi_C_AR.data" *)output m_axi_C_ARLOCK;
  (* RS_HS = "m_axi_C_AR.data" *)output [2:0] m_axi_C_ARPROT;
  (* RS_HS = "m_axi_C_AR.data" *)output [3:0] m_axi_C_ARQOS;
  (* RS_HS = "m_axi_C_AR.ready" *)input m_axi_C_ARREADY;
  (* RS_HS = "m_axi_C_AR.data" *)output [2:0] m_axi_C_ARSIZE;
  (* RS_HS = "m_axi_C_AR.valid" *)output m_axi_C_ARVALID;
  (* RS_HS = "m_axi_C_AW.data" *)output [63:0] m_axi_C_AWADDR;
  (* RS_HS = "m_axi_C_AW.data" *)output [1:0] m_axi_C_AWBURST;
  (* RS_HS = "m_axi_C_AW.data" *)output [3:0] m_axi_C_AWCACHE;
  (* RS_HS = "m_axi_C_AW.data" *)output [0:0] m_axi_C_AWID;
  (* RS_HS = "m_axi_C_AW.data" *)output [7:0] m_axi_C_AWLEN;
  (* RS_HS = "m_axi_C_AW.data" *)output m_axi_C_AWLOCK;
  (* RS_HS = "m_axi_C_AW.data" *)output [2:0] m_axi_C_AWPROT;
  (* RS_HS = "m_axi_C_AW.data" *)output [3:0] m_axi_C_AWQOS;
  (* RS_HS = "m_axi_C_AW.ready" *)input m_axi_C_AWREADY;
  (* RS_HS = "m_axi_C_AW.data" *)output [2:0] m_axi_C_AWSIZE;
  (* RS_HS = "m_axi_C_AW.valid" *)output m_axi_C_AWVALID;
  (* RS_HS = "m_axi_C_B.data" *)input [0:0] m_axi_C_BID;
  (* RS_HS = "m_axi_C_B.ready" *)output m_axi_C_BREADY;
  (* RS_HS = "m_axi_C_B.data" *)input [1:0] m_axi_C_BRESP;
  (* RS_HS = "m_axi_C_B.valid" *)input m_axi_C_BVALID;
  (* RS_HS = "m_axi_C_R.data" *)input [511:0] m_axi_C_RDATA;
  (* RS_HS = "m_axi_C_R.data" *)input [0:0] m_axi_C_RID;
  (* RS_HS = "m_axi_C_R.data" *)input m_axi_C_RLAST;
  (* RS_HS = "m_axi_C_R.ready" *)output m_axi_C_RREADY;
  (* RS_HS = "m_axi_C_R.data" *)input [1:0] m_axi_C_RRESP;
  (* RS_HS = "m_axi_C_R.valid" *)input m_axi_C_RVALID;
  (* RS_HS = "m_axi_C_W.data" *)output [511:0] m_axi_C_WDATA;
  (* RS_HS = "m_axi_C_W.data" *)output m_axi_C_WLAST;
  (* RS_HS = "m_axi_C_W.ready" *)input m_axi_C_WREADY;
  (* RS_HS = "m_axi_C_W.data" *)output [63:0] m_axi_C_WSTRB;
  (* RS_HS = "m_axi_C_W.valid" *)output m_axi_C_WVALID;
  wire ap_start;
  wire [63:0] A;
  wire [63:0] B;
  wire [63:0] C;
  wire [512:0] fifo_A_A_IO_L2_in_0__dout;
  wire fifo_A_A_IO_L2_in_0__empty_n;
  wire fifo_A_A_IO_L2_in_0__read;
  wire [512:0] fifo_A_A_IO_L2_in_0__din;
  wire fifo_A_A_IO_L2_in_0__full_n;
  wire fifo_A_A_IO_L2_in_0__write;
  wire [512:0] fifo_A_A_IO_L2_in_1__dout;
  wire fifo_A_A_IO_L2_in_1__empty_n;
  wire fifo_A_A_IO_L2_in_1__read;
  wire [512:0] fifo_A_A_IO_L2_in_1__din;
  wire fifo_A_A_IO_L2_in_1__full_n;
  wire fifo_A_A_IO_L2_in_1__write;
  wire [512:0] fifo_A_A_IO_L2_in_10__dout;
  wire fifo_A_A_IO_L2_in_10__empty_n;
  wire fifo_A_A_IO_L2_in_10__read;
  wire [512:0] fifo_A_A_IO_L2_in_10__din;
  wire fifo_A_A_IO_L2_in_10__full_n;
  wire fifo_A_A_IO_L2_in_10__write;
  wire [512:0] fifo_A_A_IO_L2_in_11__dout;
  wire fifo_A_A_IO_L2_in_11__empty_n;
  wire fifo_A_A_IO_L2_in_11__read;
  wire [512:0] fifo_A_A_IO_L2_in_11__din;
  wire fifo_A_A_IO_L2_in_11__full_n;
  wire fifo_A_A_IO_L2_in_11__write;
  wire [512:0] fifo_A_A_IO_L2_in_12__dout;
  wire fifo_A_A_IO_L2_in_12__empty_n;
  wire fifo_A_A_IO_L2_in_12__read;
  wire [512:0] fifo_A_A_IO_L2_in_12__din;
  wire fifo_A_A_IO_L2_in_12__full_n;
  wire fifo_A_A_IO_L2_in_12__write;
  wire [512:0] fifo_A_A_IO_L2_in_13__dout;
  wire fifo_A_A_IO_L2_in_13__empty_n;
  wire fifo_A_A_IO_L2_in_13__read;
  wire [512:0] fifo_A_A_IO_L2_in_13__din;
  wire fifo_A_A_IO_L2_in_13__full_n;
  wire fifo_A_A_IO_L2_in_13__write;
  wire [512:0] fifo_A_A_IO_L2_in_14__dout;
  wire fifo_A_A_IO_L2_in_14__empty_n;
  wire fifo_A_A_IO_L2_in_14__read;
  wire [512:0] fifo_A_A_IO_L2_in_14__din;
  wire fifo_A_A_IO_L2_in_14__full_n;
  wire fifo_A_A_IO_L2_in_14__write;
  wire [512:0] fifo_A_A_IO_L2_in_15__dout;
  wire fifo_A_A_IO_L2_in_15__empty_n;
  wire fifo_A_A_IO_L2_in_15__read;
  wire [512:0] fifo_A_A_IO_L2_in_15__din;
  wire fifo_A_A_IO_L2_in_15__full_n;
  wire fifo_A_A_IO_L2_in_15__write;
  wire [512:0] fifo_A_A_IO_L2_in_16__dout;
  wire fifo_A_A_IO_L2_in_16__empty_n;
  wire fifo_A_A_IO_L2_in_16__read;
  wire [512:0] fifo_A_A_IO_L2_in_16__din;
  wire fifo_A_A_IO_L2_in_16__full_n;
  wire fifo_A_A_IO_L2_in_16__write;
  wire [512:0] fifo_A_A_IO_L2_in_17__dout;
  wire fifo_A_A_IO_L2_in_17__empty_n;
  wire fifo_A_A_IO_L2_in_17__read;
  wire [512:0] fifo_A_A_IO_L2_in_17__din;
  wire fifo_A_A_IO_L2_in_17__full_n;
  wire fifo_A_A_IO_L2_in_17__write;
  wire [512:0] fifo_A_A_IO_L2_in_2__dout;
  wire fifo_A_A_IO_L2_in_2__empty_n;
  wire fifo_A_A_IO_L2_in_2__read;
  wire [512:0] fifo_A_A_IO_L2_in_2__din;
  wire fifo_A_A_IO_L2_in_2__full_n;
  wire fifo_A_A_IO_L2_in_2__write;
  wire [512:0] fifo_A_A_IO_L2_in_3__dout;
  wire fifo_A_A_IO_L2_in_3__empty_n;
  wire fifo_A_A_IO_L2_in_3__read;
  wire [512:0] fifo_A_A_IO_L2_in_3__din;
  wire fifo_A_A_IO_L2_in_3__full_n;
  wire fifo_A_A_IO_L2_in_3__write;
  wire [512:0] fifo_A_A_IO_L2_in_4__dout;
  wire fifo_A_A_IO_L2_in_4__empty_n;
  wire fifo_A_A_IO_L2_in_4__read;
  wire [512:0] fifo_A_A_IO_L2_in_4__din;
  wire fifo_A_A_IO_L2_in_4__full_n;
  wire fifo_A_A_IO_L2_in_4__write;
  wire [512:0] fifo_A_A_IO_L2_in_5__dout;
  wire fifo_A_A_IO_L2_in_5__empty_n;
  wire fifo_A_A_IO_L2_in_5__read;
  wire [512:0] fifo_A_A_IO_L2_in_5__din;
  wire fifo_A_A_IO_L2_in_5__full_n;
  wire fifo_A_A_IO_L2_in_5__write;
  wire [512:0] fifo_A_A_IO_L2_in_6__dout;
  wire fifo_A_A_IO_L2_in_6__empty_n;
  wire fifo_A_A_IO_L2_in_6__read;
  wire [512:0] fifo_A_A_IO_L2_in_6__din;
  wire fifo_A_A_IO_L2_in_6__full_n;
  wire fifo_A_A_IO_L2_in_6__write;
  wire [512:0] fifo_A_A_IO_L2_in_7__dout;
  wire fifo_A_A_IO_L2_in_7__empty_n;
  wire fifo_A_A_IO_L2_in_7__read;
  wire [512:0] fifo_A_A_IO_L2_in_7__din;
  wire fifo_A_A_IO_L2_in_7__full_n;
  wire fifo_A_A_IO_L2_in_7__write;
  wire [512:0] fifo_A_A_IO_L2_in_8__dout;
  wire fifo_A_A_IO_L2_in_8__empty_n;
  wire fifo_A_A_IO_L2_in_8__read;
  wire [512:0] fifo_A_A_IO_L2_in_8__din;
  wire fifo_A_A_IO_L2_in_8__full_n;
  wire fifo_A_A_IO_L2_in_8__write;
  wire [512:0] fifo_A_A_IO_L2_in_9__dout;
  wire fifo_A_A_IO_L2_in_9__empty_n;
  wire fifo_A_A_IO_L2_in_9__read;
  wire [512:0] fifo_A_A_IO_L2_in_9__din;
  wire fifo_A_A_IO_L2_in_9__full_n;
  wire fifo_A_A_IO_L2_in_9__write;
  wire [512:0] fifo_A_A_IO_L3_in_serialize__dout;
  wire fifo_A_A_IO_L3_in_serialize__empty_n;
  wire fifo_A_A_IO_L3_in_serialize__read;
  wire [512:0] fifo_A_A_IO_L3_in_serialize__din;
  wire fifo_A_A_IO_L3_in_serialize__full_n;
  wire fifo_A_A_IO_L3_in_serialize__write;
  wire [512:0] fifo_A_PE_0_0__dout;
  wire fifo_A_PE_0_0__empty_n;
  wire fifo_A_PE_0_0__read;
  wire [512:0] fifo_A_PE_0_0__din;
  wire fifo_A_PE_0_0__full_n;
  wire fifo_A_PE_0_0__write;
  wire [512:0] fifo_A_PE_0_1__dout;
  wire fifo_A_PE_0_1__empty_n;
  wire fifo_A_PE_0_1__read;
  wire [512:0] fifo_A_PE_0_1__din;
  wire fifo_A_PE_0_1__full_n;
  wire fifo_A_PE_0_1__write;
  wire [512:0] fifo_A_PE_0_10__dout;
  wire fifo_A_PE_0_10__empty_n;
  wire fifo_A_PE_0_10__read;
  wire [512:0] fifo_A_PE_0_10__din;
  wire fifo_A_PE_0_10__full_n;
  wire fifo_A_PE_0_10__write;
  wire [512:0] fifo_A_PE_0_11__dout;
  wire fifo_A_PE_0_11__empty_n;
  wire fifo_A_PE_0_11__read;
  wire [512:0] fifo_A_PE_0_11__din;
  wire fifo_A_PE_0_11__full_n;
  wire fifo_A_PE_0_11__write;
  wire [512:0] fifo_A_PE_0_12__dout;
  wire fifo_A_PE_0_12__empty_n;
  wire fifo_A_PE_0_12__read;
  wire [512:0] fifo_A_PE_0_12__din;
  wire fifo_A_PE_0_12__full_n;
  wire fifo_A_PE_0_12__write;
  wire [512:0] fifo_A_PE_0_13__dout;
  wire fifo_A_PE_0_13__empty_n;
  wire fifo_A_PE_0_13__read;
  wire [512:0] fifo_A_PE_0_13__din;
  wire fifo_A_PE_0_13__full_n;
  wire fifo_A_PE_0_13__write;
  wire [512:0] fifo_A_PE_0_14__dout;
  wire fifo_A_PE_0_14__empty_n;
  wire fifo_A_PE_0_14__read;
  wire [512:0] fifo_A_PE_0_14__din;
  wire fifo_A_PE_0_14__full_n;
  wire fifo_A_PE_0_14__write;
  wire [512:0] fifo_A_PE_0_15__dout;
  wire fifo_A_PE_0_15__empty_n;
  wire fifo_A_PE_0_15__read;
  wire [512:0] fifo_A_PE_0_15__din;
  wire fifo_A_PE_0_15__full_n;
  wire fifo_A_PE_0_15__write;
  wire [512:0] fifo_A_PE_0_16__dout;
  wire fifo_A_PE_0_16__empty_n;
  wire fifo_A_PE_0_16__read;
  wire [512:0] fifo_A_PE_0_16__din;
  wire fifo_A_PE_0_16__full_n;
  wire fifo_A_PE_0_16__write;
  wire [512:0] fifo_A_PE_0_17__dout;
  wire fifo_A_PE_0_17__empty_n;
  wire fifo_A_PE_0_17__read;
  wire [512:0] fifo_A_PE_0_17__din;
  wire fifo_A_PE_0_17__full_n;
  wire fifo_A_PE_0_17__write;
  wire [512:0] fifo_A_PE_0_2__dout;
  wire fifo_A_PE_0_2__empty_n;
  wire fifo_A_PE_0_2__read;
  wire [512:0] fifo_A_PE_0_2__din;
  wire fifo_A_PE_0_2__full_n;
  wire fifo_A_PE_0_2__write;
  wire [512:0] fifo_A_PE_0_3__dout;
  wire fifo_A_PE_0_3__empty_n;
  wire fifo_A_PE_0_3__read;
  wire [512:0] fifo_A_PE_0_3__din;
  wire fifo_A_PE_0_3__full_n;
  wire fifo_A_PE_0_3__write;
  wire [512:0] fifo_A_PE_0_4__dout;
  wire fifo_A_PE_0_4__empty_n;
  wire fifo_A_PE_0_4__read;
  wire [512:0] fifo_A_PE_0_4__din;
  wire fifo_A_PE_0_4__full_n;
  wire fifo_A_PE_0_4__write;
  wire [512:0] fifo_A_PE_0_5__dout;
  wire fifo_A_PE_0_5__empty_n;
  wire fifo_A_PE_0_5__read;
  wire [512:0] fifo_A_PE_0_5__din;
  wire fifo_A_PE_0_5__full_n;
  wire fifo_A_PE_0_5__write;
  wire [512:0] fifo_A_PE_0_6__dout;
  wire fifo_A_PE_0_6__empty_n;
  wire fifo_A_PE_0_6__read;
  wire [512:0] fifo_A_PE_0_6__din;
  wire fifo_A_PE_0_6__full_n;
  wire fifo_A_PE_0_6__write;
  wire [512:0] fifo_A_PE_0_7__dout;
  wire fifo_A_PE_0_7__empty_n;
  wire fifo_A_PE_0_7__read;
  wire [512:0] fifo_A_PE_0_7__din;
  wire fifo_A_PE_0_7__full_n;
  wire fifo_A_PE_0_7__write;
  wire [512:0] fifo_A_PE_0_8__dout;
  wire fifo_A_PE_0_8__empty_n;
  wire fifo_A_PE_0_8__read;
  wire [512:0] fifo_A_PE_0_8__din;
  wire fifo_A_PE_0_8__full_n;
  wire fifo_A_PE_0_8__write;
  wire [512:0] fifo_A_PE_0_9__dout;
  wire fifo_A_PE_0_9__empty_n;
  wire fifo_A_PE_0_9__read;
  wire [512:0] fifo_A_PE_0_9__din;
  wire fifo_A_PE_0_9__full_n;
  wire fifo_A_PE_0_9__write;
  wire [512:0] fifo_A_PE_10_0__dout;
  wire fifo_A_PE_10_0__empty_n;
  wire fifo_A_PE_10_0__read;
  wire [512:0] fifo_A_PE_10_0__din;
  wire fifo_A_PE_10_0__full_n;
  wire fifo_A_PE_10_0__write;
  wire [512:0] fifo_A_PE_10_1__dout;
  wire fifo_A_PE_10_1__empty_n;
  wire fifo_A_PE_10_1__read;
  wire [512:0] fifo_A_PE_10_1__din;
  wire fifo_A_PE_10_1__full_n;
  wire fifo_A_PE_10_1__write;
  wire [512:0] fifo_A_PE_10_10__dout;
  wire fifo_A_PE_10_10__empty_n;
  wire fifo_A_PE_10_10__read;
  wire [512:0] fifo_A_PE_10_10__din;
  wire fifo_A_PE_10_10__full_n;
  wire fifo_A_PE_10_10__write;
  wire [512:0] fifo_A_PE_10_11__dout;
  wire fifo_A_PE_10_11__empty_n;
  wire fifo_A_PE_10_11__read;
  wire [512:0] fifo_A_PE_10_11__din;
  wire fifo_A_PE_10_11__full_n;
  wire fifo_A_PE_10_11__write;
  wire [512:0] fifo_A_PE_10_12__dout;
  wire fifo_A_PE_10_12__empty_n;
  wire fifo_A_PE_10_12__read;
  wire [512:0] fifo_A_PE_10_12__din;
  wire fifo_A_PE_10_12__full_n;
  wire fifo_A_PE_10_12__write;
  wire [512:0] fifo_A_PE_10_13__dout;
  wire fifo_A_PE_10_13__empty_n;
  wire fifo_A_PE_10_13__read;
  wire [512:0] fifo_A_PE_10_13__din;
  wire fifo_A_PE_10_13__full_n;
  wire fifo_A_PE_10_13__write;
  wire [512:0] fifo_A_PE_10_14__dout;
  wire fifo_A_PE_10_14__empty_n;
  wire fifo_A_PE_10_14__read;
  wire [512:0] fifo_A_PE_10_14__din;
  wire fifo_A_PE_10_14__full_n;
  wire fifo_A_PE_10_14__write;
  wire [512:0] fifo_A_PE_10_15__dout;
  wire fifo_A_PE_10_15__empty_n;
  wire fifo_A_PE_10_15__read;
  wire [512:0] fifo_A_PE_10_15__din;
  wire fifo_A_PE_10_15__full_n;
  wire fifo_A_PE_10_15__write;
  wire [512:0] fifo_A_PE_10_16__dout;
  wire fifo_A_PE_10_16__empty_n;
  wire fifo_A_PE_10_16__read;
  wire [512:0] fifo_A_PE_10_16__din;
  wire fifo_A_PE_10_16__full_n;
  wire fifo_A_PE_10_16__write;
  wire [512:0] fifo_A_PE_10_17__dout;
  wire fifo_A_PE_10_17__empty_n;
  wire fifo_A_PE_10_17__read;
  wire [512:0] fifo_A_PE_10_17__din;
  wire fifo_A_PE_10_17__full_n;
  wire fifo_A_PE_10_17__write;
  wire [512:0] fifo_A_PE_10_2__dout;
  wire fifo_A_PE_10_2__empty_n;
  wire fifo_A_PE_10_2__read;
  wire [512:0] fifo_A_PE_10_2__din;
  wire fifo_A_PE_10_2__full_n;
  wire fifo_A_PE_10_2__write;
  wire [512:0] fifo_A_PE_10_3__dout;
  wire fifo_A_PE_10_3__empty_n;
  wire fifo_A_PE_10_3__read;
  wire [512:0] fifo_A_PE_10_3__din;
  wire fifo_A_PE_10_3__full_n;
  wire fifo_A_PE_10_3__write;
  wire [512:0] fifo_A_PE_10_4__dout;
  wire fifo_A_PE_10_4__empty_n;
  wire fifo_A_PE_10_4__read;
  wire [512:0] fifo_A_PE_10_4__din;
  wire fifo_A_PE_10_4__full_n;
  wire fifo_A_PE_10_4__write;
  wire [512:0] fifo_A_PE_10_5__dout;
  wire fifo_A_PE_10_5__empty_n;
  wire fifo_A_PE_10_5__read;
  wire [512:0] fifo_A_PE_10_5__din;
  wire fifo_A_PE_10_5__full_n;
  wire fifo_A_PE_10_5__write;
  wire [512:0] fifo_A_PE_10_6__dout;
  wire fifo_A_PE_10_6__empty_n;
  wire fifo_A_PE_10_6__read;
  wire [512:0] fifo_A_PE_10_6__din;
  wire fifo_A_PE_10_6__full_n;
  wire fifo_A_PE_10_6__write;
  wire [512:0] fifo_A_PE_10_7__dout;
  wire fifo_A_PE_10_7__empty_n;
  wire fifo_A_PE_10_7__read;
  wire [512:0] fifo_A_PE_10_7__din;
  wire fifo_A_PE_10_7__full_n;
  wire fifo_A_PE_10_7__write;
  wire [512:0] fifo_A_PE_10_8__dout;
  wire fifo_A_PE_10_8__empty_n;
  wire fifo_A_PE_10_8__read;
  wire [512:0] fifo_A_PE_10_8__din;
  wire fifo_A_PE_10_8__full_n;
  wire fifo_A_PE_10_8__write;
  wire [512:0] fifo_A_PE_10_9__dout;
  wire fifo_A_PE_10_9__empty_n;
  wire fifo_A_PE_10_9__read;
  wire [512:0] fifo_A_PE_10_9__din;
  wire fifo_A_PE_10_9__full_n;
  wire fifo_A_PE_10_9__write;
  wire [512:0] fifo_A_PE_11_0__dout;
  wire fifo_A_PE_11_0__empty_n;
  wire fifo_A_PE_11_0__read;
  wire [512:0] fifo_A_PE_11_0__din;
  wire fifo_A_PE_11_0__full_n;
  wire fifo_A_PE_11_0__write;
  wire [512:0] fifo_A_PE_11_1__dout;
  wire fifo_A_PE_11_1__empty_n;
  wire fifo_A_PE_11_1__read;
  wire [512:0] fifo_A_PE_11_1__din;
  wire fifo_A_PE_11_1__full_n;
  wire fifo_A_PE_11_1__write;
  wire [512:0] fifo_A_PE_11_10__dout;
  wire fifo_A_PE_11_10__empty_n;
  wire fifo_A_PE_11_10__read;
  wire [512:0] fifo_A_PE_11_10__din;
  wire fifo_A_PE_11_10__full_n;
  wire fifo_A_PE_11_10__write;
  wire [512:0] fifo_A_PE_11_11__dout;
  wire fifo_A_PE_11_11__empty_n;
  wire fifo_A_PE_11_11__read;
  wire [512:0] fifo_A_PE_11_11__din;
  wire fifo_A_PE_11_11__full_n;
  wire fifo_A_PE_11_11__write;
  wire [512:0] fifo_A_PE_11_12__dout;
  wire fifo_A_PE_11_12__empty_n;
  wire fifo_A_PE_11_12__read;
  wire [512:0] fifo_A_PE_11_12__din;
  wire fifo_A_PE_11_12__full_n;
  wire fifo_A_PE_11_12__write;
  wire [512:0] fifo_A_PE_11_13__dout;
  wire fifo_A_PE_11_13__empty_n;
  wire fifo_A_PE_11_13__read;
  wire [512:0] fifo_A_PE_11_13__din;
  wire fifo_A_PE_11_13__full_n;
  wire fifo_A_PE_11_13__write;
  wire [512:0] fifo_A_PE_11_14__dout;
  wire fifo_A_PE_11_14__empty_n;
  wire fifo_A_PE_11_14__read;
  wire [512:0] fifo_A_PE_11_14__din;
  wire fifo_A_PE_11_14__full_n;
  wire fifo_A_PE_11_14__write;
  wire [512:0] fifo_A_PE_11_15__dout;
  wire fifo_A_PE_11_15__empty_n;
  wire fifo_A_PE_11_15__read;
  wire [512:0] fifo_A_PE_11_15__din;
  wire fifo_A_PE_11_15__full_n;
  wire fifo_A_PE_11_15__write;
  wire [512:0] fifo_A_PE_11_16__dout;
  wire fifo_A_PE_11_16__empty_n;
  wire fifo_A_PE_11_16__read;
  wire [512:0] fifo_A_PE_11_16__din;
  wire fifo_A_PE_11_16__full_n;
  wire fifo_A_PE_11_16__write;
  wire [512:0] fifo_A_PE_11_17__dout;
  wire fifo_A_PE_11_17__empty_n;
  wire fifo_A_PE_11_17__read;
  wire [512:0] fifo_A_PE_11_17__din;
  wire fifo_A_PE_11_17__full_n;
  wire fifo_A_PE_11_17__write;
  wire [512:0] fifo_A_PE_11_2__dout;
  wire fifo_A_PE_11_2__empty_n;
  wire fifo_A_PE_11_2__read;
  wire [512:0] fifo_A_PE_11_2__din;
  wire fifo_A_PE_11_2__full_n;
  wire fifo_A_PE_11_2__write;
  wire [512:0] fifo_A_PE_11_3__dout;
  wire fifo_A_PE_11_3__empty_n;
  wire fifo_A_PE_11_3__read;
  wire [512:0] fifo_A_PE_11_3__din;
  wire fifo_A_PE_11_3__full_n;
  wire fifo_A_PE_11_3__write;
  wire [512:0] fifo_A_PE_11_4__dout;
  wire fifo_A_PE_11_4__empty_n;
  wire fifo_A_PE_11_4__read;
  wire [512:0] fifo_A_PE_11_4__din;
  wire fifo_A_PE_11_4__full_n;
  wire fifo_A_PE_11_4__write;
  wire [512:0] fifo_A_PE_11_5__dout;
  wire fifo_A_PE_11_5__empty_n;
  wire fifo_A_PE_11_5__read;
  wire [512:0] fifo_A_PE_11_5__din;
  wire fifo_A_PE_11_5__full_n;
  wire fifo_A_PE_11_5__write;
  wire [512:0] fifo_A_PE_11_6__dout;
  wire fifo_A_PE_11_6__empty_n;
  wire fifo_A_PE_11_6__read;
  wire [512:0] fifo_A_PE_11_6__din;
  wire fifo_A_PE_11_6__full_n;
  wire fifo_A_PE_11_6__write;
  wire [512:0] fifo_A_PE_11_7__dout;
  wire fifo_A_PE_11_7__empty_n;
  wire fifo_A_PE_11_7__read;
  wire [512:0] fifo_A_PE_11_7__din;
  wire fifo_A_PE_11_7__full_n;
  wire fifo_A_PE_11_7__write;
  wire [512:0] fifo_A_PE_11_8__dout;
  wire fifo_A_PE_11_8__empty_n;
  wire fifo_A_PE_11_8__read;
  wire [512:0] fifo_A_PE_11_8__din;
  wire fifo_A_PE_11_8__full_n;
  wire fifo_A_PE_11_8__write;
  wire [512:0] fifo_A_PE_11_9__dout;
  wire fifo_A_PE_11_9__empty_n;
  wire fifo_A_PE_11_9__read;
  wire [512:0] fifo_A_PE_11_9__din;
  wire fifo_A_PE_11_9__full_n;
  wire fifo_A_PE_11_9__write;
  wire [512:0] fifo_A_PE_12_0__dout;
  wire fifo_A_PE_12_0__empty_n;
  wire fifo_A_PE_12_0__read;
  wire [512:0] fifo_A_PE_12_0__din;
  wire fifo_A_PE_12_0__full_n;
  wire fifo_A_PE_12_0__write;
  wire [512:0] fifo_A_PE_12_1__dout;
  wire fifo_A_PE_12_1__empty_n;
  wire fifo_A_PE_12_1__read;
  wire [512:0] fifo_A_PE_12_1__din;
  wire fifo_A_PE_12_1__full_n;
  wire fifo_A_PE_12_1__write;
  wire [512:0] fifo_A_PE_12_10__dout;
  wire fifo_A_PE_12_10__empty_n;
  wire fifo_A_PE_12_10__read;
  wire [512:0] fifo_A_PE_12_10__din;
  wire fifo_A_PE_12_10__full_n;
  wire fifo_A_PE_12_10__write;
  wire [512:0] fifo_A_PE_12_11__dout;
  wire fifo_A_PE_12_11__empty_n;
  wire fifo_A_PE_12_11__read;
  wire [512:0] fifo_A_PE_12_11__din;
  wire fifo_A_PE_12_11__full_n;
  wire fifo_A_PE_12_11__write;
  wire [512:0] fifo_A_PE_12_12__dout;
  wire fifo_A_PE_12_12__empty_n;
  wire fifo_A_PE_12_12__read;
  wire [512:0] fifo_A_PE_12_12__din;
  wire fifo_A_PE_12_12__full_n;
  wire fifo_A_PE_12_12__write;
  wire [512:0] fifo_A_PE_12_13__dout;
  wire fifo_A_PE_12_13__empty_n;
  wire fifo_A_PE_12_13__read;
  wire [512:0] fifo_A_PE_12_13__din;
  wire fifo_A_PE_12_13__full_n;
  wire fifo_A_PE_12_13__write;
  wire [512:0] fifo_A_PE_12_14__dout;
  wire fifo_A_PE_12_14__empty_n;
  wire fifo_A_PE_12_14__read;
  wire [512:0] fifo_A_PE_12_14__din;
  wire fifo_A_PE_12_14__full_n;
  wire fifo_A_PE_12_14__write;
  wire [512:0] fifo_A_PE_12_15__dout;
  wire fifo_A_PE_12_15__empty_n;
  wire fifo_A_PE_12_15__read;
  wire [512:0] fifo_A_PE_12_15__din;
  wire fifo_A_PE_12_15__full_n;
  wire fifo_A_PE_12_15__write;
  wire [512:0] fifo_A_PE_12_16__dout;
  wire fifo_A_PE_12_16__empty_n;
  wire fifo_A_PE_12_16__read;
  wire [512:0] fifo_A_PE_12_16__din;
  wire fifo_A_PE_12_16__full_n;
  wire fifo_A_PE_12_16__write;
  wire [512:0] fifo_A_PE_12_17__dout;
  wire fifo_A_PE_12_17__empty_n;
  wire fifo_A_PE_12_17__read;
  wire [512:0] fifo_A_PE_12_17__din;
  wire fifo_A_PE_12_17__full_n;
  wire fifo_A_PE_12_17__write;
  wire [512:0] fifo_A_PE_12_2__dout;
  wire fifo_A_PE_12_2__empty_n;
  wire fifo_A_PE_12_2__read;
  wire [512:0] fifo_A_PE_12_2__din;
  wire fifo_A_PE_12_2__full_n;
  wire fifo_A_PE_12_2__write;
  wire [512:0] fifo_A_PE_12_3__dout;
  wire fifo_A_PE_12_3__empty_n;
  wire fifo_A_PE_12_3__read;
  wire [512:0] fifo_A_PE_12_3__din;
  wire fifo_A_PE_12_3__full_n;
  wire fifo_A_PE_12_3__write;
  wire [512:0] fifo_A_PE_12_4__dout;
  wire fifo_A_PE_12_4__empty_n;
  wire fifo_A_PE_12_4__read;
  wire [512:0] fifo_A_PE_12_4__din;
  wire fifo_A_PE_12_4__full_n;
  wire fifo_A_PE_12_4__write;
  wire [512:0] fifo_A_PE_12_5__dout;
  wire fifo_A_PE_12_5__empty_n;
  wire fifo_A_PE_12_5__read;
  wire [512:0] fifo_A_PE_12_5__din;
  wire fifo_A_PE_12_5__full_n;
  wire fifo_A_PE_12_5__write;
  wire [512:0] fifo_A_PE_12_6__dout;
  wire fifo_A_PE_12_6__empty_n;
  wire fifo_A_PE_12_6__read;
  wire [512:0] fifo_A_PE_12_6__din;
  wire fifo_A_PE_12_6__full_n;
  wire fifo_A_PE_12_6__write;
  wire [512:0] fifo_A_PE_12_7__dout;
  wire fifo_A_PE_12_7__empty_n;
  wire fifo_A_PE_12_7__read;
  wire [512:0] fifo_A_PE_12_7__din;
  wire fifo_A_PE_12_7__full_n;
  wire fifo_A_PE_12_7__write;
  wire [512:0] fifo_A_PE_12_8__dout;
  wire fifo_A_PE_12_8__empty_n;
  wire fifo_A_PE_12_8__read;
  wire [512:0] fifo_A_PE_12_8__din;
  wire fifo_A_PE_12_8__full_n;
  wire fifo_A_PE_12_8__write;
  wire [512:0] fifo_A_PE_12_9__dout;
  wire fifo_A_PE_12_9__empty_n;
  wire fifo_A_PE_12_9__read;
  wire [512:0] fifo_A_PE_12_9__din;
  wire fifo_A_PE_12_9__full_n;
  wire fifo_A_PE_12_9__write;
  wire [512:0] fifo_A_PE_13_0__dout;
  wire fifo_A_PE_13_0__empty_n;
  wire fifo_A_PE_13_0__read;
  wire [512:0] fifo_A_PE_13_0__din;
  wire fifo_A_PE_13_0__full_n;
  wire fifo_A_PE_13_0__write;
  wire [512:0] fifo_A_PE_13_1__dout;
  wire fifo_A_PE_13_1__empty_n;
  wire fifo_A_PE_13_1__read;
  wire [512:0] fifo_A_PE_13_1__din;
  wire fifo_A_PE_13_1__full_n;
  wire fifo_A_PE_13_1__write;
  wire [512:0] fifo_A_PE_13_10__dout;
  wire fifo_A_PE_13_10__empty_n;
  wire fifo_A_PE_13_10__read;
  wire [512:0] fifo_A_PE_13_10__din;
  wire fifo_A_PE_13_10__full_n;
  wire fifo_A_PE_13_10__write;
  wire [512:0] fifo_A_PE_13_11__dout;
  wire fifo_A_PE_13_11__empty_n;
  wire fifo_A_PE_13_11__read;
  wire [512:0] fifo_A_PE_13_11__din;
  wire fifo_A_PE_13_11__full_n;
  wire fifo_A_PE_13_11__write;
  wire [512:0] fifo_A_PE_13_12__dout;
  wire fifo_A_PE_13_12__empty_n;
  wire fifo_A_PE_13_12__read;
  wire [512:0] fifo_A_PE_13_12__din;
  wire fifo_A_PE_13_12__full_n;
  wire fifo_A_PE_13_12__write;
  wire [512:0] fifo_A_PE_13_13__dout;
  wire fifo_A_PE_13_13__empty_n;
  wire fifo_A_PE_13_13__read;
  wire [512:0] fifo_A_PE_13_13__din;
  wire fifo_A_PE_13_13__full_n;
  wire fifo_A_PE_13_13__write;
  wire [512:0] fifo_A_PE_13_14__dout;
  wire fifo_A_PE_13_14__empty_n;
  wire fifo_A_PE_13_14__read;
  wire [512:0] fifo_A_PE_13_14__din;
  wire fifo_A_PE_13_14__full_n;
  wire fifo_A_PE_13_14__write;
  wire [512:0] fifo_A_PE_13_15__dout;
  wire fifo_A_PE_13_15__empty_n;
  wire fifo_A_PE_13_15__read;
  wire [512:0] fifo_A_PE_13_15__din;
  wire fifo_A_PE_13_15__full_n;
  wire fifo_A_PE_13_15__write;
  wire [512:0] fifo_A_PE_13_16__dout;
  wire fifo_A_PE_13_16__empty_n;
  wire fifo_A_PE_13_16__read;
  wire [512:0] fifo_A_PE_13_16__din;
  wire fifo_A_PE_13_16__full_n;
  wire fifo_A_PE_13_16__write;
  wire [512:0] fifo_A_PE_13_17__dout;
  wire fifo_A_PE_13_17__empty_n;
  wire fifo_A_PE_13_17__read;
  wire [512:0] fifo_A_PE_13_17__din;
  wire fifo_A_PE_13_17__full_n;
  wire fifo_A_PE_13_17__write;
  wire [512:0] fifo_A_PE_13_2__dout;
  wire fifo_A_PE_13_2__empty_n;
  wire fifo_A_PE_13_2__read;
  wire [512:0] fifo_A_PE_13_2__din;
  wire fifo_A_PE_13_2__full_n;
  wire fifo_A_PE_13_2__write;
  wire [512:0] fifo_A_PE_13_3__dout;
  wire fifo_A_PE_13_3__empty_n;
  wire fifo_A_PE_13_3__read;
  wire [512:0] fifo_A_PE_13_3__din;
  wire fifo_A_PE_13_3__full_n;
  wire fifo_A_PE_13_3__write;
  wire [512:0] fifo_A_PE_13_4__dout;
  wire fifo_A_PE_13_4__empty_n;
  wire fifo_A_PE_13_4__read;
  wire [512:0] fifo_A_PE_13_4__din;
  wire fifo_A_PE_13_4__full_n;
  wire fifo_A_PE_13_4__write;
  wire [512:0] fifo_A_PE_13_5__dout;
  wire fifo_A_PE_13_5__empty_n;
  wire fifo_A_PE_13_5__read;
  wire [512:0] fifo_A_PE_13_5__din;
  wire fifo_A_PE_13_5__full_n;
  wire fifo_A_PE_13_5__write;
  wire [512:0] fifo_A_PE_13_6__dout;
  wire fifo_A_PE_13_6__empty_n;
  wire fifo_A_PE_13_6__read;
  wire [512:0] fifo_A_PE_13_6__din;
  wire fifo_A_PE_13_6__full_n;
  wire fifo_A_PE_13_6__write;
  wire [512:0] fifo_A_PE_13_7__dout;
  wire fifo_A_PE_13_7__empty_n;
  wire fifo_A_PE_13_7__read;
  wire [512:0] fifo_A_PE_13_7__din;
  wire fifo_A_PE_13_7__full_n;
  wire fifo_A_PE_13_7__write;
  wire [512:0] fifo_A_PE_13_8__dout;
  wire fifo_A_PE_13_8__empty_n;
  wire fifo_A_PE_13_8__read;
  wire [512:0] fifo_A_PE_13_8__din;
  wire fifo_A_PE_13_8__full_n;
  wire fifo_A_PE_13_8__write;
  wire [512:0] fifo_A_PE_13_9__dout;
  wire fifo_A_PE_13_9__empty_n;
  wire fifo_A_PE_13_9__read;
  wire [512:0] fifo_A_PE_13_9__din;
  wire fifo_A_PE_13_9__full_n;
  wire fifo_A_PE_13_9__write;
  wire [512:0] fifo_A_PE_14_0__dout;
  wire fifo_A_PE_14_0__empty_n;
  wire fifo_A_PE_14_0__read;
  wire [512:0] fifo_A_PE_14_0__din;
  wire fifo_A_PE_14_0__full_n;
  wire fifo_A_PE_14_0__write;
  wire [512:0] fifo_A_PE_14_1__dout;
  wire fifo_A_PE_14_1__empty_n;
  wire fifo_A_PE_14_1__read;
  wire [512:0] fifo_A_PE_14_1__din;
  wire fifo_A_PE_14_1__full_n;
  wire fifo_A_PE_14_1__write;
  wire [512:0] fifo_A_PE_14_10__dout;
  wire fifo_A_PE_14_10__empty_n;
  wire fifo_A_PE_14_10__read;
  wire [512:0] fifo_A_PE_14_10__din;
  wire fifo_A_PE_14_10__full_n;
  wire fifo_A_PE_14_10__write;
  wire [512:0] fifo_A_PE_14_11__dout;
  wire fifo_A_PE_14_11__empty_n;
  wire fifo_A_PE_14_11__read;
  wire [512:0] fifo_A_PE_14_11__din;
  wire fifo_A_PE_14_11__full_n;
  wire fifo_A_PE_14_11__write;
  wire [512:0] fifo_A_PE_14_12__dout;
  wire fifo_A_PE_14_12__empty_n;
  wire fifo_A_PE_14_12__read;
  wire [512:0] fifo_A_PE_14_12__din;
  wire fifo_A_PE_14_12__full_n;
  wire fifo_A_PE_14_12__write;
  wire [512:0] fifo_A_PE_14_13__dout;
  wire fifo_A_PE_14_13__empty_n;
  wire fifo_A_PE_14_13__read;
  wire [512:0] fifo_A_PE_14_13__din;
  wire fifo_A_PE_14_13__full_n;
  wire fifo_A_PE_14_13__write;
  wire [512:0] fifo_A_PE_14_14__dout;
  wire fifo_A_PE_14_14__empty_n;
  wire fifo_A_PE_14_14__read;
  wire [512:0] fifo_A_PE_14_14__din;
  wire fifo_A_PE_14_14__full_n;
  wire fifo_A_PE_14_14__write;
  wire [512:0] fifo_A_PE_14_15__dout;
  wire fifo_A_PE_14_15__empty_n;
  wire fifo_A_PE_14_15__read;
  wire [512:0] fifo_A_PE_14_15__din;
  wire fifo_A_PE_14_15__full_n;
  wire fifo_A_PE_14_15__write;
  wire [512:0] fifo_A_PE_14_16__dout;
  wire fifo_A_PE_14_16__empty_n;
  wire fifo_A_PE_14_16__read;
  wire [512:0] fifo_A_PE_14_16__din;
  wire fifo_A_PE_14_16__full_n;
  wire fifo_A_PE_14_16__write;
  wire [512:0] fifo_A_PE_14_17__dout;
  wire fifo_A_PE_14_17__empty_n;
  wire fifo_A_PE_14_17__read;
  wire [512:0] fifo_A_PE_14_17__din;
  wire fifo_A_PE_14_17__full_n;
  wire fifo_A_PE_14_17__write;
  wire [512:0] fifo_A_PE_14_2__dout;
  wire fifo_A_PE_14_2__empty_n;
  wire fifo_A_PE_14_2__read;
  wire [512:0] fifo_A_PE_14_2__din;
  wire fifo_A_PE_14_2__full_n;
  wire fifo_A_PE_14_2__write;
  wire [512:0] fifo_A_PE_14_3__dout;
  wire fifo_A_PE_14_3__empty_n;
  wire fifo_A_PE_14_3__read;
  wire [512:0] fifo_A_PE_14_3__din;
  wire fifo_A_PE_14_3__full_n;
  wire fifo_A_PE_14_3__write;
  wire [512:0] fifo_A_PE_14_4__dout;
  wire fifo_A_PE_14_4__empty_n;
  wire fifo_A_PE_14_4__read;
  wire [512:0] fifo_A_PE_14_4__din;
  wire fifo_A_PE_14_4__full_n;
  wire fifo_A_PE_14_4__write;
  wire [512:0] fifo_A_PE_14_5__dout;
  wire fifo_A_PE_14_5__empty_n;
  wire fifo_A_PE_14_5__read;
  wire [512:0] fifo_A_PE_14_5__din;
  wire fifo_A_PE_14_5__full_n;
  wire fifo_A_PE_14_5__write;
  wire [512:0] fifo_A_PE_14_6__dout;
  wire fifo_A_PE_14_6__empty_n;
  wire fifo_A_PE_14_6__read;
  wire [512:0] fifo_A_PE_14_6__din;
  wire fifo_A_PE_14_6__full_n;
  wire fifo_A_PE_14_6__write;
  wire [512:0] fifo_A_PE_14_7__dout;
  wire fifo_A_PE_14_7__empty_n;
  wire fifo_A_PE_14_7__read;
  wire [512:0] fifo_A_PE_14_7__din;
  wire fifo_A_PE_14_7__full_n;
  wire fifo_A_PE_14_7__write;
  wire [512:0] fifo_A_PE_14_8__dout;
  wire fifo_A_PE_14_8__empty_n;
  wire fifo_A_PE_14_8__read;
  wire [512:0] fifo_A_PE_14_8__din;
  wire fifo_A_PE_14_8__full_n;
  wire fifo_A_PE_14_8__write;
  wire [512:0] fifo_A_PE_14_9__dout;
  wire fifo_A_PE_14_9__empty_n;
  wire fifo_A_PE_14_9__read;
  wire [512:0] fifo_A_PE_14_9__din;
  wire fifo_A_PE_14_9__full_n;
  wire fifo_A_PE_14_9__write;
  wire [512:0] fifo_A_PE_15_0__dout;
  wire fifo_A_PE_15_0__empty_n;
  wire fifo_A_PE_15_0__read;
  wire [512:0] fifo_A_PE_15_0__din;
  wire fifo_A_PE_15_0__full_n;
  wire fifo_A_PE_15_0__write;
  wire [512:0] fifo_A_PE_15_1__dout;
  wire fifo_A_PE_15_1__empty_n;
  wire fifo_A_PE_15_1__read;
  wire [512:0] fifo_A_PE_15_1__din;
  wire fifo_A_PE_15_1__full_n;
  wire fifo_A_PE_15_1__write;
  wire [512:0] fifo_A_PE_15_10__dout;
  wire fifo_A_PE_15_10__empty_n;
  wire fifo_A_PE_15_10__read;
  wire [512:0] fifo_A_PE_15_10__din;
  wire fifo_A_PE_15_10__full_n;
  wire fifo_A_PE_15_10__write;
  wire [512:0] fifo_A_PE_15_11__dout;
  wire fifo_A_PE_15_11__empty_n;
  wire fifo_A_PE_15_11__read;
  wire [512:0] fifo_A_PE_15_11__din;
  wire fifo_A_PE_15_11__full_n;
  wire fifo_A_PE_15_11__write;
  wire [512:0] fifo_A_PE_15_12__dout;
  wire fifo_A_PE_15_12__empty_n;
  wire fifo_A_PE_15_12__read;
  wire [512:0] fifo_A_PE_15_12__din;
  wire fifo_A_PE_15_12__full_n;
  wire fifo_A_PE_15_12__write;
  wire [512:0] fifo_A_PE_15_13__dout;
  wire fifo_A_PE_15_13__empty_n;
  wire fifo_A_PE_15_13__read;
  wire [512:0] fifo_A_PE_15_13__din;
  wire fifo_A_PE_15_13__full_n;
  wire fifo_A_PE_15_13__write;
  wire [512:0] fifo_A_PE_15_14__dout;
  wire fifo_A_PE_15_14__empty_n;
  wire fifo_A_PE_15_14__read;
  wire [512:0] fifo_A_PE_15_14__din;
  wire fifo_A_PE_15_14__full_n;
  wire fifo_A_PE_15_14__write;
  wire [512:0] fifo_A_PE_15_15__dout;
  wire fifo_A_PE_15_15__empty_n;
  wire fifo_A_PE_15_15__read;
  wire [512:0] fifo_A_PE_15_15__din;
  wire fifo_A_PE_15_15__full_n;
  wire fifo_A_PE_15_15__write;
  wire [512:0] fifo_A_PE_15_16__dout;
  wire fifo_A_PE_15_16__empty_n;
  wire fifo_A_PE_15_16__read;
  wire [512:0] fifo_A_PE_15_16__din;
  wire fifo_A_PE_15_16__full_n;
  wire fifo_A_PE_15_16__write;
  wire [512:0] fifo_A_PE_15_17__dout;
  wire fifo_A_PE_15_17__empty_n;
  wire fifo_A_PE_15_17__read;
  wire [512:0] fifo_A_PE_15_17__din;
  wire fifo_A_PE_15_17__full_n;
  wire fifo_A_PE_15_17__write;
  wire [512:0] fifo_A_PE_15_2__dout;
  wire fifo_A_PE_15_2__empty_n;
  wire fifo_A_PE_15_2__read;
  wire [512:0] fifo_A_PE_15_2__din;
  wire fifo_A_PE_15_2__full_n;
  wire fifo_A_PE_15_2__write;
  wire [512:0] fifo_A_PE_15_3__dout;
  wire fifo_A_PE_15_3__empty_n;
  wire fifo_A_PE_15_3__read;
  wire [512:0] fifo_A_PE_15_3__din;
  wire fifo_A_PE_15_3__full_n;
  wire fifo_A_PE_15_3__write;
  wire [512:0] fifo_A_PE_15_4__dout;
  wire fifo_A_PE_15_4__empty_n;
  wire fifo_A_PE_15_4__read;
  wire [512:0] fifo_A_PE_15_4__din;
  wire fifo_A_PE_15_4__full_n;
  wire fifo_A_PE_15_4__write;
  wire [512:0] fifo_A_PE_15_5__dout;
  wire fifo_A_PE_15_5__empty_n;
  wire fifo_A_PE_15_5__read;
  wire [512:0] fifo_A_PE_15_5__din;
  wire fifo_A_PE_15_5__full_n;
  wire fifo_A_PE_15_5__write;
  wire [512:0] fifo_A_PE_15_6__dout;
  wire fifo_A_PE_15_6__empty_n;
  wire fifo_A_PE_15_6__read;
  wire [512:0] fifo_A_PE_15_6__din;
  wire fifo_A_PE_15_6__full_n;
  wire fifo_A_PE_15_6__write;
  wire [512:0] fifo_A_PE_15_7__dout;
  wire fifo_A_PE_15_7__empty_n;
  wire fifo_A_PE_15_7__read;
  wire [512:0] fifo_A_PE_15_7__din;
  wire fifo_A_PE_15_7__full_n;
  wire fifo_A_PE_15_7__write;
  wire [512:0] fifo_A_PE_15_8__dout;
  wire fifo_A_PE_15_8__empty_n;
  wire fifo_A_PE_15_8__read;
  wire [512:0] fifo_A_PE_15_8__din;
  wire fifo_A_PE_15_8__full_n;
  wire fifo_A_PE_15_8__write;
  wire [512:0] fifo_A_PE_15_9__dout;
  wire fifo_A_PE_15_9__empty_n;
  wire fifo_A_PE_15_9__read;
  wire [512:0] fifo_A_PE_15_9__din;
  wire fifo_A_PE_15_9__full_n;
  wire fifo_A_PE_15_9__write;
  wire [512:0] fifo_A_PE_16_0__dout;
  wire fifo_A_PE_16_0__empty_n;
  wire fifo_A_PE_16_0__read;
  wire [512:0] fifo_A_PE_16_0__din;
  wire fifo_A_PE_16_0__full_n;
  wire fifo_A_PE_16_0__write;
  wire [512:0] fifo_A_PE_16_1__dout;
  wire fifo_A_PE_16_1__empty_n;
  wire fifo_A_PE_16_1__read;
  wire [512:0] fifo_A_PE_16_1__din;
  wire fifo_A_PE_16_1__full_n;
  wire fifo_A_PE_16_1__write;
  wire [512:0] fifo_A_PE_16_10__dout;
  wire fifo_A_PE_16_10__empty_n;
  wire fifo_A_PE_16_10__read;
  wire [512:0] fifo_A_PE_16_10__din;
  wire fifo_A_PE_16_10__full_n;
  wire fifo_A_PE_16_10__write;
  wire [512:0] fifo_A_PE_16_11__dout;
  wire fifo_A_PE_16_11__empty_n;
  wire fifo_A_PE_16_11__read;
  wire [512:0] fifo_A_PE_16_11__din;
  wire fifo_A_PE_16_11__full_n;
  wire fifo_A_PE_16_11__write;
  wire [512:0] fifo_A_PE_16_12__dout;
  wire fifo_A_PE_16_12__empty_n;
  wire fifo_A_PE_16_12__read;
  wire [512:0] fifo_A_PE_16_12__din;
  wire fifo_A_PE_16_12__full_n;
  wire fifo_A_PE_16_12__write;
  wire [512:0] fifo_A_PE_16_13__dout;
  wire fifo_A_PE_16_13__empty_n;
  wire fifo_A_PE_16_13__read;
  wire [512:0] fifo_A_PE_16_13__din;
  wire fifo_A_PE_16_13__full_n;
  wire fifo_A_PE_16_13__write;
  wire [512:0] fifo_A_PE_16_14__dout;
  wire fifo_A_PE_16_14__empty_n;
  wire fifo_A_PE_16_14__read;
  wire [512:0] fifo_A_PE_16_14__din;
  wire fifo_A_PE_16_14__full_n;
  wire fifo_A_PE_16_14__write;
  wire [512:0] fifo_A_PE_16_15__dout;
  wire fifo_A_PE_16_15__empty_n;
  wire fifo_A_PE_16_15__read;
  wire [512:0] fifo_A_PE_16_15__din;
  wire fifo_A_PE_16_15__full_n;
  wire fifo_A_PE_16_15__write;
  wire [512:0] fifo_A_PE_16_16__dout;
  wire fifo_A_PE_16_16__empty_n;
  wire fifo_A_PE_16_16__read;
  wire [512:0] fifo_A_PE_16_16__din;
  wire fifo_A_PE_16_16__full_n;
  wire fifo_A_PE_16_16__write;
  wire [512:0] fifo_A_PE_16_17__dout;
  wire fifo_A_PE_16_17__empty_n;
  wire fifo_A_PE_16_17__read;
  wire [512:0] fifo_A_PE_16_17__din;
  wire fifo_A_PE_16_17__full_n;
  wire fifo_A_PE_16_17__write;
  wire [512:0] fifo_A_PE_16_2__dout;
  wire fifo_A_PE_16_2__empty_n;
  wire fifo_A_PE_16_2__read;
  wire [512:0] fifo_A_PE_16_2__din;
  wire fifo_A_PE_16_2__full_n;
  wire fifo_A_PE_16_2__write;
  wire [512:0] fifo_A_PE_16_3__dout;
  wire fifo_A_PE_16_3__empty_n;
  wire fifo_A_PE_16_3__read;
  wire [512:0] fifo_A_PE_16_3__din;
  wire fifo_A_PE_16_3__full_n;
  wire fifo_A_PE_16_3__write;
  wire [512:0] fifo_A_PE_16_4__dout;
  wire fifo_A_PE_16_4__empty_n;
  wire fifo_A_PE_16_4__read;
  wire [512:0] fifo_A_PE_16_4__din;
  wire fifo_A_PE_16_4__full_n;
  wire fifo_A_PE_16_4__write;
  wire [512:0] fifo_A_PE_16_5__dout;
  wire fifo_A_PE_16_5__empty_n;
  wire fifo_A_PE_16_5__read;
  wire [512:0] fifo_A_PE_16_5__din;
  wire fifo_A_PE_16_5__full_n;
  wire fifo_A_PE_16_5__write;
  wire [512:0] fifo_A_PE_16_6__dout;
  wire fifo_A_PE_16_6__empty_n;
  wire fifo_A_PE_16_6__read;
  wire [512:0] fifo_A_PE_16_6__din;
  wire fifo_A_PE_16_6__full_n;
  wire fifo_A_PE_16_6__write;
  wire [512:0] fifo_A_PE_16_7__dout;
  wire fifo_A_PE_16_7__empty_n;
  wire fifo_A_PE_16_7__read;
  wire [512:0] fifo_A_PE_16_7__din;
  wire fifo_A_PE_16_7__full_n;
  wire fifo_A_PE_16_7__write;
  wire [512:0] fifo_A_PE_16_8__dout;
  wire fifo_A_PE_16_8__empty_n;
  wire fifo_A_PE_16_8__read;
  wire [512:0] fifo_A_PE_16_8__din;
  wire fifo_A_PE_16_8__full_n;
  wire fifo_A_PE_16_8__write;
  wire [512:0] fifo_A_PE_16_9__dout;
  wire fifo_A_PE_16_9__empty_n;
  wire fifo_A_PE_16_9__read;
  wire [512:0] fifo_A_PE_16_9__din;
  wire fifo_A_PE_16_9__full_n;
  wire fifo_A_PE_16_9__write;
  wire [512:0] fifo_A_PE_17_0__dout;
  wire fifo_A_PE_17_0__empty_n;
  wire fifo_A_PE_17_0__read;
  wire [512:0] fifo_A_PE_17_0__din;
  wire fifo_A_PE_17_0__full_n;
  wire fifo_A_PE_17_0__write;
  wire [512:0] fifo_A_PE_17_1__dout;
  wire fifo_A_PE_17_1__empty_n;
  wire fifo_A_PE_17_1__read;
  wire [512:0] fifo_A_PE_17_1__din;
  wire fifo_A_PE_17_1__full_n;
  wire fifo_A_PE_17_1__write;
  wire [512:0] fifo_A_PE_17_10__dout;
  wire fifo_A_PE_17_10__empty_n;
  wire fifo_A_PE_17_10__read;
  wire [512:0] fifo_A_PE_17_10__din;
  wire fifo_A_PE_17_10__full_n;
  wire fifo_A_PE_17_10__write;
  wire [512:0] fifo_A_PE_17_11__dout;
  wire fifo_A_PE_17_11__empty_n;
  wire fifo_A_PE_17_11__read;
  wire [512:0] fifo_A_PE_17_11__din;
  wire fifo_A_PE_17_11__full_n;
  wire fifo_A_PE_17_11__write;
  wire [512:0] fifo_A_PE_17_12__dout;
  wire fifo_A_PE_17_12__empty_n;
  wire fifo_A_PE_17_12__read;
  wire [512:0] fifo_A_PE_17_12__din;
  wire fifo_A_PE_17_12__full_n;
  wire fifo_A_PE_17_12__write;
  wire [512:0] fifo_A_PE_17_13__dout;
  wire fifo_A_PE_17_13__empty_n;
  wire fifo_A_PE_17_13__read;
  wire [512:0] fifo_A_PE_17_13__din;
  wire fifo_A_PE_17_13__full_n;
  wire fifo_A_PE_17_13__write;
  wire [512:0] fifo_A_PE_17_14__dout;
  wire fifo_A_PE_17_14__empty_n;
  wire fifo_A_PE_17_14__read;
  wire [512:0] fifo_A_PE_17_14__din;
  wire fifo_A_PE_17_14__full_n;
  wire fifo_A_PE_17_14__write;
  wire [512:0] fifo_A_PE_17_15__dout;
  wire fifo_A_PE_17_15__empty_n;
  wire fifo_A_PE_17_15__read;
  wire [512:0] fifo_A_PE_17_15__din;
  wire fifo_A_PE_17_15__full_n;
  wire fifo_A_PE_17_15__write;
  wire [512:0] fifo_A_PE_17_16__dout;
  wire fifo_A_PE_17_16__empty_n;
  wire fifo_A_PE_17_16__read;
  wire [512:0] fifo_A_PE_17_16__din;
  wire fifo_A_PE_17_16__full_n;
  wire fifo_A_PE_17_16__write;
  wire [512:0] fifo_A_PE_17_17__dout;
  wire fifo_A_PE_17_17__empty_n;
  wire fifo_A_PE_17_17__read;
  wire [512:0] fifo_A_PE_17_17__din;
  wire fifo_A_PE_17_17__full_n;
  wire fifo_A_PE_17_17__write;
  wire [512:0] fifo_A_PE_17_2__dout;
  wire fifo_A_PE_17_2__empty_n;
  wire fifo_A_PE_17_2__read;
  wire [512:0] fifo_A_PE_17_2__din;
  wire fifo_A_PE_17_2__full_n;
  wire fifo_A_PE_17_2__write;
  wire [512:0] fifo_A_PE_17_3__dout;
  wire fifo_A_PE_17_3__empty_n;
  wire fifo_A_PE_17_3__read;
  wire [512:0] fifo_A_PE_17_3__din;
  wire fifo_A_PE_17_3__full_n;
  wire fifo_A_PE_17_3__write;
  wire [512:0] fifo_A_PE_17_4__dout;
  wire fifo_A_PE_17_4__empty_n;
  wire fifo_A_PE_17_4__read;
  wire [512:0] fifo_A_PE_17_4__din;
  wire fifo_A_PE_17_4__full_n;
  wire fifo_A_PE_17_4__write;
  wire [512:0] fifo_A_PE_17_5__dout;
  wire fifo_A_PE_17_5__empty_n;
  wire fifo_A_PE_17_5__read;
  wire [512:0] fifo_A_PE_17_5__din;
  wire fifo_A_PE_17_5__full_n;
  wire fifo_A_PE_17_5__write;
  wire [512:0] fifo_A_PE_17_6__dout;
  wire fifo_A_PE_17_6__empty_n;
  wire fifo_A_PE_17_6__read;
  wire [512:0] fifo_A_PE_17_6__din;
  wire fifo_A_PE_17_6__full_n;
  wire fifo_A_PE_17_6__write;
  wire [512:0] fifo_A_PE_17_7__dout;
  wire fifo_A_PE_17_7__empty_n;
  wire fifo_A_PE_17_7__read;
  wire [512:0] fifo_A_PE_17_7__din;
  wire fifo_A_PE_17_7__full_n;
  wire fifo_A_PE_17_7__write;
  wire [512:0] fifo_A_PE_17_8__dout;
  wire fifo_A_PE_17_8__empty_n;
  wire fifo_A_PE_17_8__read;
  wire [512:0] fifo_A_PE_17_8__din;
  wire fifo_A_PE_17_8__full_n;
  wire fifo_A_PE_17_8__write;
  wire [512:0] fifo_A_PE_17_9__dout;
  wire fifo_A_PE_17_9__empty_n;
  wire fifo_A_PE_17_9__read;
  wire [512:0] fifo_A_PE_17_9__din;
  wire fifo_A_PE_17_9__full_n;
  wire fifo_A_PE_17_9__write;
  wire [512:0] fifo_A_PE_1_0__dout;
  wire fifo_A_PE_1_0__empty_n;
  wire fifo_A_PE_1_0__read;
  wire [512:0] fifo_A_PE_1_0__din;
  wire fifo_A_PE_1_0__full_n;
  wire fifo_A_PE_1_0__write;
  wire [512:0] fifo_A_PE_1_1__dout;
  wire fifo_A_PE_1_1__empty_n;
  wire fifo_A_PE_1_1__read;
  wire [512:0] fifo_A_PE_1_1__din;
  wire fifo_A_PE_1_1__full_n;
  wire fifo_A_PE_1_1__write;
  wire [512:0] fifo_A_PE_1_10__dout;
  wire fifo_A_PE_1_10__empty_n;
  wire fifo_A_PE_1_10__read;
  wire [512:0] fifo_A_PE_1_10__din;
  wire fifo_A_PE_1_10__full_n;
  wire fifo_A_PE_1_10__write;
  wire [512:0] fifo_A_PE_1_11__dout;
  wire fifo_A_PE_1_11__empty_n;
  wire fifo_A_PE_1_11__read;
  wire [512:0] fifo_A_PE_1_11__din;
  wire fifo_A_PE_1_11__full_n;
  wire fifo_A_PE_1_11__write;
  wire [512:0] fifo_A_PE_1_12__dout;
  wire fifo_A_PE_1_12__empty_n;
  wire fifo_A_PE_1_12__read;
  wire [512:0] fifo_A_PE_1_12__din;
  wire fifo_A_PE_1_12__full_n;
  wire fifo_A_PE_1_12__write;
  wire [512:0] fifo_A_PE_1_13__dout;
  wire fifo_A_PE_1_13__empty_n;
  wire fifo_A_PE_1_13__read;
  wire [512:0] fifo_A_PE_1_13__din;
  wire fifo_A_PE_1_13__full_n;
  wire fifo_A_PE_1_13__write;
  wire [512:0] fifo_A_PE_1_14__dout;
  wire fifo_A_PE_1_14__empty_n;
  wire fifo_A_PE_1_14__read;
  wire [512:0] fifo_A_PE_1_14__din;
  wire fifo_A_PE_1_14__full_n;
  wire fifo_A_PE_1_14__write;
  wire [512:0] fifo_A_PE_1_15__dout;
  wire fifo_A_PE_1_15__empty_n;
  wire fifo_A_PE_1_15__read;
  wire [512:0] fifo_A_PE_1_15__din;
  wire fifo_A_PE_1_15__full_n;
  wire fifo_A_PE_1_15__write;
  wire [512:0] fifo_A_PE_1_16__dout;
  wire fifo_A_PE_1_16__empty_n;
  wire fifo_A_PE_1_16__read;
  wire [512:0] fifo_A_PE_1_16__din;
  wire fifo_A_PE_1_16__full_n;
  wire fifo_A_PE_1_16__write;
  wire [512:0] fifo_A_PE_1_17__dout;
  wire fifo_A_PE_1_17__empty_n;
  wire fifo_A_PE_1_17__read;
  wire [512:0] fifo_A_PE_1_17__din;
  wire fifo_A_PE_1_17__full_n;
  wire fifo_A_PE_1_17__write;
  wire [512:0] fifo_A_PE_1_2__dout;
  wire fifo_A_PE_1_2__empty_n;
  wire fifo_A_PE_1_2__read;
  wire [512:0] fifo_A_PE_1_2__din;
  wire fifo_A_PE_1_2__full_n;
  wire fifo_A_PE_1_2__write;
  wire [512:0] fifo_A_PE_1_3__dout;
  wire fifo_A_PE_1_3__empty_n;
  wire fifo_A_PE_1_3__read;
  wire [512:0] fifo_A_PE_1_3__din;
  wire fifo_A_PE_1_3__full_n;
  wire fifo_A_PE_1_3__write;
  wire [512:0] fifo_A_PE_1_4__dout;
  wire fifo_A_PE_1_4__empty_n;
  wire fifo_A_PE_1_4__read;
  wire [512:0] fifo_A_PE_1_4__din;
  wire fifo_A_PE_1_4__full_n;
  wire fifo_A_PE_1_4__write;
  wire [512:0] fifo_A_PE_1_5__dout;
  wire fifo_A_PE_1_5__empty_n;
  wire fifo_A_PE_1_5__read;
  wire [512:0] fifo_A_PE_1_5__din;
  wire fifo_A_PE_1_5__full_n;
  wire fifo_A_PE_1_5__write;
  wire [512:0] fifo_A_PE_1_6__dout;
  wire fifo_A_PE_1_6__empty_n;
  wire fifo_A_PE_1_6__read;
  wire [512:0] fifo_A_PE_1_6__din;
  wire fifo_A_PE_1_6__full_n;
  wire fifo_A_PE_1_6__write;
  wire [512:0] fifo_A_PE_1_7__dout;
  wire fifo_A_PE_1_7__empty_n;
  wire fifo_A_PE_1_7__read;
  wire [512:0] fifo_A_PE_1_7__din;
  wire fifo_A_PE_1_7__full_n;
  wire fifo_A_PE_1_7__write;
  wire [512:0] fifo_A_PE_1_8__dout;
  wire fifo_A_PE_1_8__empty_n;
  wire fifo_A_PE_1_8__read;
  wire [512:0] fifo_A_PE_1_8__din;
  wire fifo_A_PE_1_8__full_n;
  wire fifo_A_PE_1_8__write;
  wire [512:0] fifo_A_PE_1_9__dout;
  wire fifo_A_PE_1_9__empty_n;
  wire fifo_A_PE_1_9__read;
  wire [512:0] fifo_A_PE_1_9__din;
  wire fifo_A_PE_1_9__full_n;
  wire fifo_A_PE_1_9__write;
  wire [512:0] fifo_A_PE_2_0__dout;
  wire fifo_A_PE_2_0__empty_n;
  wire fifo_A_PE_2_0__read;
  wire [512:0] fifo_A_PE_2_0__din;
  wire fifo_A_PE_2_0__full_n;
  wire fifo_A_PE_2_0__write;
  wire [512:0] fifo_A_PE_2_1__dout;
  wire fifo_A_PE_2_1__empty_n;
  wire fifo_A_PE_2_1__read;
  wire [512:0] fifo_A_PE_2_1__din;
  wire fifo_A_PE_2_1__full_n;
  wire fifo_A_PE_2_1__write;
  wire [512:0] fifo_A_PE_2_10__dout;
  wire fifo_A_PE_2_10__empty_n;
  wire fifo_A_PE_2_10__read;
  wire [512:0] fifo_A_PE_2_10__din;
  wire fifo_A_PE_2_10__full_n;
  wire fifo_A_PE_2_10__write;
  wire [512:0] fifo_A_PE_2_11__dout;
  wire fifo_A_PE_2_11__empty_n;
  wire fifo_A_PE_2_11__read;
  wire [512:0] fifo_A_PE_2_11__din;
  wire fifo_A_PE_2_11__full_n;
  wire fifo_A_PE_2_11__write;
  wire [512:0] fifo_A_PE_2_12__dout;
  wire fifo_A_PE_2_12__empty_n;
  wire fifo_A_PE_2_12__read;
  wire [512:0] fifo_A_PE_2_12__din;
  wire fifo_A_PE_2_12__full_n;
  wire fifo_A_PE_2_12__write;
  wire [512:0] fifo_A_PE_2_13__dout;
  wire fifo_A_PE_2_13__empty_n;
  wire fifo_A_PE_2_13__read;
  wire [512:0] fifo_A_PE_2_13__din;
  wire fifo_A_PE_2_13__full_n;
  wire fifo_A_PE_2_13__write;
  wire [512:0] fifo_A_PE_2_14__dout;
  wire fifo_A_PE_2_14__empty_n;
  wire fifo_A_PE_2_14__read;
  wire [512:0] fifo_A_PE_2_14__din;
  wire fifo_A_PE_2_14__full_n;
  wire fifo_A_PE_2_14__write;
  wire [512:0] fifo_A_PE_2_15__dout;
  wire fifo_A_PE_2_15__empty_n;
  wire fifo_A_PE_2_15__read;
  wire [512:0] fifo_A_PE_2_15__din;
  wire fifo_A_PE_2_15__full_n;
  wire fifo_A_PE_2_15__write;
  wire [512:0] fifo_A_PE_2_16__dout;
  wire fifo_A_PE_2_16__empty_n;
  wire fifo_A_PE_2_16__read;
  wire [512:0] fifo_A_PE_2_16__din;
  wire fifo_A_PE_2_16__full_n;
  wire fifo_A_PE_2_16__write;
  wire [512:0] fifo_A_PE_2_17__dout;
  wire fifo_A_PE_2_17__empty_n;
  wire fifo_A_PE_2_17__read;
  wire [512:0] fifo_A_PE_2_17__din;
  wire fifo_A_PE_2_17__full_n;
  wire fifo_A_PE_2_17__write;
  wire [512:0] fifo_A_PE_2_2__dout;
  wire fifo_A_PE_2_2__empty_n;
  wire fifo_A_PE_2_2__read;
  wire [512:0] fifo_A_PE_2_2__din;
  wire fifo_A_PE_2_2__full_n;
  wire fifo_A_PE_2_2__write;
  wire [512:0] fifo_A_PE_2_3__dout;
  wire fifo_A_PE_2_3__empty_n;
  wire fifo_A_PE_2_3__read;
  wire [512:0] fifo_A_PE_2_3__din;
  wire fifo_A_PE_2_3__full_n;
  wire fifo_A_PE_2_3__write;
  wire [512:0] fifo_A_PE_2_4__dout;
  wire fifo_A_PE_2_4__empty_n;
  wire fifo_A_PE_2_4__read;
  wire [512:0] fifo_A_PE_2_4__din;
  wire fifo_A_PE_2_4__full_n;
  wire fifo_A_PE_2_4__write;
  wire [512:0] fifo_A_PE_2_5__dout;
  wire fifo_A_PE_2_5__empty_n;
  wire fifo_A_PE_2_5__read;
  wire [512:0] fifo_A_PE_2_5__din;
  wire fifo_A_PE_2_5__full_n;
  wire fifo_A_PE_2_5__write;
  wire [512:0] fifo_A_PE_2_6__dout;
  wire fifo_A_PE_2_6__empty_n;
  wire fifo_A_PE_2_6__read;
  wire [512:0] fifo_A_PE_2_6__din;
  wire fifo_A_PE_2_6__full_n;
  wire fifo_A_PE_2_6__write;
  wire [512:0] fifo_A_PE_2_7__dout;
  wire fifo_A_PE_2_7__empty_n;
  wire fifo_A_PE_2_7__read;
  wire [512:0] fifo_A_PE_2_7__din;
  wire fifo_A_PE_2_7__full_n;
  wire fifo_A_PE_2_7__write;
  wire [512:0] fifo_A_PE_2_8__dout;
  wire fifo_A_PE_2_8__empty_n;
  wire fifo_A_PE_2_8__read;
  wire [512:0] fifo_A_PE_2_8__din;
  wire fifo_A_PE_2_8__full_n;
  wire fifo_A_PE_2_8__write;
  wire [512:0] fifo_A_PE_2_9__dout;
  wire fifo_A_PE_2_9__empty_n;
  wire fifo_A_PE_2_9__read;
  wire [512:0] fifo_A_PE_2_9__din;
  wire fifo_A_PE_2_9__full_n;
  wire fifo_A_PE_2_9__write;
  wire [512:0] fifo_A_PE_3_0__dout;
  wire fifo_A_PE_3_0__empty_n;
  wire fifo_A_PE_3_0__read;
  wire [512:0] fifo_A_PE_3_0__din;
  wire fifo_A_PE_3_0__full_n;
  wire fifo_A_PE_3_0__write;
  wire [512:0] fifo_A_PE_3_1__dout;
  wire fifo_A_PE_3_1__empty_n;
  wire fifo_A_PE_3_1__read;
  wire [512:0] fifo_A_PE_3_1__din;
  wire fifo_A_PE_3_1__full_n;
  wire fifo_A_PE_3_1__write;
  wire [512:0] fifo_A_PE_3_10__dout;
  wire fifo_A_PE_3_10__empty_n;
  wire fifo_A_PE_3_10__read;
  wire [512:0] fifo_A_PE_3_10__din;
  wire fifo_A_PE_3_10__full_n;
  wire fifo_A_PE_3_10__write;
  wire [512:0] fifo_A_PE_3_11__dout;
  wire fifo_A_PE_3_11__empty_n;
  wire fifo_A_PE_3_11__read;
  wire [512:0] fifo_A_PE_3_11__din;
  wire fifo_A_PE_3_11__full_n;
  wire fifo_A_PE_3_11__write;
  wire [512:0] fifo_A_PE_3_12__dout;
  wire fifo_A_PE_3_12__empty_n;
  wire fifo_A_PE_3_12__read;
  wire [512:0] fifo_A_PE_3_12__din;
  wire fifo_A_PE_3_12__full_n;
  wire fifo_A_PE_3_12__write;
  wire [512:0] fifo_A_PE_3_13__dout;
  wire fifo_A_PE_3_13__empty_n;
  wire fifo_A_PE_3_13__read;
  wire [512:0] fifo_A_PE_3_13__din;
  wire fifo_A_PE_3_13__full_n;
  wire fifo_A_PE_3_13__write;
  wire [512:0] fifo_A_PE_3_14__dout;
  wire fifo_A_PE_3_14__empty_n;
  wire fifo_A_PE_3_14__read;
  wire [512:0] fifo_A_PE_3_14__din;
  wire fifo_A_PE_3_14__full_n;
  wire fifo_A_PE_3_14__write;
  wire [512:0] fifo_A_PE_3_15__dout;
  wire fifo_A_PE_3_15__empty_n;
  wire fifo_A_PE_3_15__read;
  wire [512:0] fifo_A_PE_3_15__din;
  wire fifo_A_PE_3_15__full_n;
  wire fifo_A_PE_3_15__write;
  wire [512:0] fifo_A_PE_3_16__dout;
  wire fifo_A_PE_3_16__empty_n;
  wire fifo_A_PE_3_16__read;
  wire [512:0] fifo_A_PE_3_16__din;
  wire fifo_A_PE_3_16__full_n;
  wire fifo_A_PE_3_16__write;
  wire [512:0] fifo_A_PE_3_17__dout;
  wire fifo_A_PE_3_17__empty_n;
  wire fifo_A_PE_3_17__read;
  wire [512:0] fifo_A_PE_3_17__din;
  wire fifo_A_PE_3_17__full_n;
  wire fifo_A_PE_3_17__write;
  wire [512:0] fifo_A_PE_3_2__dout;
  wire fifo_A_PE_3_2__empty_n;
  wire fifo_A_PE_3_2__read;
  wire [512:0] fifo_A_PE_3_2__din;
  wire fifo_A_PE_3_2__full_n;
  wire fifo_A_PE_3_2__write;
  wire [512:0] fifo_A_PE_3_3__dout;
  wire fifo_A_PE_3_3__empty_n;
  wire fifo_A_PE_3_3__read;
  wire [512:0] fifo_A_PE_3_3__din;
  wire fifo_A_PE_3_3__full_n;
  wire fifo_A_PE_3_3__write;
  wire [512:0] fifo_A_PE_3_4__dout;
  wire fifo_A_PE_3_4__empty_n;
  wire fifo_A_PE_3_4__read;
  wire [512:0] fifo_A_PE_3_4__din;
  wire fifo_A_PE_3_4__full_n;
  wire fifo_A_PE_3_4__write;
  wire [512:0] fifo_A_PE_3_5__dout;
  wire fifo_A_PE_3_5__empty_n;
  wire fifo_A_PE_3_5__read;
  wire [512:0] fifo_A_PE_3_5__din;
  wire fifo_A_PE_3_5__full_n;
  wire fifo_A_PE_3_5__write;
  wire [512:0] fifo_A_PE_3_6__dout;
  wire fifo_A_PE_3_6__empty_n;
  wire fifo_A_PE_3_6__read;
  wire [512:0] fifo_A_PE_3_6__din;
  wire fifo_A_PE_3_6__full_n;
  wire fifo_A_PE_3_6__write;
  wire [512:0] fifo_A_PE_3_7__dout;
  wire fifo_A_PE_3_7__empty_n;
  wire fifo_A_PE_3_7__read;
  wire [512:0] fifo_A_PE_3_7__din;
  wire fifo_A_PE_3_7__full_n;
  wire fifo_A_PE_3_7__write;
  wire [512:0] fifo_A_PE_3_8__dout;
  wire fifo_A_PE_3_8__empty_n;
  wire fifo_A_PE_3_8__read;
  wire [512:0] fifo_A_PE_3_8__din;
  wire fifo_A_PE_3_8__full_n;
  wire fifo_A_PE_3_8__write;
  wire [512:0] fifo_A_PE_3_9__dout;
  wire fifo_A_PE_3_9__empty_n;
  wire fifo_A_PE_3_9__read;
  wire [512:0] fifo_A_PE_3_9__din;
  wire fifo_A_PE_3_9__full_n;
  wire fifo_A_PE_3_9__write;
  wire [512:0] fifo_A_PE_4_0__dout;
  wire fifo_A_PE_4_0__empty_n;
  wire fifo_A_PE_4_0__read;
  wire [512:0] fifo_A_PE_4_0__din;
  wire fifo_A_PE_4_0__full_n;
  wire fifo_A_PE_4_0__write;
  wire [512:0] fifo_A_PE_4_1__dout;
  wire fifo_A_PE_4_1__empty_n;
  wire fifo_A_PE_4_1__read;
  wire [512:0] fifo_A_PE_4_1__din;
  wire fifo_A_PE_4_1__full_n;
  wire fifo_A_PE_4_1__write;
  wire [512:0] fifo_A_PE_4_10__dout;
  wire fifo_A_PE_4_10__empty_n;
  wire fifo_A_PE_4_10__read;
  wire [512:0] fifo_A_PE_4_10__din;
  wire fifo_A_PE_4_10__full_n;
  wire fifo_A_PE_4_10__write;
  wire [512:0] fifo_A_PE_4_11__dout;
  wire fifo_A_PE_4_11__empty_n;
  wire fifo_A_PE_4_11__read;
  wire [512:0] fifo_A_PE_4_11__din;
  wire fifo_A_PE_4_11__full_n;
  wire fifo_A_PE_4_11__write;
  wire [512:0] fifo_A_PE_4_12__dout;
  wire fifo_A_PE_4_12__empty_n;
  wire fifo_A_PE_4_12__read;
  wire [512:0] fifo_A_PE_4_12__din;
  wire fifo_A_PE_4_12__full_n;
  wire fifo_A_PE_4_12__write;
  wire [512:0] fifo_A_PE_4_13__dout;
  wire fifo_A_PE_4_13__empty_n;
  wire fifo_A_PE_4_13__read;
  wire [512:0] fifo_A_PE_4_13__din;
  wire fifo_A_PE_4_13__full_n;
  wire fifo_A_PE_4_13__write;
  wire [512:0] fifo_A_PE_4_14__dout;
  wire fifo_A_PE_4_14__empty_n;
  wire fifo_A_PE_4_14__read;
  wire [512:0] fifo_A_PE_4_14__din;
  wire fifo_A_PE_4_14__full_n;
  wire fifo_A_PE_4_14__write;
  wire [512:0] fifo_A_PE_4_15__dout;
  wire fifo_A_PE_4_15__empty_n;
  wire fifo_A_PE_4_15__read;
  wire [512:0] fifo_A_PE_4_15__din;
  wire fifo_A_PE_4_15__full_n;
  wire fifo_A_PE_4_15__write;
  wire [512:0] fifo_A_PE_4_16__dout;
  wire fifo_A_PE_4_16__empty_n;
  wire fifo_A_PE_4_16__read;
  wire [512:0] fifo_A_PE_4_16__din;
  wire fifo_A_PE_4_16__full_n;
  wire fifo_A_PE_4_16__write;
  wire [512:0] fifo_A_PE_4_17__dout;
  wire fifo_A_PE_4_17__empty_n;
  wire fifo_A_PE_4_17__read;
  wire [512:0] fifo_A_PE_4_17__din;
  wire fifo_A_PE_4_17__full_n;
  wire fifo_A_PE_4_17__write;
  wire [512:0] fifo_A_PE_4_2__dout;
  wire fifo_A_PE_4_2__empty_n;
  wire fifo_A_PE_4_2__read;
  wire [512:0] fifo_A_PE_4_2__din;
  wire fifo_A_PE_4_2__full_n;
  wire fifo_A_PE_4_2__write;
  wire [512:0] fifo_A_PE_4_3__dout;
  wire fifo_A_PE_4_3__empty_n;
  wire fifo_A_PE_4_3__read;
  wire [512:0] fifo_A_PE_4_3__din;
  wire fifo_A_PE_4_3__full_n;
  wire fifo_A_PE_4_3__write;
  wire [512:0] fifo_A_PE_4_4__dout;
  wire fifo_A_PE_4_4__empty_n;
  wire fifo_A_PE_4_4__read;
  wire [512:0] fifo_A_PE_4_4__din;
  wire fifo_A_PE_4_4__full_n;
  wire fifo_A_PE_4_4__write;
  wire [512:0] fifo_A_PE_4_5__dout;
  wire fifo_A_PE_4_5__empty_n;
  wire fifo_A_PE_4_5__read;
  wire [512:0] fifo_A_PE_4_5__din;
  wire fifo_A_PE_4_5__full_n;
  wire fifo_A_PE_4_5__write;
  wire [512:0] fifo_A_PE_4_6__dout;
  wire fifo_A_PE_4_6__empty_n;
  wire fifo_A_PE_4_6__read;
  wire [512:0] fifo_A_PE_4_6__din;
  wire fifo_A_PE_4_6__full_n;
  wire fifo_A_PE_4_6__write;
  wire [512:0] fifo_A_PE_4_7__dout;
  wire fifo_A_PE_4_7__empty_n;
  wire fifo_A_PE_4_7__read;
  wire [512:0] fifo_A_PE_4_7__din;
  wire fifo_A_PE_4_7__full_n;
  wire fifo_A_PE_4_7__write;
  wire [512:0] fifo_A_PE_4_8__dout;
  wire fifo_A_PE_4_8__empty_n;
  wire fifo_A_PE_4_8__read;
  wire [512:0] fifo_A_PE_4_8__din;
  wire fifo_A_PE_4_8__full_n;
  wire fifo_A_PE_4_8__write;
  wire [512:0] fifo_A_PE_4_9__dout;
  wire fifo_A_PE_4_9__empty_n;
  wire fifo_A_PE_4_9__read;
  wire [512:0] fifo_A_PE_4_9__din;
  wire fifo_A_PE_4_9__full_n;
  wire fifo_A_PE_4_9__write;
  wire [512:0] fifo_A_PE_5_0__dout;
  wire fifo_A_PE_5_0__empty_n;
  wire fifo_A_PE_5_0__read;
  wire [512:0] fifo_A_PE_5_0__din;
  wire fifo_A_PE_5_0__full_n;
  wire fifo_A_PE_5_0__write;
  wire [512:0] fifo_A_PE_5_1__dout;
  wire fifo_A_PE_5_1__empty_n;
  wire fifo_A_PE_5_1__read;
  wire [512:0] fifo_A_PE_5_1__din;
  wire fifo_A_PE_5_1__full_n;
  wire fifo_A_PE_5_1__write;
  wire [512:0] fifo_A_PE_5_10__dout;
  wire fifo_A_PE_5_10__empty_n;
  wire fifo_A_PE_5_10__read;
  wire [512:0] fifo_A_PE_5_10__din;
  wire fifo_A_PE_5_10__full_n;
  wire fifo_A_PE_5_10__write;
  wire [512:0] fifo_A_PE_5_11__dout;
  wire fifo_A_PE_5_11__empty_n;
  wire fifo_A_PE_5_11__read;
  wire [512:0] fifo_A_PE_5_11__din;
  wire fifo_A_PE_5_11__full_n;
  wire fifo_A_PE_5_11__write;
  wire [512:0] fifo_A_PE_5_12__dout;
  wire fifo_A_PE_5_12__empty_n;
  wire fifo_A_PE_5_12__read;
  wire [512:0] fifo_A_PE_5_12__din;
  wire fifo_A_PE_5_12__full_n;
  wire fifo_A_PE_5_12__write;
  wire [512:0] fifo_A_PE_5_13__dout;
  wire fifo_A_PE_5_13__empty_n;
  wire fifo_A_PE_5_13__read;
  wire [512:0] fifo_A_PE_5_13__din;
  wire fifo_A_PE_5_13__full_n;
  wire fifo_A_PE_5_13__write;
  wire [512:0] fifo_A_PE_5_14__dout;
  wire fifo_A_PE_5_14__empty_n;
  wire fifo_A_PE_5_14__read;
  wire [512:0] fifo_A_PE_5_14__din;
  wire fifo_A_PE_5_14__full_n;
  wire fifo_A_PE_5_14__write;
  wire [512:0] fifo_A_PE_5_15__dout;
  wire fifo_A_PE_5_15__empty_n;
  wire fifo_A_PE_5_15__read;
  wire [512:0] fifo_A_PE_5_15__din;
  wire fifo_A_PE_5_15__full_n;
  wire fifo_A_PE_5_15__write;
  wire [512:0] fifo_A_PE_5_16__dout;
  wire fifo_A_PE_5_16__empty_n;
  wire fifo_A_PE_5_16__read;
  wire [512:0] fifo_A_PE_5_16__din;
  wire fifo_A_PE_5_16__full_n;
  wire fifo_A_PE_5_16__write;
  wire [512:0] fifo_A_PE_5_17__dout;
  wire fifo_A_PE_5_17__empty_n;
  wire fifo_A_PE_5_17__read;
  wire [512:0] fifo_A_PE_5_17__din;
  wire fifo_A_PE_5_17__full_n;
  wire fifo_A_PE_5_17__write;
  wire [512:0] fifo_A_PE_5_2__dout;
  wire fifo_A_PE_5_2__empty_n;
  wire fifo_A_PE_5_2__read;
  wire [512:0] fifo_A_PE_5_2__din;
  wire fifo_A_PE_5_2__full_n;
  wire fifo_A_PE_5_2__write;
  wire [512:0] fifo_A_PE_5_3__dout;
  wire fifo_A_PE_5_3__empty_n;
  wire fifo_A_PE_5_3__read;
  wire [512:0] fifo_A_PE_5_3__din;
  wire fifo_A_PE_5_3__full_n;
  wire fifo_A_PE_5_3__write;
  wire [512:0] fifo_A_PE_5_4__dout;
  wire fifo_A_PE_5_4__empty_n;
  wire fifo_A_PE_5_4__read;
  wire [512:0] fifo_A_PE_5_4__din;
  wire fifo_A_PE_5_4__full_n;
  wire fifo_A_PE_5_4__write;
  wire [512:0] fifo_A_PE_5_5__dout;
  wire fifo_A_PE_5_5__empty_n;
  wire fifo_A_PE_5_5__read;
  wire [512:0] fifo_A_PE_5_5__din;
  wire fifo_A_PE_5_5__full_n;
  wire fifo_A_PE_5_5__write;
  wire [512:0] fifo_A_PE_5_6__dout;
  wire fifo_A_PE_5_6__empty_n;
  wire fifo_A_PE_5_6__read;
  wire [512:0] fifo_A_PE_5_6__din;
  wire fifo_A_PE_5_6__full_n;
  wire fifo_A_PE_5_6__write;
  wire [512:0] fifo_A_PE_5_7__dout;
  wire fifo_A_PE_5_7__empty_n;
  wire fifo_A_PE_5_7__read;
  wire [512:0] fifo_A_PE_5_7__din;
  wire fifo_A_PE_5_7__full_n;
  wire fifo_A_PE_5_7__write;
  wire [512:0] fifo_A_PE_5_8__dout;
  wire fifo_A_PE_5_8__empty_n;
  wire fifo_A_PE_5_8__read;
  wire [512:0] fifo_A_PE_5_8__din;
  wire fifo_A_PE_5_8__full_n;
  wire fifo_A_PE_5_8__write;
  wire [512:0] fifo_A_PE_5_9__dout;
  wire fifo_A_PE_5_9__empty_n;
  wire fifo_A_PE_5_9__read;
  wire [512:0] fifo_A_PE_5_9__din;
  wire fifo_A_PE_5_9__full_n;
  wire fifo_A_PE_5_9__write;
  wire [512:0] fifo_A_PE_6_0__dout;
  wire fifo_A_PE_6_0__empty_n;
  wire fifo_A_PE_6_0__read;
  wire [512:0] fifo_A_PE_6_0__din;
  wire fifo_A_PE_6_0__full_n;
  wire fifo_A_PE_6_0__write;
  wire [512:0] fifo_A_PE_6_1__dout;
  wire fifo_A_PE_6_1__empty_n;
  wire fifo_A_PE_6_1__read;
  wire [512:0] fifo_A_PE_6_1__din;
  wire fifo_A_PE_6_1__full_n;
  wire fifo_A_PE_6_1__write;
  wire [512:0] fifo_A_PE_6_10__dout;
  wire fifo_A_PE_6_10__empty_n;
  wire fifo_A_PE_6_10__read;
  wire [512:0] fifo_A_PE_6_10__din;
  wire fifo_A_PE_6_10__full_n;
  wire fifo_A_PE_6_10__write;
  wire [512:0] fifo_A_PE_6_11__dout;
  wire fifo_A_PE_6_11__empty_n;
  wire fifo_A_PE_6_11__read;
  wire [512:0] fifo_A_PE_6_11__din;
  wire fifo_A_PE_6_11__full_n;
  wire fifo_A_PE_6_11__write;
  wire [512:0] fifo_A_PE_6_12__dout;
  wire fifo_A_PE_6_12__empty_n;
  wire fifo_A_PE_6_12__read;
  wire [512:0] fifo_A_PE_6_12__din;
  wire fifo_A_PE_6_12__full_n;
  wire fifo_A_PE_6_12__write;
  wire [512:0] fifo_A_PE_6_13__dout;
  wire fifo_A_PE_6_13__empty_n;
  wire fifo_A_PE_6_13__read;
  wire [512:0] fifo_A_PE_6_13__din;
  wire fifo_A_PE_6_13__full_n;
  wire fifo_A_PE_6_13__write;
  wire [512:0] fifo_A_PE_6_14__dout;
  wire fifo_A_PE_6_14__empty_n;
  wire fifo_A_PE_6_14__read;
  wire [512:0] fifo_A_PE_6_14__din;
  wire fifo_A_PE_6_14__full_n;
  wire fifo_A_PE_6_14__write;
  wire [512:0] fifo_A_PE_6_15__dout;
  wire fifo_A_PE_6_15__empty_n;
  wire fifo_A_PE_6_15__read;
  wire [512:0] fifo_A_PE_6_15__din;
  wire fifo_A_PE_6_15__full_n;
  wire fifo_A_PE_6_15__write;
  wire [512:0] fifo_A_PE_6_16__dout;
  wire fifo_A_PE_6_16__empty_n;
  wire fifo_A_PE_6_16__read;
  wire [512:0] fifo_A_PE_6_16__din;
  wire fifo_A_PE_6_16__full_n;
  wire fifo_A_PE_6_16__write;
  wire [512:0] fifo_A_PE_6_17__dout;
  wire fifo_A_PE_6_17__empty_n;
  wire fifo_A_PE_6_17__read;
  wire [512:0] fifo_A_PE_6_17__din;
  wire fifo_A_PE_6_17__full_n;
  wire fifo_A_PE_6_17__write;
  wire [512:0] fifo_A_PE_6_2__dout;
  wire fifo_A_PE_6_2__empty_n;
  wire fifo_A_PE_6_2__read;
  wire [512:0] fifo_A_PE_6_2__din;
  wire fifo_A_PE_6_2__full_n;
  wire fifo_A_PE_6_2__write;
  wire [512:0] fifo_A_PE_6_3__dout;
  wire fifo_A_PE_6_3__empty_n;
  wire fifo_A_PE_6_3__read;
  wire [512:0] fifo_A_PE_6_3__din;
  wire fifo_A_PE_6_3__full_n;
  wire fifo_A_PE_6_3__write;
  wire [512:0] fifo_A_PE_6_4__dout;
  wire fifo_A_PE_6_4__empty_n;
  wire fifo_A_PE_6_4__read;
  wire [512:0] fifo_A_PE_6_4__din;
  wire fifo_A_PE_6_4__full_n;
  wire fifo_A_PE_6_4__write;
  wire [512:0] fifo_A_PE_6_5__dout;
  wire fifo_A_PE_6_5__empty_n;
  wire fifo_A_PE_6_5__read;
  wire [512:0] fifo_A_PE_6_5__din;
  wire fifo_A_PE_6_5__full_n;
  wire fifo_A_PE_6_5__write;
  wire [512:0] fifo_A_PE_6_6__dout;
  wire fifo_A_PE_6_6__empty_n;
  wire fifo_A_PE_6_6__read;
  wire [512:0] fifo_A_PE_6_6__din;
  wire fifo_A_PE_6_6__full_n;
  wire fifo_A_PE_6_6__write;
  wire [512:0] fifo_A_PE_6_7__dout;
  wire fifo_A_PE_6_7__empty_n;
  wire fifo_A_PE_6_7__read;
  wire [512:0] fifo_A_PE_6_7__din;
  wire fifo_A_PE_6_7__full_n;
  wire fifo_A_PE_6_7__write;
  wire [512:0] fifo_A_PE_6_8__dout;
  wire fifo_A_PE_6_8__empty_n;
  wire fifo_A_PE_6_8__read;
  wire [512:0] fifo_A_PE_6_8__din;
  wire fifo_A_PE_6_8__full_n;
  wire fifo_A_PE_6_8__write;
  wire [512:0] fifo_A_PE_6_9__dout;
  wire fifo_A_PE_6_9__empty_n;
  wire fifo_A_PE_6_9__read;
  wire [512:0] fifo_A_PE_6_9__din;
  wire fifo_A_PE_6_9__full_n;
  wire fifo_A_PE_6_9__write;
  wire [512:0] fifo_A_PE_7_0__dout;
  wire fifo_A_PE_7_0__empty_n;
  wire fifo_A_PE_7_0__read;
  wire [512:0] fifo_A_PE_7_0__din;
  wire fifo_A_PE_7_0__full_n;
  wire fifo_A_PE_7_0__write;
  wire [512:0] fifo_A_PE_7_1__dout;
  wire fifo_A_PE_7_1__empty_n;
  wire fifo_A_PE_7_1__read;
  wire [512:0] fifo_A_PE_7_1__din;
  wire fifo_A_PE_7_1__full_n;
  wire fifo_A_PE_7_1__write;
  wire [512:0] fifo_A_PE_7_10__dout;
  wire fifo_A_PE_7_10__empty_n;
  wire fifo_A_PE_7_10__read;
  wire [512:0] fifo_A_PE_7_10__din;
  wire fifo_A_PE_7_10__full_n;
  wire fifo_A_PE_7_10__write;
  wire [512:0] fifo_A_PE_7_11__dout;
  wire fifo_A_PE_7_11__empty_n;
  wire fifo_A_PE_7_11__read;
  wire [512:0] fifo_A_PE_7_11__din;
  wire fifo_A_PE_7_11__full_n;
  wire fifo_A_PE_7_11__write;
  wire [512:0] fifo_A_PE_7_12__dout;
  wire fifo_A_PE_7_12__empty_n;
  wire fifo_A_PE_7_12__read;
  wire [512:0] fifo_A_PE_7_12__din;
  wire fifo_A_PE_7_12__full_n;
  wire fifo_A_PE_7_12__write;
  wire [512:0] fifo_A_PE_7_13__dout;
  wire fifo_A_PE_7_13__empty_n;
  wire fifo_A_PE_7_13__read;
  wire [512:0] fifo_A_PE_7_13__din;
  wire fifo_A_PE_7_13__full_n;
  wire fifo_A_PE_7_13__write;
  wire [512:0] fifo_A_PE_7_14__dout;
  wire fifo_A_PE_7_14__empty_n;
  wire fifo_A_PE_7_14__read;
  wire [512:0] fifo_A_PE_7_14__din;
  wire fifo_A_PE_7_14__full_n;
  wire fifo_A_PE_7_14__write;
  wire [512:0] fifo_A_PE_7_15__dout;
  wire fifo_A_PE_7_15__empty_n;
  wire fifo_A_PE_7_15__read;
  wire [512:0] fifo_A_PE_7_15__din;
  wire fifo_A_PE_7_15__full_n;
  wire fifo_A_PE_7_15__write;
  wire [512:0] fifo_A_PE_7_16__dout;
  wire fifo_A_PE_7_16__empty_n;
  wire fifo_A_PE_7_16__read;
  wire [512:0] fifo_A_PE_7_16__din;
  wire fifo_A_PE_7_16__full_n;
  wire fifo_A_PE_7_16__write;
  wire [512:0] fifo_A_PE_7_17__dout;
  wire fifo_A_PE_7_17__empty_n;
  wire fifo_A_PE_7_17__read;
  wire [512:0] fifo_A_PE_7_17__din;
  wire fifo_A_PE_7_17__full_n;
  wire fifo_A_PE_7_17__write;
  wire [512:0] fifo_A_PE_7_2__dout;
  wire fifo_A_PE_7_2__empty_n;
  wire fifo_A_PE_7_2__read;
  wire [512:0] fifo_A_PE_7_2__din;
  wire fifo_A_PE_7_2__full_n;
  wire fifo_A_PE_7_2__write;
  wire [512:0] fifo_A_PE_7_3__dout;
  wire fifo_A_PE_7_3__empty_n;
  wire fifo_A_PE_7_3__read;
  wire [512:0] fifo_A_PE_7_3__din;
  wire fifo_A_PE_7_3__full_n;
  wire fifo_A_PE_7_3__write;
  wire [512:0] fifo_A_PE_7_4__dout;
  wire fifo_A_PE_7_4__empty_n;
  wire fifo_A_PE_7_4__read;
  wire [512:0] fifo_A_PE_7_4__din;
  wire fifo_A_PE_7_4__full_n;
  wire fifo_A_PE_7_4__write;
  wire [512:0] fifo_A_PE_7_5__dout;
  wire fifo_A_PE_7_5__empty_n;
  wire fifo_A_PE_7_5__read;
  wire [512:0] fifo_A_PE_7_5__din;
  wire fifo_A_PE_7_5__full_n;
  wire fifo_A_PE_7_5__write;
  wire [512:0] fifo_A_PE_7_6__dout;
  wire fifo_A_PE_7_6__empty_n;
  wire fifo_A_PE_7_6__read;
  wire [512:0] fifo_A_PE_7_6__din;
  wire fifo_A_PE_7_6__full_n;
  wire fifo_A_PE_7_6__write;
  wire [512:0] fifo_A_PE_7_7__dout;
  wire fifo_A_PE_7_7__empty_n;
  wire fifo_A_PE_7_7__read;
  wire [512:0] fifo_A_PE_7_7__din;
  wire fifo_A_PE_7_7__full_n;
  wire fifo_A_PE_7_7__write;
  wire [512:0] fifo_A_PE_7_8__dout;
  wire fifo_A_PE_7_8__empty_n;
  wire fifo_A_PE_7_8__read;
  wire [512:0] fifo_A_PE_7_8__din;
  wire fifo_A_PE_7_8__full_n;
  wire fifo_A_PE_7_8__write;
  wire [512:0] fifo_A_PE_7_9__dout;
  wire fifo_A_PE_7_9__empty_n;
  wire fifo_A_PE_7_9__read;
  wire [512:0] fifo_A_PE_7_9__din;
  wire fifo_A_PE_7_9__full_n;
  wire fifo_A_PE_7_9__write;
  wire [512:0] fifo_A_PE_8_0__dout;
  wire fifo_A_PE_8_0__empty_n;
  wire fifo_A_PE_8_0__read;
  wire [512:0] fifo_A_PE_8_0__din;
  wire fifo_A_PE_8_0__full_n;
  wire fifo_A_PE_8_0__write;
  wire [512:0] fifo_A_PE_8_1__dout;
  wire fifo_A_PE_8_1__empty_n;
  wire fifo_A_PE_8_1__read;
  wire [512:0] fifo_A_PE_8_1__din;
  wire fifo_A_PE_8_1__full_n;
  wire fifo_A_PE_8_1__write;
  wire [512:0] fifo_A_PE_8_10__dout;
  wire fifo_A_PE_8_10__empty_n;
  wire fifo_A_PE_8_10__read;
  wire [512:0] fifo_A_PE_8_10__din;
  wire fifo_A_PE_8_10__full_n;
  wire fifo_A_PE_8_10__write;
  wire [512:0] fifo_A_PE_8_11__dout;
  wire fifo_A_PE_8_11__empty_n;
  wire fifo_A_PE_8_11__read;
  wire [512:0] fifo_A_PE_8_11__din;
  wire fifo_A_PE_8_11__full_n;
  wire fifo_A_PE_8_11__write;
  wire [512:0] fifo_A_PE_8_12__dout;
  wire fifo_A_PE_8_12__empty_n;
  wire fifo_A_PE_8_12__read;
  wire [512:0] fifo_A_PE_8_12__din;
  wire fifo_A_PE_8_12__full_n;
  wire fifo_A_PE_8_12__write;
  wire [512:0] fifo_A_PE_8_13__dout;
  wire fifo_A_PE_8_13__empty_n;
  wire fifo_A_PE_8_13__read;
  wire [512:0] fifo_A_PE_8_13__din;
  wire fifo_A_PE_8_13__full_n;
  wire fifo_A_PE_8_13__write;
  wire [512:0] fifo_A_PE_8_14__dout;
  wire fifo_A_PE_8_14__empty_n;
  wire fifo_A_PE_8_14__read;
  wire [512:0] fifo_A_PE_8_14__din;
  wire fifo_A_PE_8_14__full_n;
  wire fifo_A_PE_8_14__write;
  wire [512:0] fifo_A_PE_8_15__dout;
  wire fifo_A_PE_8_15__empty_n;
  wire fifo_A_PE_8_15__read;
  wire [512:0] fifo_A_PE_8_15__din;
  wire fifo_A_PE_8_15__full_n;
  wire fifo_A_PE_8_15__write;
  wire [512:0] fifo_A_PE_8_16__dout;
  wire fifo_A_PE_8_16__empty_n;
  wire fifo_A_PE_8_16__read;
  wire [512:0] fifo_A_PE_8_16__din;
  wire fifo_A_PE_8_16__full_n;
  wire fifo_A_PE_8_16__write;
  wire [512:0] fifo_A_PE_8_17__dout;
  wire fifo_A_PE_8_17__empty_n;
  wire fifo_A_PE_8_17__read;
  wire [512:0] fifo_A_PE_8_17__din;
  wire fifo_A_PE_8_17__full_n;
  wire fifo_A_PE_8_17__write;
  wire [512:0] fifo_A_PE_8_2__dout;
  wire fifo_A_PE_8_2__empty_n;
  wire fifo_A_PE_8_2__read;
  wire [512:0] fifo_A_PE_8_2__din;
  wire fifo_A_PE_8_2__full_n;
  wire fifo_A_PE_8_2__write;
  wire [512:0] fifo_A_PE_8_3__dout;
  wire fifo_A_PE_8_3__empty_n;
  wire fifo_A_PE_8_3__read;
  wire [512:0] fifo_A_PE_8_3__din;
  wire fifo_A_PE_8_3__full_n;
  wire fifo_A_PE_8_3__write;
  wire [512:0] fifo_A_PE_8_4__dout;
  wire fifo_A_PE_8_4__empty_n;
  wire fifo_A_PE_8_4__read;
  wire [512:0] fifo_A_PE_8_4__din;
  wire fifo_A_PE_8_4__full_n;
  wire fifo_A_PE_8_4__write;
  wire [512:0] fifo_A_PE_8_5__dout;
  wire fifo_A_PE_8_5__empty_n;
  wire fifo_A_PE_8_5__read;
  wire [512:0] fifo_A_PE_8_5__din;
  wire fifo_A_PE_8_5__full_n;
  wire fifo_A_PE_8_5__write;
  wire [512:0] fifo_A_PE_8_6__dout;
  wire fifo_A_PE_8_6__empty_n;
  wire fifo_A_PE_8_6__read;
  wire [512:0] fifo_A_PE_8_6__din;
  wire fifo_A_PE_8_6__full_n;
  wire fifo_A_PE_8_6__write;
  wire [512:0] fifo_A_PE_8_7__dout;
  wire fifo_A_PE_8_7__empty_n;
  wire fifo_A_PE_8_7__read;
  wire [512:0] fifo_A_PE_8_7__din;
  wire fifo_A_PE_8_7__full_n;
  wire fifo_A_PE_8_7__write;
  wire [512:0] fifo_A_PE_8_8__dout;
  wire fifo_A_PE_8_8__empty_n;
  wire fifo_A_PE_8_8__read;
  wire [512:0] fifo_A_PE_8_8__din;
  wire fifo_A_PE_8_8__full_n;
  wire fifo_A_PE_8_8__write;
  wire [512:0] fifo_A_PE_8_9__dout;
  wire fifo_A_PE_8_9__empty_n;
  wire fifo_A_PE_8_9__read;
  wire [512:0] fifo_A_PE_8_9__din;
  wire fifo_A_PE_8_9__full_n;
  wire fifo_A_PE_8_9__write;
  wire [512:0] fifo_A_PE_9_0__dout;
  wire fifo_A_PE_9_0__empty_n;
  wire fifo_A_PE_9_0__read;
  wire [512:0] fifo_A_PE_9_0__din;
  wire fifo_A_PE_9_0__full_n;
  wire fifo_A_PE_9_0__write;
  wire [512:0] fifo_A_PE_9_1__dout;
  wire fifo_A_PE_9_1__empty_n;
  wire fifo_A_PE_9_1__read;
  wire [512:0] fifo_A_PE_9_1__din;
  wire fifo_A_PE_9_1__full_n;
  wire fifo_A_PE_9_1__write;
  wire [512:0] fifo_A_PE_9_10__dout;
  wire fifo_A_PE_9_10__empty_n;
  wire fifo_A_PE_9_10__read;
  wire [512:0] fifo_A_PE_9_10__din;
  wire fifo_A_PE_9_10__full_n;
  wire fifo_A_PE_9_10__write;
  wire [512:0] fifo_A_PE_9_11__dout;
  wire fifo_A_PE_9_11__empty_n;
  wire fifo_A_PE_9_11__read;
  wire [512:0] fifo_A_PE_9_11__din;
  wire fifo_A_PE_9_11__full_n;
  wire fifo_A_PE_9_11__write;
  wire [512:0] fifo_A_PE_9_12__dout;
  wire fifo_A_PE_9_12__empty_n;
  wire fifo_A_PE_9_12__read;
  wire [512:0] fifo_A_PE_9_12__din;
  wire fifo_A_PE_9_12__full_n;
  wire fifo_A_PE_9_12__write;
  wire [512:0] fifo_A_PE_9_13__dout;
  wire fifo_A_PE_9_13__empty_n;
  wire fifo_A_PE_9_13__read;
  wire [512:0] fifo_A_PE_9_13__din;
  wire fifo_A_PE_9_13__full_n;
  wire fifo_A_PE_9_13__write;
  wire [512:0] fifo_A_PE_9_14__dout;
  wire fifo_A_PE_9_14__empty_n;
  wire fifo_A_PE_9_14__read;
  wire [512:0] fifo_A_PE_9_14__din;
  wire fifo_A_PE_9_14__full_n;
  wire fifo_A_PE_9_14__write;
  wire [512:0] fifo_A_PE_9_15__dout;
  wire fifo_A_PE_9_15__empty_n;
  wire fifo_A_PE_9_15__read;
  wire [512:0] fifo_A_PE_9_15__din;
  wire fifo_A_PE_9_15__full_n;
  wire fifo_A_PE_9_15__write;
  wire [512:0] fifo_A_PE_9_16__dout;
  wire fifo_A_PE_9_16__empty_n;
  wire fifo_A_PE_9_16__read;
  wire [512:0] fifo_A_PE_9_16__din;
  wire fifo_A_PE_9_16__full_n;
  wire fifo_A_PE_9_16__write;
  wire [512:0] fifo_A_PE_9_17__dout;
  wire fifo_A_PE_9_17__empty_n;
  wire fifo_A_PE_9_17__read;
  wire [512:0] fifo_A_PE_9_17__din;
  wire fifo_A_PE_9_17__full_n;
  wire fifo_A_PE_9_17__write;
  wire [512:0] fifo_A_PE_9_2__dout;
  wire fifo_A_PE_9_2__empty_n;
  wire fifo_A_PE_9_2__read;
  wire [512:0] fifo_A_PE_9_2__din;
  wire fifo_A_PE_9_2__full_n;
  wire fifo_A_PE_9_2__write;
  wire [512:0] fifo_A_PE_9_3__dout;
  wire fifo_A_PE_9_3__empty_n;
  wire fifo_A_PE_9_3__read;
  wire [512:0] fifo_A_PE_9_3__din;
  wire fifo_A_PE_9_3__full_n;
  wire fifo_A_PE_9_3__write;
  wire [512:0] fifo_A_PE_9_4__dout;
  wire fifo_A_PE_9_4__empty_n;
  wire fifo_A_PE_9_4__read;
  wire [512:0] fifo_A_PE_9_4__din;
  wire fifo_A_PE_9_4__full_n;
  wire fifo_A_PE_9_4__write;
  wire [512:0] fifo_A_PE_9_5__dout;
  wire fifo_A_PE_9_5__empty_n;
  wire fifo_A_PE_9_5__read;
  wire [512:0] fifo_A_PE_9_5__din;
  wire fifo_A_PE_9_5__full_n;
  wire fifo_A_PE_9_5__write;
  wire [512:0] fifo_A_PE_9_6__dout;
  wire fifo_A_PE_9_6__empty_n;
  wire fifo_A_PE_9_6__read;
  wire [512:0] fifo_A_PE_9_6__din;
  wire fifo_A_PE_9_6__full_n;
  wire fifo_A_PE_9_6__write;
  wire [512:0] fifo_A_PE_9_7__dout;
  wire fifo_A_PE_9_7__empty_n;
  wire fifo_A_PE_9_7__read;
  wire [512:0] fifo_A_PE_9_7__din;
  wire fifo_A_PE_9_7__full_n;
  wire fifo_A_PE_9_7__write;
  wire [512:0] fifo_A_PE_9_8__dout;
  wire fifo_A_PE_9_8__empty_n;
  wire fifo_A_PE_9_8__read;
  wire [512:0] fifo_A_PE_9_8__din;
  wire fifo_A_PE_9_8__full_n;
  wire fifo_A_PE_9_8__write;
  wire [512:0] fifo_A_PE_9_9__dout;
  wire fifo_A_PE_9_9__empty_n;
  wire fifo_A_PE_9_9__read;
  wire [512:0] fifo_A_PE_9_9__din;
  wire fifo_A_PE_9_9__full_n;
  wire fifo_A_PE_9_9__write;
  wire [512:0] fifo_B_B_IO_L2_in_0__dout;
  wire fifo_B_B_IO_L2_in_0__empty_n;
  wire fifo_B_B_IO_L2_in_0__read;
  wire [512:0] fifo_B_B_IO_L2_in_0__din;
  wire fifo_B_B_IO_L2_in_0__full_n;
  wire fifo_B_B_IO_L2_in_0__write;
  wire [512:0] fifo_B_B_IO_L2_in_1__dout;
  wire fifo_B_B_IO_L2_in_1__empty_n;
  wire fifo_B_B_IO_L2_in_1__read;
  wire [512:0] fifo_B_B_IO_L2_in_1__din;
  wire fifo_B_B_IO_L2_in_1__full_n;
  wire fifo_B_B_IO_L2_in_1__write;
  wire [512:0] fifo_B_B_IO_L2_in_10__dout;
  wire fifo_B_B_IO_L2_in_10__empty_n;
  wire fifo_B_B_IO_L2_in_10__read;
  wire [512:0] fifo_B_B_IO_L2_in_10__din;
  wire fifo_B_B_IO_L2_in_10__full_n;
  wire fifo_B_B_IO_L2_in_10__write;
  wire [512:0] fifo_B_B_IO_L2_in_11__dout;
  wire fifo_B_B_IO_L2_in_11__empty_n;
  wire fifo_B_B_IO_L2_in_11__read;
  wire [512:0] fifo_B_B_IO_L2_in_11__din;
  wire fifo_B_B_IO_L2_in_11__full_n;
  wire fifo_B_B_IO_L2_in_11__write;
  wire [512:0] fifo_B_B_IO_L2_in_12__dout;
  wire fifo_B_B_IO_L2_in_12__empty_n;
  wire fifo_B_B_IO_L2_in_12__read;
  wire [512:0] fifo_B_B_IO_L2_in_12__din;
  wire fifo_B_B_IO_L2_in_12__full_n;
  wire fifo_B_B_IO_L2_in_12__write;
  wire [512:0] fifo_B_B_IO_L2_in_13__dout;
  wire fifo_B_B_IO_L2_in_13__empty_n;
  wire fifo_B_B_IO_L2_in_13__read;
  wire [512:0] fifo_B_B_IO_L2_in_13__din;
  wire fifo_B_B_IO_L2_in_13__full_n;
  wire fifo_B_B_IO_L2_in_13__write;
  wire [512:0] fifo_B_B_IO_L2_in_14__dout;
  wire fifo_B_B_IO_L2_in_14__empty_n;
  wire fifo_B_B_IO_L2_in_14__read;
  wire [512:0] fifo_B_B_IO_L2_in_14__din;
  wire fifo_B_B_IO_L2_in_14__full_n;
  wire fifo_B_B_IO_L2_in_14__write;
  wire [512:0] fifo_B_B_IO_L2_in_15__dout;
  wire fifo_B_B_IO_L2_in_15__empty_n;
  wire fifo_B_B_IO_L2_in_15__read;
  wire [512:0] fifo_B_B_IO_L2_in_15__din;
  wire fifo_B_B_IO_L2_in_15__full_n;
  wire fifo_B_B_IO_L2_in_15__write;
  wire [512:0] fifo_B_B_IO_L2_in_16__dout;
  wire fifo_B_B_IO_L2_in_16__empty_n;
  wire fifo_B_B_IO_L2_in_16__read;
  wire [512:0] fifo_B_B_IO_L2_in_16__din;
  wire fifo_B_B_IO_L2_in_16__full_n;
  wire fifo_B_B_IO_L2_in_16__write;
  wire [512:0] fifo_B_B_IO_L2_in_2__dout;
  wire fifo_B_B_IO_L2_in_2__empty_n;
  wire fifo_B_B_IO_L2_in_2__read;
  wire [512:0] fifo_B_B_IO_L2_in_2__din;
  wire fifo_B_B_IO_L2_in_2__full_n;
  wire fifo_B_B_IO_L2_in_2__write;
  wire [512:0] fifo_B_B_IO_L2_in_3__dout;
  wire fifo_B_B_IO_L2_in_3__empty_n;
  wire fifo_B_B_IO_L2_in_3__read;
  wire [512:0] fifo_B_B_IO_L2_in_3__din;
  wire fifo_B_B_IO_L2_in_3__full_n;
  wire fifo_B_B_IO_L2_in_3__write;
  wire [512:0] fifo_B_B_IO_L2_in_4__dout;
  wire fifo_B_B_IO_L2_in_4__empty_n;
  wire fifo_B_B_IO_L2_in_4__read;
  wire [512:0] fifo_B_B_IO_L2_in_4__din;
  wire fifo_B_B_IO_L2_in_4__full_n;
  wire fifo_B_B_IO_L2_in_4__write;
  wire [512:0] fifo_B_B_IO_L2_in_5__dout;
  wire fifo_B_B_IO_L2_in_5__empty_n;
  wire fifo_B_B_IO_L2_in_5__read;
  wire [512:0] fifo_B_B_IO_L2_in_5__din;
  wire fifo_B_B_IO_L2_in_5__full_n;
  wire fifo_B_B_IO_L2_in_5__write;
  wire [512:0] fifo_B_B_IO_L2_in_6__dout;
  wire fifo_B_B_IO_L2_in_6__empty_n;
  wire fifo_B_B_IO_L2_in_6__read;
  wire [512:0] fifo_B_B_IO_L2_in_6__din;
  wire fifo_B_B_IO_L2_in_6__full_n;
  wire fifo_B_B_IO_L2_in_6__write;
  wire [512:0] fifo_B_B_IO_L2_in_7__dout;
  wire fifo_B_B_IO_L2_in_7__empty_n;
  wire fifo_B_B_IO_L2_in_7__read;
  wire [512:0] fifo_B_B_IO_L2_in_7__din;
  wire fifo_B_B_IO_L2_in_7__full_n;
  wire fifo_B_B_IO_L2_in_7__write;
  wire [512:0] fifo_B_B_IO_L2_in_8__dout;
  wire fifo_B_B_IO_L2_in_8__empty_n;
  wire fifo_B_B_IO_L2_in_8__read;
  wire [512:0] fifo_B_B_IO_L2_in_8__din;
  wire fifo_B_B_IO_L2_in_8__full_n;
  wire fifo_B_B_IO_L2_in_8__write;
  wire [512:0] fifo_B_B_IO_L2_in_9__dout;
  wire fifo_B_B_IO_L2_in_9__empty_n;
  wire fifo_B_B_IO_L2_in_9__read;
  wire [512:0] fifo_B_B_IO_L2_in_9__din;
  wire fifo_B_B_IO_L2_in_9__full_n;
  wire fifo_B_B_IO_L2_in_9__write;
  wire [512:0] fifo_B_B_IO_L3_in_serialize__dout;
  wire fifo_B_B_IO_L3_in_serialize__empty_n;
  wire fifo_B_B_IO_L3_in_serialize__read;
  wire [512:0] fifo_B_B_IO_L3_in_serialize__din;
  wire fifo_B_B_IO_L3_in_serialize__full_n;
  wire fifo_B_B_IO_L3_in_serialize__write;
  wire [512:0] fifo_B_PE_0_0__dout;
  wire fifo_B_PE_0_0__empty_n;
  wire fifo_B_PE_0_0__read;
  wire [512:0] fifo_B_PE_0_0__din;
  wire fifo_B_PE_0_0__full_n;
  wire fifo_B_PE_0_0__write;
  wire [512:0] fifo_B_PE_0_1__dout;
  wire fifo_B_PE_0_1__empty_n;
  wire fifo_B_PE_0_1__read;
  wire [512:0] fifo_B_PE_0_1__din;
  wire fifo_B_PE_0_1__full_n;
  wire fifo_B_PE_0_1__write;
  wire [512:0] fifo_B_PE_0_10__dout;
  wire fifo_B_PE_0_10__empty_n;
  wire fifo_B_PE_0_10__read;
  wire [512:0] fifo_B_PE_0_10__din;
  wire fifo_B_PE_0_10__full_n;
  wire fifo_B_PE_0_10__write;
  wire [512:0] fifo_B_PE_0_11__dout;
  wire fifo_B_PE_0_11__empty_n;
  wire fifo_B_PE_0_11__read;
  wire [512:0] fifo_B_PE_0_11__din;
  wire fifo_B_PE_0_11__full_n;
  wire fifo_B_PE_0_11__write;
  wire [512:0] fifo_B_PE_0_12__dout;
  wire fifo_B_PE_0_12__empty_n;
  wire fifo_B_PE_0_12__read;
  wire [512:0] fifo_B_PE_0_12__din;
  wire fifo_B_PE_0_12__full_n;
  wire fifo_B_PE_0_12__write;
  wire [512:0] fifo_B_PE_0_13__dout;
  wire fifo_B_PE_0_13__empty_n;
  wire fifo_B_PE_0_13__read;
  wire [512:0] fifo_B_PE_0_13__din;
  wire fifo_B_PE_0_13__full_n;
  wire fifo_B_PE_0_13__write;
  wire [512:0] fifo_B_PE_0_14__dout;
  wire fifo_B_PE_0_14__empty_n;
  wire fifo_B_PE_0_14__read;
  wire [512:0] fifo_B_PE_0_14__din;
  wire fifo_B_PE_0_14__full_n;
  wire fifo_B_PE_0_14__write;
  wire [512:0] fifo_B_PE_0_15__dout;
  wire fifo_B_PE_0_15__empty_n;
  wire fifo_B_PE_0_15__read;
  wire [512:0] fifo_B_PE_0_15__din;
  wire fifo_B_PE_0_15__full_n;
  wire fifo_B_PE_0_15__write;
  wire [512:0] fifo_B_PE_0_16__dout;
  wire fifo_B_PE_0_16__empty_n;
  wire fifo_B_PE_0_16__read;
  wire [512:0] fifo_B_PE_0_16__din;
  wire fifo_B_PE_0_16__full_n;
  wire fifo_B_PE_0_16__write;
  wire [512:0] fifo_B_PE_0_2__dout;
  wire fifo_B_PE_0_2__empty_n;
  wire fifo_B_PE_0_2__read;
  wire [512:0] fifo_B_PE_0_2__din;
  wire fifo_B_PE_0_2__full_n;
  wire fifo_B_PE_0_2__write;
  wire [512:0] fifo_B_PE_0_3__dout;
  wire fifo_B_PE_0_3__empty_n;
  wire fifo_B_PE_0_3__read;
  wire [512:0] fifo_B_PE_0_3__din;
  wire fifo_B_PE_0_3__full_n;
  wire fifo_B_PE_0_3__write;
  wire [512:0] fifo_B_PE_0_4__dout;
  wire fifo_B_PE_0_4__empty_n;
  wire fifo_B_PE_0_4__read;
  wire [512:0] fifo_B_PE_0_4__din;
  wire fifo_B_PE_0_4__full_n;
  wire fifo_B_PE_0_4__write;
  wire [512:0] fifo_B_PE_0_5__dout;
  wire fifo_B_PE_0_5__empty_n;
  wire fifo_B_PE_0_5__read;
  wire [512:0] fifo_B_PE_0_5__din;
  wire fifo_B_PE_0_5__full_n;
  wire fifo_B_PE_0_5__write;
  wire [512:0] fifo_B_PE_0_6__dout;
  wire fifo_B_PE_0_6__empty_n;
  wire fifo_B_PE_0_6__read;
  wire [512:0] fifo_B_PE_0_6__din;
  wire fifo_B_PE_0_6__full_n;
  wire fifo_B_PE_0_6__write;
  wire [512:0] fifo_B_PE_0_7__dout;
  wire fifo_B_PE_0_7__empty_n;
  wire fifo_B_PE_0_7__read;
  wire [512:0] fifo_B_PE_0_7__din;
  wire fifo_B_PE_0_7__full_n;
  wire fifo_B_PE_0_7__write;
  wire [512:0] fifo_B_PE_0_8__dout;
  wire fifo_B_PE_0_8__empty_n;
  wire fifo_B_PE_0_8__read;
  wire [512:0] fifo_B_PE_0_8__din;
  wire fifo_B_PE_0_8__full_n;
  wire fifo_B_PE_0_8__write;
  wire [512:0] fifo_B_PE_0_9__dout;
  wire fifo_B_PE_0_9__empty_n;
  wire fifo_B_PE_0_9__read;
  wire [512:0] fifo_B_PE_0_9__din;
  wire fifo_B_PE_0_9__full_n;
  wire fifo_B_PE_0_9__write;
  wire [512:0] fifo_B_PE_10_0__dout;
  wire fifo_B_PE_10_0__empty_n;
  wire fifo_B_PE_10_0__read;
  wire [512:0] fifo_B_PE_10_0__din;
  wire fifo_B_PE_10_0__full_n;
  wire fifo_B_PE_10_0__write;
  wire [512:0] fifo_B_PE_10_1__dout;
  wire fifo_B_PE_10_1__empty_n;
  wire fifo_B_PE_10_1__read;
  wire [512:0] fifo_B_PE_10_1__din;
  wire fifo_B_PE_10_1__full_n;
  wire fifo_B_PE_10_1__write;
  wire [512:0] fifo_B_PE_10_10__dout;
  wire fifo_B_PE_10_10__empty_n;
  wire fifo_B_PE_10_10__read;
  wire [512:0] fifo_B_PE_10_10__din;
  wire fifo_B_PE_10_10__full_n;
  wire fifo_B_PE_10_10__write;
  wire [512:0] fifo_B_PE_10_11__dout;
  wire fifo_B_PE_10_11__empty_n;
  wire fifo_B_PE_10_11__read;
  wire [512:0] fifo_B_PE_10_11__din;
  wire fifo_B_PE_10_11__full_n;
  wire fifo_B_PE_10_11__write;
  wire [512:0] fifo_B_PE_10_12__dout;
  wire fifo_B_PE_10_12__empty_n;
  wire fifo_B_PE_10_12__read;
  wire [512:0] fifo_B_PE_10_12__din;
  wire fifo_B_PE_10_12__full_n;
  wire fifo_B_PE_10_12__write;
  wire [512:0] fifo_B_PE_10_13__dout;
  wire fifo_B_PE_10_13__empty_n;
  wire fifo_B_PE_10_13__read;
  wire [512:0] fifo_B_PE_10_13__din;
  wire fifo_B_PE_10_13__full_n;
  wire fifo_B_PE_10_13__write;
  wire [512:0] fifo_B_PE_10_14__dout;
  wire fifo_B_PE_10_14__empty_n;
  wire fifo_B_PE_10_14__read;
  wire [512:0] fifo_B_PE_10_14__din;
  wire fifo_B_PE_10_14__full_n;
  wire fifo_B_PE_10_14__write;
  wire [512:0] fifo_B_PE_10_15__dout;
  wire fifo_B_PE_10_15__empty_n;
  wire fifo_B_PE_10_15__read;
  wire [512:0] fifo_B_PE_10_15__din;
  wire fifo_B_PE_10_15__full_n;
  wire fifo_B_PE_10_15__write;
  wire [512:0] fifo_B_PE_10_16__dout;
  wire fifo_B_PE_10_16__empty_n;
  wire fifo_B_PE_10_16__read;
  wire [512:0] fifo_B_PE_10_16__din;
  wire fifo_B_PE_10_16__full_n;
  wire fifo_B_PE_10_16__write;
  wire [512:0] fifo_B_PE_10_2__dout;
  wire fifo_B_PE_10_2__empty_n;
  wire fifo_B_PE_10_2__read;
  wire [512:0] fifo_B_PE_10_2__din;
  wire fifo_B_PE_10_2__full_n;
  wire fifo_B_PE_10_2__write;
  wire [512:0] fifo_B_PE_10_3__dout;
  wire fifo_B_PE_10_3__empty_n;
  wire fifo_B_PE_10_3__read;
  wire [512:0] fifo_B_PE_10_3__din;
  wire fifo_B_PE_10_3__full_n;
  wire fifo_B_PE_10_3__write;
  wire [512:0] fifo_B_PE_10_4__dout;
  wire fifo_B_PE_10_4__empty_n;
  wire fifo_B_PE_10_4__read;
  wire [512:0] fifo_B_PE_10_4__din;
  wire fifo_B_PE_10_4__full_n;
  wire fifo_B_PE_10_4__write;
  wire [512:0] fifo_B_PE_10_5__dout;
  wire fifo_B_PE_10_5__empty_n;
  wire fifo_B_PE_10_5__read;
  wire [512:0] fifo_B_PE_10_5__din;
  wire fifo_B_PE_10_5__full_n;
  wire fifo_B_PE_10_5__write;
  wire [512:0] fifo_B_PE_10_6__dout;
  wire fifo_B_PE_10_6__empty_n;
  wire fifo_B_PE_10_6__read;
  wire [512:0] fifo_B_PE_10_6__din;
  wire fifo_B_PE_10_6__full_n;
  wire fifo_B_PE_10_6__write;
  wire [512:0] fifo_B_PE_10_7__dout;
  wire fifo_B_PE_10_7__empty_n;
  wire fifo_B_PE_10_7__read;
  wire [512:0] fifo_B_PE_10_7__din;
  wire fifo_B_PE_10_7__full_n;
  wire fifo_B_PE_10_7__write;
  wire [512:0] fifo_B_PE_10_8__dout;
  wire fifo_B_PE_10_8__empty_n;
  wire fifo_B_PE_10_8__read;
  wire [512:0] fifo_B_PE_10_8__din;
  wire fifo_B_PE_10_8__full_n;
  wire fifo_B_PE_10_8__write;
  wire [512:0] fifo_B_PE_10_9__dout;
  wire fifo_B_PE_10_9__empty_n;
  wire fifo_B_PE_10_9__read;
  wire [512:0] fifo_B_PE_10_9__din;
  wire fifo_B_PE_10_9__full_n;
  wire fifo_B_PE_10_9__write;
  wire [512:0] fifo_B_PE_11_0__dout;
  wire fifo_B_PE_11_0__empty_n;
  wire fifo_B_PE_11_0__read;
  wire [512:0] fifo_B_PE_11_0__din;
  wire fifo_B_PE_11_0__full_n;
  wire fifo_B_PE_11_0__write;
  wire [512:0] fifo_B_PE_11_1__dout;
  wire fifo_B_PE_11_1__empty_n;
  wire fifo_B_PE_11_1__read;
  wire [512:0] fifo_B_PE_11_1__din;
  wire fifo_B_PE_11_1__full_n;
  wire fifo_B_PE_11_1__write;
  wire [512:0] fifo_B_PE_11_10__dout;
  wire fifo_B_PE_11_10__empty_n;
  wire fifo_B_PE_11_10__read;
  wire [512:0] fifo_B_PE_11_10__din;
  wire fifo_B_PE_11_10__full_n;
  wire fifo_B_PE_11_10__write;
  wire [512:0] fifo_B_PE_11_11__dout;
  wire fifo_B_PE_11_11__empty_n;
  wire fifo_B_PE_11_11__read;
  wire [512:0] fifo_B_PE_11_11__din;
  wire fifo_B_PE_11_11__full_n;
  wire fifo_B_PE_11_11__write;
  wire [512:0] fifo_B_PE_11_12__dout;
  wire fifo_B_PE_11_12__empty_n;
  wire fifo_B_PE_11_12__read;
  wire [512:0] fifo_B_PE_11_12__din;
  wire fifo_B_PE_11_12__full_n;
  wire fifo_B_PE_11_12__write;
  wire [512:0] fifo_B_PE_11_13__dout;
  wire fifo_B_PE_11_13__empty_n;
  wire fifo_B_PE_11_13__read;
  wire [512:0] fifo_B_PE_11_13__din;
  wire fifo_B_PE_11_13__full_n;
  wire fifo_B_PE_11_13__write;
  wire [512:0] fifo_B_PE_11_14__dout;
  wire fifo_B_PE_11_14__empty_n;
  wire fifo_B_PE_11_14__read;
  wire [512:0] fifo_B_PE_11_14__din;
  wire fifo_B_PE_11_14__full_n;
  wire fifo_B_PE_11_14__write;
  wire [512:0] fifo_B_PE_11_15__dout;
  wire fifo_B_PE_11_15__empty_n;
  wire fifo_B_PE_11_15__read;
  wire [512:0] fifo_B_PE_11_15__din;
  wire fifo_B_PE_11_15__full_n;
  wire fifo_B_PE_11_15__write;
  wire [512:0] fifo_B_PE_11_16__dout;
  wire fifo_B_PE_11_16__empty_n;
  wire fifo_B_PE_11_16__read;
  wire [512:0] fifo_B_PE_11_16__din;
  wire fifo_B_PE_11_16__full_n;
  wire fifo_B_PE_11_16__write;
  wire [512:0] fifo_B_PE_11_2__dout;
  wire fifo_B_PE_11_2__empty_n;
  wire fifo_B_PE_11_2__read;
  wire [512:0] fifo_B_PE_11_2__din;
  wire fifo_B_PE_11_2__full_n;
  wire fifo_B_PE_11_2__write;
  wire [512:0] fifo_B_PE_11_3__dout;
  wire fifo_B_PE_11_3__empty_n;
  wire fifo_B_PE_11_3__read;
  wire [512:0] fifo_B_PE_11_3__din;
  wire fifo_B_PE_11_3__full_n;
  wire fifo_B_PE_11_3__write;
  wire [512:0] fifo_B_PE_11_4__dout;
  wire fifo_B_PE_11_4__empty_n;
  wire fifo_B_PE_11_4__read;
  wire [512:0] fifo_B_PE_11_4__din;
  wire fifo_B_PE_11_4__full_n;
  wire fifo_B_PE_11_4__write;
  wire [512:0] fifo_B_PE_11_5__dout;
  wire fifo_B_PE_11_5__empty_n;
  wire fifo_B_PE_11_5__read;
  wire [512:0] fifo_B_PE_11_5__din;
  wire fifo_B_PE_11_5__full_n;
  wire fifo_B_PE_11_5__write;
  wire [512:0] fifo_B_PE_11_6__dout;
  wire fifo_B_PE_11_6__empty_n;
  wire fifo_B_PE_11_6__read;
  wire [512:0] fifo_B_PE_11_6__din;
  wire fifo_B_PE_11_6__full_n;
  wire fifo_B_PE_11_6__write;
  wire [512:0] fifo_B_PE_11_7__dout;
  wire fifo_B_PE_11_7__empty_n;
  wire fifo_B_PE_11_7__read;
  wire [512:0] fifo_B_PE_11_7__din;
  wire fifo_B_PE_11_7__full_n;
  wire fifo_B_PE_11_7__write;
  wire [512:0] fifo_B_PE_11_8__dout;
  wire fifo_B_PE_11_8__empty_n;
  wire fifo_B_PE_11_8__read;
  wire [512:0] fifo_B_PE_11_8__din;
  wire fifo_B_PE_11_8__full_n;
  wire fifo_B_PE_11_8__write;
  wire [512:0] fifo_B_PE_11_9__dout;
  wire fifo_B_PE_11_9__empty_n;
  wire fifo_B_PE_11_9__read;
  wire [512:0] fifo_B_PE_11_9__din;
  wire fifo_B_PE_11_9__full_n;
  wire fifo_B_PE_11_9__write;
  wire [512:0] fifo_B_PE_12_0__dout;
  wire fifo_B_PE_12_0__empty_n;
  wire fifo_B_PE_12_0__read;
  wire [512:0] fifo_B_PE_12_0__din;
  wire fifo_B_PE_12_0__full_n;
  wire fifo_B_PE_12_0__write;
  wire [512:0] fifo_B_PE_12_1__dout;
  wire fifo_B_PE_12_1__empty_n;
  wire fifo_B_PE_12_1__read;
  wire [512:0] fifo_B_PE_12_1__din;
  wire fifo_B_PE_12_1__full_n;
  wire fifo_B_PE_12_1__write;
  wire [512:0] fifo_B_PE_12_10__dout;
  wire fifo_B_PE_12_10__empty_n;
  wire fifo_B_PE_12_10__read;
  wire [512:0] fifo_B_PE_12_10__din;
  wire fifo_B_PE_12_10__full_n;
  wire fifo_B_PE_12_10__write;
  wire [512:0] fifo_B_PE_12_11__dout;
  wire fifo_B_PE_12_11__empty_n;
  wire fifo_B_PE_12_11__read;
  wire [512:0] fifo_B_PE_12_11__din;
  wire fifo_B_PE_12_11__full_n;
  wire fifo_B_PE_12_11__write;
  wire [512:0] fifo_B_PE_12_12__dout;
  wire fifo_B_PE_12_12__empty_n;
  wire fifo_B_PE_12_12__read;
  wire [512:0] fifo_B_PE_12_12__din;
  wire fifo_B_PE_12_12__full_n;
  wire fifo_B_PE_12_12__write;
  wire [512:0] fifo_B_PE_12_13__dout;
  wire fifo_B_PE_12_13__empty_n;
  wire fifo_B_PE_12_13__read;
  wire [512:0] fifo_B_PE_12_13__din;
  wire fifo_B_PE_12_13__full_n;
  wire fifo_B_PE_12_13__write;
  wire [512:0] fifo_B_PE_12_14__dout;
  wire fifo_B_PE_12_14__empty_n;
  wire fifo_B_PE_12_14__read;
  wire [512:0] fifo_B_PE_12_14__din;
  wire fifo_B_PE_12_14__full_n;
  wire fifo_B_PE_12_14__write;
  wire [512:0] fifo_B_PE_12_15__dout;
  wire fifo_B_PE_12_15__empty_n;
  wire fifo_B_PE_12_15__read;
  wire [512:0] fifo_B_PE_12_15__din;
  wire fifo_B_PE_12_15__full_n;
  wire fifo_B_PE_12_15__write;
  wire [512:0] fifo_B_PE_12_16__dout;
  wire fifo_B_PE_12_16__empty_n;
  wire fifo_B_PE_12_16__read;
  wire [512:0] fifo_B_PE_12_16__din;
  wire fifo_B_PE_12_16__full_n;
  wire fifo_B_PE_12_16__write;
  wire [512:0] fifo_B_PE_12_2__dout;
  wire fifo_B_PE_12_2__empty_n;
  wire fifo_B_PE_12_2__read;
  wire [512:0] fifo_B_PE_12_2__din;
  wire fifo_B_PE_12_2__full_n;
  wire fifo_B_PE_12_2__write;
  wire [512:0] fifo_B_PE_12_3__dout;
  wire fifo_B_PE_12_3__empty_n;
  wire fifo_B_PE_12_3__read;
  wire [512:0] fifo_B_PE_12_3__din;
  wire fifo_B_PE_12_3__full_n;
  wire fifo_B_PE_12_3__write;
  wire [512:0] fifo_B_PE_12_4__dout;
  wire fifo_B_PE_12_4__empty_n;
  wire fifo_B_PE_12_4__read;
  wire [512:0] fifo_B_PE_12_4__din;
  wire fifo_B_PE_12_4__full_n;
  wire fifo_B_PE_12_4__write;
  wire [512:0] fifo_B_PE_12_5__dout;
  wire fifo_B_PE_12_5__empty_n;
  wire fifo_B_PE_12_5__read;
  wire [512:0] fifo_B_PE_12_5__din;
  wire fifo_B_PE_12_5__full_n;
  wire fifo_B_PE_12_5__write;
  wire [512:0] fifo_B_PE_12_6__dout;
  wire fifo_B_PE_12_6__empty_n;
  wire fifo_B_PE_12_6__read;
  wire [512:0] fifo_B_PE_12_6__din;
  wire fifo_B_PE_12_6__full_n;
  wire fifo_B_PE_12_6__write;
  wire [512:0] fifo_B_PE_12_7__dout;
  wire fifo_B_PE_12_7__empty_n;
  wire fifo_B_PE_12_7__read;
  wire [512:0] fifo_B_PE_12_7__din;
  wire fifo_B_PE_12_7__full_n;
  wire fifo_B_PE_12_7__write;
  wire [512:0] fifo_B_PE_12_8__dout;
  wire fifo_B_PE_12_8__empty_n;
  wire fifo_B_PE_12_8__read;
  wire [512:0] fifo_B_PE_12_8__din;
  wire fifo_B_PE_12_8__full_n;
  wire fifo_B_PE_12_8__write;
  wire [512:0] fifo_B_PE_12_9__dout;
  wire fifo_B_PE_12_9__empty_n;
  wire fifo_B_PE_12_9__read;
  wire [512:0] fifo_B_PE_12_9__din;
  wire fifo_B_PE_12_9__full_n;
  wire fifo_B_PE_12_9__write;
  wire [512:0] fifo_B_PE_13_0__dout;
  wire fifo_B_PE_13_0__empty_n;
  wire fifo_B_PE_13_0__read;
  wire [512:0] fifo_B_PE_13_0__din;
  wire fifo_B_PE_13_0__full_n;
  wire fifo_B_PE_13_0__write;
  wire [512:0] fifo_B_PE_13_1__dout;
  wire fifo_B_PE_13_1__empty_n;
  wire fifo_B_PE_13_1__read;
  wire [512:0] fifo_B_PE_13_1__din;
  wire fifo_B_PE_13_1__full_n;
  wire fifo_B_PE_13_1__write;
  wire [512:0] fifo_B_PE_13_10__dout;
  wire fifo_B_PE_13_10__empty_n;
  wire fifo_B_PE_13_10__read;
  wire [512:0] fifo_B_PE_13_10__din;
  wire fifo_B_PE_13_10__full_n;
  wire fifo_B_PE_13_10__write;
  wire [512:0] fifo_B_PE_13_11__dout;
  wire fifo_B_PE_13_11__empty_n;
  wire fifo_B_PE_13_11__read;
  wire [512:0] fifo_B_PE_13_11__din;
  wire fifo_B_PE_13_11__full_n;
  wire fifo_B_PE_13_11__write;
  wire [512:0] fifo_B_PE_13_12__dout;
  wire fifo_B_PE_13_12__empty_n;
  wire fifo_B_PE_13_12__read;
  wire [512:0] fifo_B_PE_13_12__din;
  wire fifo_B_PE_13_12__full_n;
  wire fifo_B_PE_13_12__write;
  wire [512:0] fifo_B_PE_13_13__dout;
  wire fifo_B_PE_13_13__empty_n;
  wire fifo_B_PE_13_13__read;
  wire [512:0] fifo_B_PE_13_13__din;
  wire fifo_B_PE_13_13__full_n;
  wire fifo_B_PE_13_13__write;
  wire [512:0] fifo_B_PE_13_14__dout;
  wire fifo_B_PE_13_14__empty_n;
  wire fifo_B_PE_13_14__read;
  wire [512:0] fifo_B_PE_13_14__din;
  wire fifo_B_PE_13_14__full_n;
  wire fifo_B_PE_13_14__write;
  wire [512:0] fifo_B_PE_13_15__dout;
  wire fifo_B_PE_13_15__empty_n;
  wire fifo_B_PE_13_15__read;
  wire [512:0] fifo_B_PE_13_15__din;
  wire fifo_B_PE_13_15__full_n;
  wire fifo_B_PE_13_15__write;
  wire [512:0] fifo_B_PE_13_16__dout;
  wire fifo_B_PE_13_16__empty_n;
  wire fifo_B_PE_13_16__read;
  wire [512:0] fifo_B_PE_13_16__din;
  wire fifo_B_PE_13_16__full_n;
  wire fifo_B_PE_13_16__write;
  wire [512:0] fifo_B_PE_13_2__dout;
  wire fifo_B_PE_13_2__empty_n;
  wire fifo_B_PE_13_2__read;
  wire [512:0] fifo_B_PE_13_2__din;
  wire fifo_B_PE_13_2__full_n;
  wire fifo_B_PE_13_2__write;
  wire [512:0] fifo_B_PE_13_3__dout;
  wire fifo_B_PE_13_3__empty_n;
  wire fifo_B_PE_13_3__read;
  wire [512:0] fifo_B_PE_13_3__din;
  wire fifo_B_PE_13_3__full_n;
  wire fifo_B_PE_13_3__write;
  wire [512:0] fifo_B_PE_13_4__dout;
  wire fifo_B_PE_13_4__empty_n;
  wire fifo_B_PE_13_4__read;
  wire [512:0] fifo_B_PE_13_4__din;
  wire fifo_B_PE_13_4__full_n;
  wire fifo_B_PE_13_4__write;
  wire [512:0] fifo_B_PE_13_5__dout;
  wire fifo_B_PE_13_5__empty_n;
  wire fifo_B_PE_13_5__read;
  wire [512:0] fifo_B_PE_13_5__din;
  wire fifo_B_PE_13_5__full_n;
  wire fifo_B_PE_13_5__write;
  wire [512:0] fifo_B_PE_13_6__dout;
  wire fifo_B_PE_13_6__empty_n;
  wire fifo_B_PE_13_6__read;
  wire [512:0] fifo_B_PE_13_6__din;
  wire fifo_B_PE_13_6__full_n;
  wire fifo_B_PE_13_6__write;
  wire [512:0] fifo_B_PE_13_7__dout;
  wire fifo_B_PE_13_7__empty_n;
  wire fifo_B_PE_13_7__read;
  wire [512:0] fifo_B_PE_13_7__din;
  wire fifo_B_PE_13_7__full_n;
  wire fifo_B_PE_13_7__write;
  wire [512:0] fifo_B_PE_13_8__dout;
  wire fifo_B_PE_13_8__empty_n;
  wire fifo_B_PE_13_8__read;
  wire [512:0] fifo_B_PE_13_8__din;
  wire fifo_B_PE_13_8__full_n;
  wire fifo_B_PE_13_8__write;
  wire [512:0] fifo_B_PE_13_9__dout;
  wire fifo_B_PE_13_9__empty_n;
  wire fifo_B_PE_13_9__read;
  wire [512:0] fifo_B_PE_13_9__din;
  wire fifo_B_PE_13_9__full_n;
  wire fifo_B_PE_13_9__write;
  wire [512:0] fifo_B_PE_14_0__dout;
  wire fifo_B_PE_14_0__empty_n;
  wire fifo_B_PE_14_0__read;
  wire [512:0] fifo_B_PE_14_0__din;
  wire fifo_B_PE_14_0__full_n;
  wire fifo_B_PE_14_0__write;
  wire [512:0] fifo_B_PE_14_1__dout;
  wire fifo_B_PE_14_1__empty_n;
  wire fifo_B_PE_14_1__read;
  wire [512:0] fifo_B_PE_14_1__din;
  wire fifo_B_PE_14_1__full_n;
  wire fifo_B_PE_14_1__write;
  wire [512:0] fifo_B_PE_14_10__dout;
  wire fifo_B_PE_14_10__empty_n;
  wire fifo_B_PE_14_10__read;
  wire [512:0] fifo_B_PE_14_10__din;
  wire fifo_B_PE_14_10__full_n;
  wire fifo_B_PE_14_10__write;
  wire [512:0] fifo_B_PE_14_11__dout;
  wire fifo_B_PE_14_11__empty_n;
  wire fifo_B_PE_14_11__read;
  wire [512:0] fifo_B_PE_14_11__din;
  wire fifo_B_PE_14_11__full_n;
  wire fifo_B_PE_14_11__write;
  wire [512:0] fifo_B_PE_14_12__dout;
  wire fifo_B_PE_14_12__empty_n;
  wire fifo_B_PE_14_12__read;
  wire [512:0] fifo_B_PE_14_12__din;
  wire fifo_B_PE_14_12__full_n;
  wire fifo_B_PE_14_12__write;
  wire [512:0] fifo_B_PE_14_13__dout;
  wire fifo_B_PE_14_13__empty_n;
  wire fifo_B_PE_14_13__read;
  wire [512:0] fifo_B_PE_14_13__din;
  wire fifo_B_PE_14_13__full_n;
  wire fifo_B_PE_14_13__write;
  wire [512:0] fifo_B_PE_14_14__dout;
  wire fifo_B_PE_14_14__empty_n;
  wire fifo_B_PE_14_14__read;
  wire [512:0] fifo_B_PE_14_14__din;
  wire fifo_B_PE_14_14__full_n;
  wire fifo_B_PE_14_14__write;
  wire [512:0] fifo_B_PE_14_15__dout;
  wire fifo_B_PE_14_15__empty_n;
  wire fifo_B_PE_14_15__read;
  wire [512:0] fifo_B_PE_14_15__din;
  wire fifo_B_PE_14_15__full_n;
  wire fifo_B_PE_14_15__write;
  wire [512:0] fifo_B_PE_14_16__dout;
  wire fifo_B_PE_14_16__empty_n;
  wire fifo_B_PE_14_16__read;
  wire [512:0] fifo_B_PE_14_16__din;
  wire fifo_B_PE_14_16__full_n;
  wire fifo_B_PE_14_16__write;
  wire [512:0] fifo_B_PE_14_2__dout;
  wire fifo_B_PE_14_2__empty_n;
  wire fifo_B_PE_14_2__read;
  wire [512:0] fifo_B_PE_14_2__din;
  wire fifo_B_PE_14_2__full_n;
  wire fifo_B_PE_14_2__write;
  wire [512:0] fifo_B_PE_14_3__dout;
  wire fifo_B_PE_14_3__empty_n;
  wire fifo_B_PE_14_3__read;
  wire [512:0] fifo_B_PE_14_3__din;
  wire fifo_B_PE_14_3__full_n;
  wire fifo_B_PE_14_3__write;
  wire [512:0] fifo_B_PE_14_4__dout;
  wire fifo_B_PE_14_4__empty_n;
  wire fifo_B_PE_14_4__read;
  wire [512:0] fifo_B_PE_14_4__din;
  wire fifo_B_PE_14_4__full_n;
  wire fifo_B_PE_14_4__write;
  wire [512:0] fifo_B_PE_14_5__dout;
  wire fifo_B_PE_14_5__empty_n;
  wire fifo_B_PE_14_5__read;
  wire [512:0] fifo_B_PE_14_5__din;
  wire fifo_B_PE_14_5__full_n;
  wire fifo_B_PE_14_5__write;
  wire [512:0] fifo_B_PE_14_6__dout;
  wire fifo_B_PE_14_6__empty_n;
  wire fifo_B_PE_14_6__read;
  wire [512:0] fifo_B_PE_14_6__din;
  wire fifo_B_PE_14_6__full_n;
  wire fifo_B_PE_14_6__write;
  wire [512:0] fifo_B_PE_14_7__dout;
  wire fifo_B_PE_14_7__empty_n;
  wire fifo_B_PE_14_7__read;
  wire [512:0] fifo_B_PE_14_7__din;
  wire fifo_B_PE_14_7__full_n;
  wire fifo_B_PE_14_7__write;
  wire [512:0] fifo_B_PE_14_8__dout;
  wire fifo_B_PE_14_8__empty_n;
  wire fifo_B_PE_14_8__read;
  wire [512:0] fifo_B_PE_14_8__din;
  wire fifo_B_PE_14_8__full_n;
  wire fifo_B_PE_14_8__write;
  wire [512:0] fifo_B_PE_14_9__dout;
  wire fifo_B_PE_14_9__empty_n;
  wire fifo_B_PE_14_9__read;
  wire [512:0] fifo_B_PE_14_9__din;
  wire fifo_B_PE_14_9__full_n;
  wire fifo_B_PE_14_9__write;
  wire [512:0] fifo_B_PE_15_0__dout;
  wire fifo_B_PE_15_0__empty_n;
  wire fifo_B_PE_15_0__read;
  wire [512:0] fifo_B_PE_15_0__din;
  wire fifo_B_PE_15_0__full_n;
  wire fifo_B_PE_15_0__write;
  wire [512:0] fifo_B_PE_15_1__dout;
  wire fifo_B_PE_15_1__empty_n;
  wire fifo_B_PE_15_1__read;
  wire [512:0] fifo_B_PE_15_1__din;
  wire fifo_B_PE_15_1__full_n;
  wire fifo_B_PE_15_1__write;
  wire [512:0] fifo_B_PE_15_10__dout;
  wire fifo_B_PE_15_10__empty_n;
  wire fifo_B_PE_15_10__read;
  wire [512:0] fifo_B_PE_15_10__din;
  wire fifo_B_PE_15_10__full_n;
  wire fifo_B_PE_15_10__write;
  wire [512:0] fifo_B_PE_15_11__dout;
  wire fifo_B_PE_15_11__empty_n;
  wire fifo_B_PE_15_11__read;
  wire [512:0] fifo_B_PE_15_11__din;
  wire fifo_B_PE_15_11__full_n;
  wire fifo_B_PE_15_11__write;
  wire [512:0] fifo_B_PE_15_12__dout;
  wire fifo_B_PE_15_12__empty_n;
  wire fifo_B_PE_15_12__read;
  wire [512:0] fifo_B_PE_15_12__din;
  wire fifo_B_PE_15_12__full_n;
  wire fifo_B_PE_15_12__write;
  wire [512:0] fifo_B_PE_15_13__dout;
  wire fifo_B_PE_15_13__empty_n;
  wire fifo_B_PE_15_13__read;
  wire [512:0] fifo_B_PE_15_13__din;
  wire fifo_B_PE_15_13__full_n;
  wire fifo_B_PE_15_13__write;
  wire [512:0] fifo_B_PE_15_14__dout;
  wire fifo_B_PE_15_14__empty_n;
  wire fifo_B_PE_15_14__read;
  wire [512:0] fifo_B_PE_15_14__din;
  wire fifo_B_PE_15_14__full_n;
  wire fifo_B_PE_15_14__write;
  wire [512:0] fifo_B_PE_15_15__dout;
  wire fifo_B_PE_15_15__empty_n;
  wire fifo_B_PE_15_15__read;
  wire [512:0] fifo_B_PE_15_15__din;
  wire fifo_B_PE_15_15__full_n;
  wire fifo_B_PE_15_15__write;
  wire [512:0] fifo_B_PE_15_16__dout;
  wire fifo_B_PE_15_16__empty_n;
  wire fifo_B_PE_15_16__read;
  wire [512:0] fifo_B_PE_15_16__din;
  wire fifo_B_PE_15_16__full_n;
  wire fifo_B_PE_15_16__write;
  wire [512:0] fifo_B_PE_15_2__dout;
  wire fifo_B_PE_15_2__empty_n;
  wire fifo_B_PE_15_2__read;
  wire [512:0] fifo_B_PE_15_2__din;
  wire fifo_B_PE_15_2__full_n;
  wire fifo_B_PE_15_2__write;
  wire [512:0] fifo_B_PE_15_3__dout;
  wire fifo_B_PE_15_3__empty_n;
  wire fifo_B_PE_15_3__read;
  wire [512:0] fifo_B_PE_15_3__din;
  wire fifo_B_PE_15_3__full_n;
  wire fifo_B_PE_15_3__write;
  wire [512:0] fifo_B_PE_15_4__dout;
  wire fifo_B_PE_15_4__empty_n;
  wire fifo_B_PE_15_4__read;
  wire [512:0] fifo_B_PE_15_4__din;
  wire fifo_B_PE_15_4__full_n;
  wire fifo_B_PE_15_4__write;
  wire [512:0] fifo_B_PE_15_5__dout;
  wire fifo_B_PE_15_5__empty_n;
  wire fifo_B_PE_15_5__read;
  wire [512:0] fifo_B_PE_15_5__din;
  wire fifo_B_PE_15_5__full_n;
  wire fifo_B_PE_15_5__write;
  wire [512:0] fifo_B_PE_15_6__dout;
  wire fifo_B_PE_15_6__empty_n;
  wire fifo_B_PE_15_6__read;
  wire [512:0] fifo_B_PE_15_6__din;
  wire fifo_B_PE_15_6__full_n;
  wire fifo_B_PE_15_6__write;
  wire [512:0] fifo_B_PE_15_7__dout;
  wire fifo_B_PE_15_7__empty_n;
  wire fifo_B_PE_15_7__read;
  wire [512:0] fifo_B_PE_15_7__din;
  wire fifo_B_PE_15_7__full_n;
  wire fifo_B_PE_15_7__write;
  wire [512:0] fifo_B_PE_15_8__dout;
  wire fifo_B_PE_15_8__empty_n;
  wire fifo_B_PE_15_8__read;
  wire [512:0] fifo_B_PE_15_8__din;
  wire fifo_B_PE_15_8__full_n;
  wire fifo_B_PE_15_8__write;
  wire [512:0] fifo_B_PE_15_9__dout;
  wire fifo_B_PE_15_9__empty_n;
  wire fifo_B_PE_15_9__read;
  wire [512:0] fifo_B_PE_15_9__din;
  wire fifo_B_PE_15_9__full_n;
  wire fifo_B_PE_15_9__write;
  wire [512:0] fifo_B_PE_16_0__dout;
  wire fifo_B_PE_16_0__empty_n;
  wire fifo_B_PE_16_0__read;
  wire [512:0] fifo_B_PE_16_0__din;
  wire fifo_B_PE_16_0__full_n;
  wire fifo_B_PE_16_0__write;
  wire [512:0] fifo_B_PE_16_1__dout;
  wire fifo_B_PE_16_1__empty_n;
  wire fifo_B_PE_16_1__read;
  wire [512:0] fifo_B_PE_16_1__din;
  wire fifo_B_PE_16_1__full_n;
  wire fifo_B_PE_16_1__write;
  wire [512:0] fifo_B_PE_16_10__dout;
  wire fifo_B_PE_16_10__empty_n;
  wire fifo_B_PE_16_10__read;
  wire [512:0] fifo_B_PE_16_10__din;
  wire fifo_B_PE_16_10__full_n;
  wire fifo_B_PE_16_10__write;
  wire [512:0] fifo_B_PE_16_11__dout;
  wire fifo_B_PE_16_11__empty_n;
  wire fifo_B_PE_16_11__read;
  wire [512:0] fifo_B_PE_16_11__din;
  wire fifo_B_PE_16_11__full_n;
  wire fifo_B_PE_16_11__write;
  wire [512:0] fifo_B_PE_16_12__dout;
  wire fifo_B_PE_16_12__empty_n;
  wire fifo_B_PE_16_12__read;
  wire [512:0] fifo_B_PE_16_12__din;
  wire fifo_B_PE_16_12__full_n;
  wire fifo_B_PE_16_12__write;
  wire [512:0] fifo_B_PE_16_13__dout;
  wire fifo_B_PE_16_13__empty_n;
  wire fifo_B_PE_16_13__read;
  wire [512:0] fifo_B_PE_16_13__din;
  wire fifo_B_PE_16_13__full_n;
  wire fifo_B_PE_16_13__write;
  wire [512:0] fifo_B_PE_16_14__dout;
  wire fifo_B_PE_16_14__empty_n;
  wire fifo_B_PE_16_14__read;
  wire [512:0] fifo_B_PE_16_14__din;
  wire fifo_B_PE_16_14__full_n;
  wire fifo_B_PE_16_14__write;
  wire [512:0] fifo_B_PE_16_15__dout;
  wire fifo_B_PE_16_15__empty_n;
  wire fifo_B_PE_16_15__read;
  wire [512:0] fifo_B_PE_16_15__din;
  wire fifo_B_PE_16_15__full_n;
  wire fifo_B_PE_16_15__write;
  wire [512:0] fifo_B_PE_16_16__dout;
  wire fifo_B_PE_16_16__empty_n;
  wire fifo_B_PE_16_16__read;
  wire [512:0] fifo_B_PE_16_16__din;
  wire fifo_B_PE_16_16__full_n;
  wire fifo_B_PE_16_16__write;
  wire [512:0] fifo_B_PE_16_2__dout;
  wire fifo_B_PE_16_2__empty_n;
  wire fifo_B_PE_16_2__read;
  wire [512:0] fifo_B_PE_16_2__din;
  wire fifo_B_PE_16_2__full_n;
  wire fifo_B_PE_16_2__write;
  wire [512:0] fifo_B_PE_16_3__dout;
  wire fifo_B_PE_16_3__empty_n;
  wire fifo_B_PE_16_3__read;
  wire [512:0] fifo_B_PE_16_3__din;
  wire fifo_B_PE_16_3__full_n;
  wire fifo_B_PE_16_3__write;
  wire [512:0] fifo_B_PE_16_4__dout;
  wire fifo_B_PE_16_4__empty_n;
  wire fifo_B_PE_16_4__read;
  wire [512:0] fifo_B_PE_16_4__din;
  wire fifo_B_PE_16_4__full_n;
  wire fifo_B_PE_16_4__write;
  wire [512:0] fifo_B_PE_16_5__dout;
  wire fifo_B_PE_16_5__empty_n;
  wire fifo_B_PE_16_5__read;
  wire [512:0] fifo_B_PE_16_5__din;
  wire fifo_B_PE_16_5__full_n;
  wire fifo_B_PE_16_5__write;
  wire [512:0] fifo_B_PE_16_6__dout;
  wire fifo_B_PE_16_6__empty_n;
  wire fifo_B_PE_16_6__read;
  wire [512:0] fifo_B_PE_16_6__din;
  wire fifo_B_PE_16_6__full_n;
  wire fifo_B_PE_16_6__write;
  wire [512:0] fifo_B_PE_16_7__dout;
  wire fifo_B_PE_16_7__empty_n;
  wire fifo_B_PE_16_7__read;
  wire [512:0] fifo_B_PE_16_7__din;
  wire fifo_B_PE_16_7__full_n;
  wire fifo_B_PE_16_7__write;
  wire [512:0] fifo_B_PE_16_8__dout;
  wire fifo_B_PE_16_8__empty_n;
  wire fifo_B_PE_16_8__read;
  wire [512:0] fifo_B_PE_16_8__din;
  wire fifo_B_PE_16_8__full_n;
  wire fifo_B_PE_16_8__write;
  wire [512:0] fifo_B_PE_16_9__dout;
  wire fifo_B_PE_16_9__empty_n;
  wire fifo_B_PE_16_9__read;
  wire [512:0] fifo_B_PE_16_9__din;
  wire fifo_B_PE_16_9__full_n;
  wire fifo_B_PE_16_9__write;
  wire [512:0] fifo_B_PE_17_0__dout;
  wire fifo_B_PE_17_0__empty_n;
  wire fifo_B_PE_17_0__read;
  wire [512:0] fifo_B_PE_17_0__din;
  wire fifo_B_PE_17_0__full_n;
  wire fifo_B_PE_17_0__write;
  wire [512:0] fifo_B_PE_17_1__dout;
  wire fifo_B_PE_17_1__empty_n;
  wire fifo_B_PE_17_1__read;
  wire [512:0] fifo_B_PE_17_1__din;
  wire fifo_B_PE_17_1__full_n;
  wire fifo_B_PE_17_1__write;
  wire [512:0] fifo_B_PE_17_10__dout;
  wire fifo_B_PE_17_10__empty_n;
  wire fifo_B_PE_17_10__read;
  wire [512:0] fifo_B_PE_17_10__din;
  wire fifo_B_PE_17_10__full_n;
  wire fifo_B_PE_17_10__write;
  wire [512:0] fifo_B_PE_17_11__dout;
  wire fifo_B_PE_17_11__empty_n;
  wire fifo_B_PE_17_11__read;
  wire [512:0] fifo_B_PE_17_11__din;
  wire fifo_B_PE_17_11__full_n;
  wire fifo_B_PE_17_11__write;
  wire [512:0] fifo_B_PE_17_12__dout;
  wire fifo_B_PE_17_12__empty_n;
  wire fifo_B_PE_17_12__read;
  wire [512:0] fifo_B_PE_17_12__din;
  wire fifo_B_PE_17_12__full_n;
  wire fifo_B_PE_17_12__write;
  wire [512:0] fifo_B_PE_17_13__dout;
  wire fifo_B_PE_17_13__empty_n;
  wire fifo_B_PE_17_13__read;
  wire [512:0] fifo_B_PE_17_13__din;
  wire fifo_B_PE_17_13__full_n;
  wire fifo_B_PE_17_13__write;
  wire [512:0] fifo_B_PE_17_14__dout;
  wire fifo_B_PE_17_14__empty_n;
  wire fifo_B_PE_17_14__read;
  wire [512:0] fifo_B_PE_17_14__din;
  wire fifo_B_PE_17_14__full_n;
  wire fifo_B_PE_17_14__write;
  wire [512:0] fifo_B_PE_17_15__dout;
  wire fifo_B_PE_17_15__empty_n;
  wire fifo_B_PE_17_15__read;
  wire [512:0] fifo_B_PE_17_15__din;
  wire fifo_B_PE_17_15__full_n;
  wire fifo_B_PE_17_15__write;
  wire [512:0] fifo_B_PE_17_16__dout;
  wire fifo_B_PE_17_16__empty_n;
  wire fifo_B_PE_17_16__read;
  wire [512:0] fifo_B_PE_17_16__din;
  wire fifo_B_PE_17_16__full_n;
  wire fifo_B_PE_17_16__write;
  wire [512:0] fifo_B_PE_17_2__dout;
  wire fifo_B_PE_17_2__empty_n;
  wire fifo_B_PE_17_2__read;
  wire [512:0] fifo_B_PE_17_2__din;
  wire fifo_B_PE_17_2__full_n;
  wire fifo_B_PE_17_2__write;
  wire [512:0] fifo_B_PE_17_3__dout;
  wire fifo_B_PE_17_3__empty_n;
  wire fifo_B_PE_17_3__read;
  wire [512:0] fifo_B_PE_17_3__din;
  wire fifo_B_PE_17_3__full_n;
  wire fifo_B_PE_17_3__write;
  wire [512:0] fifo_B_PE_17_4__dout;
  wire fifo_B_PE_17_4__empty_n;
  wire fifo_B_PE_17_4__read;
  wire [512:0] fifo_B_PE_17_4__din;
  wire fifo_B_PE_17_4__full_n;
  wire fifo_B_PE_17_4__write;
  wire [512:0] fifo_B_PE_17_5__dout;
  wire fifo_B_PE_17_5__empty_n;
  wire fifo_B_PE_17_5__read;
  wire [512:0] fifo_B_PE_17_5__din;
  wire fifo_B_PE_17_5__full_n;
  wire fifo_B_PE_17_5__write;
  wire [512:0] fifo_B_PE_17_6__dout;
  wire fifo_B_PE_17_6__empty_n;
  wire fifo_B_PE_17_6__read;
  wire [512:0] fifo_B_PE_17_6__din;
  wire fifo_B_PE_17_6__full_n;
  wire fifo_B_PE_17_6__write;
  wire [512:0] fifo_B_PE_17_7__dout;
  wire fifo_B_PE_17_7__empty_n;
  wire fifo_B_PE_17_7__read;
  wire [512:0] fifo_B_PE_17_7__din;
  wire fifo_B_PE_17_7__full_n;
  wire fifo_B_PE_17_7__write;
  wire [512:0] fifo_B_PE_17_8__dout;
  wire fifo_B_PE_17_8__empty_n;
  wire fifo_B_PE_17_8__read;
  wire [512:0] fifo_B_PE_17_8__din;
  wire fifo_B_PE_17_8__full_n;
  wire fifo_B_PE_17_8__write;
  wire [512:0] fifo_B_PE_17_9__dout;
  wire fifo_B_PE_17_9__empty_n;
  wire fifo_B_PE_17_9__read;
  wire [512:0] fifo_B_PE_17_9__din;
  wire fifo_B_PE_17_9__full_n;
  wire fifo_B_PE_17_9__write;
  wire [512:0] fifo_B_PE_18_0__dout;
  wire fifo_B_PE_18_0__empty_n;
  wire fifo_B_PE_18_0__read;
  wire [512:0] fifo_B_PE_18_0__din;
  wire fifo_B_PE_18_0__full_n;
  wire fifo_B_PE_18_0__write;
  wire [512:0] fifo_B_PE_18_1__dout;
  wire fifo_B_PE_18_1__empty_n;
  wire fifo_B_PE_18_1__read;
  wire [512:0] fifo_B_PE_18_1__din;
  wire fifo_B_PE_18_1__full_n;
  wire fifo_B_PE_18_1__write;
  wire [512:0] fifo_B_PE_18_10__dout;
  wire fifo_B_PE_18_10__empty_n;
  wire fifo_B_PE_18_10__read;
  wire [512:0] fifo_B_PE_18_10__din;
  wire fifo_B_PE_18_10__full_n;
  wire fifo_B_PE_18_10__write;
  wire [512:0] fifo_B_PE_18_11__dout;
  wire fifo_B_PE_18_11__empty_n;
  wire fifo_B_PE_18_11__read;
  wire [512:0] fifo_B_PE_18_11__din;
  wire fifo_B_PE_18_11__full_n;
  wire fifo_B_PE_18_11__write;
  wire [512:0] fifo_B_PE_18_12__dout;
  wire fifo_B_PE_18_12__empty_n;
  wire fifo_B_PE_18_12__read;
  wire [512:0] fifo_B_PE_18_12__din;
  wire fifo_B_PE_18_12__full_n;
  wire fifo_B_PE_18_12__write;
  wire [512:0] fifo_B_PE_18_13__dout;
  wire fifo_B_PE_18_13__empty_n;
  wire fifo_B_PE_18_13__read;
  wire [512:0] fifo_B_PE_18_13__din;
  wire fifo_B_PE_18_13__full_n;
  wire fifo_B_PE_18_13__write;
  wire [512:0] fifo_B_PE_18_14__dout;
  wire fifo_B_PE_18_14__empty_n;
  wire fifo_B_PE_18_14__read;
  wire [512:0] fifo_B_PE_18_14__din;
  wire fifo_B_PE_18_14__full_n;
  wire fifo_B_PE_18_14__write;
  wire [512:0] fifo_B_PE_18_15__dout;
  wire fifo_B_PE_18_15__empty_n;
  wire fifo_B_PE_18_15__read;
  wire [512:0] fifo_B_PE_18_15__din;
  wire fifo_B_PE_18_15__full_n;
  wire fifo_B_PE_18_15__write;
  wire [512:0] fifo_B_PE_18_16__dout;
  wire fifo_B_PE_18_16__empty_n;
  wire fifo_B_PE_18_16__read;
  wire [512:0] fifo_B_PE_18_16__din;
  wire fifo_B_PE_18_16__full_n;
  wire fifo_B_PE_18_16__write;
  wire [512:0] fifo_B_PE_18_2__dout;
  wire fifo_B_PE_18_2__empty_n;
  wire fifo_B_PE_18_2__read;
  wire [512:0] fifo_B_PE_18_2__din;
  wire fifo_B_PE_18_2__full_n;
  wire fifo_B_PE_18_2__write;
  wire [512:0] fifo_B_PE_18_3__dout;
  wire fifo_B_PE_18_3__empty_n;
  wire fifo_B_PE_18_3__read;
  wire [512:0] fifo_B_PE_18_3__din;
  wire fifo_B_PE_18_3__full_n;
  wire fifo_B_PE_18_3__write;
  wire [512:0] fifo_B_PE_18_4__dout;
  wire fifo_B_PE_18_4__empty_n;
  wire fifo_B_PE_18_4__read;
  wire [512:0] fifo_B_PE_18_4__din;
  wire fifo_B_PE_18_4__full_n;
  wire fifo_B_PE_18_4__write;
  wire [512:0] fifo_B_PE_18_5__dout;
  wire fifo_B_PE_18_5__empty_n;
  wire fifo_B_PE_18_5__read;
  wire [512:0] fifo_B_PE_18_5__din;
  wire fifo_B_PE_18_5__full_n;
  wire fifo_B_PE_18_5__write;
  wire [512:0] fifo_B_PE_18_6__dout;
  wire fifo_B_PE_18_6__empty_n;
  wire fifo_B_PE_18_6__read;
  wire [512:0] fifo_B_PE_18_6__din;
  wire fifo_B_PE_18_6__full_n;
  wire fifo_B_PE_18_6__write;
  wire [512:0] fifo_B_PE_18_7__dout;
  wire fifo_B_PE_18_7__empty_n;
  wire fifo_B_PE_18_7__read;
  wire [512:0] fifo_B_PE_18_7__din;
  wire fifo_B_PE_18_7__full_n;
  wire fifo_B_PE_18_7__write;
  wire [512:0] fifo_B_PE_18_8__dout;
  wire fifo_B_PE_18_8__empty_n;
  wire fifo_B_PE_18_8__read;
  wire [512:0] fifo_B_PE_18_8__din;
  wire fifo_B_PE_18_8__full_n;
  wire fifo_B_PE_18_8__write;
  wire [512:0] fifo_B_PE_18_9__dout;
  wire fifo_B_PE_18_9__empty_n;
  wire fifo_B_PE_18_9__read;
  wire [512:0] fifo_B_PE_18_9__din;
  wire fifo_B_PE_18_9__full_n;
  wire fifo_B_PE_18_9__write;
  wire [512:0] fifo_B_PE_1_0__dout;
  wire fifo_B_PE_1_0__empty_n;
  wire fifo_B_PE_1_0__read;
  wire [512:0] fifo_B_PE_1_0__din;
  wire fifo_B_PE_1_0__full_n;
  wire fifo_B_PE_1_0__write;
  wire [512:0] fifo_B_PE_1_1__dout;
  wire fifo_B_PE_1_1__empty_n;
  wire fifo_B_PE_1_1__read;
  wire [512:0] fifo_B_PE_1_1__din;
  wire fifo_B_PE_1_1__full_n;
  wire fifo_B_PE_1_1__write;
  wire [512:0] fifo_B_PE_1_10__dout;
  wire fifo_B_PE_1_10__empty_n;
  wire fifo_B_PE_1_10__read;
  wire [512:0] fifo_B_PE_1_10__din;
  wire fifo_B_PE_1_10__full_n;
  wire fifo_B_PE_1_10__write;
  wire [512:0] fifo_B_PE_1_11__dout;
  wire fifo_B_PE_1_11__empty_n;
  wire fifo_B_PE_1_11__read;
  wire [512:0] fifo_B_PE_1_11__din;
  wire fifo_B_PE_1_11__full_n;
  wire fifo_B_PE_1_11__write;
  wire [512:0] fifo_B_PE_1_12__dout;
  wire fifo_B_PE_1_12__empty_n;
  wire fifo_B_PE_1_12__read;
  wire [512:0] fifo_B_PE_1_12__din;
  wire fifo_B_PE_1_12__full_n;
  wire fifo_B_PE_1_12__write;
  wire [512:0] fifo_B_PE_1_13__dout;
  wire fifo_B_PE_1_13__empty_n;
  wire fifo_B_PE_1_13__read;
  wire [512:0] fifo_B_PE_1_13__din;
  wire fifo_B_PE_1_13__full_n;
  wire fifo_B_PE_1_13__write;
  wire [512:0] fifo_B_PE_1_14__dout;
  wire fifo_B_PE_1_14__empty_n;
  wire fifo_B_PE_1_14__read;
  wire [512:0] fifo_B_PE_1_14__din;
  wire fifo_B_PE_1_14__full_n;
  wire fifo_B_PE_1_14__write;
  wire [512:0] fifo_B_PE_1_15__dout;
  wire fifo_B_PE_1_15__empty_n;
  wire fifo_B_PE_1_15__read;
  wire [512:0] fifo_B_PE_1_15__din;
  wire fifo_B_PE_1_15__full_n;
  wire fifo_B_PE_1_15__write;
  wire [512:0] fifo_B_PE_1_16__dout;
  wire fifo_B_PE_1_16__empty_n;
  wire fifo_B_PE_1_16__read;
  wire [512:0] fifo_B_PE_1_16__din;
  wire fifo_B_PE_1_16__full_n;
  wire fifo_B_PE_1_16__write;
  wire [512:0] fifo_B_PE_1_2__dout;
  wire fifo_B_PE_1_2__empty_n;
  wire fifo_B_PE_1_2__read;
  wire [512:0] fifo_B_PE_1_2__din;
  wire fifo_B_PE_1_2__full_n;
  wire fifo_B_PE_1_2__write;
  wire [512:0] fifo_B_PE_1_3__dout;
  wire fifo_B_PE_1_3__empty_n;
  wire fifo_B_PE_1_3__read;
  wire [512:0] fifo_B_PE_1_3__din;
  wire fifo_B_PE_1_3__full_n;
  wire fifo_B_PE_1_3__write;
  wire [512:0] fifo_B_PE_1_4__dout;
  wire fifo_B_PE_1_4__empty_n;
  wire fifo_B_PE_1_4__read;
  wire [512:0] fifo_B_PE_1_4__din;
  wire fifo_B_PE_1_4__full_n;
  wire fifo_B_PE_1_4__write;
  wire [512:0] fifo_B_PE_1_5__dout;
  wire fifo_B_PE_1_5__empty_n;
  wire fifo_B_PE_1_5__read;
  wire [512:0] fifo_B_PE_1_5__din;
  wire fifo_B_PE_1_5__full_n;
  wire fifo_B_PE_1_5__write;
  wire [512:0] fifo_B_PE_1_6__dout;
  wire fifo_B_PE_1_6__empty_n;
  wire fifo_B_PE_1_6__read;
  wire [512:0] fifo_B_PE_1_6__din;
  wire fifo_B_PE_1_6__full_n;
  wire fifo_B_PE_1_6__write;
  wire [512:0] fifo_B_PE_1_7__dout;
  wire fifo_B_PE_1_7__empty_n;
  wire fifo_B_PE_1_7__read;
  wire [512:0] fifo_B_PE_1_7__din;
  wire fifo_B_PE_1_7__full_n;
  wire fifo_B_PE_1_7__write;
  wire [512:0] fifo_B_PE_1_8__dout;
  wire fifo_B_PE_1_8__empty_n;
  wire fifo_B_PE_1_8__read;
  wire [512:0] fifo_B_PE_1_8__din;
  wire fifo_B_PE_1_8__full_n;
  wire fifo_B_PE_1_8__write;
  wire [512:0] fifo_B_PE_1_9__dout;
  wire fifo_B_PE_1_9__empty_n;
  wire fifo_B_PE_1_9__read;
  wire [512:0] fifo_B_PE_1_9__din;
  wire fifo_B_PE_1_9__full_n;
  wire fifo_B_PE_1_9__write;
  wire [512:0] fifo_B_PE_2_0__dout;
  wire fifo_B_PE_2_0__empty_n;
  wire fifo_B_PE_2_0__read;
  wire [512:0] fifo_B_PE_2_0__din;
  wire fifo_B_PE_2_0__full_n;
  wire fifo_B_PE_2_0__write;
  wire [512:0] fifo_B_PE_2_1__dout;
  wire fifo_B_PE_2_1__empty_n;
  wire fifo_B_PE_2_1__read;
  wire [512:0] fifo_B_PE_2_1__din;
  wire fifo_B_PE_2_1__full_n;
  wire fifo_B_PE_2_1__write;
  wire [512:0] fifo_B_PE_2_10__dout;
  wire fifo_B_PE_2_10__empty_n;
  wire fifo_B_PE_2_10__read;
  wire [512:0] fifo_B_PE_2_10__din;
  wire fifo_B_PE_2_10__full_n;
  wire fifo_B_PE_2_10__write;
  wire [512:0] fifo_B_PE_2_11__dout;
  wire fifo_B_PE_2_11__empty_n;
  wire fifo_B_PE_2_11__read;
  wire [512:0] fifo_B_PE_2_11__din;
  wire fifo_B_PE_2_11__full_n;
  wire fifo_B_PE_2_11__write;
  wire [512:0] fifo_B_PE_2_12__dout;
  wire fifo_B_PE_2_12__empty_n;
  wire fifo_B_PE_2_12__read;
  wire [512:0] fifo_B_PE_2_12__din;
  wire fifo_B_PE_2_12__full_n;
  wire fifo_B_PE_2_12__write;
  wire [512:0] fifo_B_PE_2_13__dout;
  wire fifo_B_PE_2_13__empty_n;
  wire fifo_B_PE_2_13__read;
  wire [512:0] fifo_B_PE_2_13__din;
  wire fifo_B_PE_2_13__full_n;
  wire fifo_B_PE_2_13__write;
  wire [512:0] fifo_B_PE_2_14__dout;
  wire fifo_B_PE_2_14__empty_n;
  wire fifo_B_PE_2_14__read;
  wire [512:0] fifo_B_PE_2_14__din;
  wire fifo_B_PE_2_14__full_n;
  wire fifo_B_PE_2_14__write;
  wire [512:0] fifo_B_PE_2_15__dout;
  wire fifo_B_PE_2_15__empty_n;
  wire fifo_B_PE_2_15__read;
  wire [512:0] fifo_B_PE_2_15__din;
  wire fifo_B_PE_2_15__full_n;
  wire fifo_B_PE_2_15__write;
  wire [512:0] fifo_B_PE_2_16__dout;
  wire fifo_B_PE_2_16__empty_n;
  wire fifo_B_PE_2_16__read;
  wire [512:0] fifo_B_PE_2_16__din;
  wire fifo_B_PE_2_16__full_n;
  wire fifo_B_PE_2_16__write;
  wire [512:0] fifo_B_PE_2_2__dout;
  wire fifo_B_PE_2_2__empty_n;
  wire fifo_B_PE_2_2__read;
  wire [512:0] fifo_B_PE_2_2__din;
  wire fifo_B_PE_2_2__full_n;
  wire fifo_B_PE_2_2__write;
  wire [512:0] fifo_B_PE_2_3__dout;
  wire fifo_B_PE_2_3__empty_n;
  wire fifo_B_PE_2_3__read;
  wire [512:0] fifo_B_PE_2_3__din;
  wire fifo_B_PE_2_3__full_n;
  wire fifo_B_PE_2_3__write;
  wire [512:0] fifo_B_PE_2_4__dout;
  wire fifo_B_PE_2_4__empty_n;
  wire fifo_B_PE_2_4__read;
  wire [512:0] fifo_B_PE_2_4__din;
  wire fifo_B_PE_2_4__full_n;
  wire fifo_B_PE_2_4__write;
  wire [512:0] fifo_B_PE_2_5__dout;
  wire fifo_B_PE_2_5__empty_n;
  wire fifo_B_PE_2_5__read;
  wire [512:0] fifo_B_PE_2_5__din;
  wire fifo_B_PE_2_5__full_n;
  wire fifo_B_PE_2_5__write;
  wire [512:0] fifo_B_PE_2_6__dout;
  wire fifo_B_PE_2_6__empty_n;
  wire fifo_B_PE_2_6__read;
  wire [512:0] fifo_B_PE_2_6__din;
  wire fifo_B_PE_2_6__full_n;
  wire fifo_B_PE_2_6__write;
  wire [512:0] fifo_B_PE_2_7__dout;
  wire fifo_B_PE_2_7__empty_n;
  wire fifo_B_PE_2_7__read;
  wire [512:0] fifo_B_PE_2_7__din;
  wire fifo_B_PE_2_7__full_n;
  wire fifo_B_PE_2_7__write;
  wire [512:0] fifo_B_PE_2_8__dout;
  wire fifo_B_PE_2_8__empty_n;
  wire fifo_B_PE_2_8__read;
  wire [512:0] fifo_B_PE_2_8__din;
  wire fifo_B_PE_2_8__full_n;
  wire fifo_B_PE_2_8__write;
  wire [512:0] fifo_B_PE_2_9__dout;
  wire fifo_B_PE_2_9__empty_n;
  wire fifo_B_PE_2_9__read;
  wire [512:0] fifo_B_PE_2_9__din;
  wire fifo_B_PE_2_9__full_n;
  wire fifo_B_PE_2_9__write;
  wire [512:0] fifo_B_PE_3_0__dout;
  wire fifo_B_PE_3_0__empty_n;
  wire fifo_B_PE_3_0__read;
  wire [512:0] fifo_B_PE_3_0__din;
  wire fifo_B_PE_3_0__full_n;
  wire fifo_B_PE_3_0__write;
  wire [512:0] fifo_B_PE_3_1__dout;
  wire fifo_B_PE_3_1__empty_n;
  wire fifo_B_PE_3_1__read;
  wire [512:0] fifo_B_PE_3_1__din;
  wire fifo_B_PE_3_1__full_n;
  wire fifo_B_PE_3_1__write;
  wire [512:0] fifo_B_PE_3_10__dout;
  wire fifo_B_PE_3_10__empty_n;
  wire fifo_B_PE_3_10__read;
  wire [512:0] fifo_B_PE_3_10__din;
  wire fifo_B_PE_3_10__full_n;
  wire fifo_B_PE_3_10__write;
  wire [512:0] fifo_B_PE_3_11__dout;
  wire fifo_B_PE_3_11__empty_n;
  wire fifo_B_PE_3_11__read;
  wire [512:0] fifo_B_PE_3_11__din;
  wire fifo_B_PE_3_11__full_n;
  wire fifo_B_PE_3_11__write;
  wire [512:0] fifo_B_PE_3_12__dout;
  wire fifo_B_PE_3_12__empty_n;
  wire fifo_B_PE_3_12__read;
  wire [512:0] fifo_B_PE_3_12__din;
  wire fifo_B_PE_3_12__full_n;
  wire fifo_B_PE_3_12__write;
  wire [512:0] fifo_B_PE_3_13__dout;
  wire fifo_B_PE_3_13__empty_n;
  wire fifo_B_PE_3_13__read;
  wire [512:0] fifo_B_PE_3_13__din;
  wire fifo_B_PE_3_13__full_n;
  wire fifo_B_PE_3_13__write;
  wire [512:0] fifo_B_PE_3_14__dout;
  wire fifo_B_PE_3_14__empty_n;
  wire fifo_B_PE_3_14__read;
  wire [512:0] fifo_B_PE_3_14__din;
  wire fifo_B_PE_3_14__full_n;
  wire fifo_B_PE_3_14__write;
  wire [512:0] fifo_B_PE_3_15__dout;
  wire fifo_B_PE_3_15__empty_n;
  wire fifo_B_PE_3_15__read;
  wire [512:0] fifo_B_PE_3_15__din;
  wire fifo_B_PE_3_15__full_n;
  wire fifo_B_PE_3_15__write;
  wire [512:0] fifo_B_PE_3_16__dout;
  wire fifo_B_PE_3_16__empty_n;
  wire fifo_B_PE_3_16__read;
  wire [512:0] fifo_B_PE_3_16__din;
  wire fifo_B_PE_3_16__full_n;
  wire fifo_B_PE_3_16__write;
  wire [512:0] fifo_B_PE_3_2__dout;
  wire fifo_B_PE_3_2__empty_n;
  wire fifo_B_PE_3_2__read;
  wire [512:0] fifo_B_PE_3_2__din;
  wire fifo_B_PE_3_2__full_n;
  wire fifo_B_PE_3_2__write;
  wire [512:0] fifo_B_PE_3_3__dout;
  wire fifo_B_PE_3_3__empty_n;
  wire fifo_B_PE_3_3__read;
  wire [512:0] fifo_B_PE_3_3__din;
  wire fifo_B_PE_3_3__full_n;
  wire fifo_B_PE_3_3__write;
  wire [512:0] fifo_B_PE_3_4__dout;
  wire fifo_B_PE_3_4__empty_n;
  wire fifo_B_PE_3_4__read;
  wire [512:0] fifo_B_PE_3_4__din;
  wire fifo_B_PE_3_4__full_n;
  wire fifo_B_PE_3_4__write;
  wire [512:0] fifo_B_PE_3_5__dout;
  wire fifo_B_PE_3_5__empty_n;
  wire fifo_B_PE_3_5__read;
  wire [512:0] fifo_B_PE_3_5__din;
  wire fifo_B_PE_3_5__full_n;
  wire fifo_B_PE_3_5__write;
  wire [512:0] fifo_B_PE_3_6__dout;
  wire fifo_B_PE_3_6__empty_n;
  wire fifo_B_PE_3_6__read;
  wire [512:0] fifo_B_PE_3_6__din;
  wire fifo_B_PE_3_6__full_n;
  wire fifo_B_PE_3_6__write;
  wire [512:0] fifo_B_PE_3_7__dout;
  wire fifo_B_PE_3_7__empty_n;
  wire fifo_B_PE_3_7__read;
  wire [512:0] fifo_B_PE_3_7__din;
  wire fifo_B_PE_3_7__full_n;
  wire fifo_B_PE_3_7__write;
  wire [512:0] fifo_B_PE_3_8__dout;
  wire fifo_B_PE_3_8__empty_n;
  wire fifo_B_PE_3_8__read;
  wire [512:0] fifo_B_PE_3_8__din;
  wire fifo_B_PE_3_8__full_n;
  wire fifo_B_PE_3_8__write;
  wire [512:0] fifo_B_PE_3_9__dout;
  wire fifo_B_PE_3_9__empty_n;
  wire fifo_B_PE_3_9__read;
  wire [512:0] fifo_B_PE_3_9__din;
  wire fifo_B_PE_3_9__full_n;
  wire fifo_B_PE_3_9__write;
  wire [512:0] fifo_B_PE_4_0__dout;
  wire fifo_B_PE_4_0__empty_n;
  wire fifo_B_PE_4_0__read;
  wire [512:0] fifo_B_PE_4_0__din;
  wire fifo_B_PE_4_0__full_n;
  wire fifo_B_PE_4_0__write;
  wire [512:0] fifo_B_PE_4_1__dout;
  wire fifo_B_PE_4_1__empty_n;
  wire fifo_B_PE_4_1__read;
  wire [512:0] fifo_B_PE_4_1__din;
  wire fifo_B_PE_4_1__full_n;
  wire fifo_B_PE_4_1__write;
  wire [512:0] fifo_B_PE_4_10__dout;
  wire fifo_B_PE_4_10__empty_n;
  wire fifo_B_PE_4_10__read;
  wire [512:0] fifo_B_PE_4_10__din;
  wire fifo_B_PE_4_10__full_n;
  wire fifo_B_PE_4_10__write;
  wire [512:0] fifo_B_PE_4_11__dout;
  wire fifo_B_PE_4_11__empty_n;
  wire fifo_B_PE_4_11__read;
  wire [512:0] fifo_B_PE_4_11__din;
  wire fifo_B_PE_4_11__full_n;
  wire fifo_B_PE_4_11__write;
  wire [512:0] fifo_B_PE_4_12__dout;
  wire fifo_B_PE_4_12__empty_n;
  wire fifo_B_PE_4_12__read;
  wire [512:0] fifo_B_PE_4_12__din;
  wire fifo_B_PE_4_12__full_n;
  wire fifo_B_PE_4_12__write;
  wire [512:0] fifo_B_PE_4_13__dout;
  wire fifo_B_PE_4_13__empty_n;
  wire fifo_B_PE_4_13__read;
  wire [512:0] fifo_B_PE_4_13__din;
  wire fifo_B_PE_4_13__full_n;
  wire fifo_B_PE_4_13__write;
  wire [512:0] fifo_B_PE_4_14__dout;
  wire fifo_B_PE_4_14__empty_n;
  wire fifo_B_PE_4_14__read;
  wire [512:0] fifo_B_PE_4_14__din;
  wire fifo_B_PE_4_14__full_n;
  wire fifo_B_PE_4_14__write;
  wire [512:0] fifo_B_PE_4_15__dout;
  wire fifo_B_PE_4_15__empty_n;
  wire fifo_B_PE_4_15__read;
  wire [512:0] fifo_B_PE_4_15__din;
  wire fifo_B_PE_4_15__full_n;
  wire fifo_B_PE_4_15__write;
  wire [512:0] fifo_B_PE_4_16__dout;
  wire fifo_B_PE_4_16__empty_n;
  wire fifo_B_PE_4_16__read;
  wire [512:0] fifo_B_PE_4_16__din;
  wire fifo_B_PE_4_16__full_n;
  wire fifo_B_PE_4_16__write;
  wire [512:0] fifo_B_PE_4_2__dout;
  wire fifo_B_PE_4_2__empty_n;
  wire fifo_B_PE_4_2__read;
  wire [512:0] fifo_B_PE_4_2__din;
  wire fifo_B_PE_4_2__full_n;
  wire fifo_B_PE_4_2__write;
  wire [512:0] fifo_B_PE_4_3__dout;
  wire fifo_B_PE_4_3__empty_n;
  wire fifo_B_PE_4_3__read;
  wire [512:0] fifo_B_PE_4_3__din;
  wire fifo_B_PE_4_3__full_n;
  wire fifo_B_PE_4_3__write;
  wire [512:0] fifo_B_PE_4_4__dout;
  wire fifo_B_PE_4_4__empty_n;
  wire fifo_B_PE_4_4__read;
  wire [512:0] fifo_B_PE_4_4__din;
  wire fifo_B_PE_4_4__full_n;
  wire fifo_B_PE_4_4__write;
  wire [512:0] fifo_B_PE_4_5__dout;
  wire fifo_B_PE_4_5__empty_n;
  wire fifo_B_PE_4_5__read;
  wire [512:0] fifo_B_PE_4_5__din;
  wire fifo_B_PE_4_5__full_n;
  wire fifo_B_PE_4_5__write;
  wire [512:0] fifo_B_PE_4_6__dout;
  wire fifo_B_PE_4_6__empty_n;
  wire fifo_B_PE_4_6__read;
  wire [512:0] fifo_B_PE_4_6__din;
  wire fifo_B_PE_4_6__full_n;
  wire fifo_B_PE_4_6__write;
  wire [512:0] fifo_B_PE_4_7__dout;
  wire fifo_B_PE_4_7__empty_n;
  wire fifo_B_PE_4_7__read;
  wire [512:0] fifo_B_PE_4_7__din;
  wire fifo_B_PE_4_7__full_n;
  wire fifo_B_PE_4_7__write;
  wire [512:0] fifo_B_PE_4_8__dout;
  wire fifo_B_PE_4_8__empty_n;
  wire fifo_B_PE_4_8__read;
  wire [512:0] fifo_B_PE_4_8__din;
  wire fifo_B_PE_4_8__full_n;
  wire fifo_B_PE_4_8__write;
  wire [512:0] fifo_B_PE_4_9__dout;
  wire fifo_B_PE_4_9__empty_n;
  wire fifo_B_PE_4_9__read;
  wire [512:0] fifo_B_PE_4_9__din;
  wire fifo_B_PE_4_9__full_n;
  wire fifo_B_PE_4_9__write;
  wire [512:0] fifo_B_PE_5_0__dout;
  wire fifo_B_PE_5_0__empty_n;
  wire fifo_B_PE_5_0__read;
  wire [512:0] fifo_B_PE_5_0__din;
  wire fifo_B_PE_5_0__full_n;
  wire fifo_B_PE_5_0__write;
  wire [512:0] fifo_B_PE_5_1__dout;
  wire fifo_B_PE_5_1__empty_n;
  wire fifo_B_PE_5_1__read;
  wire [512:0] fifo_B_PE_5_1__din;
  wire fifo_B_PE_5_1__full_n;
  wire fifo_B_PE_5_1__write;
  wire [512:0] fifo_B_PE_5_10__dout;
  wire fifo_B_PE_5_10__empty_n;
  wire fifo_B_PE_5_10__read;
  wire [512:0] fifo_B_PE_5_10__din;
  wire fifo_B_PE_5_10__full_n;
  wire fifo_B_PE_5_10__write;
  wire [512:0] fifo_B_PE_5_11__dout;
  wire fifo_B_PE_5_11__empty_n;
  wire fifo_B_PE_5_11__read;
  wire [512:0] fifo_B_PE_5_11__din;
  wire fifo_B_PE_5_11__full_n;
  wire fifo_B_PE_5_11__write;
  wire [512:0] fifo_B_PE_5_12__dout;
  wire fifo_B_PE_5_12__empty_n;
  wire fifo_B_PE_5_12__read;
  wire [512:0] fifo_B_PE_5_12__din;
  wire fifo_B_PE_5_12__full_n;
  wire fifo_B_PE_5_12__write;
  wire [512:0] fifo_B_PE_5_13__dout;
  wire fifo_B_PE_5_13__empty_n;
  wire fifo_B_PE_5_13__read;
  wire [512:0] fifo_B_PE_5_13__din;
  wire fifo_B_PE_5_13__full_n;
  wire fifo_B_PE_5_13__write;
  wire [512:0] fifo_B_PE_5_14__dout;
  wire fifo_B_PE_5_14__empty_n;
  wire fifo_B_PE_5_14__read;
  wire [512:0] fifo_B_PE_5_14__din;
  wire fifo_B_PE_5_14__full_n;
  wire fifo_B_PE_5_14__write;
  wire [512:0] fifo_B_PE_5_15__dout;
  wire fifo_B_PE_5_15__empty_n;
  wire fifo_B_PE_5_15__read;
  wire [512:0] fifo_B_PE_5_15__din;
  wire fifo_B_PE_5_15__full_n;
  wire fifo_B_PE_5_15__write;
  wire [512:0] fifo_B_PE_5_16__dout;
  wire fifo_B_PE_5_16__empty_n;
  wire fifo_B_PE_5_16__read;
  wire [512:0] fifo_B_PE_5_16__din;
  wire fifo_B_PE_5_16__full_n;
  wire fifo_B_PE_5_16__write;
  wire [512:0] fifo_B_PE_5_2__dout;
  wire fifo_B_PE_5_2__empty_n;
  wire fifo_B_PE_5_2__read;
  wire [512:0] fifo_B_PE_5_2__din;
  wire fifo_B_PE_5_2__full_n;
  wire fifo_B_PE_5_2__write;
  wire [512:0] fifo_B_PE_5_3__dout;
  wire fifo_B_PE_5_3__empty_n;
  wire fifo_B_PE_5_3__read;
  wire [512:0] fifo_B_PE_5_3__din;
  wire fifo_B_PE_5_3__full_n;
  wire fifo_B_PE_5_3__write;
  wire [512:0] fifo_B_PE_5_4__dout;
  wire fifo_B_PE_5_4__empty_n;
  wire fifo_B_PE_5_4__read;
  wire [512:0] fifo_B_PE_5_4__din;
  wire fifo_B_PE_5_4__full_n;
  wire fifo_B_PE_5_4__write;
  wire [512:0] fifo_B_PE_5_5__dout;
  wire fifo_B_PE_5_5__empty_n;
  wire fifo_B_PE_5_5__read;
  wire [512:0] fifo_B_PE_5_5__din;
  wire fifo_B_PE_5_5__full_n;
  wire fifo_B_PE_5_5__write;
  wire [512:0] fifo_B_PE_5_6__dout;
  wire fifo_B_PE_5_6__empty_n;
  wire fifo_B_PE_5_6__read;
  wire [512:0] fifo_B_PE_5_6__din;
  wire fifo_B_PE_5_6__full_n;
  wire fifo_B_PE_5_6__write;
  wire [512:0] fifo_B_PE_5_7__dout;
  wire fifo_B_PE_5_7__empty_n;
  wire fifo_B_PE_5_7__read;
  wire [512:0] fifo_B_PE_5_7__din;
  wire fifo_B_PE_5_7__full_n;
  wire fifo_B_PE_5_7__write;
  wire [512:0] fifo_B_PE_5_8__dout;
  wire fifo_B_PE_5_8__empty_n;
  wire fifo_B_PE_5_8__read;
  wire [512:0] fifo_B_PE_5_8__din;
  wire fifo_B_PE_5_8__full_n;
  wire fifo_B_PE_5_8__write;
  wire [512:0] fifo_B_PE_5_9__dout;
  wire fifo_B_PE_5_9__empty_n;
  wire fifo_B_PE_5_9__read;
  wire [512:0] fifo_B_PE_5_9__din;
  wire fifo_B_PE_5_9__full_n;
  wire fifo_B_PE_5_9__write;
  wire [512:0] fifo_B_PE_6_0__dout;
  wire fifo_B_PE_6_0__empty_n;
  wire fifo_B_PE_6_0__read;
  wire [512:0] fifo_B_PE_6_0__din;
  wire fifo_B_PE_6_0__full_n;
  wire fifo_B_PE_6_0__write;
  wire [512:0] fifo_B_PE_6_1__dout;
  wire fifo_B_PE_6_1__empty_n;
  wire fifo_B_PE_6_1__read;
  wire [512:0] fifo_B_PE_6_1__din;
  wire fifo_B_PE_6_1__full_n;
  wire fifo_B_PE_6_1__write;
  wire [512:0] fifo_B_PE_6_10__dout;
  wire fifo_B_PE_6_10__empty_n;
  wire fifo_B_PE_6_10__read;
  wire [512:0] fifo_B_PE_6_10__din;
  wire fifo_B_PE_6_10__full_n;
  wire fifo_B_PE_6_10__write;
  wire [512:0] fifo_B_PE_6_11__dout;
  wire fifo_B_PE_6_11__empty_n;
  wire fifo_B_PE_6_11__read;
  wire [512:0] fifo_B_PE_6_11__din;
  wire fifo_B_PE_6_11__full_n;
  wire fifo_B_PE_6_11__write;
  wire [512:0] fifo_B_PE_6_12__dout;
  wire fifo_B_PE_6_12__empty_n;
  wire fifo_B_PE_6_12__read;
  wire [512:0] fifo_B_PE_6_12__din;
  wire fifo_B_PE_6_12__full_n;
  wire fifo_B_PE_6_12__write;
  wire [512:0] fifo_B_PE_6_13__dout;
  wire fifo_B_PE_6_13__empty_n;
  wire fifo_B_PE_6_13__read;
  wire [512:0] fifo_B_PE_6_13__din;
  wire fifo_B_PE_6_13__full_n;
  wire fifo_B_PE_6_13__write;
  wire [512:0] fifo_B_PE_6_14__dout;
  wire fifo_B_PE_6_14__empty_n;
  wire fifo_B_PE_6_14__read;
  wire [512:0] fifo_B_PE_6_14__din;
  wire fifo_B_PE_6_14__full_n;
  wire fifo_B_PE_6_14__write;
  wire [512:0] fifo_B_PE_6_15__dout;
  wire fifo_B_PE_6_15__empty_n;
  wire fifo_B_PE_6_15__read;
  wire [512:0] fifo_B_PE_6_15__din;
  wire fifo_B_PE_6_15__full_n;
  wire fifo_B_PE_6_15__write;
  wire [512:0] fifo_B_PE_6_16__dout;
  wire fifo_B_PE_6_16__empty_n;
  wire fifo_B_PE_6_16__read;
  wire [512:0] fifo_B_PE_6_16__din;
  wire fifo_B_PE_6_16__full_n;
  wire fifo_B_PE_6_16__write;
  wire [512:0] fifo_B_PE_6_2__dout;
  wire fifo_B_PE_6_2__empty_n;
  wire fifo_B_PE_6_2__read;
  wire [512:0] fifo_B_PE_6_2__din;
  wire fifo_B_PE_6_2__full_n;
  wire fifo_B_PE_6_2__write;
  wire [512:0] fifo_B_PE_6_3__dout;
  wire fifo_B_PE_6_3__empty_n;
  wire fifo_B_PE_6_3__read;
  wire [512:0] fifo_B_PE_6_3__din;
  wire fifo_B_PE_6_3__full_n;
  wire fifo_B_PE_6_3__write;
  wire [512:0] fifo_B_PE_6_4__dout;
  wire fifo_B_PE_6_4__empty_n;
  wire fifo_B_PE_6_4__read;
  wire [512:0] fifo_B_PE_6_4__din;
  wire fifo_B_PE_6_4__full_n;
  wire fifo_B_PE_6_4__write;
  wire [512:0] fifo_B_PE_6_5__dout;
  wire fifo_B_PE_6_5__empty_n;
  wire fifo_B_PE_6_5__read;
  wire [512:0] fifo_B_PE_6_5__din;
  wire fifo_B_PE_6_5__full_n;
  wire fifo_B_PE_6_5__write;
  wire [512:0] fifo_B_PE_6_6__dout;
  wire fifo_B_PE_6_6__empty_n;
  wire fifo_B_PE_6_6__read;
  wire [512:0] fifo_B_PE_6_6__din;
  wire fifo_B_PE_6_6__full_n;
  wire fifo_B_PE_6_6__write;
  wire [512:0] fifo_B_PE_6_7__dout;
  wire fifo_B_PE_6_7__empty_n;
  wire fifo_B_PE_6_7__read;
  wire [512:0] fifo_B_PE_6_7__din;
  wire fifo_B_PE_6_7__full_n;
  wire fifo_B_PE_6_7__write;
  wire [512:0] fifo_B_PE_6_8__dout;
  wire fifo_B_PE_6_8__empty_n;
  wire fifo_B_PE_6_8__read;
  wire [512:0] fifo_B_PE_6_8__din;
  wire fifo_B_PE_6_8__full_n;
  wire fifo_B_PE_6_8__write;
  wire [512:0] fifo_B_PE_6_9__dout;
  wire fifo_B_PE_6_9__empty_n;
  wire fifo_B_PE_6_9__read;
  wire [512:0] fifo_B_PE_6_9__din;
  wire fifo_B_PE_6_9__full_n;
  wire fifo_B_PE_6_9__write;
  wire [512:0] fifo_B_PE_7_0__dout;
  wire fifo_B_PE_7_0__empty_n;
  wire fifo_B_PE_7_0__read;
  wire [512:0] fifo_B_PE_7_0__din;
  wire fifo_B_PE_7_0__full_n;
  wire fifo_B_PE_7_0__write;
  wire [512:0] fifo_B_PE_7_1__dout;
  wire fifo_B_PE_7_1__empty_n;
  wire fifo_B_PE_7_1__read;
  wire [512:0] fifo_B_PE_7_1__din;
  wire fifo_B_PE_7_1__full_n;
  wire fifo_B_PE_7_1__write;
  wire [512:0] fifo_B_PE_7_10__dout;
  wire fifo_B_PE_7_10__empty_n;
  wire fifo_B_PE_7_10__read;
  wire [512:0] fifo_B_PE_7_10__din;
  wire fifo_B_PE_7_10__full_n;
  wire fifo_B_PE_7_10__write;
  wire [512:0] fifo_B_PE_7_11__dout;
  wire fifo_B_PE_7_11__empty_n;
  wire fifo_B_PE_7_11__read;
  wire [512:0] fifo_B_PE_7_11__din;
  wire fifo_B_PE_7_11__full_n;
  wire fifo_B_PE_7_11__write;
  wire [512:0] fifo_B_PE_7_12__dout;
  wire fifo_B_PE_7_12__empty_n;
  wire fifo_B_PE_7_12__read;
  wire [512:0] fifo_B_PE_7_12__din;
  wire fifo_B_PE_7_12__full_n;
  wire fifo_B_PE_7_12__write;
  wire [512:0] fifo_B_PE_7_13__dout;
  wire fifo_B_PE_7_13__empty_n;
  wire fifo_B_PE_7_13__read;
  wire [512:0] fifo_B_PE_7_13__din;
  wire fifo_B_PE_7_13__full_n;
  wire fifo_B_PE_7_13__write;
  wire [512:0] fifo_B_PE_7_14__dout;
  wire fifo_B_PE_7_14__empty_n;
  wire fifo_B_PE_7_14__read;
  wire [512:0] fifo_B_PE_7_14__din;
  wire fifo_B_PE_7_14__full_n;
  wire fifo_B_PE_7_14__write;
  wire [512:0] fifo_B_PE_7_15__dout;
  wire fifo_B_PE_7_15__empty_n;
  wire fifo_B_PE_7_15__read;
  wire [512:0] fifo_B_PE_7_15__din;
  wire fifo_B_PE_7_15__full_n;
  wire fifo_B_PE_7_15__write;
  wire [512:0] fifo_B_PE_7_16__dout;
  wire fifo_B_PE_7_16__empty_n;
  wire fifo_B_PE_7_16__read;
  wire [512:0] fifo_B_PE_7_16__din;
  wire fifo_B_PE_7_16__full_n;
  wire fifo_B_PE_7_16__write;
  wire [512:0] fifo_B_PE_7_2__dout;
  wire fifo_B_PE_7_2__empty_n;
  wire fifo_B_PE_7_2__read;
  wire [512:0] fifo_B_PE_7_2__din;
  wire fifo_B_PE_7_2__full_n;
  wire fifo_B_PE_7_2__write;
  wire [512:0] fifo_B_PE_7_3__dout;
  wire fifo_B_PE_7_3__empty_n;
  wire fifo_B_PE_7_3__read;
  wire [512:0] fifo_B_PE_7_3__din;
  wire fifo_B_PE_7_3__full_n;
  wire fifo_B_PE_7_3__write;
  wire [512:0] fifo_B_PE_7_4__dout;
  wire fifo_B_PE_7_4__empty_n;
  wire fifo_B_PE_7_4__read;
  wire [512:0] fifo_B_PE_7_4__din;
  wire fifo_B_PE_7_4__full_n;
  wire fifo_B_PE_7_4__write;
  wire [512:0] fifo_B_PE_7_5__dout;
  wire fifo_B_PE_7_5__empty_n;
  wire fifo_B_PE_7_5__read;
  wire [512:0] fifo_B_PE_7_5__din;
  wire fifo_B_PE_7_5__full_n;
  wire fifo_B_PE_7_5__write;
  wire [512:0] fifo_B_PE_7_6__dout;
  wire fifo_B_PE_7_6__empty_n;
  wire fifo_B_PE_7_6__read;
  wire [512:0] fifo_B_PE_7_6__din;
  wire fifo_B_PE_7_6__full_n;
  wire fifo_B_PE_7_6__write;
  wire [512:0] fifo_B_PE_7_7__dout;
  wire fifo_B_PE_7_7__empty_n;
  wire fifo_B_PE_7_7__read;
  wire [512:0] fifo_B_PE_7_7__din;
  wire fifo_B_PE_7_7__full_n;
  wire fifo_B_PE_7_7__write;
  wire [512:0] fifo_B_PE_7_8__dout;
  wire fifo_B_PE_7_8__empty_n;
  wire fifo_B_PE_7_8__read;
  wire [512:0] fifo_B_PE_7_8__din;
  wire fifo_B_PE_7_8__full_n;
  wire fifo_B_PE_7_8__write;
  wire [512:0] fifo_B_PE_7_9__dout;
  wire fifo_B_PE_7_9__empty_n;
  wire fifo_B_PE_7_9__read;
  wire [512:0] fifo_B_PE_7_9__din;
  wire fifo_B_PE_7_9__full_n;
  wire fifo_B_PE_7_9__write;
  wire [512:0] fifo_B_PE_8_0__dout;
  wire fifo_B_PE_8_0__empty_n;
  wire fifo_B_PE_8_0__read;
  wire [512:0] fifo_B_PE_8_0__din;
  wire fifo_B_PE_8_0__full_n;
  wire fifo_B_PE_8_0__write;
  wire [512:0] fifo_B_PE_8_1__dout;
  wire fifo_B_PE_8_1__empty_n;
  wire fifo_B_PE_8_1__read;
  wire [512:0] fifo_B_PE_8_1__din;
  wire fifo_B_PE_8_1__full_n;
  wire fifo_B_PE_8_1__write;
  wire [512:0] fifo_B_PE_8_10__dout;
  wire fifo_B_PE_8_10__empty_n;
  wire fifo_B_PE_8_10__read;
  wire [512:0] fifo_B_PE_8_10__din;
  wire fifo_B_PE_8_10__full_n;
  wire fifo_B_PE_8_10__write;
  wire [512:0] fifo_B_PE_8_11__dout;
  wire fifo_B_PE_8_11__empty_n;
  wire fifo_B_PE_8_11__read;
  wire [512:0] fifo_B_PE_8_11__din;
  wire fifo_B_PE_8_11__full_n;
  wire fifo_B_PE_8_11__write;
  wire [512:0] fifo_B_PE_8_12__dout;
  wire fifo_B_PE_8_12__empty_n;
  wire fifo_B_PE_8_12__read;
  wire [512:0] fifo_B_PE_8_12__din;
  wire fifo_B_PE_8_12__full_n;
  wire fifo_B_PE_8_12__write;
  wire [512:0] fifo_B_PE_8_13__dout;
  wire fifo_B_PE_8_13__empty_n;
  wire fifo_B_PE_8_13__read;
  wire [512:0] fifo_B_PE_8_13__din;
  wire fifo_B_PE_8_13__full_n;
  wire fifo_B_PE_8_13__write;
  wire [512:0] fifo_B_PE_8_14__dout;
  wire fifo_B_PE_8_14__empty_n;
  wire fifo_B_PE_8_14__read;
  wire [512:0] fifo_B_PE_8_14__din;
  wire fifo_B_PE_8_14__full_n;
  wire fifo_B_PE_8_14__write;
  wire [512:0] fifo_B_PE_8_15__dout;
  wire fifo_B_PE_8_15__empty_n;
  wire fifo_B_PE_8_15__read;
  wire [512:0] fifo_B_PE_8_15__din;
  wire fifo_B_PE_8_15__full_n;
  wire fifo_B_PE_8_15__write;
  wire [512:0] fifo_B_PE_8_16__dout;
  wire fifo_B_PE_8_16__empty_n;
  wire fifo_B_PE_8_16__read;
  wire [512:0] fifo_B_PE_8_16__din;
  wire fifo_B_PE_8_16__full_n;
  wire fifo_B_PE_8_16__write;
  wire [512:0] fifo_B_PE_8_2__dout;
  wire fifo_B_PE_8_2__empty_n;
  wire fifo_B_PE_8_2__read;
  wire [512:0] fifo_B_PE_8_2__din;
  wire fifo_B_PE_8_2__full_n;
  wire fifo_B_PE_8_2__write;
  wire [512:0] fifo_B_PE_8_3__dout;
  wire fifo_B_PE_8_3__empty_n;
  wire fifo_B_PE_8_3__read;
  wire [512:0] fifo_B_PE_8_3__din;
  wire fifo_B_PE_8_3__full_n;
  wire fifo_B_PE_8_3__write;
  wire [512:0] fifo_B_PE_8_4__dout;
  wire fifo_B_PE_8_4__empty_n;
  wire fifo_B_PE_8_4__read;
  wire [512:0] fifo_B_PE_8_4__din;
  wire fifo_B_PE_8_4__full_n;
  wire fifo_B_PE_8_4__write;
  wire [512:0] fifo_B_PE_8_5__dout;
  wire fifo_B_PE_8_5__empty_n;
  wire fifo_B_PE_8_5__read;
  wire [512:0] fifo_B_PE_8_5__din;
  wire fifo_B_PE_8_5__full_n;
  wire fifo_B_PE_8_5__write;
  wire [512:0] fifo_B_PE_8_6__dout;
  wire fifo_B_PE_8_6__empty_n;
  wire fifo_B_PE_8_6__read;
  wire [512:0] fifo_B_PE_8_6__din;
  wire fifo_B_PE_8_6__full_n;
  wire fifo_B_PE_8_6__write;
  wire [512:0] fifo_B_PE_8_7__dout;
  wire fifo_B_PE_8_7__empty_n;
  wire fifo_B_PE_8_7__read;
  wire [512:0] fifo_B_PE_8_7__din;
  wire fifo_B_PE_8_7__full_n;
  wire fifo_B_PE_8_7__write;
  wire [512:0] fifo_B_PE_8_8__dout;
  wire fifo_B_PE_8_8__empty_n;
  wire fifo_B_PE_8_8__read;
  wire [512:0] fifo_B_PE_8_8__din;
  wire fifo_B_PE_8_8__full_n;
  wire fifo_B_PE_8_8__write;
  wire [512:0] fifo_B_PE_8_9__dout;
  wire fifo_B_PE_8_9__empty_n;
  wire fifo_B_PE_8_9__read;
  wire [512:0] fifo_B_PE_8_9__din;
  wire fifo_B_PE_8_9__full_n;
  wire fifo_B_PE_8_9__write;
  wire [512:0] fifo_B_PE_9_0__dout;
  wire fifo_B_PE_9_0__empty_n;
  wire fifo_B_PE_9_0__read;
  wire [512:0] fifo_B_PE_9_0__din;
  wire fifo_B_PE_9_0__full_n;
  wire fifo_B_PE_9_0__write;
  wire [512:0] fifo_B_PE_9_1__dout;
  wire fifo_B_PE_9_1__empty_n;
  wire fifo_B_PE_9_1__read;
  wire [512:0] fifo_B_PE_9_1__din;
  wire fifo_B_PE_9_1__full_n;
  wire fifo_B_PE_9_1__write;
  wire [512:0] fifo_B_PE_9_10__dout;
  wire fifo_B_PE_9_10__empty_n;
  wire fifo_B_PE_9_10__read;
  wire [512:0] fifo_B_PE_9_10__din;
  wire fifo_B_PE_9_10__full_n;
  wire fifo_B_PE_9_10__write;
  wire [512:0] fifo_B_PE_9_11__dout;
  wire fifo_B_PE_9_11__empty_n;
  wire fifo_B_PE_9_11__read;
  wire [512:0] fifo_B_PE_9_11__din;
  wire fifo_B_PE_9_11__full_n;
  wire fifo_B_PE_9_11__write;
  wire [512:0] fifo_B_PE_9_12__dout;
  wire fifo_B_PE_9_12__empty_n;
  wire fifo_B_PE_9_12__read;
  wire [512:0] fifo_B_PE_9_12__din;
  wire fifo_B_PE_9_12__full_n;
  wire fifo_B_PE_9_12__write;
  wire [512:0] fifo_B_PE_9_13__dout;
  wire fifo_B_PE_9_13__empty_n;
  wire fifo_B_PE_9_13__read;
  wire [512:0] fifo_B_PE_9_13__din;
  wire fifo_B_PE_9_13__full_n;
  wire fifo_B_PE_9_13__write;
  wire [512:0] fifo_B_PE_9_14__dout;
  wire fifo_B_PE_9_14__empty_n;
  wire fifo_B_PE_9_14__read;
  wire [512:0] fifo_B_PE_9_14__din;
  wire fifo_B_PE_9_14__full_n;
  wire fifo_B_PE_9_14__write;
  wire [512:0] fifo_B_PE_9_15__dout;
  wire fifo_B_PE_9_15__empty_n;
  wire fifo_B_PE_9_15__read;
  wire [512:0] fifo_B_PE_9_15__din;
  wire fifo_B_PE_9_15__full_n;
  wire fifo_B_PE_9_15__write;
  wire [512:0] fifo_B_PE_9_16__dout;
  wire fifo_B_PE_9_16__empty_n;
  wire fifo_B_PE_9_16__read;
  wire [512:0] fifo_B_PE_9_16__din;
  wire fifo_B_PE_9_16__full_n;
  wire fifo_B_PE_9_16__write;
  wire [512:0] fifo_B_PE_9_2__dout;
  wire fifo_B_PE_9_2__empty_n;
  wire fifo_B_PE_9_2__read;
  wire [512:0] fifo_B_PE_9_2__din;
  wire fifo_B_PE_9_2__full_n;
  wire fifo_B_PE_9_2__write;
  wire [512:0] fifo_B_PE_9_3__dout;
  wire fifo_B_PE_9_3__empty_n;
  wire fifo_B_PE_9_3__read;
  wire [512:0] fifo_B_PE_9_3__din;
  wire fifo_B_PE_9_3__full_n;
  wire fifo_B_PE_9_3__write;
  wire [512:0] fifo_B_PE_9_4__dout;
  wire fifo_B_PE_9_4__empty_n;
  wire fifo_B_PE_9_4__read;
  wire [512:0] fifo_B_PE_9_4__din;
  wire fifo_B_PE_9_4__full_n;
  wire fifo_B_PE_9_4__write;
  wire [512:0] fifo_B_PE_9_5__dout;
  wire fifo_B_PE_9_5__empty_n;
  wire fifo_B_PE_9_5__read;
  wire [512:0] fifo_B_PE_9_5__din;
  wire fifo_B_PE_9_5__full_n;
  wire fifo_B_PE_9_5__write;
  wire [512:0] fifo_B_PE_9_6__dout;
  wire fifo_B_PE_9_6__empty_n;
  wire fifo_B_PE_9_6__read;
  wire [512:0] fifo_B_PE_9_6__din;
  wire fifo_B_PE_9_6__full_n;
  wire fifo_B_PE_9_6__write;
  wire [512:0] fifo_B_PE_9_7__dout;
  wire fifo_B_PE_9_7__empty_n;
  wire fifo_B_PE_9_7__read;
  wire [512:0] fifo_B_PE_9_7__din;
  wire fifo_B_PE_9_7__full_n;
  wire fifo_B_PE_9_7__write;
  wire [512:0] fifo_B_PE_9_8__dout;
  wire fifo_B_PE_9_8__empty_n;
  wire fifo_B_PE_9_8__read;
  wire [512:0] fifo_B_PE_9_8__din;
  wire fifo_B_PE_9_8__full_n;
  wire fifo_B_PE_9_8__write;
  wire [512:0] fifo_B_PE_9_9__dout;
  wire fifo_B_PE_9_9__empty_n;
  wire fifo_B_PE_9_9__read;
  wire [512:0] fifo_B_PE_9_9__din;
  wire fifo_B_PE_9_9__full_n;
  wire fifo_B_PE_9_9__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_0_0__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_0_0__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_0_0__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_0_0__din;
  wire fifo_C_drain_C_drain_IO_L1_out_0_0__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_0_0__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_0_1__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_0_1__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_0_1__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_0_1__din;
  wire fifo_C_drain_C_drain_IO_L1_out_0_1__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_0_1__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_0_10__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_0_10__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_0_10__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_0_10__din;
  wire fifo_C_drain_C_drain_IO_L1_out_0_10__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_0_10__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_0_11__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_0_11__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_0_11__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_0_11__din;
  wire fifo_C_drain_C_drain_IO_L1_out_0_11__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_0_11__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_0_12__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_0_12__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_0_12__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_0_12__din;
  wire fifo_C_drain_C_drain_IO_L1_out_0_12__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_0_12__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_0_13__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_0_13__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_0_13__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_0_13__din;
  wire fifo_C_drain_C_drain_IO_L1_out_0_13__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_0_13__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_0_14__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_0_14__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_0_14__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_0_14__din;
  wire fifo_C_drain_C_drain_IO_L1_out_0_14__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_0_14__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_0_15__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_0_15__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_0_15__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_0_15__din;
  wire fifo_C_drain_C_drain_IO_L1_out_0_15__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_0_15__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_0_16__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_0_16__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_0_16__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_0_16__din;
  wire fifo_C_drain_C_drain_IO_L1_out_0_16__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_0_16__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_0_17__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_0_17__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_0_17__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_0_17__din;
  wire fifo_C_drain_C_drain_IO_L1_out_0_17__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_0_17__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_0_2__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_0_2__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_0_2__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_0_2__din;
  wire fifo_C_drain_C_drain_IO_L1_out_0_2__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_0_2__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_0_3__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_0_3__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_0_3__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_0_3__din;
  wire fifo_C_drain_C_drain_IO_L1_out_0_3__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_0_3__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_0_4__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_0_4__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_0_4__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_0_4__din;
  wire fifo_C_drain_C_drain_IO_L1_out_0_4__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_0_4__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_0_5__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_0_5__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_0_5__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_0_5__din;
  wire fifo_C_drain_C_drain_IO_L1_out_0_5__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_0_5__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_0_6__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_0_6__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_0_6__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_0_6__din;
  wire fifo_C_drain_C_drain_IO_L1_out_0_6__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_0_6__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_0_7__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_0_7__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_0_7__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_0_7__din;
  wire fifo_C_drain_C_drain_IO_L1_out_0_7__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_0_7__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_0_8__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_0_8__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_0_8__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_0_8__din;
  wire fifo_C_drain_C_drain_IO_L1_out_0_8__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_0_8__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_0_9__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_0_9__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_0_9__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_0_9__din;
  wire fifo_C_drain_C_drain_IO_L1_out_0_9__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_0_9__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_10_0__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_10_0__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_10_0__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_10_0__din;
  wire fifo_C_drain_C_drain_IO_L1_out_10_0__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_10_0__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_10_1__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_10_1__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_10_1__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_10_1__din;
  wire fifo_C_drain_C_drain_IO_L1_out_10_1__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_10_1__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_10_10__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_10_10__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_10_10__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_10_10__din;
  wire fifo_C_drain_C_drain_IO_L1_out_10_10__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_10_10__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_10_11__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_10_11__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_10_11__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_10_11__din;
  wire fifo_C_drain_C_drain_IO_L1_out_10_11__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_10_11__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_10_12__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_10_12__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_10_12__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_10_12__din;
  wire fifo_C_drain_C_drain_IO_L1_out_10_12__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_10_12__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_10_13__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_10_13__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_10_13__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_10_13__din;
  wire fifo_C_drain_C_drain_IO_L1_out_10_13__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_10_13__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_10_14__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_10_14__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_10_14__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_10_14__din;
  wire fifo_C_drain_C_drain_IO_L1_out_10_14__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_10_14__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_10_15__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_10_15__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_10_15__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_10_15__din;
  wire fifo_C_drain_C_drain_IO_L1_out_10_15__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_10_15__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_10_16__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_10_16__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_10_16__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_10_16__din;
  wire fifo_C_drain_C_drain_IO_L1_out_10_16__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_10_16__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_10_17__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_10_17__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_10_17__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_10_17__din;
  wire fifo_C_drain_C_drain_IO_L1_out_10_17__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_10_17__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_10_2__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_10_2__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_10_2__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_10_2__din;
  wire fifo_C_drain_C_drain_IO_L1_out_10_2__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_10_2__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_10_3__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_10_3__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_10_3__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_10_3__din;
  wire fifo_C_drain_C_drain_IO_L1_out_10_3__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_10_3__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_10_4__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_10_4__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_10_4__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_10_4__din;
  wire fifo_C_drain_C_drain_IO_L1_out_10_4__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_10_4__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_10_5__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_10_5__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_10_5__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_10_5__din;
  wire fifo_C_drain_C_drain_IO_L1_out_10_5__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_10_5__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_10_6__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_10_6__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_10_6__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_10_6__din;
  wire fifo_C_drain_C_drain_IO_L1_out_10_6__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_10_6__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_10_7__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_10_7__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_10_7__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_10_7__din;
  wire fifo_C_drain_C_drain_IO_L1_out_10_7__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_10_7__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_10_8__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_10_8__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_10_8__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_10_8__din;
  wire fifo_C_drain_C_drain_IO_L1_out_10_8__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_10_8__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_10_9__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_10_9__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_10_9__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_10_9__din;
  wire fifo_C_drain_C_drain_IO_L1_out_10_9__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_10_9__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_11_0__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_11_0__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_11_0__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_11_0__din;
  wire fifo_C_drain_C_drain_IO_L1_out_11_0__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_11_0__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_11_1__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_11_1__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_11_1__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_11_1__din;
  wire fifo_C_drain_C_drain_IO_L1_out_11_1__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_11_1__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_11_10__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_11_10__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_11_10__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_11_10__din;
  wire fifo_C_drain_C_drain_IO_L1_out_11_10__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_11_10__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_11_11__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_11_11__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_11_11__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_11_11__din;
  wire fifo_C_drain_C_drain_IO_L1_out_11_11__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_11_11__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_11_12__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_11_12__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_11_12__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_11_12__din;
  wire fifo_C_drain_C_drain_IO_L1_out_11_12__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_11_12__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_11_13__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_11_13__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_11_13__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_11_13__din;
  wire fifo_C_drain_C_drain_IO_L1_out_11_13__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_11_13__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_11_14__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_11_14__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_11_14__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_11_14__din;
  wire fifo_C_drain_C_drain_IO_L1_out_11_14__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_11_14__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_11_15__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_11_15__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_11_15__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_11_15__din;
  wire fifo_C_drain_C_drain_IO_L1_out_11_15__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_11_15__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_11_16__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_11_16__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_11_16__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_11_16__din;
  wire fifo_C_drain_C_drain_IO_L1_out_11_16__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_11_16__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_11_17__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_11_17__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_11_17__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_11_17__din;
  wire fifo_C_drain_C_drain_IO_L1_out_11_17__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_11_17__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_11_2__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_11_2__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_11_2__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_11_2__din;
  wire fifo_C_drain_C_drain_IO_L1_out_11_2__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_11_2__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_11_3__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_11_3__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_11_3__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_11_3__din;
  wire fifo_C_drain_C_drain_IO_L1_out_11_3__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_11_3__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_11_4__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_11_4__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_11_4__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_11_4__din;
  wire fifo_C_drain_C_drain_IO_L1_out_11_4__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_11_4__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_11_5__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_11_5__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_11_5__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_11_5__din;
  wire fifo_C_drain_C_drain_IO_L1_out_11_5__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_11_5__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_11_6__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_11_6__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_11_6__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_11_6__din;
  wire fifo_C_drain_C_drain_IO_L1_out_11_6__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_11_6__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_11_7__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_11_7__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_11_7__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_11_7__din;
  wire fifo_C_drain_C_drain_IO_L1_out_11_7__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_11_7__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_11_8__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_11_8__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_11_8__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_11_8__din;
  wire fifo_C_drain_C_drain_IO_L1_out_11_8__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_11_8__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_11_9__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_11_9__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_11_9__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_11_9__din;
  wire fifo_C_drain_C_drain_IO_L1_out_11_9__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_11_9__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_12_0__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_12_0__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_12_0__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_12_0__din;
  wire fifo_C_drain_C_drain_IO_L1_out_12_0__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_12_0__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_12_1__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_12_1__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_12_1__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_12_1__din;
  wire fifo_C_drain_C_drain_IO_L1_out_12_1__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_12_1__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_12_10__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_12_10__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_12_10__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_12_10__din;
  wire fifo_C_drain_C_drain_IO_L1_out_12_10__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_12_10__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_12_11__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_12_11__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_12_11__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_12_11__din;
  wire fifo_C_drain_C_drain_IO_L1_out_12_11__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_12_11__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_12_12__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_12_12__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_12_12__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_12_12__din;
  wire fifo_C_drain_C_drain_IO_L1_out_12_12__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_12_12__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_12_13__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_12_13__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_12_13__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_12_13__din;
  wire fifo_C_drain_C_drain_IO_L1_out_12_13__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_12_13__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_12_14__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_12_14__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_12_14__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_12_14__din;
  wire fifo_C_drain_C_drain_IO_L1_out_12_14__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_12_14__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_12_15__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_12_15__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_12_15__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_12_15__din;
  wire fifo_C_drain_C_drain_IO_L1_out_12_15__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_12_15__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_12_16__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_12_16__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_12_16__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_12_16__din;
  wire fifo_C_drain_C_drain_IO_L1_out_12_16__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_12_16__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_12_17__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_12_17__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_12_17__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_12_17__din;
  wire fifo_C_drain_C_drain_IO_L1_out_12_17__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_12_17__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_12_2__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_12_2__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_12_2__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_12_2__din;
  wire fifo_C_drain_C_drain_IO_L1_out_12_2__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_12_2__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_12_3__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_12_3__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_12_3__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_12_3__din;
  wire fifo_C_drain_C_drain_IO_L1_out_12_3__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_12_3__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_12_4__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_12_4__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_12_4__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_12_4__din;
  wire fifo_C_drain_C_drain_IO_L1_out_12_4__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_12_4__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_12_5__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_12_5__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_12_5__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_12_5__din;
  wire fifo_C_drain_C_drain_IO_L1_out_12_5__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_12_5__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_12_6__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_12_6__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_12_6__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_12_6__din;
  wire fifo_C_drain_C_drain_IO_L1_out_12_6__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_12_6__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_12_7__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_12_7__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_12_7__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_12_7__din;
  wire fifo_C_drain_C_drain_IO_L1_out_12_7__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_12_7__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_12_8__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_12_8__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_12_8__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_12_8__din;
  wire fifo_C_drain_C_drain_IO_L1_out_12_8__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_12_8__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_12_9__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_12_9__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_12_9__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_12_9__din;
  wire fifo_C_drain_C_drain_IO_L1_out_12_9__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_12_9__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_13_0__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_13_0__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_13_0__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_13_0__din;
  wire fifo_C_drain_C_drain_IO_L1_out_13_0__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_13_0__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_13_1__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_13_1__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_13_1__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_13_1__din;
  wire fifo_C_drain_C_drain_IO_L1_out_13_1__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_13_1__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_13_10__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_13_10__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_13_10__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_13_10__din;
  wire fifo_C_drain_C_drain_IO_L1_out_13_10__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_13_10__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_13_11__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_13_11__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_13_11__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_13_11__din;
  wire fifo_C_drain_C_drain_IO_L1_out_13_11__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_13_11__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_13_12__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_13_12__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_13_12__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_13_12__din;
  wire fifo_C_drain_C_drain_IO_L1_out_13_12__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_13_12__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_13_13__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_13_13__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_13_13__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_13_13__din;
  wire fifo_C_drain_C_drain_IO_L1_out_13_13__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_13_13__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_13_14__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_13_14__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_13_14__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_13_14__din;
  wire fifo_C_drain_C_drain_IO_L1_out_13_14__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_13_14__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_13_15__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_13_15__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_13_15__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_13_15__din;
  wire fifo_C_drain_C_drain_IO_L1_out_13_15__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_13_15__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_13_16__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_13_16__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_13_16__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_13_16__din;
  wire fifo_C_drain_C_drain_IO_L1_out_13_16__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_13_16__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_13_17__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_13_17__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_13_17__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_13_17__din;
  wire fifo_C_drain_C_drain_IO_L1_out_13_17__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_13_17__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_13_2__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_13_2__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_13_2__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_13_2__din;
  wire fifo_C_drain_C_drain_IO_L1_out_13_2__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_13_2__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_13_3__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_13_3__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_13_3__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_13_3__din;
  wire fifo_C_drain_C_drain_IO_L1_out_13_3__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_13_3__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_13_4__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_13_4__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_13_4__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_13_4__din;
  wire fifo_C_drain_C_drain_IO_L1_out_13_4__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_13_4__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_13_5__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_13_5__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_13_5__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_13_5__din;
  wire fifo_C_drain_C_drain_IO_L1_out_13_5__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_13_5__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_13_6__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_13_6__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_13_6__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_13_6__din;
  wire fifo_C_drain_C_drain_IO_L1_out_13_6__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_13_6__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_13_7__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_13_7__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_13_7__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_13_7__din;
  wire fifo_C_drain_C_drain_IO_L1_out_13_7__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_13_7__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_13_8__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_13_8__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_13_8__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_13_8__din;
  wire fifo_C_drain_C_drain_IO_L1_out_13_8__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_13_8__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_13_9__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_13_9__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_13_9__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_13_9__din;
  wire fifo_C_drain_C_drain_IO_L1_out_13_9__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_13_9__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_14_0__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_14_0__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_14_0__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_14_0__din;
  wire fifo_C_drain_C_drain_IO_L1_out_14_0__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_14_0__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_14_1__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_14_1__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_14_1__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_14_1__din;
  wire fifo_C_drain_C_drain_IO_L1_out_14_1__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_14_1__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_14_10__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_14_10__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_14_10__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_14_10__din;
  wire fifo_C_drain_C_drain_IO_L1_out_14_10__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_14_10__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_14_11__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_14_11__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_14_11__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_14_11__din;
  wire fifo_C_drain_C_drain_IO_L1_out_14_11__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_14_11__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_14_12__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_14_12__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_14_12__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_14_12__din;
  wire fifo_C_drain_C_drain_IO_L1_out_14_12__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_14_12__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_14_13__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_14_13__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_14_13__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_14_13__din;
  wire fifo_C_drain_C_drain_IO_L1_out_14_13__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_14_13__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_14_14__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_14_14__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_14_14__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_14_14__din;
  wire fifo_C_drain_C_drain_IO_L1_out_14_14__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_14_14__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_14_15__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_14_15__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_14_15__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_14_15__din;
  wire fifo_C_drain_C_drain_IO_L1_out_14_15__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_14_15__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_14_16__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_14_16__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_14_16__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_14_16__din;
  wire fifo_C_drain_C_drain_IO_L1_out_14_16__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_14_16__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_14_17__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_14_17__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_14_17__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_14_17__din;
  wire fifo_C_drain_C_drain_IO_L1_out_14_17__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_14_17__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_14_2__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_14_2__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_14_2__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_14_2__din;
  wire fifo_C_drain_C_drain_IO_L1_out_14_2__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_14_2__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_14_3__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_14_3__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_14_3__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_14_3__din;
  wire fifo_C_drain_C_drain_IO_L1_out_14_3__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_14_3__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_14_4__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_14_4__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_14_4__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_14_4__din;
  wire fifo_C_drain_C_drain_IO_L1_out_14_4__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_14_4__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_14_5__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_14_5__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_14_5__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_14_5__din;
  wire fifo_C_drain_C_drain_IO_L1_out_14_5__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_14_5__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_14_6__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_14_6__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_14_6__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_14_6__din;
  wire fifo_C_drain_C_drain_IO_L1_out_14_6__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_14_6__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_14_7__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_14_7__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_14_7__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_14_7__din;
  wire fifo_C_drain_C_drain_IO_L1_out_14_7__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_14_7__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_14_8__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_14_8__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_14_8__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_14_8__din;
  wire fifo_C_drain_C_drain_IO_L1_out_14_8__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_14_8__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_14_9__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_14_9__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_14_9__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_14_9__din;
  wire fifo_C_drain_C_drain_IO_L1_out_14_9__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_14_9__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_15_0__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_15_0__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_15_0__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_15_0__din;
  wire fifo_C_drain_C_drain_IO_L1_out_15_0__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_15_0__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_15_1__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_15_1__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_15_1__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_15_1__din;
  wire fifo_C_drain_C_drain_IO_L1_out_15_1__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_15_1__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_15_10__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_15_10__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_15_10__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_15_10__din;
  wire fifo_C_drain_C_drain_IO_L1_out_15_10__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_15_10__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_15_11__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_15_11__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_15_11__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_15_11__din;
  wire fifo_C_drain_C_drain_IO_L1_out_15_11__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_15_11__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_15_12__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_15_12__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_15_12__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_15_12__din;
  wire fifo_C_drain_C_drain_IO_L1_out_15_12__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_15_12__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_15_13__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_15_13__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_15_13__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_15_13__din;
  wire fifo_C_drain_C_drain_IO_L1_out_15_13__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_15_13__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_15_14__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_15_14__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_15_14__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_15_14__din;
  wire fifo_C_drain_C_drain_IO_L1_out_15_14__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_15_14__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_15_15__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_15_15__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_15_15__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_15_15__din;
  wire fifo_C_drain_C_drain_IO_L1_out_15_15__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_15_15__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_15_16__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_15_16__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_15_16__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_15_16__din;
  wire fifo_C_drain_C_drain_IO_L1_out_15_16__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_15_16__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_15_17__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_15_17__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_15_17__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_15_17__din;
  wire fifo_C_drain_C_drain_IO_L1_out_15_17__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_15_17__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_15_2__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_15_2__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_15_2__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_15_2__din;
  wire fifo_C_drain_C_drain_IO_L1_out_15_2__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_15_2__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_15_3__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_15_3__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_15_3__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_15_3__din;
  wire fifo_C_drain_C_drain_IO_L1_out_15_3__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_15_3__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_15_4__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_15_4__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_15_4__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_15_4__din;
  wire fifo_C_drain_C_drain_IO_L1_out_15_4__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_15_4__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_15_5__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_15_5__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_15_5__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_15_5__din;
  wire fifo_C_drain_C_drain_IO_L1_out_15_5__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_15_5__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_15_6__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_15_6__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_15_6__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_15_6__din;
  wire fifo_C_drain_C_drain_IO_L1_out_15_6__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_15_6__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_15_7__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_15_7__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_15_7__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_15_7__din;
  wire fifo_C_drain_C_drain_IO_L1_out_15_7__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_15_7__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_15_8__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_15_8__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_15_8__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_15_8__din;
  wire fifo_C_drain_C_drain_IO_L1_out_15_8__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_15_8__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_15_9__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_15_9__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_15_9__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_15_9__din;
  wire fifo_C_drain_C_drain_IO_L1_out_15_9__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_15_9__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_16_0__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_16_0__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_16_0__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_16_0__din;
  wire fifo_C_drain_C_drain_IO_L1_out_16_0__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_16_0__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_16_1__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_16_1__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_16_1__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_16_1__din;
  wire fifo_C_drain_C_drain_IO_L1_out_16_1__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_16_1__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_16_10__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_16_10__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_16_10__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_16_10__din;
  wire fifo_C_drain_C_drain_IO_L1_out_16_10__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_16_10__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_16_11__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_16_11__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_16_11__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_16_11__din;
  wire fifo_C_drain_C_drain_IO_L1_out_16_11__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_16_11__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_16_12__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_16_12__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_16_12__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_16_12__din;
  wire fifo_C_drain_C_drain_IO_L1_out_16_12__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_16_12__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_16_13__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_16_13__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_16_13__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_16_13__din;
  wire fifo_C_drain_C_drain_IO_L1_out_16_13__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_16_13__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_16_14__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_16_14__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_16_14__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_16_14__din;
  wire fifo_C_drain_C_drain_IO_L1_out_16_14__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_16_14__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_16_15__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_16_15__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_16_15__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_16_15__din;
  wire fifo_C_drain_C_drain_IO_L1_out_16_15__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_16_15__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_16_16__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_16_16__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_16_16__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_16_16__din;
  wire fifo_C_drain_C_drain_IO_L1_out_16_16__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_16_16__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_16_17__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_16_17__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_16_17__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_16_17__din;
  wire fifo_C_drain_C_drain_IO_L1_out_16_17__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_16_17__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_16_2__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_16_2__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_16_2__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_16_2__din;
  wire fifo_C_drain_C_drain_IO_L1_out_16_2__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_16_2__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_16_3__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_16_3__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_16_3__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_16_3__din;
  wire fifo_C_drain_C_drain_IO_L1_out_16_3__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_16_3__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_16_4__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_16_4__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_16_4__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_16_4__din;
  wire fifo_C_drain_C_drain_IO_L1_out_16_4__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_16_4__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_16_5__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_16_5__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_16_5__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_16_5__din;
  wire fifo_C_drain_C_drain_IO_L1_out_16_5__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_16_5__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_16_6__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_16_6__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_16_6__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_16_6__din;
  wire fifo_C_drain_C_drain_IO_L1_out_16_6__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_16_6__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_16_7__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_16_7__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_16_7__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_16_7__din;
  wire fifo_C_drain_C_drain_IO_L1_out_16_7__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_16_7__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_16_8__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_16_8__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_16_8__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_16_8__din;
  wire fifo_C_drain_C_drain_IO_L1_out_16_8__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_16_8__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_16_9__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_16_9__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_16_9__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_16_9__din;
  wire fifo_C_drain_C_drain_IO_L1_out_16_9__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_16_9__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_1_0__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_1_0__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_1_0__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_1_0__din;
  wire fifo_C_drain_C_drain_IO_L1_out_1_0__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_1_0__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_1_1__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_1_1__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_1_1__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_1_1__din;
  wire fifo_C_drain_C_drain_IO_L1_out_1_1__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_1_1__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_1_10__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_1_10__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_1_10__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_1_10__din;
  wire fifo_C_drain_C_drain_IO_L1_out_1_10__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_1_10__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_1_11__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_1_11__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_1_11__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_1_11__din;
  wire fifo_C_drain_C_drain_IO_L1_out_1_11__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_1_11__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_1_12__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_1_12__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_1_12__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_1_12__din;
  wire fifo_C_drain_C_drain_IO_L1_out_1_12__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_1_12__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_1_13__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_1_13__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_1_13__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_1_13__din;
  wire fifo_C_drain_C_drain_IO_L1_out_1_13__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_1_13__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_1_14__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_1_14__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_1_14__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_1_14__din;
  wire fifo_C_drain_C_drain_IO_L1_out_1_14__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_1_14__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_1_15__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_1_15__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_1_15__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_1_15__din;
  wire fifo_C_drain_C_drain_IO_L1_out_1_15__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_1_15__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_1_16__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_1_16__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_1_16__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_1_16__din;
  wire fifo_C_drain_C_drain_IO_L1_out_1_16__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_1_16__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_1_17__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_1_17__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_1_17__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_1_17__din;
  wire fifo_C_drain_C_drain_IO_L1_out_1_17__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_1_17__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_1_2__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_1_2__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_1_2__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_1_2__din;
  wire fifo_C_drain_C_drain_IO_L1_out_1_2__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_1_2__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_1_3__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_1_3__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_1_3__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_1_3__din;
  wire fifo_C_drain_C_drain_IO_L1_out_1_3__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_1_3__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_1_4__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_1_4__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_1_4__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_1_4__din;
  wire fifo_C_drain_C_drain_IO_L1_out_1_4__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_1_4__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_1_5__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_1_5__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_1_5__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_1_5__din;
  wire fifo_C_drain_C_drain_IO_L1_out_1_5__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_1_5__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_1_6__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_1_6__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_1_6__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_1_6__din;
  wire fifo_C_drain_C_drain_IO_L1_out_1_6__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_1_6__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_1_7__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_1_7__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_1_7__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_1_7__din;
  wire fifo_C_drain_C_drain_IO_L1_out_1_7__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_1_7__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_1_8__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_1_8__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_1_8__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_1_8__din;
  wire fifo_C_drain_C_drain_IO_L1_out_1_8__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_1_8__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_1_9__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_1_9__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_1_9__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_1_9__din;
  wire fifo_C_drain_C_drain_IO_L1_out_1_9__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_1_9__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_2_0__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_2_0__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_2_0__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_2_0__din;
  wire fifo_C_drain_C_drain_IO_L1_out_2_0__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_2_0__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_2_1__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_2_1__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_2_1__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_2_1__din;
  wire fifo_C_drain_C_drain_IO_L1_out_2_1__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_2_1__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_2_10__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_2_10__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_2_10__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_2_10__din;
  wire fifo_C_drain_C_drain_IO_L1_out_2_10__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_2_10__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_2_11__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_2_11__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_2_11__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_2_11__din;
  wire fifo_C_drain_C_drain_IO_L1_out_2_11__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_2_11__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_2_12__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_2_12__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_2_12__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_2_12__din;
  wire fifo_C_drain_C_drain_IO_L1_out_2_12__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_2_12__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_2_13__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_2_13__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_2_13__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_2_13__din;
  wire fifo_C_drain_C_drain_IO_L1_out_2_13__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_2_13__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_2_14__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_2_14__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_2_14__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_2_14__din;
  wire fifo_C_drain_C_drain_IO_L1_out_2_14__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_2_14__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_2_15__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_2_15__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_2_15__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_2_15__din;
  wire fifo_C_drain_C_drain_IO_L1_out_2_15__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_2_15__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_2_16__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_2_16__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_2_16__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_2_16__din;
  wire fifo_C_drain_C_drain_IO_L1_out_2_16__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_2_16__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_2_17__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_2_17__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_2_17__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_2_17__din;
  wire fifo_C_drain_C_drain_IO_L1_out_2_17__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_2_17__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_2_2__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_2_2__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_2_2__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_2_2__din;
  wire fifo_C_drain_C_drain_IO_L1_out_2_2__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_2_2__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_2_3__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_2_3__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_2_3__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_2_3__din;
  wire fifo_C_drain_C_drain_IO_L1_out_2_3__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_2_3__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_2_4__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_2_4__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_2_4__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_2_4__din;
  wire fifo_C_drain_C_drain_IO_L1_out_2_4__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_2_4__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_2_5__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_2_5__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_2_5__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_2_5__din;
  wire fifo_C_drain_C_drain_IO_L1_out_2_5__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_2_5__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_2_6__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_2_6__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_2_6__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_2_6__din;
  wire fifo_C_drain_C_drain_IO_L1_out_2_6__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_2_6__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_2_7__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_2_7__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_2_7__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_2_7__din;
  wire fifo_C_drain_C_drain_IO_L1_out_2_7__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_2_7__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_2_8__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_2_8__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_2_8__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_2_8__din;
  wire fifo_C_drain_C_drain_IO_L1_out_2_8__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_2_8__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_2_9__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_2_9__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_2_9__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_2_9__din;
  wire fifo_C_drain_C_drain_IO_L1_out_2_9__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_2_9__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_3_0__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_3_0__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_3_0__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_3_0__din;
  wire fifo_C_drain_C_drain_IO_L1_out_3_0__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_3_0__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_3_1__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_3_1__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_3_1__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_3_1__din;
  wire fifo_C_drain_C_drain_IO_L1_out_3_1__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_3_1__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_3_10__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_3_10__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_3_10__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_3_10__din;
  wire fifo_C_drain_C_drain_IO_L1_out_3_10__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_3_10__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_3_11__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_3_11__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_3_11__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_3_11__din;
  wire fifo_C_drain_C_drain_IO_L1_out_3_11__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_3_11__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_3_12__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_3_12__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_3_12__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_3_12__din;
  wire fifo_C_drain_C_drain_IO_L1_out_3_12__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_3_12__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_3_13__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_3_13__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_3_13__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_3_13__din;
  wire fifo_C_drain_C_drain_IO_L1_out_3_13__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_3_13__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_3_14__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_3_14__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_3_14__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_3_14__din;
  wire fifo_C_drain_C_drain_IO_L1_out_3_14__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_3_14__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_3_15__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_3_15__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_3_15__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_3_15__din;
  wire fifo_C_drain_C_drain_IO_L1_out_3_15__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_3_15__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_3_16__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_3_16__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_3_16__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_3_16__din;
  wire fifo_C_drain_C_drain_IO_L1_out_3_16__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_3_16__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_3_17__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_3_17__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_3_17__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_3_17__din;
  wire fifo_C_drain_C_drain_IO_L1_out_3_17__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_3_17__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_3_2__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_3_2__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_3_2__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_3_2__din;
  wire fifo_C_drain_C_drain_IO_L1_out_3_2__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_3_2__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_3_3__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_3_3__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_3_3__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_3_3__din;
  wire fifo_C_drain_C_drain_IO_L1_out_3_3__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_3_3__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_3_4__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_3_4__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_3_4__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_3_4__din;
  wire fifo_C_drain_C_drain_IO_L1_out_3_4__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_3_4__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_3_5__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_3_5__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_3_5__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_3_5__din;
  wire fifo_C_drain_C_drain_IO_L1_out_3_5__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_3_5__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_3_6__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_3_6__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_3_6__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_3_6__din;
  wire fifo_C_drain_C_drain_IO_L1_out_3_6__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_3_6__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_3_7__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_3_7__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_3_7__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_3_7__din;
  wire fifo_C_drain_C_drain_IO_L1_out_3_7__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_3_7__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_3_8__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_3_8__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_3_8__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_3_8__din;
  wire fifo_C_drain_C_drain_IO_L1_out_3_8__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_3_8__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_3_9__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_3_9__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_3_9__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_3_9__din;
  wire fifo_C_drain_C_drain_IO_L1_out_3_9__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_3_9__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_4_0__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_4_0__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_4_0__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_4_0__din;
  wire fifo_C_drain_C_drain_IO_L1_out_4_0__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_4_0__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_4_1__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_4_1__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_4_1__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_4_1__din;
  wire fifo_C_drain_C_drain_IO_L1_out_4_1__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_4_1__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_4_10__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_4_10__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_4_10__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_4_10__din;
  wire fifo_C_drain_C_drain_IO_L1_out_4_10__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_4_10__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_4_11__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_4_11__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_4_11__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_4_11__din;
  wire fifo_C_drain_C_drain_IO_L1_out_4_11__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_4_11__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_4_12__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_4_12__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_4_12__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_4_12__din;
  wire fifo_C_drain_C_drain_IO_L1_out_4_12__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_4_12__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_4_13__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_4_13__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_4_13__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_4_13__din;
  wire fifo_C_drain_C_drain_IO_L1_out_4_13__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_4_13__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_4_14__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_4_14__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_4_14__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_4_14__din;
  wire fifo_C_drain_C_drain_IO_L1_out_4_14__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_4_14__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_4_15__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_4_15__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_4_15__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_4_15__din;
  wire fifo_C_drain_C_drain_IO_L1_out_4_15__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_4_15__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_4_16__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_4_16__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_4_16__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_4_16__din;
  wire fifo_C_drain_C_drain_IO_L1_out_4_16__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_4_16__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_4_17__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_4_17__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_4_17__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_4_17__din;
  wire fifo_C_drain_C_drain_IO_L1_out_4_17__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_4_17__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_4_2__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_4_2__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_4_2__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_4_2__din;
  wire fifo_C_drain_C_drain_IO_L1_out_4_2__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_4_2__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_4_3__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_4_3__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_4_3__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_4_3__din;
  wire fifo_C_drain_C_drain_IO_L1_out_4_3__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_4_3__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_4_4__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_4_4__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_4_4__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_4_4__din;
  wire fifo_C_drain_C_drain_IO_L1_out_4_4__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_4_4__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_4_5__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_4_5__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_4_5__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_4_5__din;
  wire fifo_C_drain_C_drain_IO_L1_out_4_5__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_4_5__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_4_6__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_4_6__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_4_6__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_4_6__din;
  wire fifo_C_drain_C_drain_IO_L1_out_4_6__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_4_6__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_4_7__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_4_7__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_4_7__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_4_7__din;
  wire fifo_C_drain_C_drain_IO_L1_out_4_7__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_4_7__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_4_8__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_4_8__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_4_8__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_4_8__din;
  wire fifo_C_drain_C_drain_IO_L1_out_4_8__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_4_8__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_4_9__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_4_9__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_4_9__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_4_9__din;
  wire fifo_C_drain_C_drain_IO_L1_out_4_9__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_4_9__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_5_0__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_5_0__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_5_0__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_5_0__din;
  wire fifo_C_drain_C_drain_IO_L1_out_5_0__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_5_0__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_5_1__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_5_1__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_5_1__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_5_1__din;
  wire fifo_C_drain_C_drain_IO_L1_out_5_1__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_5_1__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_5_10__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_5_10__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_5_10__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_5_10__din;
  wire fifo_C_drain_C_drain_IO_L1_out_5_10__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_5_10__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_5_11__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_5_11__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_5_11__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_5_11__din;
  wire fifo_C_drain_C_drain_IO_L1_out_5_11__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_5_11__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_5_12__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_5_12__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_5_12__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_5_12__din;
  wire fifo_C_drain_C_drain_IO_L1_out_5_12__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_5_12__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_5_13__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_5_13__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_5_13__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_5_13__din;
  wire fifo_C_drain_C_drain_IO_L1_out_5_13__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_5_13__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_5_14__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_5_14__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_5_14__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_5_14__din;
  wire fifo_C_drain_C_drain_IO_L1_out_5_14__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_5_14__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_5_15__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_5_15__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_5_15__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_5_15__din;
  wire fifo_C_drain_C_drain_IO_L1_out_5_15__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_5_15__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_5_16__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_5_16__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_5_16__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_5_16__din;
  wire fifo_C_drain_C_drain_IO_L1_out_5_16__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_5_16__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_5_17__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_5_17__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_5_17__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_5_17__din;
  wire fifo_C_drain_C_drain_IO_L1_out_5_17__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_5_17__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_5_2__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_5_2__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_5_2__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_5_2__din;
  wire fifo_C_drain_C_drain_IO_L1_out_5_2__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_5_2__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_5_3__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_5_3__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_5_3__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_5_3__din;
  wire fifo_C_drain_C_drain_IO_L1_out_5_3__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_5_3__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_5_4__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_5_4__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_5_4__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_5_4__din;
  wire fifo_C_drain_C_drain_IO_L1_out_5_4__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_5_4__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_5_5__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_5_5__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_5_5__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_5_5__din;
  wire fifo_C_drain_C_drain_IO_L1_out_5_5__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_5_5__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_5_6__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_5_6__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_5_6__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_5_6__din;
  wire fifo_C_drain_C_drain_IO_L1_out_5_6__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_5_6__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_5_7__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_5_7__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_5_7__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_5_7__din;
  wire fifo_C_drain_C_drain_IO_L1_out_5_7__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_5_7__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_5_8__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_5_8__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_5_8__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_5_8__din;
  wire fifo_C_drain_C_drain_IO_L1_out_5_8__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_5_8__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_5_9__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_5_9__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_5_9__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_5_9__din;
  wire fifo_C_drain_C_drain_IO_L1_out_5_9__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_5_9__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_6_0__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_6_0__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_6_0__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_6_0__din;
  wire fifo_C_drain_C_drain_IO_L1_out_6_0__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_6_0__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_6_1__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_6_1__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_6_1__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_6_1__din;
  wire fifo_C_drain_C_drain_IO_L1_out_6_1__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_6_1__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_6_10__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_6_10__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_6_10__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_6_10__din;
  wire fifo_C_drain_C_drain_IO_L1_out_6_10__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_6_10__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_6_11__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_6_11__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_6_11__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_6_11__din;
  wire fifo_C_drain_C_drain_IO_L1_out_6_11__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_6_11__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_6_12__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_6_12__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_6_12__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_6_12__din;
  wire fifo_C_drain_C_drain_IO_L1_out_6_12__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_6_12__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_6_13__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_6_13__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_6_13__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_6_13__din;
  wire fifo_C_drain_C_drain_IO_L1_out_6_13__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_6_13__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_6_14__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_6_14__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_6_14__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_6_14__din;
  wire fifo_C_drain_C_drain_IO_L1_out_6_14__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_6_14__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_6_15__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_6_15__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_6_15__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_6_15__din;
  wire fifo_C_drain_C_drain_IO_L1_out_6_15__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_6_15__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_6_16__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_6_16__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_6_16__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_6_16__din;
  wire fifo_C_drain_C_drain_IO_L1_out_6_16__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_6_16__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_6_17__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_6_17__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_6_17__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_6_17__din;
  wire fifo_C_drain_C_drain_IO_L1_out_6_17__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_6_17__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_6_2__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_6_2__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_6_2__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_6_2__din;
  wire fifo_C_drain_C_drain_IO_L1_out_6_2__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_6_2__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_6_3__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_6_3__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_6_3__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_6_3__din;
  wire fifo_C_drain_C_drain_IO_L1_out_6_3__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_6_3__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_6_4__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_6_4__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_6_4__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_6_4__din;
  wire fifo_C_drain_C_drain_IO_L1_out_6_4__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_6_4__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_6_5__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_6_5__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_6_5__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_6_5__din;
  wire fifo_C_drain_C_drain_IO_L1_out_6_5__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_6_5__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_6_6__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_6_6__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_6_6__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_6_6__din;
  wire fifo_C_drain_C_drain_IO_L1_out_6_6__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_6_6__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_6_7__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_6_7__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_6_7__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_6_7__din;
  wire fifo_C_drain_C_drain_IO_L1_out_6_7__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_6_7__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_6_8__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_6_8__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_6_8__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_6_8__din;
  wire fifo_C_drain_C_drain_IO_L1_out_6_8__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_6_8__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_6_9__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_6_9__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_6_9__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_6_9__din;
  wire fifo_C_drain_C_drain_IO_L1_out_6_9__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_6_9__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_7_0__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_7_0__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_7_0__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_7_0__din;
  wire fifo_C_drain_C_drain_IO_L1_out_7_0__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_7_0__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_7_1__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_7_1__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_7_1__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_7_1__din;
  wire fifo_C_drain_C_drain_IO_L1_out_7_1__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_7_1__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_7_10__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_7_10__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_7_10__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_7_10__din;
  wire fifo_C_drain_C_drain_IO_L1_out_7_10__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_7_10__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_7_11__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_7_11__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_7_11__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_7_11__din;
  wire fifo_C_drain_C_drain_IO_L1_out_7_11__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_7_11__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_7_12__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_7_12__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_7_12__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_7_12__din;
  wire fifo_C_drain_C_drain_IO_L1_out_7_12__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_7_12__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_7_13__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_7_13__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_7_13__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_7_13__din;
  wire fifo_C_drain_C_drain_IO_L1_out_7_13__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_7_13__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_7_14__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_7_14__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_7_14__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_7_14__din;
  wire fifo_C_drain_C_drain_IO_L1_out_7_14__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_7_14__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_7_15__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_7_15__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_7_15__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_7_15__din;
  wire fifo_C_drain_C_drain_IO_L1_out_7_15__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_7_15__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_7_16__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_7_16__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_7_16__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_7_16__din;
  wire fifo_C_drain_C_drain_IO_L1_out_7_16__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_7_16__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_7_17__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_7_17__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_7_17__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_7_17__din;
  wire fifo_C_drain_C_drain_IO_L1_out_7_17__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_7_17__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_7_2__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_7_2__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_7_2__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_7_2__din;
  wire fifo_C_drain_C_drain_IO_L1_out_7_2__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_7_2__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_7_3__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_7_3__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_7_3__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_7_3__din;
  wire fifo_C_drain_C_drain_IO_L1_out_7_3__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_7_3__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_7_4__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_7_4__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_7_4__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_7_4__din;
  wire fifo_C_drain_C_drain_IO_L1_out_7_4__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_7_4__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_7_5__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_7_5__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_7_5__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_7_5__din;
  wire fifo_C_drain_C_drain_IO_L1_out_7_5__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_7_5__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_7_6__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_7_6__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_7_6__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_7_6__din;
  wire fifo_C_drain_C_drain_IO_L1_out_7_6__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_7_6__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_7_7__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_7_7__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_7_7__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_7_7__din;
  wire fifo_C_drain_C_drain_IO_L1_out_7_7__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_7_7__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_7_8__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_7_8__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_7_8__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_7_8__din;
  wire fifo_C_drain_C_drain_IO_L1_out_7_8__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_7_8__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_7_9__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_7_9__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_7_9__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_7_9__din;
  wire fifo_C_drain_C_drain_IO_L1_out_7_9__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_7_9__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_8_0__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_8_0__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_8_0__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_8_0__din;
  wire fifo_C_drain_C_drain_IO_L1_out_8_0__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_8_0__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_8_1__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_8_1__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_8_1__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_8_1__din;
  wire fifo_C_drain_C_drain_IO_L1_out_8_1__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_8_1__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_8_10__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_8_10__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_8_10__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_8_10__din;
  wire fifo_C_drain_C_drain_IO_L1_out_8_10__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_8_10__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_8_11__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_8_11__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_8_11__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_8_11__din;
  wire fifo_C_drain_C_drain_IO_L1_out_8_11__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_8_11__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_8_12__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_8_12__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_8_12__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_8_12__din;
  wire fifo_C_drain_C_drain_IO_L1_out_8_12__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_8_12__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_8_13__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_8_13__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_8_13__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_8_13__din;
  wire fifo_C_drain_C_drain_IO_L1_out_8_13__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_8_13__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_8_14__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_8_14__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_8_14__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_8_14__din;
  wire fifo_C_drain_C_drain_IO_L1_out_8_14__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_8_14__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_8_15__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_8_15__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_8_15__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_8_15__din;
  wire fifo_C_drain_C_drain_IO_L1_out_8_15__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_8_15__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_8_16__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_8_16__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_8_16__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_8_16__din;
  wire fifo_C_drain_C_drain_IO_L1_out_8_16__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_8_16__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_8_17__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_8_17__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_8_17__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_8_17__din;
  wire fifo_C_drain_C_drain_IO_L1_out_8_17__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_8_17__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_8_2__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_8_2__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_8_2__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_8_2__din;
  wire fifo_C_drain_C_drain_IO_L1_out_8_2__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_8_2__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_8_3__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_8_3__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_8_3__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_8_3__din;
  wire fifo_C_drain_C_drain_IO_L1_out_8_3__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_8_3__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_8_4__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_8_4__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_8_4__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_8_4__din;
  wire fifo_C_drain_C_drain_IO_L1_out_8_4__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_8_4__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_8_5__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_8_5__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_8_5__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_8_5__din;
  wire fifo_C_drain_C_drain_IO_L1_out_8_5__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_8_5__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_8_6__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_8_6__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_8_6__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_8_6__din;
  wire fifo_C_drain_C_drain_IO_L1_out_8_6__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_8_6__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_8_7__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_8_7__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_8_7__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_8_7__din;
  wire fifo_C_drain_C_drain_IO_L1_out_8_7__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_8_7__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_8_8__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_8_8__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_8_8__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_8_8__din;
  wire fifo_C_drain_C_drain_IO_L1_out_8_8__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_8_8__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_8_9__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_8_9__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_8_9__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_8_9__din;
  wire fifo_C_drain_C_drain_IO_L1_out_8_9__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_8_9__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_9_0__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_9_0__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_9_0__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_9_0__din;
  wire fifo_C_drain_C_drain_IO_L1_out_9_0__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_9_0__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_9_1__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_9_1__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_9_1__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_9_1__din;
  wire fifo_C_drain_C_drain_IO_L1_out_9_1__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_9_1__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_9_10__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_9_10__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_9_10__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_9_10__din;
  wire fifo_C_drain_C_drain_IO_L1_out_9_10__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_9_10__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_9_11__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_9_11__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_9_11__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_9_11__din;
  wire fifo_C_drain_C_drain_IO_L1_out_9_11__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_9_11__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_9_12__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_9_12__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_9_12__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_9_12__din;
  wire fifo_C_drain_C_drain_IO_L1_out_9_12__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_9_12__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_9_13__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_9_13__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_9_13__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_9_13__din;
  wire fifo_C_drain_C_drain_IO_L1_out_9_13__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_9_13__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_9_14__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_9_14__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_9_14__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_9_14__din;
  wire fifo_C_drain_C_drain_IO_L1_out_9_14__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_9_14__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_9_15__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_9_15__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_9_15__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_9_15__din;
  wire fifo_C_drain_C_drain_IO_L1_out_9_15__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_9_15__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_9_16__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_9_16__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_9_16__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_9_16__din;
  wire fifo_C_drain_C_drain_IO_L1_out_9_16__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_9_16__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_9_17__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_9_17__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_9_17__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_9_17__din;
  wire fifo_C_drain_C_drain_IO_L1_out_9_17__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_9_17__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_9_2__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_9_2__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_9_2__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_9_2__din;
  wire fifo_C_drain_C_drain_IO_L1_out_9_2__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_9_2__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_9_3__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_9_3__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_9_3__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_9_3__din;
  wire fifo_C_drain_C_drain_IO_L1_out_9_3__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_9_3__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_9_4__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_9_4__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_9_4__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_9_4__din;
  wire fifo_C_drain_C_drain_IO_L1_out_9_4__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_9_4__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_9_5__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_9_5__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_9_5__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_9_5__din;
  wire fifo_C_drain_C_drain_IO_L1_out_9_5__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_9_5__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_9_6__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_9_6__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_9_6__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_9_6__din;
  wire fifo_C_drain_C_drain_IO_L1_out_9_6__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_9_6__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_9_7__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_9_7__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_9_7__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_9_7__din;
  wire fifo_C_drain_C_drain_IO_L1_out_9_7__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_9_7__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_9_8__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_9_8__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_9_8__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_9_8__din;
  wire fifo_C_drain_C_drain_IO_L1_out_9_8__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_9_8__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_9_9__dout;
  wire fifo_C_drain_C_drain_IO_L1_out_9_9__empty_n;
  wire fifo_C_drain_C_drain_IO_L1_out_9_9__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L1_out_9_9__din;
  wire fifo_C_drain_C_drain_IO_L1_out_9_9__full_n;
  wire fifo_C_drain_C_drain_IO_L1_out_9_9__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L2_out_0__dout;
  wire fifo_C_drain_C_drain_IO_L2_out_0__empty_n;
  wire fifo_C_drain_C_drain_IO_L2_out_0__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L2_out_0__din;
  wire fifo_C_drain_C_drain_IO_L2_out_0__full_n;
  wire fifo_C_drain_C_drain_IO_L2_out_0__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L2_out_1__dout;
  wire fifo_C_drain_C_drain_IO_L2_out_1__empty_n;
  wire fifo_C_drain_C_drain_IO_L2_out_1__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L2_out_1__din;
  wire fifo_C_drain_C_drain_IO_L2_out_1__full_n;
  wire fifo_C_drain_C_drain_IO_L2_out_1__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L2_out_10__dout;
  wire fifo_C_drain_C_drain_IO_L2_out_10__empty_n;
  wire fifo_C_drain_C_drain_IO_L2_out_10__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L2_out_10__din;
  wire fifo_C_drain_C_drain_IO_L2_out_10__full_n;
  wire fifo_C_drain_C_drain_IO_L2_out_10__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L2_out_11__dout;
  wire fifo_C_drain_C_drain_IO_L2_out_11__empty_n;
  wire fifo_C_drain_C_drain_IO_L2_out_11__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L2_out_11__din;
  wire fifo_C_drain_C_drain_IO_L2_out_11__full_n;
  wire fifo_C_drain_C_drain_IO_L2_out_11__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L2_out_12__dout;
  wire fifo_C_drain_C_drain_IO_L2_out_12__empty_n;
  wire fifo_C_drain_C_drain_IO_L2_out_12__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L2_out_12__din;
  wire fifo_C_drain_C_drain_IO_L2_out_12__full_n;
  wire fifo_C_drain_C_drain_IO_L2_out_12__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L2_out_13__dout;
  wire fifo_C_drain_C_drain_IO_L2_out_13__empty_n;
  wire fifo_C_drain_C_drain_IO_L2_out_13__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L2_out_13__din;
  wire fifo_C_drain_C_drain_IO_L2_out_13__full_n;
  wire fifo_C_drain_C_drain_IO_L2_out_13__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L2_out_14__dout;
  wire fifo_C_drain_C_drain_IO_L2_out_14__empty_n;
  wire fifo_C_drain_C_drain_IO_L2_out_14__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L2_out_14__din;
  wire fifo_C_drain_C_drain_IO_L2_out_14__full_n;
  wire fifo_C_drain_C_drain_IO_L2_out_14__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L2_out_15__dout;
  wire fifo_C_drain_C_drain_IO_L2_out_15__empty_n;
  wire fifo_C_drain_C_drain_IO_L2_out_15__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L2_out_15__din;
  wire fifo_C_drain_C_drain_IO_L2_out_15__full_n;
  wire fifo_C_drain_C_drain_IO_L2_out_15__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L2_out_16__dout;
  wire fifo_C_drain_C_drain_IO_L2_out_16__empty_n;
  wire fifo_C_drain_C_drain_IO_L2_out_16__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L2_out_16__din;
  wire fifo_C_drain_C_drain_IO_L2_out_16__full_n;
  wire fifo_C_drain_C_drain_IO_L2_out_16__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L2_out_2__dout;
  wire fifo_C_drain_C_drain_IO_L2_out_2__empty_n;
  wire fifo_C_drain_C_drain_IO_L2_out_2__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L2_out_2__din;
  wire fifo_C_drain_C_drain_IO_L2_out_2__full_n;
  wire fifo_C_drain_C_drain_IO_L2_out_2__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L2_out_3__dout;
  wire fifo_C_drain_C_drain_IO_L2_out_3__empty_n;
  wire fifo_C_drain_C_drain_IO_L2_out_3__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L2_out_3__din;
  wire fifo_C_drain_C_drain_IO_L2_out_3__full_n;
  wire fifo_C_drain_C_drain_IO_L2_out_3__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L2_out_4__dout;
  wire fifo_C_drain_C_drain_IO_L2_out_4__empty_n;
  wire fifo_C_drain_C_drain_IO_L2_out_4__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L2_out_4__din;
  wire fifo_C_drain_C_drain_IO_L2_out_4__full_n;
  wire fifo_C_drain_C_drain_IO_L2_out_4__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L2_out_5__dout;
  wire fifo_C_drain_C_drain_IO_L2_out_5__empty_n;
  wire fifo_C_drain_C_drain_IO_L2_out_5__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L2_out_5__din;
  wire fifo_C_drain_C_drain_IO_L2_out_5__full_n;
  wire fifo_C_drain_C_drain_IO_L2_out_5__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L2_out_6__dout;
  wire fifo_C_drain_C_drain_IO_L2_out_6__empty_n;
  wire fifo_C_drain_C_drain_IO_L2_out_6__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L2_out_6__din;
  wire fifo_C_drain_C_drain_IO_L2_out_6__full_n;
  wire fifo_C_drain_C_drain_IO_L2_out_6__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L2_out_7__dout;
  wire fifo_C_drain_C_drain_IO_L2_out_7__empty_n;
  wire fifo_C_drain_C_drain_IO_L2_out_7__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L2_out_7__din;
  wire fifo_C_drain_C_drain_IO_L2_out_7__full_n;
  wire fifo_C_drain_C_drain_IO_L2_out_7__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L2_out_8__dout;
  wire fifo_C_drain_C_drain_IO_L2_out_8__empty_n;
  wire fifo_C_drain_C_drain_IO_L2_out_8__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L2_out_8__din;
  wire fifo_C_drain_C_drain_IO_L2_out_8__full_n;
  wire fifo_C_drain_C_drain_IO_L2_out_8__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L2_out_9__dout;
  wire fifo_C_drain_C_drain_IO_L2_out_9__empty_n;
  wire fifo_C_drain_C_drain_IO_L2_out_9__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L2_out_9__din;
  wire fifo_C_drain_C_drain_IO_L2_out_9__full_n;
  wire fifo_C_drain_C_drain_IO_L2_out_9__write;
  wire [128:0] fifo_C_drain_C_drain_IO_L3_out_serialize__dout;
  wire fifo_C_drain_C_drain_IO_L3_out_serialize__empty_n;
  wire fifo_C_drain_C_drain_IO_L3_out_serialize__read;
  wire [128:0] fifo_C_drain_C_drain_IO_L3_out_serialize__din;
  wire fifo_C_drain_C_drain_IO_L3_out_serialize__full_n;
  wire fifo_C_drain_C_drain_IO_L3_out_serialize__write;
  wire [16:0] fifo_C_drain_PE_0_0__dout;
  wire fifo_C_drain_PE_0_0__empty_n;
  wire fifo_C_drain_PE_0_0__read;
  wire [16:0] fifo_C_drain_PE_0_0__din;
  wire fifo_C_drain_PE_0_0__full_n;
  wire fifo_C_drain_PE_0_0__write;
  wire [16:0] fifo_C_drain_PE_0_1__dout;
  wire fifo_C_drain_PE_0_1__empty_n;
  wire fifo_C_drain_PE_0_1__read;
  wire [16:0] fifo_C_drain_PE_0_1__din;
  wire fifo_C_drain_PE_0_1__full_n;
  wire fifo_C_drain_PE_0_1__write;
  wire [16:0] fifo_C_drain_PE_0_10__dout;
  wire fifo_C_drain_PE_0_10__empty_n;
  wire fifo_C_drain_PE_0_10__read;
  wire [16:0] fifo_C_drain_PE_0_10__din;
  wire fifo_C_drain_PE_0_10__full_n;
  wire fifo_C_drain_PE_0_10__write;
  wire [16:0] fifo_C_drain_PE_0_11__dout;
  wire fifo_C_drain_PE_0_11__empty_n;
  wire fifo_C_drain_PE_0_11__read;
  wire [16:0] fifo_C_drain_PE_0_11__din;
  wire fifo_C_drain_PE_0_11__full_n;
  wire fifo_C_drain_PE_0_11__write;
  wire [16:0] fifo_C_drain_PE_0_12__dout;
  wire fifo_C_drain_PE_0_12__empty_n;
  wire fifo_C_drain_PE_0_12__read;
  wire [16:0] fifo_C_drain_PE_0_12__din;
  wire fifo_C_drain_PE_0_12__full_n;
  wire fifo_C_drain_PE_0_12__write;
  wire [16:0] fifo_C_drain_PE_0_13__dout;
  wire fifo_C_drain_PE_0_13__empty_n;
  wire fifo_C_drain_PE_0_13__read;
  wire [16:0] fifo_C_drain_PE_0_13__din;
  wire fifo_C_drain_PE_0_13__full_n;
  wire fifo_C_drain_PE_0_13__write;
  wire [16:0] fifo_C_drain_PE_0_14__dout;
  wire fifo_C_drain_PE_0_14__empty_n;
  wire fifo_C_drain_PE_0_14__read;
  wire [16:0] fifo_C_drain_PE_0_14__din;
  wire fifo_C_drain_PE_0_14__full_n;
  wire fifo_C_drain_PE_0_14__write;
  wire [16:0] fifo_C_drain_PE_0_15__dout;
  wire fifo_C_drain_PE_0_15__empty_n;
  wire fifo_C_drain_PE_0_15__read;
  wire [16:0] fifo_C_drain_PE_0_15__din;
  wire fifo_C_drain_PE_0_15__full_n;
  wire fifo_C_drain_PE_0_15__write;
  wire [16:0] fifo_C_drain_PE_0_16__dout;
  wire fifo_C_drain_PE_0_16__empty_n;
  wire fifo_C_drain_PE_0_16__read;
  wire [16:0] fifo_C_drain_PE_0_16__din;
  wire fifo_C_drain_PE_0_16__full_n;
  wire fifo_C_drain_PE_0_16__write;
  wire [16:0] fifo_C_drain_PE_0_2__dout;
  wire fifo_C_drain_PE_0_2__empty_n;
  wire fifo_C_drain_PE_0_2__read;
  wire [16:0] fifo_C_drain_PE_0_2__din;
  wire fifo_C_drain_PE_0_2__full_n;
  wire fifo_C_drain_PE_0_2__write;
  wire [16:0] fifo_C_drain_PE_0_3__dout;
  wire fifo_C_drain_PE_0_3__empty_n;
  wire fifo_C_drain_PE_0_3__read;
  wire [16:0] fifo_C_drain_PE_0_3__din;
  wire fifo_C_drain_PE_0_3__full_n;
  wire fifo_C_drain_PE_0_3__write;
  wire [16:0] fifo_C_drain_PE_0_4__dout;
  wire fifo_C_drain_PE_0_4__empty_n;
  wire fifo_C_drain_PE_0_4__read;
  wire [16:0] fifo_C_drain_PE_0_4__din;
  wire fifo_C_drain_PE_0_4__full_n;
  wire fifo_C_drain_PE_0_4__write;
  wire [16:0] fifo_C_drain_PE_0_5__dout;
  wire fifo_C_drain_PE_0_5__empty_n;
  wire fifo_C_drain_PE_0_5__read;
  wire [16:0] fifo_C_drain_PE_0_5__din;
  wire fifo_C_drain_PE_0_5__full_n;
  wire fifo_C_drain_PE_0_5__write;
  wire [16:0] fifo_C_drain_PE_0_6__dout;
  wire fifo_C_drain_PE_0_6__empty_n;
  wire fifo_C_drain_PE_0_6__read;
  wire [16:0] fifo_C_drain_PE_0_6__din;
  wire fifo_C_drain_PE_0_6__full_n;
  wire fifo_C_drain_PE_0_6__write;
  wire [16:0] fifo_C_drain_PE_0_7__dout;
  wire fifo_C_drain_PE_0_7__empty_n;
  wire fifo_C_drain_PE_0_7__read;
  wire [16:0] fifo_C_drain_PE_0_7__din;
  wire fifo_C_drain_PE_0_7__full_n;
  wire fifo_C_drain_PE_0_7__write;
  wire [16:0] fifo_C_drain_PE_0_8__dout;
  wire fifo_C_drain_PE_0_8__empty_n;
  wire fifo_C_drain_PE_0_8__read;
  wire [16:0] fifo_C_drain_PE_0_8__din;
  wire fifo_C_drain_PE_0_8__full_n;
  wire fifo_C_drain_PE_0_8__write;
  wire [16:0] fifo_C_drain_PE_0_9__dout;
  wire fifo_C_drain_PE_0_9__empty_n;
  wire fifo_C_drain_PE_0_9__read;
  wire [16:0] fifo_C_drain_PE_0_9__din;
  wire fifo_C_drain_PE_0_9__full_n;
  wire fifo_C_drain_PE_0_9__write;
  wire [16:0] fifo_C_drain_PE_10_0__dout;
  wire fifo_C_drain_PE_10_0__empty_n;
  wire fifo_C_drain_PE_10_0__read;
  wire [16:0] fifo_C_drain_PE_10_0__din;
  wire fifo_C_drain_PE_10_0__full_n;
  wire fifo_C_drain_PE_10_0__write;
  wire [16:0] fifo_C_drain_PE_10_1__dout;
  wire fifo_C_drain_PE_10_1__empty_n;
  wire fifo_C_drain_PE_10_1__read;
  wire [16:0] fifo_C_drain_PE_10_1__din;
  wire fifo_C_drain_PE_10_1__full_n;
  wire fifo_C_drain_PE_10_1__write;
  wire [16:0] fifo_C_drain_PE_10_10__dout;
  wire fifo_C_drain_PE_10_10__empty_n;
  wire fifo_C_drain_PE_10_10__read;
  wire [16:0] fifo_C_drain_PE_10_10__din;
  wire fifo_C_drain_PE_10_10__full_n;
  wire fifo_C_drain_PE_10_10__write;
  wire [16:0] fifo_C_drain_PE_10_11__dout;
  wire fifo_C_drain_PE_10_11__empty_n;
  wire fifo_C_drain_PE_10_11__read;
  wire [16:0] fifo_C_drain_PE_10_11__din;
  wire fifo_C_drain_PE_10_11__full_n;
  wire fifo_C_drain_PE_10_11__write;
  wire [16:0] fifo_C_drain_PE_10_12__dout;
  wire fifo_C_drain_PE_10_12__empty_n;
  wire fifo_C_drain_PE_10_12__read;
  wire [16:0] fifo_C_drain_PE_10_12__din;
  wire fifo_C_drain_PE_10_12__full_n;
  wire fifo_C_drain_PE_10_12__write;
  wire [16:0] fifo_C_drain_PE_10_13__dout;
  wire fifo_C_drain_PE_10_13__empty_n;
  wire fifo_C_drain_PE_10_13__read;
  wire [16:0] fifo_C_drain_PE_10_13__din;
  wire fifo_C_drain_PE_10_13__full_n;
  wire fifo_C_drain_PE_10_13__write;
  wire [16:0] fifo_C_drain_PE_10_14__dout;
  wire fifo_C_drain_PE_10_14__empty_n;
  wire fifo_C_drain_PE_10_14__read;
  wire [16:0] fifo_C_drain_PE_10_14__din;
  wire fifo_C_drain_PE_10_14__full_n;
  wire fifo_C_drain_PE_10_14__write;
  wire [16:0] fifo_C_drain_PE_10_15__dout;
  wire fifo_C_drain_PE_10_15__empty_n;
  wire fifo_C_drain_PE_10_15__read;
  wire [16:0] fifo_C_drain_PE_10_15__din;
  wire fifo_C_drain_PE_10_15__full_n;
  wire fifo_C_drain_PE_10_15__write;
  wire [16:0] fifo_C_drain_PE_10_16__dout;
  wire fifo_C_drain_PE_10_16__empty_n;
  wire fifo_C_drain_PE_10_16__read;
  wire [16:0] fifo_C_drain_PE_10_16__din;
  wire fifo_C_drain_PE_10_16__full_n;
  wire fifo_C_drain_PE_10_16__write;
  wire [16:0] fifo_C_drain_PE_10_2__dout;
  wire fifo_C_drain_PE_10_2__empty_n;
  wire fifo_C_drain_PE_10_2__read;
  wire [16:0] fifo_C_drain_PE_10_2__din;
  wire fifo_C_drain_PE_10_2__full_n;
  wire fifo_C_drain_PE_10_2__write;
  wire [16:0] fifo_C_drain_PE_10_3__dout;
  wire fifo_C_drain_PE_10_3__empty_n;
  wire fifo_C_drain_PE_10_3__read;
  wire [16:0] fifo_C_drain_PE_10_3__din;
  wire fifo_C_drain_PE_10_3__full_n;
  wire fifo_C_drain_PE_10_3__write;
  wire [16:0] fifo_C_drain_PE_10_4__dout;
  wire fifo_C_drain_PE_10_4__empty_n;
  wire fifo_C_drain_PE_10_4__read;
  wire [16:0] fifo_C_drain_PE_10_4__din;
  wire fifo_C_drain_PE_10_4__full_n;
  wire fifo_C_drain_PE_10_4__write;
  wire [16:0] fifo_C_drain_PE_10_5__dout;
  wire fifo_C_drain_PE_10_5__empty_n;
  wire fifo_C_drain_PE_10_5__read;
  wire [16:0] fifo_C_drain_PE_10_5__din;
  wire fifo_C_drain_PE_10_5__full_n;
  wire fifo_C_drain_PE_10_5__write;
  wire [16:0] fifo_C_drain_PE_10_6__dout;
  wire fifo_C_drain_PE_10_6__empty_n;
  wire fifo_C_drain_PE_10_6__read;
  wire [16:0] fifo_C_drain_PE_10_6__din;
  wire fifo_C_drain_PE_10_6__full_n;
  wire fifo_C_drain_PE_10_6__write;
  wire [16:0] fifo_C_drain_PE_10_7__dout;
  wire fifo_C_drain_PE_10_7__empty_n;
  wire fifo_C_drain_PE_10_7__read;
  wire [16:0] fifo_C_drain_PE_10_7__din;
  wire fifo_C_drain_PE_10_7__full_n;
  wire fifo_C_drain_PE_10_7__write;
  wire [16:0] fifo_C_drain_PE_10_8__dout;
  wire fifo_C_drain_PE_10_8__empty_n;
  wire fifo_C_drain_PE_10_8__read;
  wire [16:0] fifo_C_drain_PE_10_8__din;
  wire fifo_C_drain_PE_10_8__full_n;
  wire fifo_C_drain_PE_10_8__write;
  wire [16:0] fifo_C_drain_PE_10_9__dout;
  wire fifo_C_drain_PE_10_9__empty_n;
  wire fifo_C_drain_PE_10_9__read;
  wire [16:0] fifo_C_drain_PE_10_9__din;
  wire fifo_C_drain_PE_10_9__full_n;
  wire fifo_C_drain_PE_10_9__write;
  wire [16:0] fifo_C_drain_PE_11_0__dout;
  wire fifo_C_drain_PE_11_0__empty_n;
  wire fifo_C_drain_PE_11_0__read;
  wire [16:0] fifo_C_drain_PE_11_0__din;
  wire fifo_C_drain_PE_11_0__full_n;
  wire fifo_C_drain_PE_11_0__write;
  wire [16:0] fifo_C_drain_PE_11_1__dout;
  wire fifo_C_drain_PE_11_1__empty_n;
  wire fifo_C_drain_PE_11_1__read;
  wire [16:0] fifo_C_drain_PE_11_1__din;
  wire fifo_C_drain_PE_11_1__full_n;
  wire fifo_C_drain_PE_11_1__write;
  wire [16:0] fifo_C_drain_PE_11_10__dout;
  wire fifo_C_drain_PE_11_10__empty_n;
  wire fifo_C_drain_PE_11_10__read;
  wire [16:0] fifo_C_drain_PE_11_10__din;
  wire fifo_C_drain_PE_11_10__full_n;
  wire fifo_C_drain_PE_11_10__write;
  wire [16:0] fifo_C_drain_PE_11_11__dout;
  wire fifo_C_drain_PE_11_11__empty_n;
  wire fifo_C_drain_PE_11_11__read;
  wire [16:0] fifo_C_drain_PE_11_11__din;
  wire fifo_C_drain_PE_11_11__full_n;
  wire fifo_C_drain_PE_11_11__write;
  wire [16:0] fifo_C_drain_PE_11_12__dout;
  wire fifo_C_drain_PE_11_12__empty_n;
  wire fifo_C_drain_PE_11_12__read;
  wire [16:0] fifo_C_drain_PE_11_12__din;
  wire fifo_C_drain_PE_11_12__full_n;
  wire fifo_C_drain_PE_11_12__write;
  wire [16:0] fifo_C_drain_PE_11_13__dout;
  wire fifo_C_drain_PE_11_13__empty_n;
  wire fifo_C_drain_PE_11_13__read;
  wire [16:0] fifo_C_drain_PE_11_13__din;
  wire fifo_C_drain_PE_11_13__full_n;
  wire fifo_C_drain_PE_11_13__write;
  wire [16:0] fifo_C_drain_PE_11_14__dout;
  wire fifo_C_drain_PE_11_14__empty_n;
  wire fifo_C_drain_PE_11_14__read;
  wire [16:0] fifo_C_drain_PE_11_14__din;
  wire fifo_C_drain_PE_11_14__full_n;
  wire fifo_C_drain_PE_11_14__write;
  wire [16:0] fifo_C_drain_PE_11_15__dout;
  wire fifo_C_drain_PE_11_15__empty_n;
  wire fifo_C_drain_PE_11_15__read;
  wire [16:0] fifo_C_drain_PE_11_15__din;
  wire fifo_C_drain_PE_11_15__full_n;
  wire fifo_C_drain_PE_11_15__write;
  wire [16:0] fifo_C_drain_PE_11_16__dout;
  wire fifo_C_drain_PE_11_16__empty_n;
  wire fifo_C_drain_PE_11_16__read;
  wire [16:0] fifo_C_drain_PE_11_16__din;
  wire fifo_C_drain_PE_11_16__full_n;
  wire fifo_C_drain_PE_11_16__write;
  wire [16:0] fifo_C_drain_PE_11_2__dout;
  wire fifo_C_drain_PE_11_2__empty_n;
  wire fifo_C_drain_PE_11_2__read;
  wire [16:0] fifo_C_drain_PE_11_2__din;
  wire fifo_C_drain_PE_11_2__full_n;
  wire fifo_C_drain_PE_11_2__write;
  wire [16:0] fifo_C_drain_PE_11_3__dout;
  wire fifo_C_drain_PE_11_3__empty_n;
  wire fifo_C_drain_PE_11_3__read;
  wire [16:0] fifo_C_drain_PE_11_3__din;
  wire fifo_C_drain_PE_11_3__full_n;
  wire fifo_C_drain_PE_11_3__write;
  wire [16:0] fifo_C_drain_PE_11_4__dout;
  wire fifo_C_drain_PE_11_4__empty_n;
  wire fifo_C_drain_PE_11_4__read;
  wire [16:0] fifo_C_drain_PE_11_4__din;
  wire fifo_C_drain_PE_11_4__full_n;
  wire fifo_C_drain_PE_11_4__write;
  wire [16:0] fifo_C_drain_PE_11_5__dout;
  wire fifo_C_drain_PE_11_5__empty_n;
  wire fifo_C_drain_PE_11_5__read;
  wire [16:0] fifo_C_drain_PE_11_5__din;
  wire fifo_C_drain_PE_11_5__full_n;
  wire fifo_C_drain_PE_11_5__write;
  wire [16:0] fifo_C_drain_PE_11_6__dout;
  wire fifo_C_drain_PE_11_6__empty_n;
  wire fifo_C_drain_PE_11_6__read;
  wire [16:0] fifo_C_drain_PE_11_6__din;
  wire fifo_C_drain_PE_11_6__full_n;
  wire fifo_C_drain_PE_11_6__write;
  wire [16:0] fifo_C_drain_PE_11_7__dout;
  wire fifo_C_drain_PE_11_7__empty_n;
  wire fifo_C_drain_PE_11_7__read;
  wire [16:0] fifo_C_drain_PE_11_7__din;
  wire fifo_C_drain_PE_11_7__full_n;
  wire fifo_C_drain_PE_11_7__write;
  wire [16:0] fifo_C_drain_PE_11_8__dout;
  wire fifo_C_drain_PE_11_8__empty_n;
  wire fifo_C_drain_PE_11_8__read;
  wire [16:0] fifo_C_drain_PE_11_8__din;
  wire fifo_C_drain_PE_11_8__full_n;
  wire fifo_C_drain_PE_11_8__write;
  wire [16:0] fifo_C_drain_PE_11_9__dout;
  wire fifo_C_drain_PE_11_9__empty_n;
  wire fifo_C_drain_PE_11_9__read;
  wire [16:0] fifo_C_drain_PE_11_9__din;
  wire fifo_C_drain_PE_11_9__full_n;
  wire fifo_C_drain_PE_11_9__write;
  wire [16:0] fifo_C_drain_PE_12_0__dout;
  wire fifo_C_drain_PE_12_0__empty_n;
  wire fifo_C_drain_PE_12_0__read;
  wire [16:0] fifo_C_drain_PE_12_0__din;
  wire fifo_C_drain_PE_12_0__full_n;
  wire fifo_C_drain_PE_12_0__write;
  wire [16:0] fifo_C_drain_PE_12_1__dout;
  wire fifo_C_drain_PE_12_1__empty_n;
  wire fifo_C_drain_PE_12_1__read;
  wire [16:0] fifo_C_drain_PE_12_1__din;
  wire fifo_C_drain_PE_12_1__full_n;
  wire fifo_C_drain_PE_12_1__write;
  wire [16:0] fifo_C_drain_PE_12_10__dout;
  wire fifo_C_drain_PE_12_10__empty_n;
  wire fifo_C_drain_PE_12_10__read;
  wire [16:0] fifo_C_drain_PE_12_10__din;
  wire fifo_C_drain_PE_12_10__full_n;
  wire fifo_C_drain_PE_12_10__write;
  wire [16:0] fifo_C_drain_PE_12_11__dout;
  wire fifo_C_drain_PE_12_11__empty_n;
  wire fifo_C_drain_PE_12_11__read;
  wire [16:0] fifo_C_drain_PE_12_11__din;
  wire fifo_C_drain_PE_12_11__full_n;
  wire fifo_C_drain_PE_12_11__write;
  wire [16:0] fifo_C_drain_PE_12_12__dout;
  wire fifo_C_drain_PE_12_12__empty_n;
  wire fifo_C_drain_PE_12_12__read;
  wire [16:0] fifo_C_drain_PE_12_12__din;
  wire fifo_C_drain_PE_12_12__full_n;
  wire fifo_C_drain_PE_12_12__write;
  wire [16:0] fifo_C_drain_PE_12_13__dout;
  wire fifo_C_drain_PE_12_13__empty_n;
  wire fifo_C_drain_PE_12_13__read;
  wire [16:0] fifo_C_drain_PE_12_13__din;
  wire fifo_C_drain_PE_12_13__full_n;
  wire fifo_C_drain_PE_12_13__write;
  wire [16:0] fifo_C_drain_PE_12_14__dout;
  wire fifo_C_drain_PE_12_14__empty_n;
  wire fifo_C_drain_PE_12_14__read;
  wire [16:0] fifo_C_drain_PE_12_14__din;
  wire fifo_C_drain_PE_12_14__full_n;
  wire fifo_C_drain_PE_12_14__write;
  wire [16:0] fifo_C_drain_PE_12_15__dout;
  wire fifo_C_drain_PE_12_15__empty_n;
  wire fifo_C_drain_PE_12_15__read;
  wire [16:0] fifo_C_drain_PE_12_15__din;
  wire fifo_C_drain_PE_12_15__full_n;
  wire fifo_C_drain_PE_12_15__write;
  wire [16:0] fifo_C_drain_PE_12_16__dout;
  wire fifo_C_drain_PE_12_16__empty_n;
  wire fifo_C_drain_PE_12_16__read;
  wire [16:0] fifo_C_drain_PE_12_16__din;
  wire fifo_C_drain_PE_12_16__full_n;
  wire fifo_C_drain_PE_12_16__write;
  wire [16:0] fifo_C_drain_PE_12_2__dout;
  wire fifo_C_drain_PE_12_2__empty_n;
  wire fifo_C_drain_PE_12_2__read;
  wire [16:0] fifo_C_drain_PE_12_2__din;
  wire fifo_C_drain_PE_12_2__full_n;
  wire fifo_C_drain_PE_12_2__write;
  wire [16:0] fifo_C_drain_PE_12_3__dout;
  wire fifo_C_drain_PE_12_3__empty_n;
  wire fifo_C_drain_PE_12_3__read;
  wire [16:0] fifo_C_drain_PE_12_3__din;
  wire fifo_C_drain_PE_12_3__full_n;
  wire fifo_C_drain_PE_12_3__write;
  wire [16:0] fifo_C_drain_PE_12_4__dout;
  wire fifo_C_drain_PE_12_4__empty_n;
  wire fifo_C_drain_PE_12_4__read;
  wire [16:0] fifo_C_drain_PE_12_4__din;
  wire fifo_C_drain_PE_12_4__full_n;
  wire fifo_C_drain_PE_12_4__write;
  wire [16:0] fifo_C_drain_PE_12_5__dout;
  wire fifo_C_drain_PE_12_5__empty_n;
  wire fifo_C_drain_PE_12_5__read;
  wire [16:0] fifo_C_drain_PE_12_5__din;
  wire fifo_C_drain_PE_12_5__full_n;
  wire fifo_C_drain_PE_12_5__write;
  wire [16:0] fifo_C_drain_PE_12_6__dout;
  wire fifo_C_drain_PE_12_6__empty_n;
  wire fifo_C_drain_PE_12_6__read;
  wire [16:0] fifo_C_drain_PE_12_6__din;
  wire fifo_C_drain_PE_12_6__full_n;
  wire fifo_C_drain_PE_12_6__write;
  wire [16:0] fifo_C_drain_PE_12_7__dout;
  wire fifo_C_drain_PE_12_7__empty_n;
  wire fifo_C_drain_PE_12_7__read;
  wire [16:0] fifo_C_drain_PE_12_7__din;
  wire fifo_C_drain_PE_12_7__full_n;
  wire fifo_C_drain_PE_12_7__write;
  wire [16:0] fifo_C_drain_PE_12_8__dout;
  wire fifo_C_drain_PE_12_8__empty_n;
  wire fifo_C_drain_PE_12_8__read;
  wire [16:0] fifo_C_drain_PE_12_8__din;
  wire fifo_C_drain_PE_12_8__full_n;
  wire fifo_C_drain_PE_12_8__write;
  wire [16:0] fifo_C_drain_PE_12_9__dout;
  wire fifo_C_drain_PE_12_9__empty_n;
  wire fifo_C_drain_PE_12_9__read;
  wire [16:0] fifo_C_drain_PE_12_9__din;
  wire fifo_C_drain_PE_12_9__full_n;
  wire fifo_C_drain_PE_12_9__write;
  wire [16:0] fifo_C_drain_PE_13_0__dout;
  wire fifo_C_drain_PE_13_0__empty_n;
  wire fifo_C_drain_PE_13_0__read;
  wire [16:0] fifo_C_drain_PE_13_0__din;
  wire fifo_C_drain_PE_13_0__full_n;
  wire fifo_C_drain_PE_13_0__write;
  wire [16:0] fifo_C_drain_PE_13_1__dout;
  wire fifo_C_drain_PE_13_1__empty_n;
  wire fifo_C_drain_PE_13_1__read;
  wire [16:0] fifo_C_drain_PE_13_1__din;
  wire fifo_C_drain_PE_13_1__full_n;
  wire fifo_C_drain_PE_13_1__write;
  wire [16:0] fifo_C_drain_PE_13_10__dout;
  wire fifo_C_drain_PE_13_10__empty_n;
  wire fifo_C_drain_PE_13_10__read;
  wire [16:0] fifo_C_drain_PE_13_10__din;
  wire fifo_C_drain_PE_13_10__full_n;
  wire fifo_C_drain_PE_13_10__write;
  wire [16:0] fifo_C_drain_PE_13_11__dout;
  wire fifo_C_drain_PE_13_11__empty_n;
  wire fifo_C_drain_PE_13_11__read;
  wire [16:0] fifo_C_drain_PE_13_11__din;
  wire fifo_C_drain_PE_13_11__full_n;
  wire fifo_C_drain_PE_13_11__write;
  wire [16:0] fifo_C_drain_PE_13_12__dout;
  wire fifo_C_drain_PE_13_12__empty_n;
  wire fifo_C_drain_PE_13_12__read;
  wire [16:0] fifo_C_drain_PE_13_12__din;
  wire fifo_C_drain_PE_13_12__full_n;
  wire fifo_C_drain_PE_13_12__write;
  wire [16:0] fifo_C_drain_PE_13_13__dout;
  wire fifo_C_drain_PE_13_13__empty_n;
  wire fifo_C_drain_PE_13_13__read;
  wire [16:0] fifo_C_drain_PE_13_13__din;
  wire fifo_C_drain_PE_13_13__full_n;
  wire fifo_C_drain_PE_13_13__write;
  wire [16:0] fifo_C_drain_PE_13_14__dout;
  wire fifo_C_drain_PE_13_14__empty_n;
  wire fifo_C_drain_PE_13_14__read;
  wire [16:0] fifo_C_drain_PE_13_14__din;
  wire fifo_C_drain_PE_13_14__full_n;
  wire fifo_C_drain_PE_13_14__write;
  wire [16:0] fifo_C_drain_PE_13_15__dout;
  wire fifo_C_drain_PE_13_15__empty_n;
  wire fifo_C_drain_PE_13_15__read;
  wire [16:0] fifo_C_drain_PE_13_15__din;
  wire fifo_C_drain_PE_13_15__full_n;
  wire fifo_C_drain_PE_13_15__write;
  wire [16:0] fifo_C_drain_PE_13_16__dout;
  wire fifo_C_drain_PE_13_16__empty_n;
  wire fifo_C_drain_PE_13_16__read;
  wire [16:0] fifo_C_drain_PE_13_16__din;
  wire fifo_C_drain_PE_13_16__full_n;
  wire fifo_C_drain_PE_13_16__write;
  wire [16:0] fifo_C_drain_PE_13_2__dout;
  wire fifo_C_drain_PE_13_2__empty_n;
  wire fifo_C_drain_PE_13_2__read;
  wire [16:0] fifo_C_drain_PE_13_2__din;
  wire fifo_C_drain_PE_13_2__full_n;
  wire fifo_C_drain_PE_13_2__write;
  wire [16:0] fifo_C_drain_PE_13_3__dout;
  wire fifo_C_drain_PE_13_3__empty_n;
  wire fifo_C_drain_PE_13_3__read;
  wire [16:0] fifo_C_drain_PE_13_3__din;
  wire fifo_C_drain_PE_13_3__full_n;
  wire fifo_C_drain_PE_13_3__write;
  wire [16:0] fifo_C_drain_PE_13_4__dout;
  wire fifo_C_drain_PE_13_4__empty_n;
  wire fifo_C_drain_PE_13_4__read;
  wire [16:0] fifo_C_drain_PE_13_4__din;
  wire fifo_C_drain_PE_13_4__full_n;
  wire fifo_C_drain_PE_13_4__write;
  wire [16:0] fifo_C_drain_PE_13_5__dout;
  wire fifo_C_drain_PE_13_5__empty_n;
  wire fifo_C_drain_PE_13_5__read;
  wire [16:0] fifo_C_drain_PE_13_5__din;
  wire fifo_C_drain_PE_13_5__full_n;
  wire fifo_C_drain_PE_13_5__write;
  wire [16:0] fifo_C_drain_PE_13_6__dout;
  wire fifo_C_drain_PE_13_6__empty_n;
  wire fifo_C_drain_PE_13_6__read;
  wire [16:0] fifo_C_drain_PE_13_6__din;
  wire fifo_C_drain_PE_13_6__full_n;
  wire fifo_C_drain_PE_13_6__write;
  wire [16:0] fifo_C_drain_PE_13_7__dout;
  wire fifo_C_drain_PE_13_7__empty_n;
  wire fifo_C_drain_PE_13_7__read;
  wire [16:0] fifo_C_drain_PE_13_7__din;
  wire fifo_C_drain_PE_13_7__full_n;
  wire fifo_C_drain_PE_13_7__write;
  wire [16:0] fifo_C_drain_PE_13_8__dout;
  wire fifo_C_drain_PE_13_8__empty_n;
  wire fifo_C_drain_PE_13_8__read;
  wire [16:0] fifo_C_drain_PE_13_8__din;
  wire fifo_C_drain_PE_13_8__full_n;
  wire fifo_C_drain_PE_13_8__write;
  wire [16:0] fifo_C_drain_PE_13_9__dout;
  wire fifo_C_drain_PE_13_9__empty_n;
  wire fifo_C_drain_PE_13_9__read;
  wire [16:0] fifo_C_drain_PE_13_9__din;
  wire fifo_C_drain_PE_13_9__full_n;
  wire fifo_C_drain_PE_13_9__write;
  wire [16:0] fifo_C_drain_PE_14_0__dout;
  wire fifo_C_drain_PE_14_0__empty_n;
  wire fifo_C_drain_PE_14_0__read;
  wire [16:0] fifo_C_drain_PE_14_0__din;
  wire fifo_C_drain_PE_14_0__full_n;
  wire fifo_C_drain_PE_14_0__write;
  wire [16:0] fifo_C_drain_PE_14_1__dout;
  wire fifo_C_drain_PE_14_1__empty_n;
  wire fifo_C_drain_PE_14_1__read;
  wire [16:0] fifo_C_drain_PE_14_1__din;
  wire fifo_C_drain_PE_14_1__full_n;
  wire fifo_C_drain_PE_14_1__write;
  wire [16:0] fifo_C_drain_PE_14_10__dout;
  wire fifo_C_drain_PE_14_10__empty_n;
  wire fifo_C_drain_PE_14_10__read;
  wire [16:0] fifo_C_drain_PE_14_10__din;
  wire fifo_C_drain_PE_14_10__full_n;
  wire fifo_C_drain_PE_14_10__write;
  wire [16:0] fifo_C_drain_PE_14_11__dout;
  wire fifo_C_drain_PE_14_11__empty_n;
  wire fifo_C_drain_PE_14_11__read;
  wire [16:0] fifo_C_drain_PE_14_11__din;
  wire fifo_C_drain_PE_14_11__full_n;
  wire fifo_C_drain_PE_14_11__write;
  wire [16:0] fifo_C_drain_PE_14_12__dout;
  wire fifo_C_drain_PE_14_12__empty_n;
  wire fifo_C_drain_PE_14_12__read;
  wire [16:0] fifo_C_drain_PE_14_12__din;
  wire fifo_C_drain_PE_14_12__full_n;
  wire fifo_C_drain_PE_14_12__write;
  wire [16:0] fifo_C_drain_PE_14_13__dout;
  wire fifo_C_drain_PE_14_13__empty_n;
  wire fifo_C_drain_PE_14_13__read;
  wire [16:0] fifo_C_drain_PE_14_13__din;
  wire fifo_C_drain_PE_14_13__full_n;
  wire fifo_C_drain_PE_14_13__write;
  wire [16:0] fifo_C_drain_PE_14_14__dout;
  wire fifo_C_drain_PE_14_14__empty_n;
  wire fifo_C_drain_PE_14_14__read;
  wire [16:0] fifo_C_drain_PE_14_14__din;
  wire fifo_C_drain_PE_14_14__full_n;
  wire fifo_C_drain_PE_14_14__write;
  wire [16:0] fifo_C_drain_PE_14_15__dout;
  wire fifo_C_drain_PE_14_15__empty_n;
  wire fifo_C_drain_PE_14_15__read;
  wire [16:0] fifo_C_drain_PE_14_15__din;
  wire fifo_C_drain_PE_14_15__full_n;
  wire fifo_C_drain_PE_14_15__write;
  wire [16:0] fifo_C_drain_PE_14_16__dout;
  wire fifo_C_drain_PE_14_16__empty_n;
  wire fifo_C_drain_PE_14_16__read;
  wire [16:0] fifo_C_drain_PE_14_16__din;
  wire fifo_C_drain_PE_14_16__full_n;
  wire fifo_C_drain_PE_14_16__write;
  wire [16:0] fifo_C_drain_PE_14_2__dout;
  wire fifo_C_drain_PE_14_2__empty_n;
  wire fifo_C_drain_PE_14_2__read;
  wire [16:0] fifo_C_drain_PE_14_2__din;
  wire fifo_C_drain_PE_14_2__full_n;
  wire fifo_C_drain_PE_14_2__write;
  wire [16:0] fifo_C_drain_PE_14_3__dout;
  wire fifo_C_drain_PE_14_3__empty_n;
  wire fifo_C_drain_PE_14_3__read;
  wire [16:0] fifo_C_drain_PE_14_3__din;
  wire fifo_C_drain_PE_14_3__full_n;
  wire fifo_C_drain_PE_14_3__write;
  wire [16:0] fifo_C_drain_PE_14_4__dout;
  wire fifo_C_drain_PE_14_4__empty_n;
  wire fifo_C_drain_PE_14_4__read;
  wire [16:0] fifo_C_drain_PE_14_4__din;
  wire fifo_C_drain_PE_14_4__full_n;
  wire fifo_C_drain_PE_14_4__write;
  wire [16:0] fifo_C_drain_PE_14_5__dout;
  wire fifo_C_drain_PE_14_5__empty_n;
  wire fifo_C_drain_PE_14_5__read;
  wire [16:0] fifo_C_drain_PE_14_5__din;
  wire fifo_C_drain_PE_14_5__full_n;
  wire fifo_C_drain_PE_14_5__write;
  wire [16:0] fifo_C_drain_PE_14_6__dout;
  wire fifo_C_drain_PE_14_6__empty_n;
  wire fifo_C_drain_PE_14_6__read;
  wire [16:0] fifo_C_drain_PE_14_6__din;
  wire fifo_C_drain_PE_14_6__full_n;
  wire fifo_C_drain_PE_14_6__write;
  wire [16:0] fifo_C_drain_PE_14_7__dout;
  wire fifo_C_drain_PE_14_7__empty_n;
  wire fifo_C_drain_PE_14_7__read;
  wire [16:0] fifo_C_drain_PE_14_7__din;
  wire fifo_C_drain_PE_14_7__full_n;
  wire fifo_C_drain_PE_14_7__write;
  wire [16:0] fifo_C_drain_PE_14_8__dout;
  wire fifo_C_drain_PE_14_8__empty_n;
  wire fifo_C_drain_PE_14_8__read;
  wire [16:0] fifo_C_drain_PE_14_8__din;
  wire fifo_C_drain_PE_14_8__full_n;
  wire fifo_C_drain_PE_14_8__write;
  wire [16:0] fifo_C_drain_PE_14_9__dout;
  wire fifo_C_drain_PE_14_9__empty_n;
  wire fifo_C_drain_PE_14_9__read;
  wire [16:0] fifo_C_drain_PE_14_9__din;
  wire fifo_C_drain_PE_14_9__full_n;
  wire fifo_C_drain_PE_14_9__write;
  wire [16:0] fifo_C_drain_PE_15_0__dout;
  wire fifo_C_drain_PE_15_0__empty_n;
  wire fifo_C_drain_PE_15_0__read;
  wire [16:0] fifo_C_drain_PE_15_0__din;
  wire fifo_C_drain_PE_15_0__full_n;
  wire fifo_C_drain_PE_15_0__write;
  wire [16:0] fifo_C_drain_PE_15_1__dout;
  wire fifo_C_drain_PE_15_1__empty_n;
  wire fifo_C_drain_PE_15_1__read;
  wire [16:0] fifo_C_drain_PE_15_1__din;
  wire fifo_C_drain_PE_15_1__full_n;
  wire fifo_C_drain_PE_15_1__write;
  wire [16:0] fifo_C_drain_PE_15_10__dout;
  wire fifo_C_drain_PE_15_10__empty_n;
  wire fifo_C_drain_PE_15_10__read;
  wire [16:0] fifo_C_drain_PE_15_10__din;
  wire fifo_C_drain_PE_15_10__full_n;
  wire fifo_C_drain_PE_15_10__write;
  wire [16:0] fifo_C_drain_PE_15_11__dout;
  wire fifo_C_drain_PE_15_11__empty_n;
  wire fifo_C_drain_PE_15_11__read;
  wire [16:0] fifo_C_drain_PE_15_11__din;
  wire fifo_C_drain_PE_15_11__full_n;
  wire fifo_C_drain_PE_15_11__write;
  wire [16:0] fifo_C_drain_PE_15_12__dout;
  wire fifo_C_drain_PE_15_12__empty_n;
  wire fifo_C_drain_PE_15_12__read;
  wire [16:0] fifo_C_drain_PE_15_12__din;
  wire fifo_C_drain_PE_15_12__full_n;
  wire fifo_C_drain_PE_15_12__write;
  wire [16:0] fifo_C_drain_PE_15_13__dout;
  wire fifo_C_drain_PE_15_13__empty_n;
  wire fifo_C_drain_PE_15_13__read;
  wire [16:0] fifo_C_drain_PE_15_13__din;
  wire fifo_C_drain_PE_15_13__full_n;
  wire fifo_C_drain_PE_15_13__write;
  wire [16:0] fifo_C_drain_PE_15_14__dout;
  wire fifo_C_drain_PE_15_14__empty_n;
  wire fifo_C_drain_PE_15_14__read;
  wire [16:0] fifo_C_drain_PE_15_14__din;
  wire fifo_C_drain_PE_15_14__full_n;
  wire fifo_C_drain_PE_15_14__write;
  wire [16:0] fifo_C_drain_PE_15_15__dout;
  wire fifo_C_drain_PE_15_15__empty_n;
  wire fifo_C_drain_PE_15_15__read;
  wire [16:0] fifo_C_drain_PE_15_15__din;
  wire fifo_C_drain_PE_15_15__full_n;
  wire fifo_C_drain_PE_15_15__write;
  wire [16:0] fifo_C_drain_PE_15_16__dout;
  wire fifo_C_drain_PE_15_16__empty_n;
  wire fifo_C_drain_PE_15_16__read;
  wire [16:0] fifo_C_drain_PE_15_16__din;
  wire fifo_C_drain_PE_15_16__full_n;
  wire fifo_C_drain_PE_15_16__write;
  wire [16:0] fifo_C_drain_PE_15_2__dout;
  wire fifo_C_drain_PE_15_2__empty_n;
  wire fifo_C_drain_PE_15_2__read;
  wire [16:0] fifo_C_drain_PE_15_2__din;
  wire fifo_C_drain_PE_15_2__full_n;
  wire fifo_C_drain_PE_15_2__write;
  wire [16:0] fifo_C_drain_PE_15_3__dout;
  wire fifo_C_drain_PE_15_3__empty_n;
  wire fifo_C_drain_PE_15_3__read;
  wire [16:0] fifo_C_drain_PE_15_3__din;
  wire fifo_C_drain_PE_15_3__full_n;
  wire fifo_C_drain_PE_15_3__write;
  wire [16:0] fifo_C_drain_PE_15_4__dout;
  wire fifo_C_drain_PE_15_4__empty_n;
  wire fifo_C_drain_PE_15_4__read;
  wire [16:0] fifo_C_drain_PE_15_4__din;
  wire fifo_C_drain_PE_15_4__full_n;
  wire fifo_C_drain_PE_15_4__write;
  wire [16:0] fifo_C_drain_PE_15_5__dout;
  wire fifo_C_drain_PE_15_5__empty_n;
  wire fifo_C_drain_PE_15_5__read;
  wire [16:0] fifo_C_drain_PE_15_5__din;
  wire fifo_C_drain_PE_15_5__full_n;
  wire fifo_C_drain_PE_15_5__write;
  wire [16:0] fifo_C_drain_PE_15_6__dout;
  wire fifo_C_drain_PE_15_6__empty_n;
  wire fifo_C_drain_PE_15_6__read;
  wire [16:0] fifo_C_drain_PE_15_6__din;
  wire fifo_C_drain_PE_15_6__full_n;
  wire fifo_C_drain_PE_15_6__write;
  wire [16:0] fifo_C_drain_PE_15_7__dout;
  wire fifo_C_drain_PE_15_7__empty_n;
  wire fifo_C_drain_PE_15_7__read;
  wire [16:0] fifo_C_drain_PE_15_7__din;
  wire fifo_C_drain_PE_15_7__full_n;
  wire fifo_C_drain_PE_15_7__write;
  wire [16:0] fifo_C_drain_PE_15_8__dout;
  wire fifo_C_drain_PE_15_8__empty_n;
  wire fifo_C_drain_PE_15_8__read;
  wire [16:0] fifo_C_drain_PE_15_8__din;
  wire fifo_C_drain_PE_15_8__full_n;
  wire fifo_C_drain_PE_15_8__write;
  wire [16:0] fifo_C_drain_PE_15_9__dout;
  wire fifo_C_drain_PE_15_9__empty_n;
  wire fifo_C_drain_PE_15_9__read;
  wire [16:0] fifo_C_drain_PE_15_9__din;
  wire fifo_C_drain_PE_15_9__full_n;
  wire fifo_C_drain_PE_15_9__write;
  wire [16:0] fifo_C_drain_PE_16_0__dout;
  wire fifo_C_drain_PE_16_0__empty_n;
  wire fifo_C_drain_PE_16_0__read;
  wire [16:0] fifo_C_drain_PE_16_0__din;
  wire fifo_C_drain_PE_16_0__full_n;
  wire fifo_C_drain_PE_16_0__write;
  wire [16:0] fifo_C_drain_PE_16_1__dout;
  wire fifo_C_drain_PE_16_1__empty_n;
  wire fifo_C_drain_PE_16_1__read;
  wire [16:0] fifo_C_drain_PE_16_1__din;
  wire fifo_C_drain_PE_16_1__full_n;
  wire fifo_C_drain_PE_16_1__write;
  wire [16:0] fifo_C_drain_PE_16_10__dout;
  wire fifo_C_drain_PE_16_10__empty_n;
  wire fifo_C_drain_PE_16_10__read;
  wire [16:0] fifo_C_drain_PE_16_10__din;
  wire fifo_C_drain_PE_16_10__full_n;
  wire fifo_C_drain_PE_16_10__write;
  wire [16:0] fifo_C_drain_PE_16_11__dout;
  wire fifo_C_drain_PE_16_11__empty_n;
  wire fifo_C_drain_PE_16_11__read;
  wire [16:0] fifo_C_drain_PE_16_11__din;
  wire fifo_C_drain_PE_16_11__full_n;
  wire fifo_C_drain_PE_16_11__write;
  wire [16:0] fifo_C_drain_PE_16_12__dout;
  wire fifo_C_drain_PE_16_12__empty_n;
  wire fifo_C_drain_PE_16_12__read;
  wire [16:0] fifo_C_drain_PE_16_12__din;
  wire fifo_C_drain_PE_16_12__full_n;
  wire fifo_C_drain_PE_16_12__write;
  wire [16:0] fifo_C_drain_PE_16_13__dout;
  wire fifo_C_drain_PE_16_13__empty_n;
  wire fifo_C_drain_PE_16_13__read;
  wire [16:0] fifo_C_drain_PE_16_13__din;
  wire fifo_C_drain_PE_16_13__full_n;
  wire fifo_C_drain_PE_16_13__write;
  wire [16:0] fifo_C_drain_PE_16_14__dout;
  wire fifo_C_drain_PE_16_14__empty_n;
  wire fifo_C_drain_PE_16_14__read;
  wire [16:0] fifo_C_drain_PE_16_14__din;
  wire fifo_C_drain_PE_16_14__full_n;
  wire fifo_C_drain_PE_16_14__write;
  wire [16:0] fifo_C_drain_PE_16_15__dout;
  wire fifo_C_drain_PE_16_15__empty_n;
  wire fifo_C_drain_PE_16_15__read;
  wire [16:0] fifo_C_drain_PE_16_15__din;
  wire fifo_C_drain_PE_16_15__full_n;
  wire fifo_C_drain_PE_16_15__write;
  wire [16:0] fifo_C_drain_PE_16_16__dout;
  wire fifo_C_drain_PE_16_16__empty_n;
  wire fifo_C_drain_PE_16_16__read;
  wire [16:0] fifo_C_drain_PE_16_16__din;
  wire fifo_C_drain_PE_16_16__full_n;
  wire fifo_C_drain_PE_16_16__write;
  wire [16:0] fifo_C_drain_PE_16_2__dout;
  wire fifo_C_drain_PE_16_2__empty_n;
  wire fifo_C_drain_PE_16_2__read;
  wire [16:0] fifo_C_drain_PE_16_2__din;
  wire fifo_C_drain_PE_16_2__full_n;
  wire fifo_C_drain_PE_16_2__write;
  wire [16:0] fifo_C_drain_PE_16_3__dout;
  wire fifo_C_drain_PE_16_3__empty_n;
  wire fifo_C_drain_PE_16_3__read;
  wire [16:0] fifo_C_drain_PE_16_3__din;
  wire fifo_C_drain_PE_16_3__full_n;
  wire fifo_C_drain_PE_16_3__write;
  wire [16:0] fifo_C_drain_PE_16_4__dout;
  wire fifo_C_drain_PE_16_4__empty_n;
  wire fifo_C_drain_PE_16_4__read;
  wire [16:0] fifo_C_drain_PE_16_4__din;
  wire fifo_C_drain_PE_16_4__full_n;
  wire fifo_C_drain_PE_16_4__write;
  wire [16:0] fifo_C_drain_PE_16_5__dout;
  wire fifo_C_drain_PE_16_5__empty_n;
  wire fifo_C_drain_PE_16_5__read;
  wire [16:0] fifo_C_drain_PE_16_5__din;
  wire fifo_C_drain_PE_16_5__full_n;
  wire fifo_C_drain_PE_16_5__write;
  wire [16:0] fifo_C_drain_PE_16_6__dout;
  wire fifo_C_drain_PE_16_6__empty_n;
  wire fifo_C_drain_PE_16_6__read;
  wire [16:0] fifo_C_drain_PE_16_6__din;
  wire fifo_C_drain_PE_16_6__full_n;
  wire fifo_C_drain_PE_16_6__write;
  wire [16:0] fifo_C_drain_PE_16_7__dout;
  wire fifo_C_drain_PE_16_7__empty_n;
  wire fifo_C_drain_PE_16_7__read;
  wire [16:0] fifo_C_drain_PE_16_7__din;
  wire fifo_C_drain_PE_16_7__full_n;
  wire fifo_C_drain_PE_16_7__write;
  wire [16:0] fifo_C_drain_PE_16_8__dout;
  wire fifo_C_drain_PE_16_8__empty_n;
  wire fifo_C_drain_PE_16_8__read;
  wire [16:0] fifo_C_drain_PE_16_8__din;
  wire fifo_C_drain_PE_16_8__full_n;
  wire fifo_C_drain_PE_16_8__write;
  wire [16:0] fifo_C_drain_PE_16_9__dout;
  wire fifo_C_drain_PE_16_9__empty_n;
  wire fifo_C_drain_PE_16_9__read;
  wire [16:0] fifo_C_drain_PE_16_9__din;
  wire fifo_C_drain_PE_16_9__full_n;
  wire fifo_C_drain_PE_16_9__write;
  wire [16:0] fifo_C_drain_PE_17_0__dout;
  wire fifo_C_drain_PE_17_0__empty_n;
  wire fifo_C_drain_PE_17_0__read;
  wire [16:0] fifo_C_drain_PE_17_0__din;
  wire fifo_C_drain_PE_17_0__full_n;
  wire fifo_C_drain_PE_17_0__write;
  wire [16:0] fifo_C_drain_PE_17_1__dout;
  wire fifo_C_drain_PE_17_1__empty_n;
  wire fifo_C_drain_PE_17_1__read;
  wire [16:0] fifo_C_drain_PE_17_1__din;
  wire fifo_C_drain_PE_17_1__full_n;
  wire fifo_C_drain_PE_17_1__write;
  wire [16:0] fifo_C_drain_PE_17_10__dout;
  wire fifo_C_drain_PE_17_10__empty_n;
  wire fifo_C_drain_PE_17_10__read;
  wire [16:0] fifo_C_drain_PE_17_10__din;
  wire fifo_C_drain_PE_17_10__full_n;
  wire fifo_C_drain_PE_17_10__write;
  wire [16:0] fifo_C_drain_PE_17_11__dout;
  wire fifo_C_drain_PE_17_11__empty_n;
  wire fifo_C_drain_PE_17_11__read;
  wire [16:0] fifo_C_drain_PE_17_11__din;
  wire fifo_C_drain_PE_17_11__full_n;
  wire fifo_C_drain_PE_17_11__write;
  wire [16:0] fifo_C_drain_PE_17_12__dout;
  wire fifo_C_drain_PE_17_12__empty_n;
  wire fifo_C_drain_PE_17_12__read;
  wire [16:0] fifo_C_drain_PE_17_12__din;
  wire fifo_C_drain_PE_17_12__full_n;
  wire fifo_C_drain_PE_17_12__write;
  wire [16:0] fifo_C_drain_PE_17_13__dout;
  wire fifo_C_drain_PE_17_13__empty_n;
  wire fifo_C_drain_PE_17_13__read;
  wire [16:0] fifo_C_drain_PE_17_13__din;
  wire fifo_C_drain_PE_17_13__full_n;
  wire fifo_C_drain_PE_17_13__write;
  wire [16:0] fifo_C_drain_PE_17_14__dout;
  wire fifo_C_drain_PE_17_14__empty_n;
  wire fifo_C_drain_PE_17_14__read;
  wire [16:0] fifo_C_drain_PE_17_14__din;
  wire fifo_C_drain_PE_17_14__full_n;
  wire fifo_C_drain_PE_17_14__write;
  wire [16:0] fifo_C_drain_PE_17_15__dout;
  wire fifo_C_drain_PE_17_15__empty_n;
  wire fifo_C_drain_PE_17_15__read;
  wire [16:0] fifo_C_drain_PE_17_15__din;
  wire fifo_C_drain_PE_17_15__full_n;
  wire fifo_C_drain_PE_17_15__write;
  wire [16:0] fifo_C_drain_PE_17_16__dout;
  wire fifo_C_drain_PE_17_16__empty_n;
  wire fifo_C_drain_PE_17_16__read;
  wire [16:0] fifo_C_drain_PE_17_16__din;
  wire fifo_C_drain_PE_17_16__full_n;
  wire fifo_C_drain_PE_17_16__write;
  wire [16:0] fifo_C_drain_PE_17_2__dout;
  wire fifo_C_drain_PE_17_2__empty_n;
  wire fifo_C_drain_PE_17_2__read;
  wire [16:0] fifo_C_drain_PE_17_2__din;
  wire fifo_C_drain_PE_17_2__full_n;
  wire fifo_C_drain_PE_17_2__write;
  wire [16:0] fifo_C_drain_PE_17_3__dout;
  wire fifo_C_drain_PE_17_3__empty_n;
  wire fifo_C_drain_PE_17_3__read;
  wire [16:0] fifo_C_drain_PE_17_3__din;
  wire fifo_C_drain_PE_17_3__full_n;
  wire fifo_C_drain_PE_17_3__write;
  wire [16:0] fifo_C_drain_PE_17_4__dout;
  wire fifo_C_drain_PE_17_4__empty_n;
  wire fifo_C_drain_PE_17_4__read;
  wire [16:0] fifo_C_drain_PE_17_4__din;
  wire fifo_C_drain_PE_17_4__full_n;
  wire fifo_C_drain_PE_17_4__write;
  wire [16:0] fifo_C_drain_PE_17_5__dout;
  wire fifo_C_drain_PE_17_5__empty_n;
  wire fifo_C_drain_PE_17_5__read;
  wire [16:0] fifo_C_drain_PE_17_5__din;
  wire fifo_C_drain_PE_17_5__full_n;
  wire fifo_C_drain_PE_17_5__write;
  wire [16:0] fifo_C_drain_PE_17_6__dout;
  wire fifo_C_drain_PE_17_6__empty_n;
  wire fifo_C_drain_PE_17_6__read;
  wire [16:0] fifo_C_drain_PE_17_6__din;
  wire fifo_C_drain_PE_17_6__full_n;
  wire fifo_C_drain_PE_17_6__write;
  wire [16:0] fifo_C_drain_PE_17_7__dout;
  wire fifo_C_drain_PE_17_7__empty_n;
  wire fifo_C_drain_PE_17_7__read;
  wire [16:0] fifo_C_drain_PE_17_7__din;
  wire fifo_C_drain_PE_17_7__full_n;
  wire fifo_C_drain_PE_17_7__write;
  wire [16:0] fifo_C_drain_PE_17_8__dout;
  wire fifo_C_drain_PE_17_8__empty_n;
  wire fifo_C_drain_PE_17_8__read;
  wire [16:0] fifo_C_drain_PE_17_8__din;
  wire fifo_C_drain_PE_17_8__full_n;
  wire fifo_C_drain_PE_17_8__write;
  wire [16:0] fifo_C_drain_PE_17_9__dout;
  wire fifo_C_drain_PE_17_9__empty_n;
  wire fifo_C_drain_PE_17_9__read;
  wire [16:0] fifo_C_drain_PE_17_9__din;
  wire fifo_C_drain_PE_17_9__full_n;
  wire fifo_C_drain_PE_17_9__write;
  wire [16:0] fifo_C_drain_PE_1_0__dout;
  wire fifo_C_drain_PE_1_0__empty_n;
  wire fifo_C_drain_PE_1_0__read;
  wire [16:0] fifo_C_drain_PE_1_0__din;
  wire fifo_C_drain_PE_1_0__full_n;
  wire fifo_C_drain_PE_1_0__write;
  wire [16:0] fifo_C_drain_PE_1_1__dout;
  wire fifo_C_drain_PE_1_1__empty_n;
  wire fifo_C_drain_PE_1_1__read;
  wire [16:0] fifo_C_drain_PE_1_1__din;
  wire fifo_C_drain_PE_1_1__full_n;
  wire fifo_C_drain_PE_1_1__write;
  wire [16:0] fifo_C_drain_PE_1_10__dout;
  wire fifo_C_drain_PE_1_10__empty_n;
  wire fifo_C_drain_PE_1_10__read;
  wire [16:0] fifo_C_drain_PE_1_10__din;
  wire fifo_C_drain_PE_1_10__full_n;
  wire fifo_C_drain_PE_1_10__write;
  wire [16:0] fifo_C_drain_PE_1_11__dout;
  wire fifo_C_drain_PE_1_11__empty_n;
  wire fifo_C_drain_PE_1_11__read;
  wire [16:0] fifo_C_drain_PE_1_11__din;
  wire fifo_C_drain_PE_1_11__full_n;
  wire fifo_C_drain_PE_1_11__write;
  wire [16:0] fifo_C_drain_PE_1_12__dout;
  wire fifo_C_drain_PE_1_12__empty_n;
  wire fifo_C_drain_PE_1_12__read;
  wire [16:0] fifo_C_drain_PE_1_12__din;
  wire fifo_C_drain_PE_1_12__full_n;
  wire fifo_C_drain_PE_1_12__write;
  wire [16:0] fifo_C_drain_PE_1_13__dout;
  wire fifo_C_drain_PE_1_13__empty_n;
  wire fifo_C_drain_PE_1_13__read;
  wire [16:0] fifo_C_drain_PE_1_13__din;
  wire fifo_C_drain_PE_1_13__full_n;
  wire fifo_C_drain_PE_1_13__write;
  wire [16:0] fifo_C_drain_PE_1_14__dout;
  wire fifo_C_drain_PE_1_14__empty_n;
  wire fifo_C_drain_PE_1_14__read;
  wire [16:0] fifo_C_drain_PE_1_14__din;
  wire fifo_C_drain_PE_1_14__full_n;
  wire fifo_C_drain_PE_1_14__write;
  wire [16:0] fifo_C_drain_PE_1_15__dout;
  wire fifo_C_drain_PE_1_15__empty_n;
  wire fifo_C_drain_PE_1_15__read;
  wire [16:0] fifo_C_drain_PE_1_15__din;
  wire fifo_C_drain_PE_1_15__full_n;
  wire fifo_C_drain_PE_1_15__write;
  wire [16:0] fifo_C_drain_PE_1_16__dout;
  wire fifo_C_drain_PE_1_16__empty_n;
  wire fifo_C_drain_PE_1_16__read;
  wire [16:0] fifo_C_drain_PE_1_16__din;
  wire fifo_C_drain_PE_1_16__full_n;
  wire fifo_C_drain_PE_1_16__write;
  wire [16:0] fifo_C_drain_PE_1_2__dout;
  wire fifo_C_drain_PE_1_2__empty_n;
  wire fifo_C_drain_PE_1_2__read;
  wire [16:0] fifo_C_drain_PE_1_2__din;
  wire fifo_C_drain_PE_1_2__full_n;
  wire fifo_C_drain_PE_1_2__write;
  wire [16:0] fifo_C_drain_PE_1_3__dout;
  wire fifo_C_drain_PE_1_3__empty_n;
  wire fifo_C_drain_PE_1_3__read;
  wire [16:0] fifo_C_drain_PE_1_3__din;
  wire fifo_C_drain_PE_1_3__full_n;
  wire fifo_C_drain_PE_1_3__write;
  wire [16:0] fifo_C_drain_PE_1_4__dout;
  wire fifo_C_drain_PE_1_4__empty_n;
  wire fifo_C_drain_PE_1_4__read;
  wire [16:0] fifo_C_drain_PE_1_4__din;
  wire fifo_C_drain_PE_1_4__full_n;
  wire fifo_C_drain_PE_1_4__write;
  wire [16:0] fifo_C_drain_PE_1_5__dout;
  wire fifo_C_drain_PE_1_5__empty_n;
  wire fifo_C_drain_PE_1_5__read;
  wire [16:0] fifo_C_drain_PE_1_5__din;
  wire fifo_C_drain_PE_1_5__full_n;
  wire fifo_C_drain_PE_1_5__write;
  wire [16:0] fifo_C_drain_PE_1_6__dout;
  wire fifo_C_drain_PE_1_6__empty_n;
  wire fifo_C_drain_PE_1_6__read;
  wire [16:0] fifo_C_drain_PE_1_6__din;
  wire fifo_C_drain_PE_1_6__full_n;
  wire fifo_C_drain_PE_1_6__write;
  wire [16:0] fifo_C_drain_PE_1_7__dout;
  wire fifo_C_drain_PE_1_7__empty_n;
  wire fifo_C_drain_PE_1_7__read;
  wire [16:0] fifo_C_drain_PE_1_7__din;
  wire fifo_C_drain_PE_1_7__full_n;
  wire fifo_C_drain_PE_1_7__write;
  wire [16:0] fifo_C_drain_PE_1_8__dout;
  wire fifo_C_drain_PE_1_8__empty_n;
  wire fifo_C_drain_PE_1_8__read;
  wire [16:0] fifo_C_drain_PE_1_8__din;
  wire fifo_C_drain_PE_1_8__full_n;
  wire fifo_C_drain_PE_1_8__write;
  wire [16:0] fifo_C_drain_PE_1_9__dout;
  wire fifo_C_drain_PE_1_9__empty_n;
  wire fifo_C_drain_PE_1_9__read;
  wire [16:0] fifo_C_drain_PE_1_9__din;
  wire fifo_C_drain_PE_1_9__full_n;
  wire fifo_C_drain_PE_1_9__write;
  wire [16:0] fifo_C_drain_PE_2_0__dout;
  wire fifo_C_drain_PE_2_0__empty_n;
  wire fifo_C_drain_PE_2_0__read;
  wire [16:0] fifo_C_drain_PE_2_0__din;
  wire fifo_C_drain_PE_2_0__full_n;
  wire fifo_C_drain_PE_2_0__write;
  wire [16:0] fifo_C_drain_PE_2_1__dout;
  wire fifo_C_drain_PE_2_1__empty_n;
  wire fifo_C_drain_PE_2_1__read;
  wire [16:0] fifo_C_drain_PE_2_1__din;
  wire fifo_C_drain_PE_2_1__full_n;
  wire fifo_C_drain_PE_2_1__write;
  wire [16:0] fifo_C_drain_PE_2_10__dout;
  wire fifo_C_drain_PE_2_10__empty_n;
  wire fifo_C_drain_PE_2_10__read;
  wire [16:0] fifo_C_drain_PE_2_10__din;
  wire fifo_C_drain_PE_2_10__full_n;
  wire fifo_C_drain_PE_2_10__write;
  wire [16:0] fifo_C_drain_PE_2_11__dout;
  wire fifo_C_drain_PE_2_11__empty_n;
  wire fifo_C_drain_PE_2_11__read;
  wire [16:0] fifo_C_drain_PE_2_11__din;
  wire fifo_C_drain_PE_2_11__full_n;
  wire fifo_C_drain_PE_2_11__write;
  wire [16:0] fifo_C_drain_PE_2_12__dout;
  wire fifo_C_drain_PE_2_12__empty_n;
  wire fifo_C_drain_PE_2_12__read;
  wire [16:0] fifo_C_drain_PE_2_12__din;
  wire fifo_C_drain_PE_2_12__full_n;
  wire fifo_C_drain_PE_2_12__write;
  wire [16:0] fifo_C_drain_PE_2_13__dout;
  wire fifo_C_drain_PE_2_13__empty_n;
  wire fifo_C_drain_PE_2_13__read;
  wire [16:0] fifo_C_drain_PE_2_13__din;
  wire fifo_C_drain_PE_2_13__full_n;
  wire fifo_C_drain_PE_2_13__write;
  wire [16:0] fifo_C_drain_PE_2_14__dout;
  wire fifo_C_drain_PE_2_14__empty_n;
  wire fifo_C_drain_PE_2_14__read;
  wire [16:0] fifo_C_drain_PE_2_14__din;
  wire fifo_C_drain_PE_2_14__full_n;
  wire fifo_C_drain_PE_2_14__write;
  wire [16:0] fifo_C_drain_PE_2_15__dout;
  wire fifo_C_drain_PE_2_15__empty_n;
  wire fifo_C_drain_PE_2_15__read;
  wire [16:0] fifo_C_drain_PE_2_15__din;
  wire fifo_C_drain_PE_2_15__full_n;
  wire fifo_C_drain_PE_2_15__write;
  wire [16:0] fifo_C_drain_PE_2_16__dout;
  wire fifo_C_drain_PE_2_16__empty_n;
  wire fifo_C_drain_PE_2_16__read;
  wire [16:0] fifo_C_drain_PE_2_16__din;
  wire fifo_C_drain_PE_2_16__full_n;
  wire fifo_C_drain_PE_2_16__write;
  wire [16:0] fifo_C_drain_PE_2_2__dout;
  wire fifo_C_drain_PE_2_2__empty_n;
  wire fifo_C_drain_PE_2_2__read;
  wire [16:0] fifo_C_drain_PE_2_2__din;
  wire fifo_C_drain_PE_2_2__full_n;
  wire fifo_C_drain_PE_2_2__write;
  wire [16:0] fifo_C_drain_PE_2_3__dout;
  wire fifo_C_drain_PE_2_3__empty_n;
  wire fifo_C_drain_PE_2_3__read;
  wire [16:0] fifo_C_drain_PE_2_3__din;
  wire fifo_C_drain_PE_2_3__full_n;
  wire fifo_C_drain_PE_2_3__write;
  wire [16:0] fifo_C_drain_PE_2_4__dout;
  wire fifo_C_drain_PE_2_4__empty_n;
  wire fifo_C_drain_PE_2_4__read;
  wire [16:0] fifo_C_drain_PE_2_4__din;
  wire fifo_C_drain_PE_2_4__full_n;
  wire fifo_C_drain_PE_2_4__write;
  wire [16:0] fifo_C_drain_PE_2_5__dout;
  wire fifo_C_drain_PE_2_5__empty_n;
  wire fifo_C_drain_PE_2_5__read;
  wire [16:0] fifo_C_drain_PE_2_5__din;
  wire fifo_C_drain_PE_2_5__full_n;
  wire fifo_C_drain_PE_2_5__write;
  wire [16:0] fifo_C_drain_PE_2_6__dout;
  wire fifo_C_drain_PE_2_6__empty_n;
  wire fifo_C_drain_PE_2_6__read;
  wire [16:0] fifo_C_drain_PE_2_6__din;
  wire fifo_C_drain_PE_2_6__full_n;
  wire fifo_C_drain_PE_2_6__write;
  wire [16:0] fifo_C_drain_PE_2_7__dout;
  wire fifo_C_drain_PE_2_7__empty_n;
  wire fifo_C_drain_PE_2_7__read;
  wire [16:0] fifo_C_drain_PE_2_7__din;
  wire fifo_C_drain_PE_2_7__full_n;
  wire fifo_C_drain_PE_2_7__write;
  wire [16:0] fifo_C_drain_PE_2_8__dout;
  wire fifo_C_drain_PE_2_8__empty_n;
  wire fifo_C_drain_PE_2_8__read;
  wire [16:0] fifo_C_drain_PE_2_8__din;
  wire fifo_C_drain_PE_2_8__full_n;
  wire fifo_C_drain_PE_2_8__write;
  wire [16:0] fifo_C_drain_PE_2_9__dout;
  wire fifo_C_drain_PE_2_9__empty_n;
  wire fifo_C_drain_PE_2_9__read;
  wire [16:0] fifo_C_drain_PE_2_9__din;
  wire fifo_C_drain_PE_2_9__full_n;
  wire fifo_C_drain_PE_2_9__write;
  wire [16:0] fifo_C_drain_PE_3_0__dout;
  wire fifo_C_drain_PE_3_0__empty_n;
  wire fifo_C_drain_PE_3_0__read;
  wire [16:0] fifo_C_drain_PE_3_0__din;
  wire fifo_C_drain_PE_3_0__full_n;
  wire fifo_C_drain_PE_3_0__write;
  wire [16:0] fifo_C_drain_PE_3_1__dout;
  wire fifo_C_drain_PE_3_1__empty_n;
  wire fifo_C_drain_PE_3_1__read;
  wire [16:0] fifo_C_drain_PE_3_1__din;
  wire fifo_C_drain_PE_3_1__full_n;
  wire fifo_C_drain_PE_3_1__write;
  wire [16:0] fifo_C_drain_PE_3_10__dout;
  wire fifo_C_drain_PE_3_10__empty_n;
  wire fifo_C_drain_PE_3_10__read;
  wire [16:0] fifo_C_drain_PE_3_10__din;
  wire fifo_C_drain_PE_3_10__full_n;
  wire fifo_C_drain_PE_3_10__write;
  wire [16:0] fifo_C_drain_PE_3_11__dout;
  wire fifo_C_drain_PE_3_11__empty_n;
  wire fifo_C_drain_PE_3_11__read;
  wire [16:0] fifo_C_drain_PE_3_11__din;
  wire fifo_C_drain_PE_3_11__full_n;
  wire fifo_C_drain_PE_3_11__write;
  wire [16:0] fifo_C_drain_PE_3_12__dout;
  wire fifo_C_drain_PE_3_12__empty_n;
  wire fifo_C_drain_PE_3_12__read;
  wire [16:0] fifo_C_drain_PE_3_12__din;
  wire fifo_C_drain_PE_3_12__full_n;
  wire fifo_C_drain_PE_3_12__write;
  wire [16:0] fifo_C_drain_PE_3_13__dout;
  wire fifo_C_drain_PE_3_13__empty_n;
  wire fifo_C_drain_PE_3_13__read;
  wire [16:0] fifo_C_drain_PE_3_13__din;
  wire fifo_C_drain_PE_3_13__full_n;
  wire fifo_C_drain_PE_3_13__write;
  wire [16:0] fifo_C_drain_PE_3_14__dout;
  wire fifo_C_drain_PE_3_14__empty_n;
  wire fifo_C_drain_PE_3_14__read;
  wire [16:0] fifo_C_drain_PE_3_14__din;
  wire fifo_C_drain_PE_3_14__full_n;
  wire fifo_C_drain_PE_3_14__write;
  wire [16:0] fifo_C_drain_PE_3_15__dout;
  wire fifo_C_drain_PE_3_15__empty_n;
  wire fifo_C_drain_PE_3_15__read;
  wire [16:0] fifo_C_drain_PE_3_15__din;
  wire fifo_C_drain_PE_3_15__full_n;
  wire fifo_C_drain_PE_3_15__write;
  wire [16:0] fifo_C_drain_PE_3_16__dout;
  wire fifo_C_drain_PE_3_16__empty_n;
  wire fifo_C_drain_PE_3_16__read;
  wire [16:0] fifo_C_drain_PE_3_16__din;
  wire fifo_C_drain_PE_3_16__full_n;
  wire fifo_C_drain_PE_3_16__write;
  wire [16:0] fifo_C_drain_PE_3_2__dout;
  wire fifo_C_drain_PE_3_2__empty_n;
  wire fifo_C_drain_PE_3_2__read;
  wire [16:0] fifo_C_drain_PE_3_2__din;
  wire fifo_C_drain_PE_3_2__full_n;
  wire fifo_C_drain_PE_3_2__write;
  wire [16:0] fifo_C_drain_PE_3_3__dout;
  wire fifo_C_drain_PE_3_3__empty_n;
  wire fifo_C_drain_PE_3_3__read;
  wire [16:0] fifo_C_drain_PE_3_3__din;
  wire fifo_C_drain_PE_3_3__full_n;
  wire fifo_C_drain_PE_3_3__write;
  wire [16:0] fifo_C_drain_PE_3_4__dout;
  wire fifo_C_drain_PE_3_4__empty_n;
  wire fifo_C_drain_PE_3_4__read;
  wire [16:0] fifo_C_drain_PE_3_4__din;
  wire fifo_C_drain_PE_3_4__full_n;
  wire fifo_C_drain_PE_3_4__write;
  wire [16:0] fifo_C_drain_PE_3_5__dout;
  wire fifo_C_drain_PE_3_5__empty_n;
  wire fifo_C_drain_PE_3_5__read;
  wire [16:0] fifo_C_drain_PE_3_5__din;
  wire fifo_C_drain_PE_3_5__full_n;
  wire fifo_C_drain_PE_3_5__write;
  wire [16:0] fifo_C_drain_PE_3_6__dout;
  wire fifo_C_drain_PE_3_6__empty_n;
  wire fifo_C_drain_PE_3_6__read;
  wire [16:0] fifo_C_drain_PE_3_6__din;
  wire fifo_C_drain_PE_3_6__full_n;
  wire fifo_C_drain_PE_3_6__write;
  wire [16:0] fifo_C_drain_PE_3_7__dout;
  wire fifo_C_drain_PE_3_7__empty_n;
  wire fifo_C_drain_PE_3_7__read;
  wire [16:0] fifo_C_drain_PE_3_7__din;
  wire fifo_C_drain_PE_3_7__full_n;
  wire fifo_C_drain_PE_3_7__write;
  wire [16:0] fifo_C_drain_PE_3_8__dout;
  wire fifo_C_drain_PE_3_8__empty_n;
  wire fifo_C_drain_PE_3_8__read;
  wire [16:0] fifo_C_drain_PE_3_8__din;
  wire fifo_C_drain_PE_3_8__full_n;
  wire fifo_C_drain_PE_3_8__write;
  wire [16:0] fifo_C_drain_PE_3_9__dout;
  wire fifo_C_drain_PE_3_9__empty_n;
  wire fifo_C_drain_PE_3_9__read;
  wire [16:0] fifo_C_drain_PE_3_9__din;
  wire fifo_C_drain_PE_3_9__full_n;
  wire fifo_C_drain_PE_3_9__write;
  wire [16:0] fifo_C_drain_PE_4_0__dout;
  wire fifo_C_drain_PE_4_0__empty_n;
  wire fifo_C_drain_PE_4_0__read;
  wire [16:0] fifo_C_drain_PE_4_0__din;
  wire fifo_C_drain_PE_4_0__full_n;
  wire fifo_C_drain_PE_4_0__write;
  wire [16:0] fifo_C_drain_PE_4_1__dout;
  wire fifo_C_drain_PE_4_1__empty_n;
  wire fifo_C_drain_PE_4_1__read;
  wire [16:0] fifo_C_drain_PE_4_1__din;
  wire fifo_C_drain_PE_4_1__full_n;
  wire fifo_C_drain_PE_4_1__write;
  wire [16:0] fifo_C_drain_PE_4_10__dout;
  wire fifo_C_drain_PE_4_10__empty_n;
  wire fifo_C_drain_PE_4_10__read;
  wire [16:0] fifo_C_drain_PE_4_10__din;
  wire fifo_C_drain_PE_4_10__full_n;
  wire fifo_C_drain_PE_4_10__write;
  wire [16:0] fifo_C_drain_PE_4_11__dout;
  wire fifo_C_drain_PE_4_11__empty_n;
  wire fifo_C_drain_PE_4_11__read;
  wire [16:0] fifo_C_drain_PE_4_11__din;
  wire fifo_C_drain_PE_4_11__full_n;
  wire fifo_C_drain_PE_4_11__write;
  wire [16:0] fifo_C_drain_PE_4_12__dout;
  wire fifo_C_drain_PE_4_12__empty_n;
  wire fifo_C_drain_PE_4_12__read;
  wire [16:0] fifo_C_drain_PE_4_12__din;
  wire fifo_C_drain_PE_4_12__full_n;
  wire fifo_C_drain_PE_4_12__write;
  wire [16:0] fifo_C_drain_PE_4_13__dout;
  wire fifo_C_drain_PE_4_13__empty_n;
  wire fifo_C_drain_PE_4_13__read;
  wire [16:0] fifo_C_drain_PE_4_13__din;
  wire fifo_C_drain_PE_4_13__full_n;
  wire fifo_C_drain_PE_4_13__write;
  wire [16:0] fifo_C_drain_PE_4_14__dout;
  wire fifo_C_drain_PE_4_14__empty_n;
  wire fifo_C_drain_PE_4_14__read;
  wire [16:0] fifo_C_drain_PE_4_14__din;
  wire fifo_C_drain_PE_4_14__full_n;
  wire fifo_C_drain_PE_4_14__write;
  wire [16:0] fifo_C_drain_PE_4_15__dout;
  wire fifo_C_drain_PE_4_15__empty_n;
  wire fifo_C_drain_PE_4_15__read;
  wire [16:0] fifo_C_drain_PE_4_15__din;
  wire fifo_C_drain_PE_4_15__full_n;
  wire fifo_C_drain_PE_4_15__write;
  wire [16:0] fifo_C_drain_PE_4_16__dout;
  wire fifo_C_drain_PE_4_16__empty_n;
  wire fifo_C_drain_PE_4_16__read;
  wire [16:0] fifo_C_drain_PE_4_16__din;
  wire fifo_C_drain_PE_4_16__full_n;
  wire fifo_C_drain_PE_4_16__write;
  wire [16:0] fifo_C_drain_PE_4_2__dout;
  wire fifo_C_drain_PE_4_2__empty_n;
  wire fifo_C_drain_PE_4_2__read;
  wire [16:0] fifo_C_drain_PE_4_2__din;
  wire fifo_C_drain_PE_4_2__full_n;
  wire fifo_C_drain_PE_4_2__write;
  wire [16:0] fifo_C_drain_PE_4_3__dout;
  wire fifo_C_drain_PE_4_3__empty_n;
  wire fifo_C_drain_PE_4_3__read;
  wire [16:0] fifo_C_drain_PE_4_3__din;
  wire fifo_C_drain_PE_4_3__full_n;
  wire fifo_C_drain_PE_4_3__write;
  wire [16:0] fifo_C_drain_PE_4_4__dout;
  wire fifo_C_drain_PE_4_4__empty_n;
  wire fifo_C_drain_PE_4_4__read;
  wire [16:0] fifo_C_drain_PE_4_4__din;
  wire fifo_C_drain_PE_4_4__full_n;
  wire fifo_C_drain_PE_4_4__write;
  wire [16:0] fifo_C_drain_PE_4_5__dout;
  wire fifo_C_drain_PE_4_5__empty_n;
  wire fifo_C_drain_PE_4_5__read;
  wire [16:0] fifo_C_drain_PE_4_5__din;
  wire fifo_C_drain_PE_4_5__full_n;
  wire fifo_C_drain_PE_4_5__write;
  wire [16:0] fifo_C_drain_PE_4_6__dout;
  wire fifo_C_drain_PE_4_6__empty_n;
  wire fifo_C_drain_PE_4_6__read;
  wire [16:0] fifo_C_drain_PE_4_6__din;
  wire fifo_C_drain_PE_4_6__full_n;
  wire fifo_C_drain_PE_4_6__write;
  wire [16:0] fifo_C_drain_PE_4_7__dout;
  wire fifo_C_drain_PE_4_7__empty_n;
  wire fifo_C_drain_PE_4_7__read;
  wire [16:0] fifo_C_drain_PE_4_7__din;
  wire fifo_C_drain_PE_4_7__full_n;
  wire fifo_C_drain_PE_4_7__write;
  wire [16:0] fifo_C_drain_PE_4_8__dout;
  wire fifo_C_drain_PE_4_8__empty_n;
  wire fifo_C_drain_PE_4_8__read;
  wire [16:0] fifo_C_drain_PE_4_8__din;
  wire fifo_C_drain_PE_4_8__full_n;
  wire fifo_C_drain_PE_4_8__write;
  wire [16:0] fifo_C_drain_PE_4_9__dout;
  wire fifo_C_drain_PE_4_9__empty_n;
  wire fifo_C_drain_PE_4_9__read;
  wire [16:0] fifo_C_drain_PE_4_9__din;
  wire fifo_C_drain_PE_4_9__full_n;
  wire fifo_C_drain_PE_4_9__write;
  wire [16:0] fifo_C_drain_PE_5_0__dout;
  wire fifo_C_drain_PE_5_0__empty_n;
  wire fifo_C_drain_PE_5_0__read;
  wire [16:0] fifo_C_drain_PE_5_0__din;
  wire fifo_C_drain_PE_5_0__full_n;
  wire fifo_C_drain_PE_5_0__write;
  wire [16:0] fifo_C_drain_PE_5_1__dout;
  wire fifo_C_drain_PE_5_1__empty_n;
  wire fifo_C_drain_PE_5_1__read;
  wire [16:0] fifo_C_drain_PE_5_1__din;
  wire fifo_C_drain_PE_5_1__full_n;
  wire fifo_C_drain_PE_5_1__write;
  wire [16:0] fifo_C_drain_PE_5_10__dout;
  wire fifo_C_drain_PE_5_10__empty_n;
  wire fifo_C_drain_PE_5_10__read;
  wire [16:0] fifo_C_drain_PE_5_10__din;
  wire fifo_C_drain_PE_5_10__full_n;
  wire fifo_C_drain_PE_5_10__write;
  wire [16:0] fifo_C_drain_PE_5_11__dout;
  wire fifo_C_drain_PE_5_11__empty_n;
  wire fifo_C_drain_PE_5_11__read;
  wire [16:0] fifo_C_drain_PE_5_11__din;
  wire fifo_C_drain_PE_5_11__full_n;
  wire fifo_C_drain_PE_5_11__write;
  wire [16:0] fifo_C_drain_PE_5_12__dout;
  wire fifo_C_drain_PE_5_12__empty_n;
  wire fifo_C_drain_PE_5_12__read;
  wire [16:0] fifo_C_drain_PE_5_12__din;
  wire fifo_C_drain_PE_5_12__full_n;
  wire fifo_C_drain_PE_5_12__write;
  wire [16:0] fifo_C_drain_PE_5_13__dout;
  wire fifo_C_drain_PE_5_13__empty_n;
  wire fifo_C_drain_PE_5_13__read;
  wire [16:0] fifo_C_drain_PE_5_13__din;
  wire fifo_C_drain_PE_5_13__full_n;
  wire fifo_C_drain_PE_5_13__write;
  wire [16:0] fifo_C_drain_PE_5_14__dout;
  wire fifo_C_drain_PE_5_14__empty_n;
  wire fifo_C_drain_PE_5_14__read;
  wire [16:0] fifo_C_drain_PE_5_14__din;
  wire fifo_C_drain_PE_5_14__full_n;
  wire fifo_C_drain_PE_5_14__write;
  wire [16:0] fifo_C_drain_PE_5_15__dout;
  wire fifo_C_drain_PE_5_15__empty_n;
  wire fifo_C_drain_PE_5_15__read;
  wire [16:0] fifo_C_drain_PE_5_15__din;
  wire fifo_C_drain_PE_5_15__full_n;
  wire fifo_C_drain_PE_5_15__write;
  wire [16:0] fifo_C_drain_PE_5_16__dout;
  wire fifo_C_drain_PE_5_16__empty_n;
  wire fifo_C_drain_PE_5_16__read;
  wire [16:0] fifo_C_drain_PE_5_16__din;
  wire fifo_C_drain_PE_5_16__full_n;
  wire fifo_C_drain_PE_5_16__write;
  wire [16:0] fifo_C_drain_PE_5_2__dout;
  wire fifo_C_drain_PE_5_2__empty_n;
  wire fifo_C_drain_PE_5_2__read;
  wire [16:0] fifo_C_drain_PE_5_2__din;
  wire fifo_C_drain_PE_5_2__full_n;
  wire fifo_C_drain_PE_5_2__write;
  wire [16:0] fifo_C_drain_PE_5_3__dout;
  wire fifo_C_drain_PE_5_3__empty_n;
  wire fifo_C_drain_PE_5_3__read;
  wire [16:0] fifo_C_drain_PE_5_3__din;
  wire fifo_C_drain_PE_5_3__full_n;
  wire fifo_C_drain_PE_5_3__write;
  wire [16:0] fifo_C_drain_PE_5_4__dout;
  wire fifo_C_drain_PE_5_4__empty_n;
  wire fifo_C_drain_PE_5_4__read;
  wire [16:0] fifo_C_drain_PE_5_4__din;
  wire fifo_C_drain_PE_5_4__full_n;
  wire fifo_C_drain_PE_5_4__write;
  wire [16:0] fifo_C_drain_PE_5_5__dout;
  wire fifo_C_drain_PE_5_5__empty_n;
  wire fifo_C_drain_PE_5_5__read;
  wire [16:0] fifo_C_drain_PE_5_5__din;
  wire fifo_C_drain_PE_5_5__full_n;
  wire fifo_C_drain_PE_5_5__write;
  wire [16:0] fifo_C_drain_PE_5_6__dout;
  wire fifo_C_drain_PE_5_6__empty_n;
  wire fifo_C_drain_PE_5_6__read;
  wire [16:0] fifo_C_drain_PE_5_6__din;
  wire fifo_C_drain_PE_5_6__full_n;
  wire fifo_C_drain_PE_5_6__write;
  wire [16:0] fifo_C_drain_PE_5_7__dout;
  wire fifo_C_drain_PE_5_7__empty_n;
  wire fifo_C_drain_PE_5_7__read;
  wire [16:0] fifo_C_drain_PE_5_7__din;
  wire fifo_C_drain_PE_5_7__full_n;
  wire fifo_C_drain_PE_5_7__write;
  wire [16:0] fifo_C_drain_PE_5_8__dout;
  wire fifo_C_drain_PE_5_8__empty_n;
  wire fifo_C_drain_PE_5_8__read;
  wire [16:0] fifo_C_drain_PE_5_8__din;
  wire fifo_C_drain_PE_5_8__full_n;
  wire fifo_C_drain_PE_5_8__write;
  wire [16:0] fifo_C_drain_PE_5_9__dout;
  wire fifo_C_drain_PE_5_9__empty_n;
  wire fifo_C_drain_PE_5_9__read;
  wire [16:0] fifo_C_drain_PE_5_9__din;
  wire fifo_C_drain_PE_5_9__full_n;
  wire fifo_C_drain_PE_5_9__write;
  wire [16:0] fifo_C_drain_PE_6_0__dout;
  wire fifo_C_drain_PE_6_0__empty_n;
  wire fifo_C_drain_PE_6_0__read;
  wire [16:0] fifo_C_drain_PE_6_0__din;
  wire fifo_C_drain_PE_6_0__full_n;
  wire fifo_C_drain_PE_6_0__write;
  wire [16:0] fifo_C_drain_PE_6_1__dout;
  wire fifo_C_drain_PE_6_1__empty_n;
  wire fifo_C_drain_PE_6_1__read;
  wire [16:0] fifo_C_drain_PE_6_1__din;
  wire fifo_C_drain_PE_6_1__full_n;
  wire fifo_C_drain_PE_6_1__write;
  wire [16:0] fifo_C_drain_PE_6_10__dout;
  wire fifo_C_drain_PE_6_10__empty_n;
  wire fifo_C_drain_PE_6_10__read;
  wire [16:0] fifo_C_drain_PE_6_10__din;
  wire fifo_C_drain_PE_6_10__full_n;
  wire fifo_C_drain_PE_6_10__write;
  wire [16:0] fifo_C_drain_PE_6_11__dout;
  wire fifo_C_drain_PE_6_11__empty_n;
  wire fifo_C_drain_PE_6_11__read;
  wire [16:0] fifo_C_drain_PE_6_11__din;
  wire fifo_C_drain_PE_6_11__full_n;
  wire fifo_C_drain_PE_6_11__write;
  wire [16:0] fifo_C_drain_PE_6_12__dout;
  wire fifo_C_drain_PE_6_12__empty_n;
  wire fifo_C_drain_PE_6_12__read;
  wire [16:0] fifo_C_drain_PE_6_12__din;
  wire fifo_C_drain_PE_6_12__full_n;
  wire fifo_C_drain_PE_6_12__write;
  wire [16:0] fifo_C_drain_PE_6_13__dout;
  wire fifo_C_drain_PE_6_13__empty_n;
  wire fifo_C_drain_PE_6_13__read;
  wire [16:0] fifo_C_drain_PE_6_13__din;
  wire fifo_C_drain_PE_6_13__full_n;
  wire fifo_C_drain_PE_6_13__write;
  wire [16:0] fifo_C_drain_PE_6_14__dout;
  wire fifo_C_drain_PE_6_14__empty_n;
  wire fifo_C_drain_PE_6_14__read;
  wire [16:0] fifo_C_drain_PE_6_14__din;
  wire fifo_C_drain_PE_6_14__full_n;
  wire fifo_C_drain_PE_6_14__write;
  wire [16:0] fifo_C_drain_PE_6_15__dout;
  wire fifo_C_drain_PE_6_15__empty_n;
  wire fifo_C_drain_PE_6_15__read;
  wire [16:0] fifo_C_drain_PE_6_15__din;
  wire fifo_C_drain_PE_6_15__full_n;
  wire fifo_C_drain_PE_6_15__write;
  wire [16:0] fifo_C_drain_PE_6_16__dout;
  wire fifo_C_drain_PE_6_16__empty_n;
  wire fifo_C_drain_PE_6_16__read;
  wire [16:0] fifo_C_drain_PE_6_16__din;
  wire fifo_C_drain_PE_6_16__full_n;
  wire fifo_C_drain_PE_6_16__write;
  wire [16:0] fifo_C_drain_PE_6_2__dout;
  wire fifo_C_drain_PE_6_2__empty_n;
  wire fifo_C_drain_PE_6_2__read;
  wire [16:0] fifo_C_drain_PE_6_2__din;
  wire fifo_C_drain_PE_6_2__full_n;
  wire fifo_C_drain_PE_6_2__write;
  wire [16:0] fifo_C_drain_PE_6_3__dout;
  wire fifo_C_drain_PE_6_3__empty_n;
  wire fifo_C_drain_PE_6_3__read;
  wire [16:0] fifo_C_drain_PE_6_3__din;
  wire fifo_C_drain_PE_6_3__full_n;
  wire fifo_C_drain_PE_6_3__write;
  wire [16:0] fifo_C_drain_PE_6_4__dout;
  wire fifo_C_drain_PE_6_4__empty_n;
  wire fifo_C_drain_PE_6_4__read;
  wire [16:0] fifo_C_drain_PE_6_4__din;
  wire fifo_C_drain_PE_6_4__full_n;
  wire fifo_C_drain_PE_6_4__write;
  wire [16:0] fifo_C_drain_PE_6_5__dout;
  wire fifo_C_drain_PE_6_5__empty_n;
  wire fifo_C_drain_PE_6_5__read;
  wire [16:0] fifo_C_drain_PE_6_5__din;
  wire fifo_C_drain_PE_6_5__full_n;
  wire fifo_C_drain_PE_6_5__write;
  wire [16:0] fifo_C_drain_PE_6_6__dout;
  wire fifo_C_drain_PE_6_6__empty_n;
  wire fifo_C_drain_PE_6_6__read;
  wire [16:0] fifo_C_drain_PE_6_6__din;
  wire fifo_C_drain_PE_6_6__full_n;
  wire fifo_C_drain_PE_6_6__write;
  wire [16:0] fifo_C_drain_PE_6_7__dout;
  wire fifo_C_drain_PE_6_7__empty_n;
  wire fifo_C_drain_PE_6_7__read;
  wire [16:0] fifo_C_drain_PE_6_7__din;
  wire fifo_C_drain_PE_6_7__full_n;
  wire fifo_C_drain_PE_6_7__write;
  wire [16:0] fifo_C_drain_PE_6_8__dout;
  wire fifo_C_drain_PE_6_8__empty_n;
  wire fifo_C_drain_PE_6_8__read;
  wire [16:0] fifo_C_drain_PE_6_8__din;
  wire fifo_C_drain_PE_6_8__full_n;
  wire fifo_C_drain_PE_6_8__write;
  wire [16:0] fifo_C_drain_PE_6_9__dout;
  wire fifo_C_drain_PE_6_9__empty_n;
  wire fifo_C_drain_PE_6_9__read;
  wire [16:0] fifo_C_drain_PE_6_9__din;
  wire fifo_C_drain_PE_6_9__full_n;
  wire fifo_C_drain_PE_6_9__write;
  wire [16:0] fifo_C_drain_PE_7_0__dout;
  wire fifo_C_drain_PE_7_0__empty_n;
  wire fifo_C_drain_PE_7_0__read;
  wire [16:0] fifo_C_drain_PE_7_0__din;
  wire fifo_C_drain_PE_7_0__full_n;
  wire fifo_C_drain_PE_7_0__write;
  wire [16:0] fifo_C_drain_PE_7_1__dout;
  wire fifo_C_drain_PE_7_1__empty_n;
  wire fifo_C_drain_PE_7_1__read;
  wire [16:0] fifo_C_drain_PE_7_1__din;
  wire fifo_C_drain_PE_7_1__full_n;
  wire fifo_C_drain_PE_7_1__write;
  wire [16:0] fifo_C_drain_PE_7_10__dout;
  wire fifo_C_drain_PE_7_10__empty_n;
  wire fifo_C_drain_PE_7_10__read;
  wire [16:0] fifo_C_drain_PE_7_10__din;
  wire fifo_C_drain_PE_7_10__full_n;
  wire fifo_C_drain_PE_7_10__write;
  wire [16:0] fifo_C_drain_PE_7_11__dout;
  wire fifo_C_drain_PE_7_11__empty_n;
  wire fifo_C_drain_PE_7_11__read;
  wire [16:0] fifo_C_drain_PE_7_11__din;
  wire fifo_C_drain_PE_7_11__full_n;
  wire fifo_C_drain_PE_7_11__write;
  wire [16:0] fifo_C_drain_PE_7_12__dout;
  wire fifo_C_drain_PE_7_12__empty_n;
  wire fifo_C_drain_PE_7_12__read;
  wire [16:0] fifo_C_drain_PE_7_12__din;
  wire fifo_C_drain_PE_7_12__full_n;
  wire fifo_C_drain_PE_7_12__write;
  wire [16:0] fifo_C_drain_PE_7_13__dout;
  wire fifo_C_drain_PE_7_13__empty_n;
  wire fifo_C_drain_PE_7_13__read;
  wire [16:0] fifo_C_drain_PE_7_13__din;
  wire fifo_C_drain_PE_7_13__full_n;
  wire fifo_C_drain_PE_7_13__write;
  wire [16:0] fifo_C_drain_PE_7_14__dout;
  wire fifo_C_drain_PE_7_14__empty_n;
  wire fifo_C_drain_PE_7_14__read;
  wire [16:0] fifo_C_drain_PE_7_14__din;
  wire fifo_C_drain_PE_7_14__full_n;
  wire fifo_C_drain_PE_7_14__write;
  wire [16:0] fifo_C_drain_PE_7_15__dout;
  wire fifo_C_drain_PE_7_15__empty_n;
  wire fifo_C_drain_PE_7_15__read;
  wire [16:0] fifo_C_drain_PE_7_15__din;
  wire fifo_C_drain_PE_7_15__full_n;
  wire fifo_C_drain_PE_7_15__write;
  wire [16:0] fifo_C_drain_PE_7_16__dout;
  wire fifo_C_drain_PE_7_16__empty_n;
  wire fifo_C_drain_PE_7_16__read;
  wire [16:0] fifo_C_drain_PE_7_16__din;
  wire fifo_C_drain_PE_7_16__full_n;
  wire fifo_C_drain_PE_7_16__write;
  wire [16:0] fifo_C_drain_PE_7_2__dout;
  wire fifo_C_drain_PE_7_2__empty_n;
  wire fifo_C_drain_PE_7_2__read;
  wire [16:0] fifo_C_drain_PE_7_2__din;
  wire fifo_C_drain_PE_7_2__full_n;
  wire fifo_C_drain_PE_7_2__write;
  wire [16:0] fifo_C_drain_PE_7_3__dout;
  wire fifo_C_drain_PE_7_3__empty_n;
  wire fifo_C_drain_PE_7_3__read;
  wire [16:0] fifo_C_drain_PE_7_3__din;
  wire fifo_C_drain_PE_7_3__full_n;
  wire fifo_C_drain_PE_7_3__write;
  wire [16:0] fifo_C_drain_PE_7_4__dout;
  wire fifo_C_drain_PE_7_4__empty_n;
  wire fifo_C_drain_PE_7_4__read;
  wire [16:0] fifo_C_drain_PE_7_4__din;
  wire fifo_C_drain_PE_7_4__full_n;
  wire fifo_C_drain_PE_7_4__write;
  wire [16:0] fifo_C_drain_PE_7_5__dout;
  wire fifo_C_drain_PE_7_5__empty_n;
  wire fifo_C_drain_PE_7_5__read;
  wire [16:0] fifo_C_drain_PE_7_5__din;
  wire fifo_C_drain_PE_7_5__full_n;
  wire fifo_C_drain_PE_7_5__write;
  wire [16:0] fifo_C_drain_PE_7_6__dout;
  wire fifo_C_drain_PE_7_6__empty_n;
  wire fifo_C_drain_PE_7_6__read;
  wire [16:0] fifo_C_drain_PE_7_6__din;
  wire fifo_C_drain_PE_7_6__full_n;
  wire fifo_C_drain_PE_7_6__write;
  wire [16:0] fifo_C_drain_PE_7_7__dout;
  wire fifo_C_drain_PE_7_7__empty_n;
  wire fifo_C_drain_PE_7_7__read;
  wire [16:0] fifo_C_drain_PE_7_7__din;
  wire fifo_C_drain_PE_7_7__full_n;
  wire fifo_C_drain_PE_7_7__write;
  wire [16:0] fifo_C_drain_PE_7_8__dout;
  wire fifo_C_drain_PE_7_8__empty_n;
  wire fifo_C_drain_PE_7_8__read;
  wire [16:0] fifo_C_drain_PE_7_8__din;
  wire fifo_C_drain_PE_7_8__full_n;
  wire fifo_C_drain_PE_7_8__write;
  wire [16:0] fifo_C_drain_PE_7_9__dout;
  wire fifo_C_drain_PE_7_9__empty_n;
  wire fifo_C_drain_PE_7_9__read;
  wire [16:0] fifo_C_drain_PE_7_9__din;
  wire fifo_C_drain_PE_7_9__full_n;
  wire fifo_C_drain_PE_7_9__write;
  wire [16:0] fifo_C_drain_PE_8_0__dout;
  wire fifo_C_drain_PE_8_0__empty_n;
  wire fifo_C_drain_PE_8_0__read;
  wire [16:0] fifo_C_drain_PE_8_0__din;
  wire fifo_C_drain_PE_8_0__full_n;
  wire fifo_C_drain_PE_8_0__write;
  wire [16:0] fifo_C_drain_PE_8_1__dout;
  wire fifo_C_drain_PE_8_1__empty_n;
  wire fifo_C_drain_PE_8_1__read;
  wire [16:0] fifo_C_drain_PE_8_1__din;
  wire fifo_C_drain_PE_8_1__full_n;
  wire fifo_C_drain_PE_8_1__write;
  wire [16:0] fifo_C_drain_PE_8_10__dout;
  wire fifo_C_drain_PE_8_10__empty_n;
  wire fifo_C_drain_PE_8_10__read;
  wire [16:0] fifo_C_drain_PE_8_10__din;
  wire fifo_C_drain_PE_8_10__full_n;
  wire fifo_C_drain_PE_8_10__write;
  wire [16:0] fifo_C_drain_PE_8_11__dout;
  wire fifo_C_drain_PE_8_11__empty_n;
  wire fifo_C_drain_PE_8_11__read;
  wire [16:0] fifo_C_drain_PE_8_11__din;
  wire fifo_C_drain_PE_8_11__full_n;
  wire fifo_C_drain_PE_8_11__write;
  wire [16:0] fifo_C_drain_PE_8_12__dout;
  wire fifo_C_drain_PE_8_12__empty_n;
  wire fifo_C_drain_PE_8_12__read;
  wire [16:0] fifo_C_drain_PE_8_12__din;
  wire fifo_C_drain_PE_8_12__full_n;
  wire fifo_C_drain_PE_8_12__write;
  wire [16:0] fifo_C_drain_PE_8_13__dout;
  wire fifo_C_drain_PE_8_13__empty_n;
  wire fifo_C_drain_PE_8_13__read;
  wire [16:0] fifo_C_drain_PE_8_13__din;
  wire fifo_C_drain_PE_8_13__full_n;
  wire fifo_C_drain_PE_8_13__write;
  wire [16:0] fifo_C_drain_PE_8_14__dout;
  wire fifo_C_drain_PE_8_14__empty_n;
  wire fifo_C_drain_PE_8_14__read;
  wire [16:0] fifo_C_drain_PE_8_14__din;
  wire fifo_C_drain_PE_8_14__full_n;
  wire fifo_C_drain_PE_8_14__write;
  wire [16:0] fifo_C_drain_PE_8_15__dout;
  wire fifo_C_drain_PE_8_15__empty_n;
  wire fifo_C_drain_PE_8_15__read;
  wire [16:0] fifo_C_drain_PE_8_15__din;
  wire fifo_C_drain_PE_8_15__full_n;
  wire fifo_C_drain_PE_8_15__write;
  wire [16:0] fifo_C_drain_PE_8_16__dout;
  wire fifo_C_drain_PE_8_16__empty_n;
  wire fifo_C_drain_PE_8_16__read;
  wire [16:0] fifo_C_drain_PE_8_16__din;
  wire fifo_C_drain_PE_8_16__full_n;
  wire fifo_C_drain_PE_8_16__write;
  wire [16:0] fifo_C_drain_PE_8_2__dout;
  wire fifo_C_drain_PE_8_2__empty_n;
  wire fifo_C_drain_PE_8_2__read;
  wire [16:0] fifo_C_drain_PE_8_2__din;
  wire fifo_C_drain_PE_8_2__full_n;
  wire fifo_C_drain_PE_8_2__write;
  wire [16:0] fifo_C_drain_PE_8_3__dout;
  wire fifo_C_drain_PE_8_3__empty_n;
  wire fifo_C_drain_PE_8_3__read;
  wire [16:0] fifo_C_drain_PE_8_3__din;
  wire fifo_C_drain_PE_8_3__full_n;
  wire fifo_C_drain_PE_8_3__write;
  wire [16:0] fifo_C_drain_PE_8_4__dout;
  wire fifo_C_drain_PE_8_4__empty_n;
  wire fifo_C_drain_PE_8_4__read;
  wire [16:0] fifo_C_drain_PE_8_4__din;
  wire fifo_C_drain_PE_8_4__full_n;
  wire fifo_C_drain_PE_8_4__write;
  wire [16:0] fifo_C_drain_PE_8_5__dout;
  wire fifo_C_drain_PE_8_5__empty_n;
  wire fifo_C_drain_PE_8_5__read;
  wire [16:0] fifo_C_drain_PE_8_5__din;
  wire fifo_C_drain_PE_8_5__full_n;
  wire fifo_C_drain_PE_8_5__write;
  wire [16:0] fifo_C_drain_PE_8_6__dout;
  wire fifo_C_drain_PE_8_6__empty_n;
  wire fifo_C_drain_PE_8_6__read;
  wire [16:0] fifo_C_drain_PE_8_6__din;
  wire fifo_C_drain_PE_8_6__full_n;
  wire fifo_C_drain_PE_8_6__write;
  wire [16:0] fifo_C_drain_PE_8_7__dout;
  wire fifo_C_drain_PE_8_7__empty_n;
  wire fifo_C_drain_PE_8_7__read;
  wire [16:0] fifo_C_drain_PE_8_7__din;
  wire fifo_C_drain_PE_8_7__full_n;
  wire fifo_C_drain_PE_8_7__write;
  wire [16:0] fifo_C_drain_PE_8_8__dout;
  wire fifo_C_drain_PE_8_8__empty_n;
  wire fifo_C_drain_PE_8_8__read;
  wire [16:0] fifo_C_drain_PE_8_8__din;
  wire fifo_C_drain_PE_8_8__full_n;
  wire fifo_C_drain_PE_8_8__write;
  wire [16:0] fifo_C_drain_PE_8_9__dout;
  wire fifo_C_drain_PE_8_9__empty_n;
  wire fifo_C_drain_PE_8_9__read;
  wire [16:0] fifo_C_drain_PE_8_9__din;
  wire fifo_C_drain_PE_8_9__full_n;
  wire fifo_C_drain_PE_8_9__write;
  wire [16:0] fifo_C_drain_PE_9_0__dout;
  wire fifo_C_drain_PE_9_0__empty_n;
  wire fifo_C_drain_PE_9_0__read;
  wire [16:0] fifo_C_drain_PE_9_0__din;
  wire fifo_C_drain_PE_9_0__full_n;
  wire fifo_C_drain_PE_9_0__write;
  wire [16:0] fifo_C_drain_PE_9_1__dout;
  wire fifo_C_drain_PE_9_1__empty_n;
  wire fifo_C_drain_PE_9_1__read;
  wire [16:0] fifo_C_drain_PE_9_1__din;
  wire fifo_C_drain_PE_9_1__full_n;
  wire fifo_C_drain_PE_9_1__write;
  wire [16:0] fifo_C_drain_PE_9_10__dout;
  wire fifo_C_drain_PE_9_10__empty_n;
  wire fifo_C_drain_PE_9_10__read;
  wire [16:0] fifo_C_drain_PE_9_10__din;
  wire fifo_C_drain_PE_9_10__full_n;
  wire fifo_C_drain_PE_9_10__write;
  wire [16:0] fifo_C_drain_PE_9_11__dout;
  wire fifo_C_drain_PE_9_11__empty_n;
  wire fifo_C_drain_PE_9_11__read;
  wire [16:0] fifo_C_drain_PE_9_11__din;
  wire fifo_C_drain_PE_9_11__full_n;
  wire fifo_C_drain_PE_9_11__write;
  wire [16:0] fifo_C_drain_PE_9_12__dout;
  wire fifo_C_drain_PE_9_12__empty_n;
  wire fifo_C_drain_PE_9_12__read;
  wire [16:0] fifo_C_drain_PE_9_12__din;
  wire fifo_C_drain_PE_9_12__full_n;
  wire fifo_C_drain_PE_9_12__write;
  wire [16:0] fifo_C_drain_PE_9_13__dout;
  wire fifo_C_drain_PE_9_13__empty_n;
  wire fifo_C_drain_PE_9_13__read;
  wire [16:0] fifo_C_drain_PE_9_13__din;
  wire fifo_C_drain_PE_9_13__full_n;
  wire fifo_C_drain_PE_9_13__write;
  wire [16:0] fifo_C_drain_PE_9_14__dout;
  wire fifo_C_drain_PE_9_14__empty_n;
  wire fifo_C_drain_PE_9_14__read;
  wire [16:0] fifo_C_drain_PE_9_14__din;
  wire fifo_C_drain_PE_9_14__full_n;
  wire fifo_C_drain_PE_9_14__write;
  wire [16:0] fifo_C_drain_PE_9_15__dout;
  wire fifo_C_drain_PE_9_15__empty_n;
  wire fifo_C_drain_PE_9_15__read;
  wire [16:0] fifo_C_drain_PE_9_15__din;
  wire fifo_C_drain_PE_9_15__full_n;
  wire fifo_C_drain_PE_9_15__write;
  wire [16:0] fifo_C_drain_PE_9_16__dout;
  wire fifo_C_drain_PE_9_16__empty_n;
  wire fifo_C_drain_PE_9_16__read;
  wire [16:0] fifo_C_drain_PE_9_16__din;
  wire fifo_C_drain_PE_9_16__full_n;
  wire fifo_C_drain_PE_9_16__write;
  wire [16:0] fifo_C_drain_PE_9_2__dout;
  wire fifo_C_drain_PE_9_2__empty_n;
  wire fifo_C_drain_PE_9_2__read;
  wire [16:0] fifo_C_drain_PE_9_2__din;
  wire fifo_C_drain_PE_9_2__full_n;
  wire fifo_C_drain_PE_9_2__write;
  wire [16:0] fifo_C_drain_PE_9_3__dout;
  wire fifo_C_drain_PE_9_3__empty_n;
  wire fifo_C_drain_PE_9_3__read;
  wire [16:0] fifo_C_drain_PE_9_3__din;
  wire fifo_C_drain_PE_9_3__full_n;
  wire fifo_C_drain_PE_9_3__write;
  wire [16:0] fifo_C_drain_PE_9_4__dout;
  wire fifo_C_drain_PE_9_4__empty_n;
  wire fifo_C_drain_PE_9_4__read;
  wire [16:0] fifo_C_drain_PE_9_4__din;
  wire fifo_C_drain_PE_9_4__full_n;
  wire fifo_C_drain_PE_9_4__write;
  wire [16:0] fifo_C_drain_PE_9_5__dout;
  wire fifo_C_drain_PE_9_5__empty_n;
  wire fifo_C_drain_PE_9_5__read;
  wire [16:0] fifo_C_drain_PE_9_5__din;
  wire fifo_C_drain_PE_9_5__full_n;
  wire fifo_C_drain_PE_9_5__write;
  wire [16:0] fifo_C_drain_PE_9_6__dout;
  wire fifo_C_drain_PE_9_6__empty_n;
  wire fifo_C_drain_PE_9_6__read;
  wire [16:0] fifo_C_drain_PE_9_6__din;
  wire fifo_C_drain_PE_9_6__full_n;
  wire fifo_C_drain_PE_9_6__write;
  wire [16:0] fifo_C_drain_PE_9_7__dout;
  wire fifo_C_drain_PE_9_7__empty_n;
  wire fifo_C_drain_PE_9_7__read;
  wire [16:0] fifo_C_drain_PE_9_7__din;
  wire fifo_C_drain_PE_9_7__full_n;
  wire fifo_C_drain_PE_9_7__write;
  wire [16:0] fifo_C_drain_PE_9_8__dout;
  wire fifo_C_drain_PE_9_8__empty_n;
  wire fifo_C_drain_PE_9_8__read;
  wire [16:0] fifo_C_drain_PE_9_8__din;
  wire fifo_C_drain_PE_9_8__full_n;
  wire fifo_C_drain_PE_9_8__write;
  wire [16:0] fifo_C_drain_PE_9_9__dout;
  wire fifo_C_drain_PE_9_9__empty_n;
  wire fifo_C_drain_PE_9_9__read;
  wire [16:0] fifo_C_drain_PE_9_9__din;
  wire fifo_C_drain_PE_9_9__full_n;
  wire fifo_C_drain_PE_9_9__write;
  wire A_IO_L2_in_0__ap_start;
  wire A_IO_L2_in_0__ap_ready;
  wire A_IO_L2_in_0__ap_done;
  wire A_IO_L2_in_0__ap_idle;
  wire A_IO_L2_in_1__ap_start;
  wire A_IO_L2_in_1__ap_ready;
  wire A_IO_L2_in_1__ap_done;
  wire A_IO_L2_in_1__ap_idle;
  wire A_IO_L2_in_2__ap_start;
  wire A_IO_L2_in_2__ap_ready;
  wire A_IO_L2_in_2__ap_done;
  wire A_IO_L2_in_2__ap_idle;
  wire A_IO_L2_in_3__ap_start;
  wire A_IO_L2_in_3__ap_ready;
  wire A_IO_L2_in_3__ap_done;
  wire A_IO_L2_in_3__ap_idle;
  wire A_IO_L2_in_4__ap_start;
  wire A_IO_L2_in_4__ap_ready;
  wire A_IO_L2_in_4__ap_done;
  wire A_IO_L2_in_4__ap_idle;
  wire A_IO_L2_in_5__ap_start;
  wire A_IO_L2_in_5__ap_ready;
  wire A_IO_L2_in_5__ap_done;
  wire A_IO_L2_in_5__ap_idle;
  wire A_IO_L2_in_6__ap_start;
  wire A_IO_L2_in_6__ap_ready;
  wire A_IO_L2_in_6__ap_done;
  wire A_IO_L2_in_6__ap_idle;
  wire A_IO_L2_in_7__ap_start;
  wire A_IO_L2_in_7__ap_ready;
  wire A_IO_L2_in_7__ap_done;
  wire A_IO_L2_in_7__ap_idle;
  wire A_IO_L2_in_8__ap_start;
  wire A_IO_L2_in_8__ap_ready;
  wire A_IO_L2_in_8__ap_done;
  wire A_IO_L2_in_8__ap_idle;
  wire A_IO_L2_in_9__ap_start;
  wire A_IO_L2_in_9__ap_ready;
  wire A_IO_L2_in_9__ap_done;
  wire A_IO_L2_in_9__ap_idle;
  wire A_IO_L2_in_10__ap_start;
  wire A_IO_L2_in_10__ap_ready;
  wire A_IO_L2_in_10__ap_done;
  wire A_IO_L2_in_10__ap_idle;
  wire A_IO_L2_in_11__ap_start;
  wire A_IO_L2_in_11__ap_ready;
  wire A_IO_L2_in_11__ap_done;
  wire A_IO_L2_in_11__ap_idle;
  wire A_IO_L2_in_12__ap_start;
  wire A_IO_L2_in_12__ap_ready;
  wire A_IO_L2_in_12__ap_done;
  wire A_IO_L2_in_12__ap_idle;
  wire A_IO_L2_in_13__ap_start;
  wire A_IO_L2_in_13__ap_ready;
  wire A_IO_L2_in_13__ap_done;
  wire A_IO_L2_in_13__ap_idle;
  wire A_IO_L2_in_14__ap_start;
  wire A_IO_L2_in_14__ap_ready;
  wire A_IO_L2_in_14__ap_done;
  wire A_IO_L2_in_14__ap_idle;
  wire A_IO_L2_in_15__ap_start;
  wire A_IO_L2_in_15__ap_ready;
  wire A_IO_L2_in_15__ap_done;
  wire A_IO_L2_in_15__ap_idle;
  wire A_IO_L2_in_16__ap_start;
  wire A_IO_L2_in_16__ap_ready;
  wire A_IO_L2_in_16__ap_done;
  wire A_IO_L2_in_16__ap_idle;
  wire A_IO_L2_in_boundary_0__ap_start;
  wire A_IO_L2_in_boundary_0__ap_ready;
  wire A_IO_L2_in_boundary_0__ap_done;
  wire A_IO_L2_in_boundary_0__ap_idle;
  wire A_IO_L3_in_0__ap_start;
  wire A_IO_L3_in_0__ap_ready;
  wire A_IO_L3_in_0__ap_done;
  wire A_IO_L3_in_0__ap_idle;
  wire [63:0] A_IO_L3_in_serialize_0___A__q0;
  wire A_IO_L3_in_serialize_0__ap_start;
  wire A_IO_L3_in_serialize_0__ap_ready;
  wire A_IO_L3_in_serialize_0__ap_done;
  wire A_IO_L3_in_serialize_0__ap_idle;
  wire A_PE_dummy_in_0__ap_start;
  wire A_PE_dummy_in_0__ap_ready;
  wire A_PE_dummy_in_0__ap_done;
  wire A_PE_dummy_in_0__ap_idle;
  wire A_PE_dummy_in_1__ap_start;
  wire A_PE_dummy_in_1__ap_ready;
  wire A_PE_dummy_in_1__ap_done;
  wire A_PE_dummy_in_1__ap_idle;
  wire A_PE_dummy_in_2__ap_start;
  wire A_PE_dummy_in_2__ap_ready;
  wire A_PE_dummy_in_2__ap_done;
  wire A_PE_dummy_in_2__ap_idle;
  wire A_PE_dummy_in_3__ap_start;
  wire A_PE_dummy_in_3__ap_ready;
  wire A_PE_dummy_in_3__ap_done;
  wire A_PE_dummy_in_3__ap_idle;
  wire A_PE_dummy_in_4__ap_start;
  wire A_PE_dummy_in_4__ap_ready;
  wire A_PE_dummy_in_4__ap_done;
  wire A_PE_dummy_in_4__ap_idle;
  wire A_PE_dummy_in_5__ap_start;
  wire A_PE_dummy_in_5__ap_ready;
  wire A_PE_dummy_in_5__ap_done;
  wire A_PE_dummy_in_5__ap_idle;
  wire A_PE_dummy_in_6__ap_start;
  wire A_PE_dummy_in_6__ap_ready;
  wire A_PE_dummy_in_6__ap_done;
  wire A_PE_dummy_in_6__ap_idle;
  wire A_PE_dummy_in_7__ap_start;
  wire A_PE_dummy_in_7__ap_ready;
  wire A_PE_dummy_in_7__ap_done;
  wire A_PE_dummy_in_7__ap_idle;
  wire A_PE_dummy_in_8__ap_start;
  wire A_PE_dummy_in_8__ap_ready;
  wire A_PE_dummy_in_8__ap_done;
  wire A_PE_dummy_in_8__ap_idle;
  wire A_PE_dummy_in_9__ap_start;
  wire A_PE_dummy_in_9__ap_ready;
  wire A_PE_dummy_in_9__ap_done;
  wire A_PE_dummy_in_9__ap_idle;
  wire A_PE_dummy_in_10__ap_start;
  wire A_PE_dummy_in_10__ap_ready;
  wire A_PE_dummy_in_10__ap_done;
  wire A_PE_dummy_in_10__ap_idle;
  wire A_PE_dummy_in_11__ap_start;
  wire A_PE_dummy_in_11__ap_ready;
  wire A_PE_dummy_in_11__ap_done;
  wire A_PE_dummy_in_11__ap_idle;
  wire A_PE_dummy_in_12__ap_start;
  wire A_PE_dummy_in_12__ap_ready;
  wire A_PE_dummy_in_12__ap_done;
  wire A_PE_dummy_in_12__ap_idle;
  wire A_PE_dummy_in_13__ap_start;
  wire A_PE_dummy_in_13__ap_ready;
  wire A_PE_dummy_in_13__ap_done;
  wire A_PE_dummy_in_13__ap_idle;
  wire A_PE_dummy_in_14__ap_start;
  wire A_PE_dummy_in_14__ap_ready;
  wire A_PE_dummy_in_14__ap_done;
  wire A_PE_dummy_in_14__ap_idle;
  wire A_PE_dummy_in_15__ap_start;
  wire A_PE_dummy_in_15__ap_ready;
  wire A_PE_dummy_in_15__ap_done;
  wire A_PE_dummy_in_15__ap_idle;
  wire A_PE_dummy_in_16__ap_start;
  wire A_PE_dummy_in_16__ap_ready;
  wire A_PE_dummy_in_16__ap_done;
  wire A_PE_dummy_in_16__ap_idle;
  wire A_PE_dummy_in_17__ap_start;
  wire A_PE_dummy_in_17__ap_ready;
  wire A_PE_dummy_in_17__ap_done;
  wire A_PE_dummy_in_17__ap_idle;
  wire B_IO_L2_in_0__ap_start;
  wire B_IO_L2_in_0__ap_ready;
  wire B_IO_L2_in_0__ap_done;
  wire B_IO_L2_in_0__ap_idle;
  wire B_IO_L2_in_1__ap_start;
  wire B_IO_L2_in_1__ap_ready;
  wire B_IO_L2_in_1__ap_done;
  wire B_IO_L2_in_1__ap_idle;
  wire B_IO_L2_in_2__ap_start;
  wire B_IO_L2_in_2__ap_ready;
  wire B_IO_L2_in_2__ap_done;
  wire B_IO_L2_in_2__ap_idle;
  wire B_IO_L2_in_3__ap_start;
  wire B_IO_L2_in_3__ap_ready;
  wire B_IO_L2_in_3__ap_done;
  wire B_IO_L2_in_3__ap_idle;
  wire B_IO_L2_in_4__ap_start;
  wire B_IO_L2_in_4__ap_ready;
  wire B_IO_L2_in_4__ap_done;
  wire B_IO_L2_in_4__ap_idle;
  wire B_IO_L2_in_5__ap_start;
  wire B_IO_L2_in_5__ap_ready;
  wire B_IO_L2_in_5__ap_done;
  wire B_IO_L2_in_5__ap_idle;
  wire B_IO_L2_in_6__ap_start;
  wire B_IO_L2_in_6__ap_ready;
  wire B_IO_L2_in_6__ap_done;
  wire B_IO_L2_in_6__ap_idle;
  wire B_IO_L2_in_7__ap_start;
  wire B_IO_L2_in_7__ap_ready;
  wire B_IO_L2_in_7__ap_done;
  wire B_IO_L2_in_7__ap_idle;
  wire B_IO_L2_in_8__ap_start;
  wire B_IO_L2_in_8__ap_ready;
  wire B_IO_L2_in_8__ap_done;
  wire B_IO_L2_in_8__ap_idle;
  wire B_IO_L2_in_9__ap_start;
  wire B_IO_L2_in_9__ap_ready;
  wire B_IO_L2_in_9__ap_done;
  wire B_IO_L2_in_9__ap_idle;
  wire B_IO_L2_in_10__ap_start;
  wire B_IO_L2_in_10__ap_ready;
  wire B_IO_L2_in_10__ap_done;
  wire B_IO_L2_in_10__ap_idle;
  wire B_IO_L2_in_11__ap_start;
  wire B_IO_L2_in_11__ap_ready;
  wire B_IO_L2_in_11__ap_done;
  wire B_IO_L2_in_11__ap_idle;
  wire B_IO_L2_in_12__ap_start;
  wire B_IO_L2_in_12__ap_ready;
  wire B_IO_L2_in_12__ap_done;
  wire B_IO_L2_in_12__ap_idle;
  wire B_IO_L2_in_13__ap_start;
  wire B_IO_L2_in_13__ap_ready;
  wire B_IO_L2_in_13__ap_done;
  wire B_IO_L2_in_13__ap_idle;
  wire B_IO_L2_in_14__ap_start;
  wire B_IO_L2_in_14__ap_ready;
  wire B_IO_L2_in_14__ap_done;
  wire B_IO_L2_in_14__ap_idle;
  wire B_IO_L2_in_15__ap_start;
  wire B_IO_L2_in_15__ap_ready;
  wire B_IO_L2_in_15__ap_done;
  wire B_IO_L2_in_15__ap_idle;
  wire B_IO_L2_in_boundary_0__ap_start;
  wire B_IO_L2_in_boundary_0__ap_ready;
  wire B_IO_L2_in_boundary_0__ap_done;
  wire B_IO_L2_in_boundary_0__ap_idle;
  wire B_IO_L3_in_0__ap_start;
  wire B_IO_L3_in_0__ap_ready;
  wire B_IO_L3_in_0__ap_done;
  wire B_IO_L3_in_0__ap_idle;
  wire [63:0] B_IO_L3_in_serialize_0___B__q0;
  wire B_IO_L3_in_serialize_0__ap_start;
  wire B_IO_L3_in_serialize_0__ap_ready;
  wire B_IO_L3_in_serialize_0__ap_done;
  wire B_IO_L3_in_serialize_0__ap_idle;
  wire B_PE_dummy_in_0__ap_start;
  wire B_PE_dummy_in_0__ap_ready;
  wire B_PE_dummy_in_0__ap_done;
  wire B_PE_dummy_in_0__ap_idle;
  wire B_PE_dummy_in_1__ap_start;
  wire B_PE_dummy_in_1__ap_ready;
  wire B_PE_dummy_in_1__ap_done;
  wire B_PE_dummy_in_1__ap_idle;
  wire B_PE_dummy_in_2__ap_start;
  wire B_PE_dummy_in_2__ap_ready;
  wire B_PE_dummy_in_2__ap_done;
  wire B_PE_dummy_in_2__ap_idle;
  wire B_PE_dummy_in_3__ap_start;
  wire B_PE_dummy_in_3__ap_ready;
  wire B_PE_dummy_in_3__ap_done;
  wire B_PE_dummy_in_3__ap_idle;
  wire B_PE_dummy_in_4__ap_start;
  wire B_PE_dummy_in_4__ap_ready;
  wire B_PE_dummy_in_4__ap_done;
  wire B_PE_dummy_in_4__ap_idle;
  wire B_PE_dummy_in_5__ap_start;
  wire B_PE_dummy_in_5__ap_ready;
  wire B_PE_dummy_in_5__ap_done;
  wire B_PE_dummy_in_5__ap_idle;
  wire B_PE_dummy_in_6__ap_start;
  wire B_PE_dummy_in_6__ap_ready;
  wire B_PE_dummy_in_6__ap_done;
  wire B_PE_dummy_in_6__ap_idle;
  wire B_PE_dummy_in_7__ap_start;
  wire B_PE_dummy_in_7__ap_ready;
  wire B_PE_dummy_in_7__ap_done;
  wire B_PE_dummy_in_7__ap_idle;
  wire B_PE_dummy_in_8__ap_start;
  wire B_PE_dummy_in_8__ap_ready;
  wire B_PE_dummy_in_8__ap_done;
  wire B_PE_dummy_in_8__ap_idle;
  wire B_PE_dummy_in_9__ap_start;
  wire B_PE_dummy_in_9__ap_ready;
  wire B_PE_dummy_in_9__ap_done;
  wire B_PE_dummy_in_9__ap_idle;
  wire B_PE_dummy_in_10__ap_start;
  wire B_PE_dummy_in_10__ap_ready;
  wire B_PE_dummy_in_10__ap_done;
  wire B_PE_dummy_in_10__ap_idle;
  wire B_PE_dummy_in_11__ap_start;
  wire B_PE_dummy_in_11__ap_ready;
  wire B_PE_dummy_in_11__ap_done;
  wire B_PE_dummy_in_11__ap_idle;
  wire B_PE_dummy_in_12__ap_start;
  wire B_PE_dummy_in_12__ap_ready;
  wire B_PE_dummy_in_12__ap_done;
  wire B_PE_dummy_in_12__ap_idle;
  wire B_PE_dummy_in_13__ap_start;
  wire B_PE_dummy_in_13__ap_ready;
  wire B_PE_dummy_in_13__ap_done;
  wire B_PE_dummy_in_13__ap_idle;
  wire B_PE_dummy_in_14__ap_start;
  wire B_PE_dummy_in_14__ap_ready;
  wire B_PE_dummy_in_14__ap_done;
  wire B_PE_dummy_in_14__ap_idle;
  wire B_PE_dummy_in_15__ap_start;
  wire B_PE_dummy_in_15__ap_ready;
  wire B_PE_dummy_in_15__ap_done;
  wire B_PE_dummy_in_15__ap_idle;
  wire B_PE_dummy_in_16__ap_start;
  wire B_PE_dummy_in_16__ap_ready;
  wire B_PE_dummy_in_16__ap_done;
  wire B_PE_dummy_in_16__ap_idle;
  wire C_drain_IO_L1_out_boundary_wrapper_0__ap_start;
  wire C_drain_IO_L1_out_boundary_wrapper_0__ap_ready;
  wire C_drain_IO_L1_out_boundary_wrapper_0__ap_done;
  wire C_drain_IO_L1_out_boundary_wrapper_0__ap_idle;
  wire C_drain_IO_L1_out_boundary_wrapper_1__ap_start;
  wire C_drain_IO_L1_out_boundary_wrapper_1__ap_ready;
  wire C_drain_IO_L1_out_boundary_wrapper_1__ap_done;
  wire C_drain_IO_L1_out_boundary_wrapper_1__ap_idle;
  wire C_drain_IO_L1_out_boundary_wrapper_2__ap_start;
  wire C_drain_IO_L1_out_boundary_wrapper_2__ap_ready;
  wire C_drain_IO_L1_out_boundary_wrapper_2__ap_done;
  wire C_drain_IO_L1_out_boundary_wrapper_2__ap_idle;
  wire C_drain_IO_L1_out_boundary_wrapper_3__ap_start;
  wire C_drain_IO_L1_out_boundary_wrapper_3__ap_ready;
  wire C_drain_IO_L1_out_boundary_wrapper_3__ap_done;
  wire C_drain_IO_L1_out_boundary_wrapper_3__ap_idle;
  wire C_drain_IO_L1_out_boundary_wrapper_4__ap_start;
  wire C_drain_IO_L1_out_boundary_wrapper_4__ap_ready;
  wire C_drain_IO_L1_out_boundary_wrapper_4__ap_done;
  wire C_drain_IO_L1_out_boundary_wrapper_4__ap_idle;
  wire C_drain_IO_L1_out_boundary_wrapper_5__ap_start;
  wire C_drain_IO_L1_out_boundary_wrapper_5__ap_ready;
  wire C_drain_IO_L1_out_boundary_wrapper_5__ap_done;
  wire C_drain_IO_L1_out_boundary_wrapper_5__ap_idle;
  wire C_drain_IO_L1_out_boundary_wrapper_6__ap_start;
  wire C_drain_IO_L1_out_boundary_wrapper_6__ap_ready;
  wire C_drain_IO_L1_out_boundary_wrapper_6__ap_done;
  wire C_drain_IO_L1_out_boundary_wrapper_6__ap_idle;
  wire C_drain_IO_L1_out_boundary_wrapper_7__ap_start;
  wire C_drain_IO_L1_out_boundary_wrapper_7__ap_ready;
  wire C_drain_IO_L1_out_boundary_wrapper_7__ap_done;
  wire C_drain_IO_L1_out_boundary_wrapper_7__ap_idle;
  wire C_drain_IO_L1_out_boundary_wrapper_8__ap_start;
  wire C_drain_IO_L1_out_boundary_wrapper_8__ap_ready;
  wire C_drain_IO_L1_out_boundary_wrapper_8__ap_done;
  wire C_drain_IO_L1_out_boundary_wrapper_8__ap_idle;
  wire C_drain_IO_L1_out_boundary_wrapper_9__ap_start;
  wire C_drain_IO_L1_out_boundary_wrapper_9__ap_ready;
  wire C_drain_IO_L1_out_boundary_wrapper_9__ap_done;
  wire C_drain_IO_L1_out_boundary_wrapper_9__ap_idle;
  wire C_drain_IO_L1_out_boundary_wrapper_10__ap_start;
  wire C_drain_IO_L1_out_boundary_wrapper_10__ap_ready;
  wire C_drain_IO_L1_out_boundary_wrapper_10__ap_done;
  wire C_drain_IO_L1_out_boundary_wrapper_10__ap_idle;
  wire C_drain_IO_L1_out_boundary_wrapper_11__ap_start;
  wire C_drain_IO_L1_out_boundary_wrapper_11__ap_ready;
  wire C_drain_IO_L1_out_boundary_wrapper_11__ap_done;
  wire C_drain_IO_L1_out_boundary_wrapper_11__ap_idle;
  wire C_drain_IO_L1_out_boundary_wrapper_12__ap_start;
  wire C_drain_IO_L1_out_boundary_wrapper_12__ap_ready;
  wire C_drain_IO_L1_out_boundary_wrapper_12__ap_done;
  wire C_drain_IO_L1_out_boundary_wrapper_12__ap_idle;
  wire C_drain_IO_L1_out_boundary_wrapper_13__ap_start;
  wire C_drain_IO_L1_out_boundary_wrapper_13__ap_ready;
  wire C_drain_IO_L1_out_boundary_wrapper_13__ap_done;
  wire C_drain_IO_L1_out_boundary_wrapper_13__ap_idle;
  wire C_drain_IO_L1_out_boundary_wrapper_14__ap_start;
  wire C_drain_IO_L1_out_boundary_wrapper_14__ap_ready;
  wire C_drain_IO_L1_out_boundary_wrapper_14__ap_done;
  wire C_drain_IO_L1_out_boundary_wrapper_14__ap_idle;
  wire C_drain_IO_L1_out_boundary_wrapper_15__ap_start;
  wire C_drain_IO_L1_out_boundary_wrapper_15__ap_ready;
  wire C_drain_IO_L1_out_boundary_wrapper_15__ap_done;
  wire C_drain_IO_L1_out_boundary_wrapper_15__ap_idle;
  wire C_drain_IO_L1_out_boundary_wrapper_16__ap_start;
  wire C_drain_IO_L1_out_boundary_wrapper_16__ap_ready;
  wire C_drain_IO_L1_out_boundary_wrapper_16__ap_done;
  wire C_drain_IO_L1_out_boundary_wrapper_16__ap_idle;
  wire C_drain_IO_L1_out_wrapper_0__ap_start;
  wire C_drain_IO_L1_out_wrapper_0__ap_ready;
  wire C_drain_IO_L1_out_wrapper_0__ap_done;
  wire C_drain_IO_L1_out_wrapper_0__ap_idle;
  wire C_drain_IO_L1_out_wrapper_1__ap_start;
  wire C_drain_IO_L1_out_wrapper_1__ap_ready;
  wire C_drain_IO_L1_out_wrapper_1__ap_done;
  wire C_drain_IO_L1_out_wrapper_1__ap_idle;
  wire C_drain_IO_L1_out_wrapper_2__ap_start;
  wire C_drain_IO_L1_out_wrapper_2__ap_ready;
  wire C_drain_IO_L1_out_wrapper_2__ap_done;
  wire C_drain_IO_L1_out_wrapper_2__ap_idle;
  wire C_drain_IO_L1_out_wrapper_3__ap_start;
  wire C_drain_IO_L1_out_wrapper_3__ap_ready;
  wire C_drain_IO_L1_out_wrapper_3__ap_done;
  wire C_drain_IO_L1_out_wrapper_3__ap_idle;
  wire C_drain_IO_L1_out_wrapper_4__ap_start;
  wire C_drain_IO_L1_out_wrapper_4__ap_ready;
  wire C_drain_IO_L1_out_wrapper_4__ap_done;
  wire C_drain_IO_L1_out_wrapper_4__ap_idle;
  wire C_drain_IO_L1_out_wrapper_5__ap_start;
  wire C_drain_IO_L1_out_wrapper_5__ap_ready;
  wire C_drain_IO_L1_out_wrapper_5__ap_done;
  wire C_drain_IO_L1_out_wrapper_5__ap_idle;
  wire C_drain_IO_L1_out_wrapper_6__ap_start;
  wire C_drain_IO_L1_out_wrapper_6__ap_ready;
  wire C_drain_IO_L1_out_wrapper_6__ap_done;
  wire C_drain_IO_L1_out_wrapper_6__ap_idle;
  wire C_drain_IO_L1_out_wrapper_7__ap_start;
  wire C_drain_IO_L1_out_wrapper_7__ap_ready;
  wire C_drain_IO_L1_out_wrapper_7__ap_done;
  wire C_drain_IO_L1_out_wrapper_7__ap_idle;
  wire C_drain_IO_L1_out_wrapper_8__ap_start;
  wire C_drain_IO_L1_out_wrapper_8__ap_ready;
  wire C_drain_IO_L1_out_wrapper_8__ap_done;
  wire C_drain_IO_L1_out_wrapper_8__ap_idle;
  wire C_drain_IO_L1_out_wrapper_9__ap_start;
  wire C_drain_IO_L1_out_wrapper_9__ap_ready;
  wire C_drain_IO_L1_out_wrapper_9__ap_done;
  wire C_drain_IO_L1_out_wrapper_9__ap_idle;
  wire C_drain_IO_L1_out_wrapper_10__ap_start;
  wire C_drain_IO_L1_out_wrapper_10__ap_ready;
  wire C_drain_IO_L1_out_wrapper_10__ap_done;
  wire C_drain_IO_L1_out_wrapper_10__ap_idle;
  wire C_drain_IO_L1_out_wrapper_11__ap_start;
  wire C_drain_IO_L1_out_wrapper_11__ap_ready;
  wire C_drain_IO_L1_out_wrapper_11__ap_done;
  wire C_drain_IO_L1_out_wrapper_11__ap_idle;
  wire C_drain_IO_L1_out_wrapper_12__ap_start;
  wire C_drain_IO_L1_out_wrapper_12__ap_ready;
  wire C_drain_IO_L1_out_wrapper_12__ap_done;
  wire C_drain_IO_L1_out_wrapper_12__ap_idle;
  wire C_drain_IO_L1_out_wrapper_13__ap_start;
  wire C_drain_IO_L1_out_wrapper_13__ap_ready;
  wire C_drain_IO_L1_out_wrapper_13__ap_done;
  wire C_drain_IO_L1_out_wrapper_13__ap_idle;
  wire C_drain_IO_L1_out_wrapper_14__ap_start;
  wire C_drain_IO_L1_out_wrapper_14__ap_ready;
  wire C_drain_IO_L1_out_wrapper_14__ap_done;
  wire C_drain_IO_L1_out_wrapper_14__ap_idle;
  wire C_drain_IO_L1_out_wrapper_15__ap_start;
  wire C_drain_IO_L1_out_wrapper_15__ap_ready;
  wire C_drain_IO_L1_out_wrapper_15__ap_done;
  wire C_drain_IO_L1_out_wrapper_15__ap_idle;
  wire C_drain_IO_L1_out_wrapper_16__ap_start;
  wire C_drain_IO_L1_out_wrapper_16__ap_ready;
  wire C_drain_IO_L1_out_wrapper_16__ap_done;
  wire C_drain_IO_L1_out_wrapper_16__ap_idle;
  wire C_drain_IO_L1_out_wrapper_17__ap_start;
  wire C_drain_IO_L1_out_wrapper_17__ap_ready;
  wire C_drain_IO_L1_out_wrapper_17__ap_done;
  wire C_drain_IO_L1_out_wrapper_17__ap_idle;
  wire C_drain_IO_L1_out_wrapper_18__ap_start;
  wire C_drain_IO_L1_out_wrapper_18__ap_ready;
  wire C_drain_IO_L1_out_wrapper_18__ap_done;
  wire C_drain_IO_L1_out_wrapper_18__ap_idle;
  wire C_drain_IO_L1_out_wrapper_19__ap_start;
  wire C_drain_IO_L1_out_wrapper_19__ap_ready;
  wire C_drain_IO_L1_out_wrapper_19__ap_done;
  wire C_drain_IO_L1_out_wrapper_19__ap_idle;
  wire C_drain_IO_L1_out_wrapper_20__ap_start;
  wire C_drain_IO_L1_out_wrapper_20__ap_ready;
  wire C_drain_IO_L1_out_wrapper_20__ap_done;
  wire C_drain_IO_L1_out_wrapper_20__ap_idle;
  wire C_drain_IO_L1_out_wrapper_21__ap_start;
  wire C_drain_IO_L1_out_wrapper_21__ap_ready;
  wire C_drain_IO_L1_out_wrapper_21__ap_done;
  wire C_drain_IO_L1_out_wrapper_21__ap_idle;
  wire C_drain_IO_L1_out_wrapper_22__ap_start;
  wire C_drain_IO_L1_out_wrapper_22__ap_ready;
  wire C_drain_IO_L1_out_wrapper_22__ap_done;
  wire C_drain_IO_L1_out_wrapper_22__ap_idle;
  wire C_drain_IO_L1_out_wrapper_23__ap_start;
  wire C_drain_IO_L1_out_wrapper_23__ap_ready;
  wire C_drain_IO_L1_out_wrapper_23__ap_done;
  wire C_drain_IO_L1_out_wrapper_23__ap_idle;
  wire C_drain_IO_L1_out_wrapper_24__ap_start;
  wire C_drain_IO_L1_out_wrapper_24__ap_ready;
  wire C_drain_IO_L1_out_wrapper_24__ap_done;
  wire C_drain_IO_L1_out_wrapper_24__ap_idle;
  wire C_drain_IO_L1_out_wrapper_25__ap_start;
  wire C_drain_IO_L1_out_wrapper_25__ap_ready;
  wire C_drain_IO_L1_out_wrapper_25__ap_done;
  wire C_drain_IO_L1_out_wrapper_25__ap_idle;
  wire C_drain_IO_L1_out_wrapper_26__ap_start;
  wire C_drain_IO_L1_out_wrapper_26__ap_ready;
  wire C_drain_IO_L1_out_wrapper_26__ap_done;
  wire C_drain_IO_L1_out_wrapper_26__ap_idle;
  wire C_drain_IO_L1_out_wrapper_27__ap_start;
  wire C_drain_IO_L1_out_wrapper_27__ap_ready;
  wire C_drain_IO_L1_out_wrapper_27__ap_done;
  wire C_drain_IO_L1_out_wrapper_27__ap_idle;
  wire C_drain_IO_L1_out_wrapper_28__ap_start;
  wire C_drain_IO_L1_out_wrapper_28__ap_ready;
  wire C_drain_IO_L1_out_wrapper_28__ap_done;
  wire C_drain_IO_L1_out_wrapper_28__ap_idle;
  wire C_drain_IO_L1_out_wrapper_29__ap_start;
  wire C_drain_IO_L1_out_wrapper_29__ap_ready;
  wire C_drain_IO_L1_out_wrapper_29__ap_done;
  wire C_drain_IO_L1_out_wrapper_29__ap_idle;
  wire C_drain_IO_L1_out_wrapper_30__ap_start;
  wire C_drain_IO_L1_out_wrapper_30__ap_ready;
  wire C_drain_IO_L1_out_wrapper_30__ap_done;
  wire C_drain_IO_L1_out_wrapper_30__ap_idle;
  wire C_drain_IO_L1_out_wrapper_31__ap_start;
  wire C_drain_IO_L1_out_wrapper_31__ap_ready;
  wire C_drain_IO_L1_out_wrapper_31__ap_done;
  wire C_drain_IO_L1_out_wrapper_31__ap_idle;
  wire C_drain_IO_L1_out_wrapper_32__ap_start;
  wire C_drain_IO_L1_out_wrapper_32__ap_ready;
  wire C_drain_IO_L1_out_wrapper_32__ap_done;
  wire C_drain_IO_L1_out_wrapper_32__ap_idle;
  wire C_drain_IO_L1_out_wrapper_33__ap_start;
  wire C_drain_IO_L1_out_wrapper_33__ap_ready;
  wire C_drain_IO_L1_out_wrapper_33__ap_done;
  wire C_drain_IO_L1_out_wrapper_33__ap_idle;
  wire C_drain_IO_L1_out_wrapper_34__ap_start;
  wire C_drain_IO_L1_out_wrapper_34__ap_ready;
  wire C_drain_IO_L1_out_wrapper_34__ap_done;
  wire C_drain_IO_L1_out_wrapper_34__ap_idle;
  wire C_drain_IO_L1_out_wrapper_35__ap_start;
  wire C_drain_IO_L1_out_wrapper_35__ap_ready;
  wire C_drain_IO_L1_out_wrapper_35__ap_done;
  wire C_drain_IO_L1_out_wrapper_35__ap_idle;
  wire C_drain_IO_L1_out_wrapper_36__ap_start;
  wire C_drain_IO_L1_out_wrapper_36__ap_ready;
  wire C_drain_IO_L1_out_wrapper_36__ap_done;
  wire C_drain_IO_L1_out_wrapper_36__ap_idle;
  wire C_drain_IO_L1_out_wrapper_37__ap_start;
  wire C_drain_IO_L1_out_wrapper_37__ap_ready;
  wire C_drain_IO_L1_out_wrapper_37__ap_done;
  wire C_drain_IO_L1_out_wrapper_37__ap_idle;
  wire C_drain_IO_L1_out_wrapper_38__ap_start;
  wire C_drain_IO_L1_out_wrapper_38__ap_ready;
  wire C_drain_IO_L1_out_wrapper_38__ap_done;
  wire C_drain_IO_L1_out_wrapper_38__ap_idle;
  wire C_drain_IO_L1_out_wrapper_39__ap_start;
  wire C_drain_IO_L1_out_wrapper_39__ap_ready;
  wire C_drain_IO_L1_out_wrapper_39__ap_done;
  wire C_drain_IO_L1_out_wrapper_39__ap_idle;
  wire C_drain_IO_L1_out_wrapper_40__ap_start;
  wire C_drain_IO_L1_out_wrapper_40__ap_ready;
  wire C_drain_IO_L1_out_wrapper_40__ap_done;
  wire C_drain_IO_L1_out_wrapper_40__ap_idle;
  wire C_drain_IO_L1_out_wrapper_41__ap_start;
  wire C_drain_IO_L1_out_wrapper_41__ap_ready;
  wire C_drain_IO_L1_out_wrapper_41__ap_done;
  wire C_drain_IO_L1_out_wrapper_41__ap_idle;
  wire C_drain_IO_L1_out_wrapper_42__ap_start;
  wire C_drain_IO_L1_out_wrapper_42__ap_ready;
  wire C_drain_IO_L1_out_wrapper_42__ap_done;
  wire C_drain_IO_L1_out_wrapper_42__ap_idle;
  wire C_drain_IO_L1_out_wrapper_43__ap_start;
  wire C_drain_IO_L1_out_wrapper_43__ap_ready;
  wire C_drain_IO_L1_out_wrapper_43__ap_done;
  wire C_drain_IO_L1_out_wrapper_43__ap_idle;
  wire C_drain_IO_L1_out_wrapper_44__ap_start;
  wire C_drain_IO_L1_out_wrapper_44__ap_ready;
  wire C_drain_IO_L1_out_wrapper_44__ap_done;
  wire C_drain_IO_L1_out_wrapper_44__ap_idle;
  wire C_drain_IO_L1_out_wrapper_45__ap_start;
  wire C_drain_IO_L1_out_wrapper_45__ap_ready;
  wire C_drain_IO_L1_out_wrapper_45__ap_done;
  wire C_drain_IO_L1_out_wrapper_45__ap_idle;
  wire C_drain_IO_L1_out_wrapper_46__ap_start;
  wire C_drain_IO_L1_out_wrapper_46__ap_ready;
  wire C_drain_IO_L1_out_wrapper_46__ap_done;
  wire C_drain_IO_L1_out_wrapper_46__ap_idle;
  wire C_drain_IO_L1_out_wrapper_47__ap_start;
  wire C_drain_IO_L1_out_wrapper_47__ap_ready;
  wire C_drain_IO_L1_out_wrapper_47__ap_done;
  wire C_drain_IO_L1_out_wrapper_47__ap_idle;
  wire C_drain_IO_L1_out_wrapper_48__ap_start;
  wire C_drain_IO_L1_out_wrapper_48__ap_ready;
  wire C_drain_IO_L1_out_wrapper_48__ap_done;
  wire C_drain_IO_L1_out_wrapper_48__ap_idle;
  wire C_drain_IO_L1_out_wrapper_49__ap_start;
  wire C_drain_IO_L1_out_wrapper_49__ap_ready;
  wire C_drain_IO_L1_out_wrapper_49__ap_done;
  wire C_drain_IO_L1_out_wrapper_49__ap_idle;
  wire C_drain_IO_L1_out_wrapper_50__ap_start;
  wire C_drain_IO_L1_out_wrapper_50__ap_ready;
  wire C_drain_IO_L1_out_wrapper_50__ap_done;
  wire C_drain_IO_L1_out_wrapper_50__ap_idle;
  wire C_drain_IO_L1_out_wrapper_51__ap_start;
  wire C_drain_IO_L1_out_wrapper_51__ap_ready;
  wire C_drain_IO_L1_out_wrapper_51__ap_done;
  wire C_drain_IO_L1_out_wrapper_51__ap_idle;
  wire C_drain_IO_L1_out_wrapper_52__ap_start;
  wire C_drain_IO_L1_out_wrapper_52__ap_ready;
  wire C_drain_IO_L1_out_wrapper_52__ap_done;
  wire C_drain_IO_L1_out_wrapper_52__ap_idle;
  wire C_drain_IO_L1_out_wrapper_53__ap_start;
  wire C_drain_IO_L1_out_wrapper_53__ap_ready;
  wire C_drain_IO_L1_out_wrapper_53__ap_done;
  wire C_drain_IO_L1_out_wrapper_53__ap_idle;
  wire C_drain_IO_L1_out_wrapper_54__ap_start;
  wire C_drain_IO_L1_out_wrapper_54__ap_ready;
  wire C_drain_IO_L1_out_wrapper_54__ap_done;
  wire C_drain_IO_L1_out_wrapper_54__ap_idle;
  wire C_drain_IO_L1_out_wrapper_55__ap_start;
  wire C_drain_IO_L1_out_wrapper_55__ap_ready;
  wire C_drain_IO_L1_out_wrapper_55__ap_done;
  wire C_drain_IO_L1_out_wrapper_55__ap_idle;
  wire C_drain_IO_L1_out_wrapper_56__ap_start;
  wire C_drain_IO_L1_out_wrapper_56__ap_ready;
  wire C_drain_IO_L1_out_wrapper_56__ap_done;
  wire C_drain_IO_L1_out_wrapper_56__ap_idle;
  wire C_drain_IO_L1_out_wrapper_57__ap_start;
  wire C_drain_IO_L1_out_wrapper_57__ap_ready;
  wire C_drain_IO_L1_out_wrapper_57__ap_done;
  wire C_drain_IO_L1_out_wrapper_57__ap_idle;
  wire C_drain_IO_L1_out_wrapper_58__ap_start;
  wire C_drain_IO_L1_out_wrapper_58__ap_ready;
  wire C_drain_IO_L1_out_wrapper_58__ap_done;
  wire C_drain_IO_L1_out_wrapper_58__ap_idle;
  wire C_drain_IO_L1_out_wrapper_59__ap_start;
  wire C_drain_IO_L1_out_wrapper_59__ap_ready;
  wire C_drain_IO_L1_out_wrapper_59__ap_done;
  wire C_drain_IO_L1_out_wrapper_59__ap_idle;
  wire C_drain_IO_L1_out_wrapper_60__ap_start;
  wire C_drain_IO_L1_out_wrapper_60__ap_ready;
  wire C_drain_IO_L1_out_wrapper_60__ap_done;
  wire C_drain_IO_L1_out_wrapper_60__ap_idle;
  wire C_drain_IO_L1_out_wrapper_61__ap_start;
  wire C_drain_IO_L1_out_wrapper_61__ap_ready;
  wire C_drain_IO_L1_out_wrapper_61__ap_done;
  wire C_drain_IO_L1_out_wrapper_61__ap_idle;
  wire C_drain_IO_L1_out_wrapper_62__ap_start;
  wire C_drain_IO_L1_out_wrapper_62__ap_ready;
  wire C_drain_IO_L1_out_wrapper_62__ap_done;
  wire C_drain_IO_L1_out_wrapper_62__ap_idle;
  wire C_drain_IO_L1_out_wrapper_63__ap_start;
  wire C_drain_IO_L1_out_wrapper_63__ap_ready;
  wire C_drain_IO_L1_out_wrapper_63__ap_done;
  wire C_drain_IO_L1_out_wrapper_63__ap_idle;
  wire C_drain_IO_L1_out_wrapper_64__ap_start;
  wire C_drain_IO_L1_out_wrapper_64__ap_ready;
  wire C_drain_IO_L1_out_wrapper_64__ap_done;
  wire C_drain_IO_L1_out_wrapper_64__ap_idle;
  wire C_drain_IO_L1_out_wrapper_65__ap_start;
  wire C_drain_IO_L1_out_wrapper_65__ap_ready;
  wire C_drain_IO_L1_out_wrapper_65__ap_done;
  wire C_drain_IO_L1_out_wrapper_65__ap_idle;
  wire C_drain_IO_L1_out_wrapper_66__ap_start;
  wire C_drain_IO_L1_out_wrapper_66__ap_ready;
  wire C_drain_IO_L1_out_wrapper_66__ap_done;
  wire C_drain_IO_L1_out_wrapper_66__ap_idle;
  wire C_drain_IO_L1_out_wrapper_67__ap_start;
  wire C_drain_IO_L1_out_wrapper_67__ap_ready;
  wire C_drain_IO_L1_out_wrapper_67__ap_done;
  wire C_drain_IO_L1_out_wrapper_67__ap_idle;
  wire C_drain_IO_L1_out_wrapper_68__ap_start;
  wire C_drain_IO_L1_out_wrapper_68__ap_ready;
  wire C_drain_IO_L1_out_wrapper_68__ap_done;
  wire C_drain_IO_L1_out_wrapper_68__ap_idle;
  wire C_drain_IO_L1_out_wrapper_69__ap_start;
  wire C_drain_IO_L1_out_wrapper_69__ap_ready;
  wire C_drain_IO_L1_out_wrapper_69__ap_done;
  wire C_drain_IO_L1_out_wrapper_69__ap_idle;
  wire C_drain_IO_L1_out_wrapper_70__ap_start;
  wire C_drain_IO_L1_out_wrapper_70__ap_ready;
  wire C_drain_IO_L1_out_wrapper_70__ap_done;
  wire C_drain_IO_L1_out_wrapper_70__ap_idle;
  wire C_drain_IO_L1_out_wrapper_71__ap_start;
  wire C_drain_IO_L1_out_wrapper_71__ap_ready;
  wire C_drain_IO_L1_out_wrapper_71__ap_done;
  wire C_drain_IO_L1_out_wrapper_71__ap_idle;
  wire C_drain_IO_L1_out_wrapper_72__ap_start;
  wire C_drain_IO_L1_out_wrapper_72__ap_ready;
  wire C_drain_IO_L1_out_wrapper_72__ap_done;
  wire C_drain_IO_L1_out_wrapper_72__ap_idle;
  wire C_drain_IO_L1_out_wrapper_73__ap_start;
  wire C_drain_IO_L1_out_wrapper_73__ap_ready;
  wire C_drain_IO_L1_out_wrapper_73__ap_done;
  wire C_drain_IO_L1_out_wrapper_73__ap_idle;
  wire C_drain_IO_L1_out_wrapper_74__ap_start;
  wire C_drain_IO_L1_out_wrapper_74__ap_ready;
  wire C_drain_IO_L1_out_wrapper_74__ap_done;
  wire C_drain_IO_L1_out_wrapper_74__ap_idle;
  wire C_drain_IO_L1_out_wrapper_75__ap_start;
  wire C_drain_IO_L1_out_wrapper_75__ap_ready;
  wire C_drain_IO_L1_out_wrapper_75__ap_done;
  wire C_drain_IO_L1_out_wrapper_75__ap_idle;
  wire C_drain_IO_L1_out_wrapper_76__ap_start;
  wire C_drain_IO_L1_out_wrapper_76__ap_ready;
  wire C_drain_IO_L1_out_wrapper_76__ap_done;
  wire C_drain_IO_L1_out_wrapper_76__ap_idle;
  wire C_drain_IO_L1_out_wrapper_77__ap_start;
  wire C_drain_IO_L1_out_wrapper_77__ap_ready;
  wire C_drain_IO_L1_out_wrapper_77__ap_done;
  wire C_drain_IO_L1_out_wrapper_77__ap_idle;
  wire C_drain_IO_L1_out_wrapper_78__ap_start;
  wire C_drain_IO_L1_out_wrapper_78__ap_ready;
  wire C_drain_IO_L1_out_wrapper_78__ap_done;
  wire C_drain_IO_L1_out_wrapper_78__ap_idle;
  wire C_drain_IO_L1_out_wrapper_79__ap_start;
  wire C_drain_IO_L1_out_wrapper_79__ap_ready;
  wire C_drain_IO_L1_out_wrapper_79__ap_done;
  wire C_drain_IO_L1_out_wrapper_79__ap_idle;
  wire C_drain_IO_L1_out_wrapper_80__ap_start;
  wire C_drain_IO_L1_out_wrapper_80__ap_ready;
  wire C_drain_IO_L1_out_wrapper_80__ap_done;
  wire C_drain_IO_L1_out_wrapper_80__ap_idle;
  wire C_drain_IO_L1_out_wrapper_81__ap_start;
  wire C_drain_IO_L1_out_wrapper_81__ap_ready;
  wire C_drain_IO_L1_out_wrapper_81__ap_done;
  wire C_drain_IO_L1_out_wrapper_81__ap_idle;
  wire C_drain_IO_L1_out_wrapper_82__ap_start;
  wire C_drain_IO_L1_out_wrapper_82__ap_ready;
  wire C_drain_IO_L1_out_wrapper_82__ap_done;
  wire C_drain_IO_L1_out_wrapper_82__ap_idle;
  wire C_drain_IO_L1_out_wrapper_83__ap_start;
  wire C_drain_IO_L1_out_wrapper_83__ap_ready;
  wire C_drain_IO_L1_out_wrapper_83__ap_done;
  wire C_drain_IO_L1_out_wrapper_83__ap_idle;
  wire C_drain_IO_L1_out_wrapper_84__ap_start;
  wire C_drain_IO_L1_out_wrapper_84__ap_ready;
  wire C_drain_IO_L1_out_wrapper_84__ap_done;
  wire C_drain_IO_L1_out_wrapper_84__ap_idle;
  wire C_drain_IO_L1_out_wrapper_85__ap_start;
  wire C_drain_IO_L1_out_wrapper_85__ap_ready;
  wire C_drain_IO_L1_out_wrapper_85__ap_done;
  wire C_drain_IO_L1_out_wrapper_85__ap_idle;
  wire C_drain_IO_L1_out_wrapper_86__ap_start;
  wire C_drain_IO_L1_out_wrapper_86__ap_ready;
  wire C_drain_IO_L1_out_wrapper_86__ap_done;
  wire C_drain_IO_L1_out_wrapper_86__ap_idle;
  wire C_drain_IO_L1_out_wrapper_87__ap_start;
  wire C_drain_IO_L1_out_wrapper_87__ap_ready;
  wire C_drain_IO_L1_out_wrapper_87__ap_done;
  wire C_drain_IO_L1_out_wrapper_87__ap_idle;
  wire C_drain_IO_L1_out_wrapper_88__ap_start;
  wire C_drain_IO_L1_out_wrapper_88__ap_ready;
  wire C_drain_IO_L1_out_wrapper_88__ap_done;
  wire C_drain_IO_L1_out_wrapper_88__ap_idle;
  wire C_drain_IO_L1_out_wrapper_89__ap_start;
  wire C_drain_IO_L1_out_wrapper_89__ap_ready;
  wire C_drain_IO_L1_out_wrapper_89__ap_done;
  wire C_drain_IO_L1_out_wrapper_89__ap_idle;
  wire C_drain_IO_L1_out_wrapper_90__ap_start;
  wire C_drain_IO_L1_out_wrapper_90__ap_ready;
  wire C_drain_IO_L1_out_wrapper_90__ap_done;
  wire C_drain_IO_L1_out_wrapper_90__ap_idle;
  wire C_drain_IO_L1_out_wrapper_91__ap_start;
  wire C_drain_IO_L1_out_wrapper_91__ap_ready;
  wire C_drain_IO_L1_out_wrapper_91__ap_done;
  wire C_drain_IO_L1_out_wrapper_91__ap_idle;
  wire C_drain_IO_L1_out_wrapper_92__ap_start;
  wire C_drain_IO_L1_out_wrapper_92__ap_ready;
  wire C_drain_IO_L1_out_wrapper_92__ap_done;
  wire C_drain_IO_L1_out_wrapper_92__ap_idle;
  wire C_drain_IO_L1_out_wrapper_93__ap_start;
  wire C_drain_IO_L1_out_wrapper_93__ap_ready;
  wire C_drain_IO_L1_out_wrapper_93__ap_done;
  wire C_drain_IO_L1_out_wrapper_93__ap_idle;
  wire C_drain_IO_L1_out_wrapper_94__ap_start;
  wire C_drain_IO_L1_out_wrapper_94__ap_ready;
  wire C_drain_IO_L1_out_wrapper_94__ap_done;
  wire C_drain_IO_L1_out_wrapper_94__ap_idle;
  wire C_drain_IO_L1_out_wrapper_95__ap_start;
  wire C_drain_IO_L1_out_wrapper_95__ap_ready;
  wire C_drain_IO_L1_out_wrapper_95__ap_done;
  wire C_drain_IO_L1_out_wrapper_95__ap_idle;
  wire C_drain_IO_L1_out_wrapper_96__ap_start;
  wire C_drain_IO_L1_out_wrapper_96__ap_ready;
  wire C_drain_IO_L1_out_wrapper_96__ap_done;
  wire C_drain_IO_L1_out_wrapper_96__ap_idle;
  wire C_drain_IO_L1_out_wrapper_97__ap_start;
  wire C_drain_IO_L1_out_wrapper_97__ap_ready;
  wire C_drain_IO_L1_out_wrapper_97__ap_done;
  wire C_drain_IO_L1_out_wrapper_97__ap_idle;
  wire C_drain_IO_L1_out_wrapper_98__ap_start;
  wire C_drain_IO_L1_out_wrapper_98__ap_ready;
  wire C_drain_IO_L1_out_wrapper_98__ap_done;
  wire C_drain_IO_L1_out_wrapper_98__ap_idle;
  wire C_drain_IO_L1_out_wrapper_99__ap_start;
  wire C_drain_IO_L1_out_wrapper_99__ap_ready;
  wire C_drain_IO_L1_out_wrapper_99__ap_done;
  wire C_drain_IO_L1_out_wrapper_99__ap_idle;
  wire C_drain_IO_L1_out_wrapper_100__ap_start;
  wire C_drain_IO_L1_out_wrapper_100__ap_ready;
  wire C_drain_IO_L1_out_wrapper_100__ap_done;
  wire C_drain_IO_L1_out_wrapper_100__ap_idle;
  wire C_drain_IO_L1_out_wrapper_101__ap_start;
  wire C_drain_IO_L1_out_wrapper_101__ap_ready;
  wire C_drain_IO_L1_out_wrapper_101__ap_done;
  wire C_drain_IO_L1_out_wrapper_101__ap_idle;
  wire C_drain_IO_L1_out_wrapper_102__ap_start;
  wire C_drain_IO_L1_out_wrapper_102__ap_ready;
  wire C_drain_IO_L1_out_wrapper_102__ap_done;
  wire C_drain_IO_L1_out_wrapper_102__ap_idle;
  wire C_drain_IO_L1_out_wrapper_103__ap_start;
  wire C_drain_IO_L1_out_wrapper_103__ap_ready;
  wire C_drain_IO_L1_out_wrapper_103__ap_done;
  wire C_drain_IO_L1_out_wrapper_103__ap_idle;
  wire C_drain_IO_L1_out_wrapper_104__ap_start;
  wire C_drain_IO_L1_out_wrapper_104__ap_ready;
  wire C_drain_IO_L1_out_wrapper_104__ap_done;
  wire C_drain_IO_L1_out_wrapper_104__ap_idle;
  wire C_drain_IO_L1_out_wrapper_105__ap_start;
  wire C_drain_IO_L1_out_wrapper_105__ap_ready;
  wire C_drain_IO_L1_out_wrapper_105__ap_done;
  wire C_drain_IO_L1_out_wrapper_105__ap_idle;
  wire C_drain_IO_L1_out_wrapper_106__ap_start;
  wire C_drain_IO_L1_out_wrapper_106__ap_ready;
  wire C_drain_IO_L1_out_wrapper_106__ap_done;
  wire C_drain_IO_L1_out_wrapper_106__ap_idle;
  wire C_drain_IO_L1_out_wrapper_107__ap_start;
  wire C_drain_IO_L1_out_wrapper_107__ap_ready;
  wire C_drain_IO_L1_out_wrapper_107__ap_done;
  wire C_drain_IO_L1_out_wrapper_107__ap_idle;
  wire C_drain_IO_L1_out_wrapper_108__ap_start;
  wire C_drain_IO_L1_out_wrapper_108__ap_ready;
  wire C_drain_IO_L1_out_wrapper_108__ap_done;
  wire C_drain_IO_L1_out_wrapper_108__ap_idle;
  wire C_drain_IO_L1_out_wrapper_109__ap_start;
  wire C_drain_IO_L1_out_wrapper_109__ap_ready;
  wire C_drain_IO_L1_out_wrapper_109__ap_done;
  wire C_drain_IO_L1_out_wrapper_109__ap_idle;
  wire C_drain_IO_L1_out_wrapper_110__ap_start;
  wire C_drain_IO_L1_out_wrapper_110__ap_ready;
  wire C_drain_IO_L1_out_wrapper_110__ap_done;
  wire C_drain_IO_L1_out_wrapper_110__ap_idle;
  wire C_drain_IO_L1_out_wrapper_111__ap_start;
  wire C_drain_IO_L1_out_wrapper_111__ap_ready;
  wire C_drain_IO_L1_out_wrapper_111__ap_done;
  wire C_drain_IO_L1_out_wrapper_111__ap_idle;
  wire C_drain_IO_L1_out_wrapper_112__ap_start;
  wire C_drain_IO_L1_out_wrapper_112__ap_ready;
  wire C_drain_IO_L1_out_wrapper_112__ap_done;
  wire C_drain_IO_L1_out_wrapper_112__ap_idle;
  wire C_drain_IO_L1_out_wrapper_113__ap_start;
  wire C_drain_IO_L1_out_wrapper_113__ap_ready;
  wire C_drain_IO_L1_out_wrapper_113__ap_done;
  wire C_drain_IO_L1_out_wrapper_113__ap_idle;
  wire C_drain_IO_L1_out_wrapper_114__ap_start;
  wire C_drain_IO_L1_out_wrapper_114__ap_ready;
  wire C_drain_IO_L1_out_wrapper_114__ap_done;
  wire C_drain_IO_L1_out_wrapper_114__ap_idle;
  wire C_drain_IO_L1_out_wrapper_115__ap_start;
  wire C_drain_IO_L1_out_wrapper_115__ap_ready;
  wire C_drain_IO_L1_out_wrapper_115__ap_done;
  wire C_drain_IO_L1_out_wrapper_115__ap_idle;
  wire C_drain_IO_L1_out_wrapper_116__ap_start;
  wire C_drain_IO_L1_out_wrapper_116__ap_ready;
  wire C_drain_IO_L1_out_wrapper_116__ap_done;
  wire C_drain_IO_L1_out_wrapper_116__ap_idle;
  wire C_drain_IO_L1_out_wrapper_117__ap_start;
  wire C_drain_IO_L1_out_wrapper_117__ap_ready;
  wire C_drain_IO_L1_out_wrapper_117__ap_done;
  wire C_drain_IO_L1_out_wrapper_117__ap_idle;
  wire C_drain_IO_L1_out_wrapper_118__ap_start;
  wire C_drain_IO_L1_out_wrapper_118__ap_ready;
  wire C_drain_IO_L1_out_wrapper_118__ap_done;
  wire C_drain_IO_L1_out_wrapper_118__ap_idle;
  wire C_drain_IO_L1_out_wrapper_119__ap_start;
  wire C_drain_IO_L1_out_wrapper_119__ap_ready;
  wire C_drain_IO_L1_out_wrapper_119__ap_done;
  wire C_drain_IO_L1_out_wrapper_119__ap_idle;
  wire C_drain_IO_L1_out_wrapper_120__ap_start;
  wire C_drain_IO_L1_out_wrapper_120__ap_ready;
  wire C_drain_IO_L1_out_wrapper_120__ap_done;
  wire C_drain_IO_L1_out_wrapper_120__ap_idle;
  wire C_drain_IO_L1_out_wrapper_121__ap_start;
  wire C_drain_IO_L1_out_wrapper_121__ap_ready;
  wire C_drain_IO_L1_out_wrapper_121__ap_done;
  wire C_drain_IO_L1_out_wrapper_121__ap_idle;
  wire C_drain_IO_L1_out_wrapper_122__ap_start;
  wire C_drain_IO_L1_out_wrapper_122__ap_ready;
  wire C_drain_IO_L1_out_wrapper_122__ap_done;
  wire C_drain_IO_L1_out_wrapper_122__ap_idle;
  wire C_drain_IO_L1_out_wrapper_123__ap_start;
  wire C_drain_IO_L1_out_wrapper_123__ap_ready;
  wire C_drain_IO_L1_out_wrapper_123__ap_done;
  wire C_drain_IO_L1_out_wrapper_123__ap_idle;
  wire C_drain_IO_L1_out_wrapper_124__ap_start;
  wire C_drain_IO_L1_out_wrapper_124__ap_ready;
  wire C_drain_IO_L1_out_wrapper_124__ap_done;
  wire C_drain_IO_L1_out_wrapper_124__ap_idle;
  wire C_drain_IO_L1_out_wrapper_125__ap_start;
  wire C_drain_IO_L1_out_wrapper_125__ap_ready;
  wire C_drain_IO_L1_out_wrapper_125__ap_done;
  wire C_drain_IO_L1_out_wrapper_125__ap_idle;
  wire C_drain_IO_L1_out_wrapper_126__ap_start;
  wire C_drain_IO_L1_out_wrapper_126__ap_ready;
  wire C_drain_IO_L1_out_wrapper_126__ap_done;
  wire C_drain_IO_L1_out_wrapper_126__ap_idle;
  wire C_drain_IO_L1_out_wrapper_127__ap_start;
  wire C_drain_IO_L1_out_wrapper_127__ap_ready;
  wire C_drain_IO_L1_out_wrapper_127__ap_done;
  wire C_drain_IO_L1_out_wrapper_127__ap_idle;
  wire C_drain_IO_L1_out_wrapper_128__ap_start;
  wire C_drain_IO_L1_out_wrapper_128__ap_ready;
  wire C_drain_IO_L1_out_wrapper_128__ap_done;
  wire C_drain_IO_L1_out_wrapper_128__ap_idle;
  wire C_drain_IO_L1_out_wrapper_129__ap_start;
  wire C_drain_IO_L1_out_wrapper_129__ap_ready;
  wire C_drain_IO_L1_out_wrapper_129__ap_done;
  wire C_drain_IO_L1_out_wrapper_129__ap_idle;
  wire C_drain_IO_L1_out_wrapper_130__ap_start;
  wire C_drain_IO_L1_out_wrapper_130__ap_ready;
  wire C_drain_IO_L1_out_wrapper_130__ap_done;
  wire C_drain_IO_L1_out_wrapper_130__ap_idle;
  wire C_drain_IO_L1_out_wrapper_131__ap_start;
  wire C_drain_IO_L1_out_wrapper_131__ap_ready;
  wire C_drain_IO_L1_out_wrapper_131__ap_done;
  wire C_drain_IO_L1_out_wrapper_131__ap_idle;
  wire C_drain_IO_L1_out_wrapper_132__ap_start;
  wire C_drain_IO_L1_out_wrapper_132__ap_ready;
  wire C_drain_IO_L1_out_wrapper_132__ap_done;
  wire C_drain_IO_L1_out_wrapper_132__ap_idle;
  wire C_drain_IO_L1_out_wrapper_133__ap_start;
  wire C_drain_IO_L1_out_wrapper_133__ap_ready;
  wire C_drain_IO_L1_out_wrapper_133__ap_done;
  wire C_drain_IO_L1_out_wrapper_133__ap_idle;
  wire C_drain_IO_L1_out_wrapper_134__ap_start;
  wire C_drain_IO_L1_out_wrapper_134__ap_ready;
  wire C_drain_IO_L1_out_wrapper_134__ap_done;
  wire C_drain_IO_L1_out_wrapper_134__ap_idle;
  wire C_drain_IO_L1_out_wrapper_135__ap_start;
  wire C_drain_IO_L1_out_wrapper_135__ap_ready;
  wire C_drain_IO_L1_out_wrapper_135__ap_done;
  wire C_drain_IO_L1_out_wrapper_135__ap_idle;
  wire C_drain_IO_L1_out_wrapper_136__ap_start;
  wire C_drain_IO_L1_out_wrapper_136__ap_ready;
  wire C_drain_IO_L1_out_wrapper_136__ap_done;
  wire C_drain_IO_L1_out_wrapper_136__ap_idle;
  wire C_drain_IO_L1_out_wrapper_137__ap_start;
  wire C_drain_IO_L1_out_wrapper_137__ap_ready;
  wire C_drain_IO_L1_out_wrapper_137__ap_done;
  wire C_drain_IO_L1_out_wrapper_137__ap_idle;
  wire C_drain_IO_L1_out_wrapper_138__ap_start;
  wire C_drain_IO_L1_out_wrapper_138__ap_ready;
  wire C_drain_IO_L1_out_wrapper_138__ap_done;
  wire C_drain_IO_L1_out_wrapper_138__ap_idle;
  wire C_drain_IO_L1_out_wrapper_139__ap_start;
  wire C_drain_IO_L1_out_wrapper_139__ap_ready;
  wire C_drain_IO_L1_out_wrapper_139__ap_done;
  wire C_drain_IO_L1_out_wrapper_139__ap_idle;
  wire C_drain_IO_L1_out_wrapper_140__ap_start;
  wire C_drain_IO_L1_out_wrapper_140__ap_ready;
  wire C_drain_IO_L1_out_wrapper_140__ap_done;
  wire C_drain_IO_L1_out_wrapper_140__ap_idle;
  wire C_drain_IO_L1_out_wrapper_141__ap_start;
  wire C_drain_IO_L1_out_wrapper_141__ap_ready;
  wire C_drain_IO_L1_out_wrapper_141__ap_done;
  wire C_drain_IO_L1_out_wrapper_141__ap_idle;
  wire C_drain_IO_L1_out_wrapper_142__ap_start;
  wire C_drain_IO_L1_out_wrapper_142__ap_ready;
  wire C_drain_IO_L1_out_wrapper_142__ap_done;
  wire C_drain_IO_L1_out_wrapper_142__ap_idle;
  wire C_drain_IO_L1_out_wrapper_143__ap_start;
  wire C_drain_IO_L1_out_wrapper_143__ap_ready;
  wire C_drain_IO_L1_out_wrapper_143__ap_done;
  wire C_drain_IO_L1_out_wrapper_143__ap_idle;
  wire C_drain_IO_L1_out_wrapper_144__ap_start;
  wire C_drain_IO_L1_out_wrapper_144__ap_ready;
  wire C_drain_IO_L1_out_wrapper_144__ap_done;
  wire C_drain_IO_L1_out_wrapper_144__ap_idle;
  wire C_drain_IO_L1_out_wrapper_145__ap_start;
  wire C_drain_IO_L1_out_wrapper_145__ap_ready;
  wire C_drain_IO_L1_out_wrapper_145__ap_done;
  wire C_drain_IO_L1_out_wrapper_145__ap_idle;
  wire C_drain_IO_L1_out_wrapper_146__ap_start;
  wire C_drain_IO_L1_out_wrapper_146__ap_ready;
  wire C_drain_IO_L1_out_wrapper_146__ap_done;
  wire C_drain_IO_L1_out_wrapper_146__ap_idle;
  wire C_drain_IO_L1_out_wrapper_147__ap_start;
  wire C_drain_IO_L1_out_wrapper_147__ap_ready;
  wire C_drain_IO_L1_out_wrapper_147__ap_done;
  wire C_drain_IO_L1_out_wrapper_147__ap_idle;
  wire C_drain_IO_L1_out_wrapper_148__ap_start;
  wire C_drain_IO_L1_out_wrapper_148__ap_ready;
  wire C_drain_IO_L1_out_wrapper_148__ap_done;
  wire C_drain_IO_L1_out_wrapper_148__ap_idle;
  wire C_drain_IO_L1_out_wrapper_149__ap_start;
  wire C_drain_IO_L1_out_wrapper_149__ap_ready;
  wire C_drain_IO_L1_out_wrapper_149__ap_done;
  wire C_drain_IO_L1_out_wrapper_149__ap_idle;
  wire C_drain_IO_L1_out_wrapper_150__ap_start;
  wire C_drain_IO_L1_out_wrapper_150__ap_ready;
  wire C_drain_IO_L1_out_wrapper_150__ap_done;
  wire C_drain_IO_L1_out_wrapper_150__ap_idle;
  wire C_drain_IO_L1_out_wrapper_151__ap_start;
  wire C_drain_IO_L1_out_wrapper_151__ap_ready;
  wire C_drain_IO_L1_out_wrapper_151__ap_done;
  wire C_drain_IO_L1_out_wrapper_151__ap_idle;
  wire C_drain_IO_L1_out_wrapper_152__ap_start;
  wire C_drain_IO_L1_out_wrapper_152__ap_ready;
  wire C_drain_IO_L1_out_wrapper_152__ap_done;
  wire C_drain_IO_L1_out_wrapper_152__ap_idle;
  wire C_drain_IO_L1_out_wrapper_153__ap_start;
  wire C_drain_IO_L1_out_wrapper_153__ap_ready;
  wire C_drain_IO_L1_out_wrapper_153__ap_done;
  wire C_drain_IO_L1_out_wrapper_153__ap_idle;
  wire C_drain_IO_L1_out_wrapper_154__ap_start;
  wire C_drain_IO_L1_out_wrapper_154__ap_ready;
  wire C_drain_IO_L1_out_wrapper_154__ap_done;
  wire C_drain_IO_L1_out_wrapper_154__ap_idle;
  wire C_drain_IO_L1_out_wrapper_155__ap_start;
  wire C_drain_IO_L1_out_wrapper_155__ap_ready;
  wire C_drain_IO_L1_out_wrapper_155__ap_done;
  wire C_drain_IO_L1_out_wrapper_155__ap_idle;
  wire C_drain_IO_L1_out_wrapper_156__ap_start;
  wire C_drain_IO_L1_out_wrapper_156__ap_ready;
  wire C_drain_IO_L1_out_wrapper_156__ap_done;
  wire C_drain_IO_L1_out_wrapper_156__ap_idle;
  wire C_drain_IO_L1_out_wrapper_157__ap_start;
  wire C_drain_IO_L1_out_wrapper_157__ap_ready;
  wire C_drain_IO_L1_out_wrapper_157__ap_done;
  wire C_drain_IO_L1_out_wrapper_157__ap_idle;
  wire C_drain_IO_L1_out_wrapper_158__ap_start;
  wire C_drain_IO_L1_out_wrapper_158__ap_ready;
  wire C_drain_IO_L1_out_wrapper_158__ap_done;
  wire C_drain_IO_L1_out_wrapper_158__ap_idle;
  wire C_drain_IO_L1_out_wrapper_159__ap_start;
  wire C_drain_IO_L1_out_wrapper_159__ap_ready;
  wire C_drain_IO_L1_out_wrapper_159__ap_done;
  wire C_drain_IO_L1_out_wrapper_159__ap_idle;
  wire C_drain_IO_L1_out_wrapper_160__ap_start;
  wire C_drain_IO_L1_out_wrapper_160__ap_ready;
  wire C_drain_IO_L1_out_wrapper_160__ap_done;
  wire C_drain_IO_L1_out_wrapper_160__ap_idle;
  wire C_drain_IO_L1_out_wrapper_161__ap_start;
  wire C_drain_IO_L1_out_wrapper_161__ap_ready;
  wire C_drain_IO_L1_out_wrapper_161__ap_done;
  wire C_drain_IO_L1_out_wrapper_161__ap_idle;
  wire C_drain_IO_L1_out_wrapper_162__ap_start;
  wire C_drain_IO_L1_out_wrapper_162__ap_ready;
  wire C_drain_IO_L1_out_wrapper_162__ap_done;
  wire C_drain_IO_L1_out_wrapper_162__ap_idle;
  wire C_drain_IO_L1_out_wrapper_163__ap_start;
  wire C_drain_IO_L1_out_wrapper_163__ap_ready;
  wire C_drain_IO_L1_out_wrapper_163__ap_done;
  wire C_drain_IO_L1_out_wrapper_163__ap_idle;
  wire C_drain_IO_L1_out_wrapper_164__ap_start;
  wire C_drain_IO_L1_out_wrapper_164__ap_ready;
  wire C_drain_IO_L1_out_wrapper_164__ap_done;
  wire C_drain_IO_L1_out_wrapper_164__ap_idle;
  wire C_drain_IO_L1_out_wrapper_165__ap_start;
  wire C_drain_IO_L1_out_wrapper_165__ap_ready;
  wire C_drain_IO_L1_out_wrapper_165__ap_done;
  wire C_drain_IO_L1_out_wrapper_165__ap_idle;
  wire C_drain_IO_L1_out_wrapper_166__ap_start;
  wire C_drain_IO_L1_out_wrapper_166__ap_ready;
  wire C_drain_IO_L1_out_wrapper_166__ap_done;
  wire C_drain_IO_L1_out_wrapper_166__ap_idle;
  wire C_drain_IO_L1_out_wrapper_167__ap_start;
  wire C_drain_IO_L1_out_wrapper_167__ap_ready;
  wire C_drain_IO_L1_out_wrapper_167__ap_done;
  wire C_drain_IO_L1_out_wrapper_167__ap_idle;
  wire C_drain_IO_L1_out_wrapper_168__ap_start;
  wire C_drain_IO_L1_out_wrapper_168__ap_ready;
  wire C_drain_IO_L1_out_wrapper_168__ap_done;
  wire C_drain_IO_L1_out_wrapper_168__ap_idle;
  wire C_drain_IO_L1_out_wrapper_169__ap_start;
  wire C_drain_IO_L1_out_wrapper_169__ap_ready;
  wire C_drain_IO_L1_out_wrapper_169__ap_done;
  wire C_drain_IO_L1_out_wrapper_169__ap_idle;
  wire C_drain_IO_L1_out_wrapper_170__ap_start;
  wire C_drain_IO_L1_out_wrapper_170__ap_ready;
  wire C_drain_IO_L1_out_wrapper_170__ap_done;
  wire C_drain_IO_L1_out_wrapper_170__ap_idle;
  wire C_drain_IO_L1_out_wrapper_171__ap_start;
  wire C_drain_IO_L1_out_wrapper_171__ap_ready;
  wire C_drain_IO_L1_out_wrapper_171__ap_done;
  wire C_drain_IO_L1_out_wrapper_171__ap_idle;
  wire C_drain_IO_L1_out_wrapper_172__ap_start;
  wire C_drain_IO_L1_out_wrapper_172__ap_ready;
  wire C_drain_IO_L1_out_wrapper_172__ap_done;
  wire C_drain_IO_L1_out_wrapper_172__ap_idle;
  wire C_drain_IO_L1_out_wrapper_173__ap_start;
  wire C_drain_IO_L1_out_wrapper_173__ap_ready;
  wire C_drain_IO_L1_out_wrapper_173__ap_done;
  wire C_drain_IO_L1_out_wrapper_173__ap_idle;
  wire C_drain_IO_L1_out_wrapper_174__ap_start;
  wire C_drain_IO_L1_out_wrapper_174__ap_ready;
  wire C_drain_IO_L1_out_wrapper_174__ap_done;
  wire C_drain_IO_L1_out_wrapper_174__ap_idle;
  wire C_drain_IO_L1_out_wrapper_175__ap_start;
  wire C_drain_IO_L1_out_wrapper_175__ap_ready;
  wire C_drain_IO_L1_out_wrapper_175__ap_done;
  wire C_drain_IO_L1_out_wrapper_175__ap_idle;
  wire C_drain_IO_L1_out_wrapper_176__ap_start;
  wire C_drain_IO_L1_out_wrapper_176__ap_ready;
  wire C_drain_IO_L1_out_wrapper_176__ap_done;
  wire C_drain_IO_L1_out_wrapper_176__ap_idle;
  wire C_drain_IO_L1_out_wrapper_177__ap_start;
  wire C_drain_IO_L1_out_wrapper_177__ap_ready;
  wire C_drain_IO_L1_out_wrapper_177__ap_done;
  wire C_drain_IO_L1_out_wrapper_177__ap_idle;
  wire C_drain_IO_L1_out_wrapper_178__ap_start;
  wire C_drain_IO_L1_out_wrapper_178__ap_ready;
  wire C_drain_IO_L1_out_wrapper_178__ap_done;
  wire C_drain_IO_L1_out_wrapper_178__ap_idle;
  wire C_drain_IO_L1_out_wrapper_179__ap_start;
  wire C_drain_IO_L1_out_wrapper_179__ap_ready;
  wire C_drain_IO_L1_out_wrapper_179__ap_done;
  wire C_drain_IO_L1_out_wrapper_179__ap_idle;
  wire C_drain_IO_L1_out_wrapper_180__ap_start;
  wire C_drain_IO_L1_out_wrapper_180__ap_ready;
  wire C_drain_IO_L1_out_wrapper_180__ap_done;
  wire C_drain_IO_L1_out_wrapper_180__ap_idle;
  wire C_drain_IO_L1_out_wrapper_181__ap_start;
  wire C_drain_IO_L1_out_wrapper_181__ap_ready;
  wire C_drain_IO_L1_out_wrapper_181__ap_done;
  wire C_drain_IO_L1_out_wrapper_181__ap_idle;
  wire C_drain_IO_L1_out_wrapper_182__ap_start;
  wire C_drain_IO_L1_out_wrapper_182__ap_ready;
  wire C_drain_IO_L1_out_wrapper_182__ap_done;
  wire C_drain_IO_L1_out_wrapper_182__ap_idle;
  wire C_drain_IO_L1_out_wrapper_183__ap_start;
  wire C_drain_IO_L1_out_wrapper_183__ap_ready;
  wire C_drain_IO_L1_out_wrapper_183__ap_done;
  wire C_drain_IO_L1_out_wrapper_183__ap_idle;
  wire C_drain_IO_L1_out_wrapper_184__ap_start;
  wire C_drain_IO_L1_out_wrapper_184__ap_ready;
  wire C_drain_IO_L1_out_wrapper_184__ap_done;
  wire C_drain_IO_L1_out_wrapper_184__ap_idle;
  wire C_drain_IO_L1_out_wrapper_185__ap_start;
  wire C_drain_IO_L1_out_wrapper_185__ap_ready;
  wire C_drain_IO_L1_out_wrapper_185__ap_done;
  wire C_drain_IO_L1_out_wrapper_185__ap_idle;
  wire C_drain_IO_L1_out_wrapper_186__ap_start;
  wire C_drain_IO_L1_out_wrapper_186__ap_ready;
  wire C_drain_IO_L1_out_wrapper_186__ap_done;
  wire C_drain_IO_L1_out_wrapper_186__ap_idle;
  wire C_drain_IO_L1_out_wrapper_187__ap_start;
  wire C_drain_IO_L1_out_wrapper_187__ap_ready;
  wire C_drain_IO_L1_out_wrapper_187__ap_done;
  wire C_drain_IO_L1_out_wrapper_187__ap_idle;
  wire C_drain_IO_L1_out_wrapper_188__ap_start;
  wire C_drain_IO_L1_out_wrapper_188__ap_ready;
  wire C_drain_IO_L1_out_wrapper_188__ap_done;
  wire C_drain_IO_L1_out_wrapper_188__ap_idle;
  wire C_drain_IO_L1_out_wrapper_189__ap_start;
  wire C_drain_IO_L1_out_wrapper_189__ap_ready;
  wire C_drain_IO_L1_out_wrapper_189__ap_done;
  wire C_drain_IO_L1_out_wrapper_189__ap_idle;
  wire C_drain_IO_L1_out_wrapper_190__ap_start;
  wire C_drain_IO_L1_out_wrapper_190__ap_ready;
  wire C_drain_IO_L1_out_wrapper_190__ap_done;
  wire C_drain_IO_L1_out_wrapper_190__ap_idle;
  wire C_drain_IO_L1_out_wrapper_191__ap_start;
  wire C_drain_IO_L1_out_wrapper_191__ap_ready;
  wire C_drain_IO_L1_out_wrapper_191__ap_done;
  wire C_drain_IO_L1_out_wrapper_191__ap_idle;
  wire C_drain_IO_L1_out_wrapper_192__ap_start;
  wire C_drain_IO_L1_out_wrapper_192__ap_ready;
  wire C_drain_IO_L1_out_wrapper_192__ap_done;
  wire C_drain_IO_L1_out_wrapper_192__ap_idle;
  wire C_drain_IO_L1_out_wrapper_193__ap_start;
  wire C_drain_IO_L1_out_wrapper_193__ap_ready;
  wire C_drain_IO_L1_out_wrapper_193__ap_done;
  wire C_drain_IO_L1_out_wrapper_193__ap_idle;
  wire C_drain_IO_L1_out_wrapper_194__ap_start;
  wire C_drain_IO_L1_out_wrapper_194__ap_ready;
  wire C_drain_IO_L1_out_wrapper_194__ap_done;
  wire C_drain_IO_L1_out_wrapper_194__ap_idle;
  wire C_drain_IO_L1_out_wrapper_195__ap_start;
  wire C_drain_IO_L1_out_wrapper_195__ap_ready;
  wire C_drain_IO_L1_out_wrapper_195__ap_done;
  wire C_drain_IO_L1_out_wrapper_195__ap_idle;
  wire C_drain_IO_L1_out_wrapper_196__ap_start;
  wire C_drain_IO_L1_out_wrapper_196__ap_ready;
  wire C_drain_IO_L1_out_wrapper_196__ap_done;
  wire C_drain_IO_L1_out_wrapper_196__ap_idle;
  wire C_drain_IO_L1_out_wrapper_197__ap_start;
  wire C_drain_IO_L1_out_wrapper_197__ap_ready;
  wire C_drain_IO_L1_out_wrapper_197__ap_done;
  wire C_drain_IO_L1_out_wrapper_197__ap_idle;
  wire C_drain_IO_L1_out_wrapper_198__ap_start;
  wire C_drain_IO_L1_out_wrapper_198__ap_ready;
  wire C_drain_IO_L1_out_wrapper_198__ap_done;
  wire C_drain_IO_L1_out_wrapper_198__ap_idle;
  wire C_drain_IO_L1_out_wrapper_199__ap_start;
  wire C_drain_IO_L1_out_wrapper_199__ap_ready;
  wire C_drain_IO_L1_out_wrapper_199__ap_done;
  wire C_drain_IO_L1_out_wrapper_199__ap_idle;
  wire C_drain_IO_L1_out_wrapper_200__ap_start;
  wire C_drain_IO_L1_out_wrapper_200__ap_ready;
  wire C_drain_IO_L1_out_wrapper_200__ap_done;
  wire C_drain_IO_L1_out_wrapper_200__ap_idle;
  wire C_drain_IO_L1_out_wrapper_201__ap_start;
  wire C_drain_IO_L1_out_wrapper_201__ap_ready;
  wire C_drain_IO_L1_out_wrapper_201__ap_done;
  wire C_drain_IO_L1_out_wrapper_201__ap_idle;
  wire C_drain_IO_L1_out_wrapper_202__ap_start;
  wire C_drain_IO_L1_out_wrapper_202__ap_ready;
  wire C_drain_IO_L1_out_wrapper_202__ap_done;
  wire C_drain_IO_L1_out_wrapper_202__ap_idle;
  wire C_drain_IO_L1_out_wrapper_203__ap_start;
  wire C_drain_IO_L1_out_wrapper_203__ap_ready;
  wire C_drain_IO_L1_out_wrapper_203__ap_done;
  wire C_drain_IO_L1_out_wrapper_203__ap_idle;
  wire C_drain_IO_L1_out_wrapper_204__ap_start;
  wire C_drain_IO_L1_out_wrapper_204__ap_ready;
  wire C_drain_IO_L1_out_wrapper_204__ap_done;
  wire C_drain_IO_L1_out_wrapper_204__ap_idle;
  wire C_drain_IO_L1_out_wrapper_205__ap_start;
  wire C_drain_IO_L1_out_wrapper_205__ap_ready;
  wire C_drain_IO_L1_out_wrapper_205__ap_done;
  wire C_drain_IO_L1_out_wrapper_205__ap_idle;
  wire C_drain_IO_L1_out_wrapper_206__ap_start;
  wire C_drain_IO_L1_out_wrapper_206__ap_ready;
  wire C_drain_IO_L1_out_wrapper_206__ap_done;
  wire C_drain_IO_L1_out_wrapper_206__ap_idle;
  wire C_drain_IO_L1_out_wrapper_207__ap_start;
  wire C_drain_IO_L1_out_wrapper_207__ap_ready;
  wire C_drain_IO_L1_out_wrapper_207__ap_done;
  wire C_drain_IO_L1_out_wrapper_207__ap_idle;
  wire C_drain_IO_L1_out_wrapper_208__ap_start;
  wire C_drain_IO_L1_out_wrapper_208__ap_ready;
  wire C_drain_IO_L1_out_wrapper_208__ap_done;
  wire C_drain_IO_L1_out_wrapper_208__ap_idle;
  wire C_drain_IO_L1_out_wrapper_209__ap_start;
  wire C_drain_IO_L1_out_wrapper_209__ap_ready;
  wire C_drain_IO_L1_out_wrapper_209__ap_done;
  wire C_drain_IO_L1_out_wrapper_209__ap_idle;
  wire C_drain_IO_L1_out_wrapper_210__ap_start;
  wire C_drain_IO_L1_out_wrapper_210__ap_ready;
  wire C_drain_IO_L1_out_wrapper_210__ap_done;
  wire C_drain_IO_L1_out_wrapper_210__ap_idle;
  wire C_drain_IO_L1_out_wrapper_211__ap_start;
  wire C_drain_IO_L1_out_wrapper_211__ap_ready;
  wire C_drain_IO_L1_out_wrapper_211__ap_done;
  wire C_drain_IO_L1_out_wrapper_211__ap_idle;
  wire C_drain_IO_L1_out_wrapper_212__ap_start;
  wire C_drain_IO_L1_out_wrapper_212__ap_ready;
  wire C_drain_IO_L1_out_wrapper_212__ap_done;
  wire C_drain_IO_L1_out_wrapper_212__ap_idle;
  wire C_drain_IO_L1_out_wrapper_213__ap_start;
  wire C_drain_IO_L1_out_wrapper_213__ap_ready;
  wire C_drain_IO_L1_out_wrapper_213__ap_done;
  wire C_drain_IO_L1_out_wrapper_213__ap_idle;
  wire C_drain_IO_L1_out_wrapper_214__ap_start;
  wire C_drain_IO_L1_out_wrapper_214__ap_ready;
  wire C_drain_IO_L1_out_wrapper_214__ap_done;
  wire C_drain_IO_L1_out_wrapper_214__ap_idle;
  wire C_drain_IO_L1_out_wrapper_215__ap_start;
  wire C_drain_IO_L1_out_wrapper_215__ap_ready;
  wire C_drain_IO_L1_out_wrapper_215__ap_done;
  wire C_drain_IO_L1_out_wrapper_215__ap_idle;
  wire C_drain_IO_L1_out_wrapper_216__ap_start;
  wire C_drain_IO_L1_out_wrapper_216__ap_ready;
  wire C_drain_IO_L1_out_wrapper_216__ap_done;
  wire C_drain_IO_L1_out_wrapper_216__ap_idle;
  wire C_drain_IO_L1_out_wrapper_217__ap_start;
  wire C_drain_IO_L1_out_wrapper_217__ap_ready;
  wire C_drain_IO_L1_out_wrapper_217__ap_done;
  wire C_drain_IO_L1_out_wrapper_217__ap_idle;
  wire C_drain_IO_L1_out_wrapper_218__ap_start;
  wire C_drain_IO_L1_out_wrapper_218__ap_ready;
  wire C_drain_IO_L1_out_wrapper_218__ap_done;
  wire C_drain_IO_L1_out_wrapper_218__ap_idle;
  wire C_drain_IO_L1_out_wrapper_219__ap_start;
  wire C_drain_IO_L1_out_wrapper_219__ap_ready;
  wire C_drain_IO_L1_out_wrapper_219__ap_done;
  wire C_drain_IO_L1_out_wrapper_219__ap_idle;
  wire C_drain_IO_L1_out_wrapper_220__ap_start;
  wire C_drain_IO_L1_out_wrapper_220__ap_ready;
  wire C_drain_IO_L1_out_wrapper_220__ap_done;
  wire C_drain_IO_L1_out_wrapper_220__ap_idle;
  wire C_drain_IO_L1_out_wrapper_221__ap_start;
  wire C_drain_IO_L1_out_wrapper_221__ap_ready;
  wire C_drain_IO_L1_out_wrapper_221__ap_done;
  wire C_drain_IO_L1_out_wrapper_221__ap_idle;
  wire C_drain_IO_L1_out_wrapper_222__ap_start;
  wire C_drain_IO_L1_out_wrapper_222__ap_ready;
  wire C_drain_IO_L1_out_wrapper_222__ap_done;
  wire C_drain_IO_L1_out_wrapper_222__ap_idle;
  wire C_drain_IO_L1_out_wrapper_223__ap_start;
  wire C_drain_IO_L1_out_wrapper_223__ap_ready;
  wire C_drain_IO_L1_out_wrapper_223__ap_done;
  wire C_drain_IO_L1_out_wrapper_223__ap_idle;
  wire C_drain_IO_L1_out_wrapper_224__ap_start;
  wire C_drain_IO_L1_out_wrapper_224__ap_ready;
  wire C_drain_IO_L1_out_wrapper_224__ap_done;
  wire C_drain_IO_L1_out_wrapper_224__ap_idle;
  wire C_drain_IO_L1_out_wrapper_225__ap_start;
  wire C_drain_IO_L1_out_wrapper_225__ap_ready;
  wire C_drain_IO_L1_out_wrapper_225__ap_done;
  wire C_drain_IO_L1_out_wrapper_225__ap_idle;
  wire C_drain_IO_L1_out_wrapper_226__ap_start;
  wire C_drain_IO_L1_out_wrapper_226__ap_ready;
  wire C_drain_IO_L1_out_wrapper_226__ap_done;
  wire C_drain_IO_L1_out_wrapper_226__ap_idle;
  wire C_drain_IO_L1_out_wrapper_227__ap_start;
  wire C_drain_IO_L1_out_wrapper_227__ap_ready;
  wire C_drain_IO_L1_out_wrapper_227__ap_done;
  wire C_drain_IO_L1_out_wrapper_227__ap_idle;
  wire C_drain_IO_L1_out_wrapper_228__ap_start;
  wire C_drain_IO_L1_out_wrapper_228__ap_ready;
  wire C_drain_IO_L1_out_wrapper_228__ap_done;
  wire C_drain_IO_L1_out_wrapper_228__ap_idle;
  wire C_drain_IO_L1_out_wrapper_229__ap_start;
  wire C_drain_IO_L1_out_wrapper_229__ap_ready;
  wire C_drain_IO_L1_out_wrapper_229__ap_done;
  wire C_drain_IO_L1_out_wrapper_229__ap_idle;
  wire C_drain_IO_L1_out_wrapper_230__ap_start;
  wire C_drain_IO_L1_out_wrapper_230__ap_ready;
  wire C_drain_IO_L1_out_wrapper_230__ap_done;
  wire C_drain_IO_L1_out_wrapper_230__ap_idle;
  wire C_drain_IO_L1_out_wrapper_231__ap_start;
  wire C_drain_IO_L1_out_wrapper_231__ap_ready;
  wire C_drain_IO_L1_out_wrapper_231__ap_done;
  wire C_drain_IO_L1_out_wrapper_231__ap_idle;
  wire C_drain_IO_L1_out_wrapper_232__ap_start;
  wire C_drain_IO_L1_out_wrapper_232__ap_ready;
  wire C_drain_IO_L1_out_wrapper_232__ap_done;
  wire C_drain_IO_L1_out_wrapper_232__ap_idle;
  wire C_drain_IO_L1_out_wrapper_233__ap_start;
  wire C_drain_IO_L1_out_wrapper_233__ap_ready;
  wire C_drain_IO_L1_out_wrapper_233__ap_done;
  wire C_drain_IO_L1_out_wrapper_233__ap_idle;
  wire C_drain_IO_L1_out_wrapper_234__ap_start;
  wire C_drain_IO_L1_out_wrapper_234__ap_ready;
  wire C_drain_IO_L1_out_wrapper_234__ap_done;
  wire C_drain_IO_L1_out_wrapper_234__ap_idle;
  wire C_drain_IO_L1_out_wrapper_235__ap_start;
  wire C_drain_IO_L1_out_wrapper_235__ap_ready;
  wire C_drain_IO_L1_out_wrapper_235__ap_done;
  wire C_drain_IO_L1_out_wrapper_235__ap_idle;
  wire C_drain_IO_L1_out_wrapper_236__ap_start;
  wire C_drain_IO_L1_out_wrapper_236__ap_ready;
  wire C_drain_IO_L1_out_wrapper_236__ap_done;
  wire C_drain_IO_L1_out_wrapper_236__ap_idle;
  wire C_drain_IO_L1_out_wrapper_237__ap_start;
  wire C_drain_IO_L1_out_wrapper_237__ap_ready;
  wire C_drain_IO_L1_out_wrapper_237__ap_done;
  wire C_drain_IO_L1_out_wrapper_237__ap_idle;
  wire C_drain_IO_L1_out_wrapper_238__ap_start;
  wire C_drain_IO_L1_out_wrapper_238__ap_ready;
  wire C_drain_IO_L1_out_wrapper_238__ap_done;
  wire C_drain_IO_L1_out_wrapper_238__ap_idle;
  wire C_drain_IO_L1_out_wrapper_239__ap_start;
  wire C_drain_IO_L1_out_wrapper_239__ap_ready;
  wire C_drain_IO_L1_out_wrapper_239__ap_done;
  wire C_drain_IO_L1_out_wrapper_239__ap_idle;
  wire C_drain_IO_L1_out_wrapper_240__ap_start;
  wire C_drain_IO_L1_out_wrapper_240__ap_ready;
  wire C_drain_IO_L1_out_wrapper_240__ap_done;
  wire C_drain_IO_L1_out_wrapper_240__ap_idle;
  wire C_drain_IO_L1_out_wrapper_241__ap_start;
  wire C_drain_IO_L1_out_wrapper_241__ap_ready;
  wire C_drain_IO_L1_out_wrapper_241__ap_done;
  wire C_drain_IO_L1_out_wrapper_241__ap_idle;
  wire C_drain_IO_L1_out_wrapper_242__ap_start;
  wire C_drain_IO_L1_out_wrapper_242__ap_ready;
  wire C_drain_IO_L1_out_wrapper_242__ap_done;
  wire C_drain_IO_L1_out_wrapper_242__ap_idle;
  wire C_drain_IO_L1_out_wrapper_243__ap_start;
  wire C_drain_IO_L1_out_wrapper_243__ap_ready;
  wire C_drain_IO_L1_out_wrapper_243__ap_done;
  wire C_drain_IO_L1_out_wrapper_243__ap_idle;
  wire C_drain_IO_L1_out_wrapper_244__ap_start;
  wire C_drain_IO_L1_out_wrapper_244__ap_ready;
  wire C_drain_IO_L1_out_wrapper_244__ap_done;
  wire C_drain_IO_L1_out_wrapper_244__ap_idle;
  wire C_drain_IO_L1_out_wrapper_245__ap_start;
  wire C_drain_IO_L1_out_wrapper_245__ap_ready;
  wire C_drain_IO_L1_out_wrapper_245__ap_done;
  wire C_drain_IO_L1_out_wrapper_245__ap_idle;
  wire C_drain_IO_L1_out_wrapper_246__ap_start;
  wire C_drain_IO_L1_out_wrapper_246__ap_ready;
  wire C_drain_IO_L1_out_wrapper_246__ap_done;
  wire C_drain_IO_L1_out_wrapper_246__ap_idle;
  wire C_drain_IO_L1_out_wrapper_247__ap_start;
  wire C_drain_IO_L1_out_wrapper_247__ap_ready;
  wire C_drain_IO_L1_out_wrapper_247__ap_done;
  wire C_drain_IO_L1_out_wrapper_247__ap_idle;
  wire C_drain_IO_L1_out_wrapper_248__ap_start;
  wire C_drain_IO_L1_out_wrapper_248__ap_ready;
  wire C_drain_IO_L1_out_wrapper_248__ap_done;
  wire C_drain_IO_L1_out_wrapper_248__ap_idle;
  wire C_drain_IO_L1_out_wrapper_249__ap_start;
  wire C_drain_IO_L1_out_wrapper_249__ap_ready;
  wire C_drain_IO_L1_out_wrapper_249__ap_done;
  wire C_drain_IO_L1_out_wrapper_249__ap_idle;
  wire C_drain_IO_L1_out_wrapper_250__ap_start;
  wire C_drain_IO_L1_out_wrapper_250__ap_ready;
  wire C_drain_IO_L1_out_wrapper_250__ap_done;
  wire C_drain_IO_L1_out_wrapper_250__ap_idle;
  wire C_drain_IO_L1_out_wrapper_251__ap_start;
  wire C_drain_IO_L1_out_wrapper_251__ap_ready;
  wire C_drain_IO_L1_out_wrapper_251__ap_done;
  wire C_drain_IO_L1_out_wrapper_251__ap_idle;
  wire C_drain_IO_L1_out_wrapper_252__ap_start;
  wire C_drain_IO_L1_out_wrapper_252__ap_ready;
  wire C_drain_IO_L1_out_wrapper_252__ap_done;
  wire C_drain_IO_L1_out_wrapper_252__ap_idle;
  wire C_drain_IO_L1_out_wrapper_253__ap_start;
  wire C_drain_IO_L1_out_wrapper_253__ap_ready;
  wire C_drain_IO_L1_out_wrapper_253__ap_done;
  wire C_drain_IO_L1_out_wrapper_253__ap_idle;
  wire C_drain_IO_L1_out_wrapper_254__ap_start;
  wire C_drain_IO_L1_out_wrapper_254__ap_ready;
  wire C_drain_IO_L1_out_wrapper_254__ap_done;
  wire C_drain_IO_L1_out_wrapper_254__ap_idle;
  wire C_drain_IO_L1_out_wrapper_255__ap_start;
  wire C_drain_IO_L1_out_wrapper_255__ap_ready;
  wire C_drain_IO_L1_out_wrapper_255__ap_done;
  wire C_drain_IO_L1_out_wrapper_255__ap_idle;
  wire C_drain_IO_L1_out_wrapper_256__ap_start;
  wire C_drain_IO_L1_out_wrapper_256__ap_ready;
  wire C_drain_IO_L1_out_wrapper_256__ap_done;
  wire C_drain_IO_L1_out_wrapper_256__ap_idle;
  wire C_drain_IO_L1_out_wrapper_257__ap_start;
  wire C_drain_IO_L1_out_wrapper_257__ap_ready;
  wire C_drain_IO_L1_out_wrapper_257__ap_done;
  wire C_drain_IO_L1_out_wrapper_257__ap_idle;
  wire C_drain_IO_L1_out_wrapper_258__ap_start;
  wire C_drain_IO_L1_out_wrapper_258__ap_ready;
  wire C_drain_IO_L1_out_wrapper_258__ap_done;
  wire C_drain_IO_L1_out_wrapper_258__ap_idle;
  wire C_drain_IO_L1_out_wrapper_259__ap_start;
  wire C_drain_IO_L1_out_wrapper_259__ap_ready;
  wire C_drain_IO_L1_out_wrapper_259__ap_done;
  wire C_drain_IO_L1_out_wrapper_259__ap_idle;
  wire C_drain_IO_L1_out_wrapper_260__ap_start;
  wire C_drain_IO_L1_out_wrapper_260__ap_ready;
  wire C_drain_IO_L1_out_wrapper_260__ap_done;
  wire C_drain_IO_L1_out_wrapper_260__ap_idle;
  wire C_drain_IO_L1_out_wrapper_261__ap_start;
  wire C_drain_IO_L1_out_wrapper_261__ap_ready;
  wire C_drain_IO_L1_out_wrapper_261__ap_done;
  wire C_drain_IO_L1_out_wrapper_261__ap_idle;
  wire C_drain_IO_L1_out_wrapper_262__ap_start;
  wire C_drain_IO_L1_out_wrapper_262__ap_ready;
  wire C_drain_IO_L1_out_wrapper_262__ap_done;
  wire C_drain_IO_L1_out_wrapper_262__ap_idle;
  wire C_drain_IO_L1_out_wrapper_263__ap_start;
  wire C_drain_IO_L1_out_wrapper_263__ap_ready;
  wire C_drain_IO_L1_out_wrapper_263__ap_done;
  wire C_drain_IO_L1_out_wrapper_263__ap_idle;
  wire C_drain_IO_L1_out_wrapper_264__ap_start;
  wire C_drain_IO_L1_out_wrapper_264__ap_ready;
  wire C_drain_IO_L1_out_wrapper_264__ap_done;
  wire C_drain_IO_L1_out_wrapper_264__ap_idle;
  wire C_drain_IO_L1_out_wrapper_265__ap_start;
  wire C_drain_IO_L1_out_wrapper_265__ap_ready;
  wire C_drain_IO_L1_out_wrapper_265__ap_done;
  wire C_drain_IO_L1_out_wrapper_265__ap_idle;
  wire C_drain_IO_L1_out_wrapper_266__ap_start;
  wire C_drain_IO_L1_out_wrapper_266__ap_ready;
  wire C_drain_IO_L1_out_wrapper_266__ap_done;
  wire C_drain_IO_L1_out_wrapper_266__ap_idle;
  wire C_drain_IO_L1_out_wrapper_267__ap_start;
  wire C_drain_IO_L1_out_wrapper_267__ap_ready;
  wire C_drain_IO_L1_out_wrapper_267__ap_done;
  wire C_drain_IO_L1_out_wrapper_267__ap_idle;
  wire C_drain_IO_L1_out_wrapper_268__ap_start;
  wire C_drain_IO_L1_out_wrapper_268__ap_ready;
  wire C_drain_IO_L1_out_wrapper_268__ap_done;
  wire C_drain_IO_L1_out_wrapper_268__ap_idle;
  wire C_drain_IO_L1_out_wrapper_269__ap_start;
  wire C_drain_IO_L1_out_wrapper_269__ap_ready;
  wire C_drain_IO_L1_out_wrapper_269__ap_done;
  wire C_drain_IO_L1_out_wrapper_269__ap_idle;
  wire C_drain_IO_L1_out_wrapper_270__ap_start;
  wire C_drain_IO_L1_out_wrapper_270__ap_ready;
  wire C_drain_IO_L1_out_wrapper_270__ap_done;
  wire C_drain_IO_L1_out_wrapper_270__ap_idle;
  wire C_drain_IO_L1_out_wrapper_271__ap_start;
  wire C_drain_IO_L1_out_wrapper_271__ap_ready;
  wire C_drain_IO_L1_out_wrapper_271__ap_done;
  wire C_drain_IO_L1_out_wrapper_271__ap_idle;
  wire C_drain_IO_L1_out_wrapper_272__ap_start;
  wire C_drain_IO_L1_out_wrapper_272__ap_ready;
  wire C_drain_IO_L1_out_wrapper_272__ap_done;
  wire C_drain_IO_L1_out_wrapper_272__ap_idle;
  wire C_drain_IO_L1_out_wrapper_273__ap_start;
  wire C_drain_IO_L1_out_wrapper_273__ap_ready;
  wire C_drain_IO_L1_out_wrapper_273__ap_done;
  wire C_drain_IO_L1_out_wrapper_273__ap_idle;
  wire C_drain_IO_L1_out_wrapper_274__ap_start;
  wire C_drain_IO_L1_out_wrapper_274__ap_ready;
  wire C_drain_IO_L1_out_wrapper_274__ap_done;
  wire C_drain_IO_L1_out_wrapper_274__ap_idle;
  wire C_drain_IO_L1_out_wrapper_275__ap_start;
  wire C_drain_IO_L1_out_wrapper_275__ap_ready;
  wire C_drain_IO_L1_out_wrapper_275__ap_done;
  wire C_drain_IO_L1_out_wrapper_275__ap_idle;
  wire C_drain_IO_L1_out_wrapper_276__ap_start;
  wire C_drain_IO_L1_out_wrapper_276__ap_ready;
  wire C_drain_IO_L1_out_wrapper_276__ap_done;
  wire C_drain_IO_L1_out_wrapper_276__ap_idle;
  wire C_drain_IO_L1_out_wrapper_277__ap_start;
  wire C_drain_IO_L1_out_wrapper_277__ap_ready;
  wire C_drain_IO_L1_out_wrapper_277__ap_done;
  wire C_drain_IO_L1_out_wrapper_277__ap_idle;
  wire C_drain_IO_L1_out_wrapper_278__ap_start;
  wire C_drain_IO_L1_out_wrapper_278__ap_ready;
  wire C_drain_IO_L1_out_wrapper_278__ap_done;
  wire C_drain_IO_L1_out_wrapper_278__ap_idle;
  wire C_drain_IO_L1_out_wrapper_279__ap_start;
  wire C_drain_IO_L1_out_wrapper_279__ap_ready;
  wire C_drain_IO_L1_out_wrapper_279__ap_done;
  wire C_drain_IO_L1_out_wrapper_279__ap_idle;
  wire C_drain_IO_L1_out_wrapper_280__ap_start;
  wire C_drain_IO_L1_out_wrapper_280__ap_ready;
  wire C_drain_IO_L1_out_wrapper_280__ap_done;
  wire C_drain_IO_L1_out_wrapper_280__ap_idle;
  wire C_drain_IO_L1_out_wrapper_281__ap_start;
  wire C_drain_IO_L1_out_wrapper_281__ap_ready;
  wire C_drain_IO_L1_out_wrapper_281__ap_done;
  wire C_drain_IO_L1_out_wrapper_281__ap_idle;
  wire C_drain_IO_L1_out_wrapper_282__ap_start;
  wire C_drain_IO_L1_out_wrapper_282__ap_ready;
  wire C_drain_IO_L1_out_wrapper_282__ap_done;
  wire C_drain_IO_L1_out_wrapper_282__ap_idle;
  wire C_drain_IO_L1_out_wrapper_283__ap_start;
  wire C_drain_IO_L1_out_wrapper_283__ap_ready;
  wire C_drain_IO_L1_out_wrapper_283__ap_done;
  wire C_drain_IO_L1_out_wrapper_283__ap_idle;
  wire C_drain_IO_L1_out_wrapper_284__ap_start;
  wire C_drain_IO_L1_out_wrapper_284__ap_ready;
  wire C_drain_IO_L1_out_wrapper_284__ap_done;
  wire C_drain_IO_L1_out_wrapper_284__ap_idle;
  wire C_drain_IO_L1_out_wrapper_285__ap_start;
  wire C_drain_IO_L1_out_wrapper_285__ap_ready;
  wire C_drain_IO_L1_out_wrapper_285__ap_done;
  wire C_drain_IO_L1_out_wrapper_285__ap_idle;
  wire C_drain_IO_L1_out_wrapper_286__ap_start;
  wire C_drain_IO_L1_out_wrapper_286__ap_ready;
  wire C_drain_IO_L1_out_wrapper_286__ap_done;
  wire C_drain_IO_L1_out_wrapper_286__ap_idle;
  wire C_drain_IO_L1_out_wrapper_287__ap_start;
  wire C_drain_IO_L1_out_wrapper_287__ap_ready;
  wire C_drain_IO_L1_out_wrapper_287__ap_done;
  wire C_drain_IO_L1_out_wrapper_287__ap_idle;
  wire C_drain_IO_L1_out_wrapper_288__ap_start;
  wire C_drain_IO_L1_out_wrapper_288__ap_ready;
  wire C_drain_IO_L1_out_wrapper_288__ap_done;
  wire C_drain_IO_L1_out_wrapper_288__ap_idle;
  wire C_drain_IO_L2_out_0__ap_start;
  wire C_drain_IO_L2_out_0__ap_ready;
  wire C_drain_IO_L2_out_0__ap_done;
  wire C_drain_IO_L2_out_0__ap_idle;
  wire C_drain_IO_L2_out_1__ap_start;
  wire C_drain_IO_L2_out_1__ap_ready;
  wire C_drain_IO_L2_out_1__ap_done;
  wire C_drain_IO_L2_out_1__ap_idle;
  wire C_drain_IO_L2_out_2__ap_start;
  wire C_drain_IO_L2_out_2__ap_ready;
  wire C_drain_IO_L2_out_2__ap_done;
  wire C_drain_IO_L2_out_2__ap_idle;
  wire C_drain_IO_L2_out_3__ap_start;
  wire C_drain_IO_L2_out_3__ap_ready;
  wire C_drain_IO_L2_out_3__ap_done;
  wire C_drain_IO_L2_out_3__ap_idle;
  wire C_drain_IO_L2_out_4__ap_start;
  wire C_drain_IO_L2_out_4__ap_ready;
  wire C_drain_IO_L2_out_4__ap_done;
  wire C_drain_IO_L2_out_4__ap_idle;
  wire C_drain_IO_L2_out_5__ap_start;
  wire C_drain_IO_L2_out_5__ap_ready;
  wire C_drain_IO_L2_out_5__ap_done;
  wire C_drain_IO_L2_out_5__ap_idle;
  wire C_drain_IO_L2_out_6__ap_start;
  wire C_drain_IO_L2_out_6__ap_ready;
  wire C_drain_IO_L2_out_6__ap_done;
  wire C_drain_IO_L2_out_6__ap_idle;
  wire C_drain_IO_L2_out_7__ap_start;
  wire C_drain_IO_L2_out_7__ap_ready;
  wire C_drain_IO_L2_out_7__ap_done;
  wire C_drain_IO_L2_out_7__ap_idle;
  wire C_drain_IO_L2_out_8__ap_start;
  wire C_drain_IO_L2_out_8__ap_ready;
  wire C_drain_IO_L2_out_8__ap_done;
  wire C_drain_IO_L2_out_8__ap_idle;
  wire C_drain_IO_L2_out_9__ap_start;
  wire C_drain_IO_L2_out_9__ap_ready;
  wire C_drain_IO_L2_out_9__ap_done;
  wire C_drain_IO_L2_out_9__ap_idle;
  wire C_drain_IO_L2_out_10__ap_start;
  wire C_drain_IO_L2_out_10__ap_ready;
  wire C_drain_IO_L2_out_10__ap_done;
  wire C_drain_IO_L2_out_10__ap_idle;
  wire C_drain_IO_L2_out_11__ap_start;
  wire C_drain_IO_L2_out_11__ap_ready;
  wire C_drain_IO_L2_out_11__ap_done;
  wire C_drain_IO_L2_out_11__ap_idle;
  wire C_drain_IO_L2_out_12__ap_start;
  wire C_drain_IO_L2_out_12__ap_ready;
  wire C_drain_IO_L2_out_12__ap_done;
  wire C_drain_IO_L2_out_12__ap_idle;
  wire C_drain_IO_L2_out_13__ap_start;
  wire C_drain_IO_L2_out_13__ap_ready;
  wire C_drain_IO_L2_out_13__ap_done;
  wire C_drain_IO_L2_out_13__ap_idle;
  wire C_drain_IO_L2_out_14__ap_start;
  wire C_drain_IO_L2_out_14__ap_ready;
  wire C_drain_IO_L2_out_14__ap_done;
  wire C_drain_IO_L2_out_14__ap_idle;
  wire C_drain_IO_L2_out_15__ap_start;
  wire C_drain_IO_L2_out_15__ap_ready;
  wire C_drain_IO_L2_out_15__ap_done;
  wire C_drain_IO_L2_out_15__ap_idle;
  wire C_drain_IO_L2_out_boundary_0__ap_start;
  wire C_drain_IO_L2_out_boundary_0__ap_ready;
  wire C_drain_IO_L2_out_boundary_0__ap_done;
  wire C_drain_IO_L2_out_boundary_0__ap_idle;
  wire C_drain_IO_L3_out_0__ap_start;
  wire C_drain_IO_L3_out_0__ap_ready;
  wire C_drain_IO_L3_out_0__ap_done;
  wire C_drain_IO_L3_out_0__ap_idle;
  wire [63:0] C_drain_IO_L3_out_serialize_0___C__q0;
  wire C_drain_IO_L3_out_serialize_0__ap_start;
  wire C_drain_IO_L3_out_serialize_0__ap_ready;
  wire C_drain_IO_L3_out_serialize_0__ap_done;
  wire C_drain_IO_L3_out_serialize_0__ap_idle;
  wire PE_wrapper_0__ap_start;
  wire PE_wrapper_0__ap_ready;
  wire PE_wrapper_0__ap_done;
  wire PE_wrapper_0__ap_idle;
  wire PE_wrapper_1__ap_start;
  wire PE_wrapper_1__ap_ready;
  wire PE_wrapper_1__ap_done;
  wire PE_wrapper_1__ap_idle;
  wire PE_wrapper_2__ap_start;
  wire PE_wrapper_2__ap_ready;
  wire PE_wrapper_2__ap_done;
  wire PE_wrapper_2__ap_idle;
  wire PE_wrapper_3__ap_start;
  wire PE_wrapper_3__ap_ready;
  wire PE_wrapper_3__ap_done;
  wire PE_wrapper_3__ap_idle;
  wire PE_wrapper_4__ap_start;
  wire PE_wrapper_4__ap_ready;
  wire PE_wrapper_4__ap_done;
  wire PE_wrapper_4__ap_idle;
  wire PE_wrapper_5__ap_start;
  wire PE_wrapper_5__ap_ready;
  wire PE_wrapper_5__ap_done;
  wire PE_wrapper_5__ap_idle;
  wire PE_wrapper_6__ap_start;
  wire PE_wrapper_6__ap_ready;
  wire PE_wrapper_6__ap_done;
  wire PE_wrapper_6__ap_idle;
  wire PE_wrapper_7__ap_start;
  wire PE_wrapper_7__ap_ready;
  wire PE_wrapper_7__ap_done;
  wire PE_wrapper_7__ap_idle;
  wire PE_wrapper_8__ap_start;
  wire PE_wrapper_8__ap_ready;
  wire PE_wrapper_8__ap_done;
  wire PE_wrapper_8__ap_idle;
  wire PE_wrapper_9__ap_start;
  wire PE_wrapper_9__ap_ready;
  wire PE_wrapper_9__ap_done;
  wire PE_wrapper_9__ap_idle;
  wire PE_wrapper_10__ap_start;
  wire PE_wrapper_10__ap_ready;
  wire PE_wrapper_10__ap_done;
  wire PE_wrapper_10__ap_idle;
  wire PE_wrapper_11__ap_start;
  wire PE_wrapper_11__ap_ready;
  wire PE_wrapper_11__ap_done;
  wire PE_wrapper_11__ap_idle;
  wire PE_wrapper_12__ap_start;
  wire PE_wrapper_12__ap_ready;
  wire PE_wrapper_12__ap_done;
  wire PE_wrapper_12__ap_idle;
  wire PE_wrapper_13__ap_start;
  wire PE_wrapper_13__ap_ready;
  wire PE_wrapper_13__ap_done;
  wire PE_wrapper_13__ap_idle;
  wire PE_wrapper_14__ap_start;
  wire PE_wrapper_14__ap_ready;
  wire PE_wrapper_14__ap_done;
  wire PE_wrapper_14__ap_idle;
  wire PE_wrapper_15__ap_start;
  wire PE_wrapper_15__ap_ready;
  wire PE_wrapper_15__ap_done;
  wire PE_wrapper_15__ap_idle;
  wire PE_wrapper_16__ap_start;
  wire PE_wrapper_16__ap_ready;
  wire PE_wrapper_16__ap_done;
  wire PE_wrapper_16__ap_idle;
  wire PE_wrapper_17__ap_start;
  wire PE_wrapper_17__ap_ready;
  wire PE_wrapper_17__ap_done;
  wire PE_wrapper_17__ap_idle;
  wire PE_wrapper_18__ap_start;
  wire PE_wrapper_18__ap_ready;
  wire PE_wrapper_18__ap_done;
  wire PE_wrapper_18__ap_idle;
  wire PE_wrapper_19__ap_start;
  wire PE_wrapper_19__ap_ready;
  wire PE_wrapper_19__ap_done;
  wire PE_wrapper_19__ap_idle;
  wire PE_wrapper_20__ap_start;
  wire PE_wrapper_20__ap_ready;
  wire PE_wrapper_20__ap_done;
  wire PE_wrapper_20__ap_idle;
  wire PE_wrapper_21__ap_start;
  wire PE_wrapper_21__ap_ready;
  wire PE_wrapper_21__ap_done;
  wire PE_wrapper_21__ap_idle;
  wire PE_wrapper_22__ap_start;
  wire PE_wrapper_22__ap_ready;
  wire PE_wrapper_22__ap_done;
  wire PE_wrapper_22__ap_idle;
  wire PE_wrapper_23__ap_start;
  wire PE_wrapper_23__ap_ready;
  wire PE_wrapper_23__ap_done;
  wire PE_wrapper_23__ap_idle;
  wire PE_wrapper_24__ap_start;
  wire PE_wrapper_24__ap_ready;
  wire PE_wrapper_24__ap_done;
  wire PE_wrapper_24__ap_idle;
  wire PE_wrapper_25__ap_start;
  wire PE_wrapper_25__ap_ready;
  wire PE_wrapper_25__ap_done;
  wire PE_wrapper_25__ap_idle;
  wire PE_wrapper_26__ap_start;
  wire PE_wrapper_26__ap_ready;
  wire PE_wrapper_26__ap_done;
  wire PE_wrapper_26__ap_idle;
  wire PE_wrapper_27__ap_start;
  wire PE_wrapper_27__ap_ready;
  wire PE_wrapper_27__ap_done;
  wire PE_wrapper_27__ap_idle;
  wire PE_wrapper_28__ap_start;
  wire PE_wrapper_28__ap_ready;
  wire PE_wrapper_28__ap_done;
  wire PE_wrapper_28__ap_idle;
  wire PE_wrapper_29__ap_start;
  wire PE_wrapper_29__ap_ready;
  wire PE_wrapper_29__ap_done;
  wire PE_wrapper_29__ap_idle;
  wire PE_wrapper_30__ap_start;
  wire PE_wrapper_30__ap_ready;
  wire PE_wrapper_30__ap_done;
  wire PE_wrapper_30__ap_idle;
  wire PE_wrapper_31__ap_start;
  wire PE_wrapper_31__ap_ready;
  wire PE_wrapper_31__ap_done;
  wire PE_wrapper_31__ap_idle;
  wire PE_wrapper_32__ap_start;
  wire PE_wrapper_32__ap_ready;
  wire PE_wrapper_32__ap_done;
  wire PE_wrapper_32__ap_idle;
  wire PE_wrapper_33__ap_start;
  wire PE_wrapper_33__ap_ready;
  wire PE_wrapper_33__ap_done;
  wire PE_wrapper_33__ap_idle;
  wire PE_wrapper_34__ap_start;
  wire PE_wrapper_34__ap_ready;
  wire PE_wrapper_34__ap_done;
  wire PE_wrapper_34__ap_idle;
  wire PE_wrapper_35__ap_start;
  wire PE_wrapper_35__ap_ready;
  wire PE_wrapper_35__ap_done;
  wire PE_wrapper_35__ap_idle;
  wire PE_wrapper_36__ap_start;
  wire PE_wrapper_36__ap_ready;
  wire PE_wrapper_36__ap_done;
  wire PE_wrapper_36__ap_idle;
  wire PE_wrapper_37__ap_start;
  wire PE_wrapper_37__ap_ready;
  wire PE_wrapper_37__ap_done;
  wire PE_wrapper_37__ap_idle;
  wire PE_wrapper_38__ap_start;
  wire PE_wrapper_38__ap_ready;
  wire PE_wrapper_38__ap_done;
  wire PE_wrapper_38__ap_idle;
  wire PE_wrapper_39__ap_start;
  wire PE_wrapper_39__ap_ready;
  wire PE_wrapper_39__ap_done;
  wire PE_wrapper_39__ap_idle;
  wire PE_wrapper_40__ap_start;
  wire PE_wrapper_40__ap_ready;
  wire PE_wrapper_40__ap_done;
  wire PE_wrapper_40__ap_idle;
  wire PE_wrapper_41__ap_start;
  wire PE_wrapper_41__ap_ready;
  wire PE_wrapper_41__ap_done;
  wire PE_wrapper_41__ap_idle;
  wire PE_wrapper_42__ap_start;
  wire PE_wrapper_42__ap_ready;
  wire PE_wrapper_42__ap_done;
  wire PE_wrapper_42__ap_idle;
  wire PE_wrapper_43__ap_start;
  wire PE_wrapper_43__ap_ready;
  wire PE_wrapper_43__ap_done;
  wire PE_wrapper_43__ap_idle;
  wire PE_wrapper_44__ap_start;
  wire PE_wrapper_44__ap_ready;
  wire PE_wrapper_44__ap_done;
  wire PE_wrapper_44__ap_idle;
  wire PE_wrapper_45__ap_start;
  wire PE_wrapper_45__ap_ready;
  wire PE_wrapper_45__ap_done;
  wire PE_wrapper_45__ap_idle;
  wire PE_wrapper_46__ap_start;
  wire PE_wrapper_46__ap_ready;
  wire PE_wrapper_46__ap_done;
  wire PE_wrapper_46__ap_idle;
  wire PE_wrapper_47__ap_start;
  wire PE_wrapper_47__ap_ready;
  wire PE_wrapper_47__ap_done;
  wire PE_wrapper_47__ap_idle;
  wire PE_wrapper_48__ap_start;
  wire PE_wrapper_48__ap_ready;
  wire PE_wrapper_48__ap_done;
  wire PE_wrapper_48__ap_idle;
  wire PE_wrapper_49__ap_start;
  wire PE_wrapper_49__ap_ready;
  wire PE_wrapper_49__ap_done;
  wire PE_wrapper_49__ap_idle;
  wire PE_wrapper_50__ap_start;
  wire PE_wrapper_50__ap_ready;
  wire PE_wrapper_50__ap_done;
  wire PE_wrapper_50__ap_idle;
  wire PE_wrapper_51__ap_start;
  wire PE_wrapper_51__ap_ready;
  wire PE_wrapper_51__ap_done;
  wire PE_wrapper_51__ap_idle;
  wire PE_wrapper_52__ap_start;
  wire PE_wrapper_52__ap_ready;
  wire PE_wrapper_52__ap_done;
  wire PE_wrapper_52__ap_idle;
  wire PE_wrapper_53__ap_start;
  wire PE_wrapper_53__ap_ready;
  wire PE_wrapper_53__ap_done;
  wire PE_wrapper_53__ap_idle;
  wire PE_wrapper_54__ap_start;
  wire PE_wrapper_54__ap_ready;
  wire PE_wrapper_54__ap_done;
  wire PE_wrapper_54__ap_idle;
  wire PE_wrapper_55__ap_start;
  wire PE_wrapper_55__ap_ready;
  wire PE_wrapper_55__ap_done;
  wire PE_wrapper_55__ap_idle;
  wire PE_wrapper_56__ap_start;
  wire PE_wrapper_56__ap_ready;
  wire PE_wrapper_56__ap_done;
  wire PE_wrapper_56__ap_idle;
  wire PE_wrapper_57__ap_start;
  wire PE_wrapper_57__ap_ready;
  wire PE_wrapper_57__ap_done;
  wire PE_wrapper_57__ap_idle;
  wire PE_wrapper_58__ap_start;
  wire PE_wrapper_58__ap_ready;
  wire PE_wrapper_58__ap_done;
  wire PE_wrapper_58__ap_idle;
  wire PE_wrapper_59__ap_start;
  wire PE_wrapper_59__ap_ready;
  wire PE_wrapper_59__ap_done;
  wire PE_wrapper_59__ap_idle;
  wire PE_wrapper_60__ap_start;
  wire PE_wrapper_60__ap_ready;
  wire PE_wrapper_60__ap_done;
  wire PE_wrapper_60__ap_idle;
  wire PE_wrapper_61__ap_start;
  wire PE_wrapper_61__ap_ready;
  wire PE_wrapper_61__ap_done;
  wire PE_wrapper_61__ap_idle;
  wire PE_wrapper_62__ap_start;
  wire PE_wrapper_62__ap_ready;
  wire PE_wrapper_62__ap_done;
  wire PE_wrapper_62__ap_idle;
  wire PE_wrapper_63__ap_start;
  wire PE_wrapper_63__ap_ready;
  wire PE_wrapper_63__ap_done;
  wire PE_wrapper_63__ap_idle;
  wire PE_wrapper_64__ap_start;
  wire PE_wrapper_64__ap_ready;
  wire PE_wrapper_64__ap_done;
  wire PE_wrapper_64__ap_idle;
  wire PE_wrapper_65__ap_start;
  wire PE_wrapper_65__ap_ready;
  wire PE_wrapper_65__ap_done;
  wire PE_wrapper_65__ap_idle;
  wire PE_wrapper_66__ap_start;
  wire PE_wrapper_66__ap_ready;
  wire PE_wrapper_66__ap_done;
  wire PE_wrapper_66__ap_idle;
  wire PE_wrapper_67__ap_start;
  wire PE_wrapper_67__ap_ready;
  wire PE_wrapper_67__ap_done;
  wire PE_wrapper_67__ap_idle;
  wire PE_wrapper_68__ap_start;
  wire PE_wrapper_68__ap_ready;
  wire PE_wrapper_68__ap_done;
  wire PE_wrapper_68__ap_idle;
  wire PE_wrapper_69__ap_start;
  wire PE_wrapper_69__ap_ready;
  wire PE_wrapper_69__ap_done;
  wire PE_wrapper_69__ap_idle;
  wire PE_wrapper_70__ap_start;
  wire PE_wrapper_70__ap_ready;
  wire PE_wrapper_70__ap_done;
  wire PE_wrapper_70__ap_idle;
  wire PE_wrapper_71__ap_start;
  wire PE_wrapper_71__ap_ready;
  wire PE_wrapper_71__ap_done;
  wire PE_wrapper_71__ap_idle;
  wire PE_wrapper_72__ap_start;
  wire PE_wrapper_72__ap_ready;
  wire PE_wrapper_72__ap_done;
  wire PE_wrapper_72__ap_idle;
  wire PE_wrapper_73__ap_start;
  wire PE_wrapper_73__ap_ready;
  wire PE_wrapper_73__ap_done;
  wire PE_wrapper_73__ap_idle;
  wire PE_wrapper_74__ap_start;
  wire PE_wrapper_74__ap_ready;
  wire PE_wrapper_74__ap_done;
  wire PE_wrapper_74__ap_idle;
  wire PE_wrapper_75__ap_start;
  wire PE_wrapper_75__ap_ready;
  wire PE_wrapper_75__ap_done;
  wire PE_wrapper_75__ap_idle;
  wire PE_wrapper_76__ap_start;
  wire PE_wrapper_76__ap_ready;
  wire PE_wrapper_76__ap_done;
  wire PE_wrapper_76__ap_idle;
  wire PE_wrapper_77__ap_start;
  wire PE_wrapper_77__ap_ready;
  wire PE_wrapper_77__ap_done;
  wire PE_wrapper_77__ap_idle;
  wire PE_wrapper_78__ap_start;
  wire PE_wrapper_78__ap_ready;
  wire PE_wrapper_78__ap_done;
  wire PE_wrapper_78__ap_idle;
  wire PE_wrapper_79__ap_start;
  wire PE_wrapper_79__ap_ready;
  wire PE_wrapper_79__ap_done;
  wire PE_wrapper_79__ap_idle;
  wire PE_wrapper_80__ap_start;
  wire PE_wrapper_80__ap_ready;
  wire PE_wrapper_80__ap_done;
  wire PE_wrapper_80__ap_idle;
  wire PE_wrapper_81__ap_start;
  wire PE_wrapper_81__ap_ready;
  wire PE_wrapper_81__ap_done;
  wire PE_wrapper_81__ap_idle;
  wire PE_wrapper_82__ap_start;
  wire PE_wrapper_82__ap_ready;
  wire PE_wrapper_82__ap_done;
  wire PE_wrapper_82__ap_idle;
  wire PE_wrapper_83__ap_start;
  wire PE_wrapper_83__ap_ready;
  wire PE_wrapper_83__ap_done;
  wire PE_wrapper_83__ap_idle;
  wire PE_wrapper_84__ap_start;
  wire PE_wrapper_84__ap_ready;
  wire PE_wrapper_84__ap_done;
  wire PE_wrapper_84__ap_idle;
  wire PE_wrapper_85__ap_start;
  wire PE_wrapper_85__ap_ready;
  wire PE_wrapper_85__ap_done;
  wire PE_wrapper_85__ap_idle;
  wire PE_wrapper_86__ap_start;
  wire PE_wrapper_86__ap_ready;
  wire PE_wrapper_86__ap_done;
  wire PE_wrapper_86__ap_idle;
  wire PE_wrapper_87__ap_start;
  wire PE_wrapper_87__ap_ready;
  wire PE_wrapper_87__ap_done;
  wire PE_wrapper_87__ap_idle;
  wire PE_wrapper_88__ap_start;
  wire PE_wrapper_88__ap_ready;
  wire PE_wrapper_88__ap_done;
  wire PE_wrapper_88__ap_idle;
  wire PE_wrapper_89__ap_start;
  wire PE_wrapper_89__ap_ready;
  wire PE_wrapper_89__ap_done;
  wire PE_wrapper_89__ap_idle;
  wire PE_wrapper_90__ap_start;
  wire PE_wrapper_90__ap_ready;
  wire PE_wrapper_90__ap_done;
  wire PE_wrapper_90__ap_idle;
  wire PE_wrapper_91__ap_start;
  wire PE_wrapper_91__ap_ready;
  wire PE_wrapper_91__ap_done;
  wire PE_wrapper_91__ap_idle;
  wire PE_wrapper_92__ap_start;
  wire PE_wrapper_92__ap_ready;
  wire PE_wrapper_92__ap_done;
  wire PE_wrapper_92__ap_idle;
  wire PE_wrapper_93__ap_start;
  wire PE_wrapper_93__ap_ready;
  wire PE_wrapper_93__ap_done;
  wire PE_wrapper_93__ap_idle;
  wire PE_wrapper_94__ap_start;
  wire PE_wrapper_94__ap_ready;
  wire PE_wrapper_94__ap_done;
  wire PE_wrapper_94__ap_idle;
  wire PE_wrapper_95__ap_start;
  wire PE_wrapper_95__ap_ready;
  wire PE_wrapper_95__ap_done;
  wire PE_wrapper_95__ap_idle;
  wire PE_wrapper_96__ap_start;
  wire PE_wrapper_96__ap_ready;
  wire PE_wrapper_96__ap_done;
  wire PE_wrapper_96__ap_idle;
  wire PE_wrapper_97__ap_start;
  wire PE_wrapper_97__ap_ready;
  wire PE_wrapper_97__ap_done;
  wire PE_wrapper_97__ap_idle;
  wire PE_wrapper_98__ap_start;
  wire PE_wrapper_98__ap_ready;
  wire PE_wrapper_98__ap_done;
  wire PE_wrapper_98__ap_idle;
  wire PE_wrapper_99__ap_start;
  wire PE_wrapper_99__ap_ready;
  wire PE_wrapper_99__ap_done;
  wire PE_wrapper_99__ap_idle;
  wire PE_wrapper_100__ap_start;
  wire PE_wrapper_100__ap_ready;
  wire PE_wrapper_100__ap_done;
  wire PE_wrapper_100__ap_idle;
  wire PE_wrapper_101__ap_start;
  wire PE_wrapper_101__ap_ready;
  wire PE_wrapper_101__ap_done;
  wire PE_wrapper_101__ap_idle;
  wire PE_wrapper_102__ap_start;
  wire PE_wrapper_102__ap_ready;
  wire PE_wrapper_102__ap_done;
  wire PE_wrapper_102__ap_idle;
  wire PE_wrapper_103__ap_start;
  wire PE_wrapper_103__ap_ready;
  wire PE_wrapper_103__ap_done;
  wire PE_wrapper_103__ap_idle;
  wire PE_wrapper_104__ap_start;
  wire PE_wrapper_104__ap_ready;
  wire PE_wrapper_104__ap_done;
  wire PE_wrapper_104__ap_idle;
  wire PE_wrapper_105__ap_start;
  wire PE_wrapper_105__ap_ready;
  wire PE_wrapper_105__ap_done;
  wire PE_wrapper_105__ap_idle;
  wire PE_wrapper_106__ap_start;
  wire PE_wrapper_106__ap_ready;
  wire PE_wrapper_106__ap_done;
  wire PE_wrapper_106__ap_idle;
  wire PE_wrapper_107__ap_start;
  wire PE_wrapper_107__ap_ready;
  wire PE_wrapper_107__ap_done;
  wire PE_wrapper_107__ap_idle;
  wire PE_wrapper_108__ap_start;
  wire PE_wrapper_108__ap_ready;
  wire PE_wrapper_108__ap_done;
  wire PE_wrapper_108__ap_idle;
  wire PE_wrapper_109__ap_start;
  wire PE_wrapper_109__ap_ready;
  wire PE_wrapper_109__ap_done;
  wire PE_wrapper_109__ap_idle;
  wire PE_wrapper_110__ap_start;
  wire PE_wrapper_110__ap_ready;
  wire PE_wrapper_110__ap_done;
  wire PE_wrapper_110__ap_idle;
  wire PE_wrapper_111__ap_start;
  wire PE_wrapper_111__ap_ready;
  wire PE_wrapper_111__ap_done;
  wire PE_wrapper_111__ap_idle;
  wire PE_wrapper_112__ap_start;
  wire PE_wrapper_112__ap_ready;
  wire PE_wrapper_112__ap_done;
  wire PE_wrapper_112__ap_idle;
  wire PE_wrapper_113__ap_start;
  wire PE_wrapper_113__ap_ready;
  wire PE_wrapper_113__ap_done;
  wire PE_wrapper_113__ap_idle;
  wire PE_wrapper_114__ap_start;
  wire PE_wrapper_114__ap_ready;
  wire PE_wrapper_114__ap_done;
  wire PE_wrapper_114__ap_idle;
  wire PE_wrapper_115__ap_start;
  wire PE_wrapper_115__ap_ready;
  wire PE_wrapper_115__ap_done;
  wire PE_wrapper_115__ap_idle;
  wire PE_wrapper_116__ap_start;
  wire PE_wrapper_116__ap_ready;
  wire PE_wrapper_116__ap_done;
  wire PE_wrapper_116__ap_idle;
  wire PE_wrapper_117__ap_start;
  wire PE_wrapper_117__ap_ready;
  wire PE_wrapper_117__ap_done;
  wire PE_wrapper_117__ap_idle;
  wire PE_wrapper_118__ap_start;
  wire PE_wrapper_118__ap_ready;
  wire PE_wrapper_118__ap_done;
  wire PE_wrapper_118__ap_idle;
  wire PE_wrapper_119__ap_start;
  wire PE_wrapper_119__ap_ready;
  wire PE_wrapper_119__ap_done;
  wire PE_wrapper_119__ap_idle;
  wire PE_wrapper_120__ap_start;
  wire PE_wrapper_120__ap_ready;
  wire PE_wrapper_120__ap_done;
  wire PE_wrapper_120__ap_idle;
  wire PE_wrapper_121__ap_start;
  wire PE_wrapper_121__ap_ready;
  wire PE_wrapper_121__ap_done;
  wire PE_wrapper_121__ap_idle;
  wire PE_wrapper_122__ap_start;
  wire PE_wrapper_122__ap_ready;
  wire PE_wrapper_122__ap_done;
  wire PE_wrapper_122__ap_idle;
  wire PE_wrapper_123__ap_start;
  wire PE_wrapper_123__ap_ready;
  wire PE_wrapper_123__ap_done;
  wire PE_wrapper_123__ap_idle;
  wire PE_wrapper_124__ap_start;
  wire PE_wrapper_124__ap_ready;
  wire PE_wrapper_124__ap_done;
  wire PE_wrapper_124__ap_idle;
  wire PE_wrapper_125__ap_start;
  wire PE_wrapper_125__ap_ready;
  wire PE_wrapper_125__ap_done;
  wire PE_wrapper_125__ap_idle;
  wire PE_wrapper_126__ap_start;
  wire PE_wrapper_126__ap_ready;
  wire PE_wrapper_126__ap_done;
  wire PE_wrapper_126__ap_idle;
  wire PE_wrapper_127__ap_start;
  wire PE_wrapper_127__ap_ready;
  wire PE_wrapper_127__ap_done;
  wire PE_wrapper_127__ap_idle;
  wire PE_wrapper_128__ap_start;
  wire PE_wrapper_128__ap_ready;
  wire PE_wrapper_128__ap_done;
  wire PE_wrapper_128__ap_idle;
  wire PE_wrapper_129__ap_start;
  wire PE_wrapper_129__ap_ready;
  wire PE_wrapper_129__ap_done;
  wire PE_wrapper_129__ap_idle;
  wire PE_wrapper_130__ap_start;
  wire PE_wrapper_130__ap_ready;
  wire PE_wrapper_130__ap_done;
  wire PE_wrapper_130__ap_idle;
  wire PE_wrapper_131__ap_start;
  wire PE_wrapper_131__ap_ready;
  wire PE_wrapper_131__ap_done;
  wire PE_wrapper_131__ap_idle;
  wire PE_wrapper_132__ap_start;
  wire PE_wrapper_132__ap_ready;
  wire PE_wrapper_132__ap_done;
  wire PE_wrapper_132__ap_idle;
  wire PE_wrapper_133__ap_start;
  wire PE_wrapper_133__ap_ready;
  wire PE_wrapper_133__ap_done;
  wire PE_wrapper_133__ap_idle;
  wire PE_wrapper_134__ap_start;
  wire PE_wrapper_134__ap_ready;
  wire PE_wrapper_134__ap_done;
  wire PE_wrapper_134__ap_idle;
  wire PE_wrapper_135__ap_start;
  wire PE_wrapper_135__ap_ready;
  wire PE_wrapper_135__ap_done;
  wire PE_wrapper_135__ap_idle;
  wire PE_wrapper_136__ap_start;
  wire PE_wrapper_136__ap_ready;
  wire PE_wrapper_136__ap_done;
  wire PE_wrapper_136__ap_idle;
  wire PE_wrapper_137__ap_start;
  wire PE_wrapper_137__ap_ready;
  wire PE_wrapper_137__ap_done;
  wire PE_wrapper_137__ap_idle;
  wire PE_wrapper_138__ap_start;
  wire PE_wrapper_138__ap_ready;
  wire PE_wrapper_138__ap_done;
  wire PE_wrapper_138__ap_idle;
  wire PE_wrapper_139__ap_start;
  wire PE_wrapper_139__ap_ready;
  wire PE_wrapper_139__ap_done;
  wire PE_wrapper_139__ap_idle;
  wire PE_wrapper_140__ap_start;
  wire PE_wrapper_140__ap_ready;
  wire PE_wrapper_140__ap_done;
  wire PE_wrapper_140__ap_idle;
  wire PE_wrapper_141__ap_start;
  wire PE_wrapper_141__ap_ready;
  wire PE_wrapper_141__ap_done;
  wire PE_wrapper_141__ap_idle;
  wire PE_wrapper_142__ap_start;
  wire PE_wrapper_142__ap_ready;
  wire PE_wrapper_142__ap_done;
  wire PE_wrapper_142__ap_idle;
  wire PE_wrapper_143__ap_start;
  wire PE_wrapper_143__ap_ready;
  wire PE_wrapper_143__ap_done;
  wire PE_wrapper_143__ap_idle;
  wire PE_wrapper_144__ap_start;
  wire PE_wrapper_144__ap_ready;
  wire PE_wrapper_144__ap_done;
  wire PE_wrapper_144__ap_idle;
  wire PE_wrapper_145__ap_start;
  wire PE_wrapper_145__ap_ready;
  wire PE_wrapper_145__ap_done;
  wire PE_wrapper_145__ap_idle;
  wire PE_wrapper_146__ap_start;
  wire PE_wrapper_146__ap_ready;
  wire PE_wrapper_146__ap_done;
  wire PE_wrapper_146__ap_idle;
  wire PE_wrapper_147__ap_start;
  wire PE_wrapper_147__ap_ready;
  wire PE_wrapper_147__ap_done;
  wire PE_wrapper_147__ap_idle;
  wire PE_wrapper_148__ap_start;
  wire PE_wrapper_148__ap_ready;
  wire PE_wrapper_148__ap_done;
  wire PE_wrapper_148__ap_idle;
  wire PE_wrapper_149__ap_start;
  wire PE_wrapper_149__ap_ready;
  wire PE_wrapper_149__ap_done;
  wire PE_wrapper_149__ap_idle;
  wire PE_wrapper_150__ap_start;
  wire PE_wrapper_150__ap_ready;
  wire PE_wrapper_150__ap_done;
  wire PE_wrapper_150__ap_idle;
  wire PE_wrapper_151__ap_start;
  wire PE_wrapper_151__ap_ready;
  wire PE_wrapper_151__ap_done;
  wire PE_wrapper_151__ap_idle;
  wire PE_wrapper_152__ap_start;
  wire PE_wrapper_152__ap_ready;
  wire PE_wrapper_152__ap_done;
  wire PE_wrapper_152__ap_idle;
  wire PE_wrapper_153__ap_start;
  wire PE_wrapper_153__ap_ready;
  wire PE_wrapper_153__ap_done;
  wire PE_wrapper_153__ap_idle;
  wire PE_wrapper_154__ap_start;
  wire PE_wrapper_154__ap_ready;
  wire PE_wrapper_154__ap_done;
  wire PE_wrapper_154__ap_idle;
  wire PE_wrapper_155__ap_start;
  wire PE_wrapper_155__ap_ready;
  wire PE_wrapper_155__ap_done;
  wire PE_wrapper_155__ap_idle;
  wire PE_wrapper_156__ap_start;
  wire PE_wrapper_156__ap_ready;
  wire PE_wrapper_156__ap_done;
  wire PE_wrapper_156__ap_idle;
  wire PE_wrapper_157__ap_start;
  wire PE_wrapper_157__ap_ready;
  wire PE_wrapper_157__ap_done;
  wire PE_wrapper_157__ap_idle;
  wire PE_wrapper_158__ap_start;
  wire PE_wrapper_158__ap_ready;
  wire PE_wrapper_158__ap_done;
  wire PE_wrapper_158__ap_idle;
  wire PE_wrapper_159__ap_start;
  wire PE_wrapper_159__ap_ready;
  wire PE_wrapper_159__ap_done;
  wire PE_wrapper_159__ap_idle;
  wire PE_wrapper_160__ap_start;
  wire PE_wrapper_160__ap_ready;
  wire PE_wrapper_160__ap_done;
  wire PE_wrapper_160__ap_idle;
  wire PE_wrapper_161__ap_start;
  wire PE_wrapper_161__ap_ready;
  wire PE_wrapper_161__ap_done;
  wire PE_wrapper_161__ap_idle;
  wire PE_wrapper_162__ap_start;
  wire PE_wrapper_162__ap_ready;
  wire PE_wrapper_162__ap_done;
  wire PE_wrapper_162__ap_idle;
  wire PE_wrapper_163__ap_start;
  wire PE_wrapper_163__ap_ready;
  wire PE_wrapper_163__ap_done;
  wire PE_wrapper_163__ap_idle;
  wire PE_wrapper_164__ap_start;
  wire PE_wrapper_164__ap_ready;
  wire PE_wrapper_164__ap_done;
  wire PE_wrapper_164__ap_idle;
  wire PE_wrapper_165__ap_start;
  wire PE_wrapper_165__ap_ready;
  wire PE_wrapper_165__ap_done;
  wire PE_wrapper_165__ap_idle;
  wire PE_wrapper_166__ap_start;
  wire PE_wrapper_166__ap_ready;
  wire PE_wrapper_166__ap_done;
  wire PE_wrapper_166__ap_idle;
  wire PE_wrapper_167__ap_start;
  wire PE_wrapper_167__ap_ready;
  wire PE_wrapper_167__ap_done;
  wire PE_wrapper_167__ap_idle;
  wire PE_wrapper_168__ap_start;
  wire PE_wrapper_168__ap_ready;
  wire PE_wrapper_168__ap_done;
  wire PE_wrapper_168__ap_idle;
  wire PE_wrapper_169__ap_start;
  wire PE_wrapper_169__ap_ready;
  wire PE_wrapper_169__ap_done;
  wire PE_wrapper_169__ap_idle;
  wire PE_wrapper_170__ap_start;
  wire PE_wrapper_170__ap_ready;
  wire PE_wrapper_170__ap_done;
  wire PE_wrapper_170__ap_idle;
  wire PE_wrapper_171__ap_start;
  wire PE_wrapper_171__ap_ready;
  wire PE_wrapper_171__ap_done;
  wire PE_wrapper_171__ap_idle;
  wire PE_wrapper_172__ap_start;
  wire PE_wrapper_172__ap_ready;
  wire PE_wrapper_172__ap_done;
  wire PE_wrapper_172__ap_idle;
  wire PE_wrapper_173__ap_start;
  wire PE_wrapper_173__ap_ready;
  wire PE_wrapper_173__ap_done;
  wire PE_wrapper_173__ap_idle;
  wire PE_wrapper_174__ap_start;
  wire PE_wrapper_174__ap_ready;
  wire PE_wrapper_174__ap_done;
  wire PE_wrapper_174__ap_idle;
  wire PE_wrapper_175__ap_start;
  wire PE_wrapper_175__ap_ready;
  wire PE_wrapper_175__ap_done;
  wire PE_wrapper_175__ap_idle;
  wire PE_wrapper_176__ap_start;
  wire PE_wrapper_176__ap_ready;
  wire PE_wrapper_176__ap_done;
  wire PE_wrapper_176__ap_idle;
  wire PE_wrapper_177__ap_start;
  wire PE_wrapper_177__ap_ready;
  wire PE_wrapper_177__ap_done;
  wire PE_wrapper_177__ap_idle;
  wire PE_wrapper_178__ap_start;
  wire PE_wrapper_178__ap_ready;
  wire PE_wrapper_178__ap_done;
  wire PE_wrapper_178__ap_idle;
  wire PE_wrapper_179__ap_start;
  wire PE_wrapper_179__ap_ready;
  wire PE_wrapper_179__ap_done;
  wire PE_wrapper_179__ap_idle;
  wire PE_wrapper_180__ap_start;
  wire PE_wrapper_180__ap_ready;
  wire PE_wrapper_180__ap_done;
  wire PE_wrapper_180__ap_idle;
  wire PE_wrapper_181__ap_start;
  wire PE_wrapper_181__ap_ready;
  wire PE_wrapper_181__ap_done;
  wire PE_wrapper_181__ap_idle;
  wire PE_wrapper_182__ap_start;
  wire PE_wrapper_182__ap_ready;
  wire PE_wrapper_182__ap_done;
  wire PE_wrapper_182__ap_idle;
  wire PE_wrapper_183__ap_start;
  wire PE_wrapper_183__ap_ready;
  wire PE_wrapper_183__ap_done;
  wire PE_wrapper_183__ap_idle;
  wire PE_wrapper_184__ap_start;
  wire PE_wrapper_184__ap_ready;
  wire PE_wrapper_184__ap_done;
  wire PE_wrapper_184__ap_idle;
  wire PE_wrapper_185__ap_start;
  wire PE_wrapper_185__ap_ready;
  wire PE_wrapper_185__ap_done;
  wire PE_wrapper_185__ap_idle;
  wire PE_wrapper_186__ap_start;
  wire PE_wrapper_186__ap_ready;
  wire PE_wrapper_186__ap_done;
  wire PE_wrapper_186__ap_idle;
  wire PE_wrapper_187__ap_start;
  wire PE_wrapper_187__ap_ready;
  wire PE_wrapper_187__ap_done;
  wire PE_wrapper_187__ap_idle;
  wire PE_wrapper_188__ap_start;
  wire PE_wrapper_188__ap_ready;
  wire PE_wrapper_188__ap_done;
  wire PE_wrapper_188__ap_idle;
  wire PE_wrapper_189__ap_start;
  wire PE_wrapper_189__ap_ready;
  wire PE_wrapper_189__ap_done;
  wire PE_wrapper_189__ap_idle;
  wire PE_wrapper_190__ap_start;
  wire PE_wrapper_190__ap_ready;
  wire PE_wrapper_190__ap_done;
  wire PE_wrapper_190__ap_idle;
  wire PE_wrapper_191__ap_start;
  wire PE_wrapper_191__ap_ready;
  wire PE_wrapper_191__ap_done;
  wire PE_wrapper_191__ap_idle;
  wire PE_wrapper_192__ap_start;
  wire PE_wrapper_192__ap_ready;
  wire PE_wrapper_192__ap_done;
  wire PE_wrapper_192__ap_idle;
  wire PE_wrapper_193__ap_start;
  wire PE_wrapper_193__ap_ready;
  wire PE_wrapper_193__ap_done;
  wire PE_wrapper_193__ap_idle;
  wire PE_wrapper_194__ap_start;
  wire PE_wrapper_194__ap_ready;
  wire PE_wrapper_194__ap_done;
  wire PE_wrapper_194__ap_idle;
  wire PE_wrapper_195__ap_start;
  wire PE_wrapper_195__ap_ready;
  wire PE_wrapper_195__ap_done;
  wire PE_wrapper_195__ap_idle;
  wire PE_wrapper_196__ap_start;
  wire PE_wrapper_196__ap_ready;
  wire PE_wrapper_196__ap_done;
  wire PE_wrapper_196__ap_idle;
  wire PE_wrapper_197__ap_start;
  wire PE_wrapper_197__ap_ready;
  wire PE_wrapper_197__ap_done;
  wire PE_wrapper_197__ap_idle;
  wire PE_wrapper_198__ap_start;
  wire PE_wrapper_198__ap_ready;
  wire PE_wrapper_198__ap_done;
  wire PE_wrapper_198__ap_idle;
  wire PE_wrapper_199__ap_start;
  wire PE_wrapper_199__ap_ready;
  wire PE_wrapper_199__ap_done;
  wire PE_wrapper_199__ap_idle;
  wire PE_wrapper_200__ap_start;
  wire PE_wrapper_200__ap_ready;
  wire PE_wrapper_200__ap_done;
  wire PE_wrapper_200__ap_idle;
  wire PE_wrapper_201__ap_start;
  wire PE_wrapper_201__ap_ready;
  wire PE_wrapper_201__ap_done;
  wire PE_wrapper_201__ap_idle;
  wire PE_wrapper_202__ap_start;
  wire PE_wrapper_202__ap_ready;
  wire PE_wrapper_202__ap_done;
  wire PE_wrapper_202__ap_idle;
  wire PE_wrapper_203__ap_start;
  wire PE_wrapper_203__ap_ready;
  wire PE_wrapper_203__ap_done;
  wire PE_wrapper_203__ap_idle;
  wire PE_wrapper_204__ap_start;
  wire PE_wrapper_204__ap_ready;
  wire PE_wrapper_204__ap_done;
  wire PE_wrapper_204__ap_idle;
  wire PE_wrapper_205__ap_start;
  wire PE_wrapper_205__ap_ready;
  wire PE_wrapper_205__ap_done;
  wire PE_wrapper_205__ap_idle;
  wire PE_wrapper_206__ap_start;
  wire PE_wrapper_206__ap_ready;
  wire PE_wrapper_206__ap_done;
  wire PE_wrapper_206__ap_idle;
  wire PE_wrapper_207__ap_start;
  wire PE_wrapper_207__ap_ready;
  wire PE_wrapper_207__ap_done;
  wire PE_wrapper_207__ap_idle;
  wire PE_wrapper_208__ap_start;
  wire PE_wrapper_208__ap_ready;
  wire PE_wrapper_208__ap_done;
  wire PE_wrapper_208__ap_idle;
  wire PE_wrapper_209__ap_start;
  wire PE_wrapper_209__ap_ready;
  wire PE_wrapper_209__ap_done;
  wire PE_wrapper_209__ap_idle;
  wire PE_wrapper_210__ap_start;
  wire PE_wrapper_210__ap_ready;
  wire PE_wrapper_210__ap_done;
  wire PE_wrapper_210__ap_idle;
  wire PE_wrapper_211__ap_start;
  wire PE_wrapper_211__ap_ready;
  wire PE_wrapper_211__ap_done;
  wire PE_wrapper_211__ap_idle;
  wire PE_wrapper_212__ap_start;
  wire PE_wrapper_212__ap_ready;
  wire PE_wrapper_212__ap_done;
  wire PE_wrapper_212__ap_idle;
  wire PE_wrapper_213__ap_start;
  wire PE_wrapper_213__ap_ready;
  wire PE_wrapper_213__ap_done;
  wire PE_wrapper_213__ap_idle;
  wire PE_wrapper_214__ap_start;
  wire PE_wrapper_214__ap_ready;
  wire PE_wrapper_214__ap_done;
  wire PE_wrapper_214__ap_idle;
  wire PE_wrapper_215__ap_start;
  wire PE_wrapper_215__ap_ready;
  wire PE_wrapper_215__ap_done;
  wire PE_wrapper_215__ap_idle;
  wire PE_wrapper_216__ap_start;
  wire PE_wrapper_216__ap_ready;
  wire PE_wrapper_216__ap_done;
  wire PE_wrapper_216__ap_idle;
  wire PE_wrapper_217__ap_start;
  wire PE_wrapper_217__ap_ready;
  wire PE_wrapper_217__ap_done;
  wire PE_wrapper_217__ap_idle;
  wire PE_wrapper_218__ap_start;
  wire PE_wrapper_218__ap_ready;
  wire PE_wrapper_218__ap_done;
  wire PE_wrapper_218__ap_idle;
  wire PE_wrapper_219__ap_start;
  wire PE_wrapper_219__ap_ready;
  wire PE_wrapper_219__ap_done;
  wire PE_wrapper_219__ap_idle;
  wire PE_wrapper_220__ap_start;
  wire PE_wrapper_220__ap_ready;
  wire PE_wrapper_220__ap_done;
  wire PE_wrapper_220__ap_idle;
  wire PE_wrapper_221__ap_start;
  wire PE_wrapper_221__ap_ready;
  wire PE_wrapper_221__ap_done;
  wire PE_wrapper_221__ap_idle;
  wire PE_wrapper_222__ap_start;
  wire PE_wrapper_222__ap_ready;
  wire PE_wrapper_222__ap_done;
  wire PE_wrapper_222__ap_idle;
  wire PE_wrapper_223__ap_start;
  wire PE_wrapper_223__ap_ready;
  wire PE_wrapper_223__ap_done;
  wire PE_wrapper_223__ap_idle;
  wire PE_wrapper_224__ap_start;
  wire PE_wrapper_224__ap_ready;
  wire PE_wrapper_224__ap_done;
  wire PE_wrapper_224__ap_idle;
  wire PE_wrapper_225__ap_start;
  wire PE_wrapper_225__ap_ready;
  wire PE_wrapper_225__ap_done;
  wire PE_wrapper_225__ap_idle;
  wire PE_wrapper_226__ap_start;
  wire PE_wrapper_226__ap_ready;
  wire PE_wrapper_226__ap_done;
  wire PE_wrapper_226__ap_idle;
  wire PE_wrapper_227__ap_start;
  wire PE_wrapper_227__ap_ready;
  wire PE_wrapper_227__ap_done;
  wire PE_wrapper_227__ap_idle;
  wire PE_wrapper_228__ap_start;
  wire PE_wrapper_228__ap_ready;
  wire PE_wrapper_228__ap_done;
  wire PE_wrapper_228__ap_idle;
  wire PE_wrapper_229__ap_start;
  wire PE_wrapper_229__ap_ready;
  wire PE_wrapper_229__ap_done;
  wire PE_wrapper_229__ap_idle;
  wire PE_wrapper_230__ap_start;
  wire PE_wrapper_230__ap_ready;
  wire PE_wrapper_230__ap_done;
  wire PE_wrapper_230__ap_idle;
  wire PE_wrapper_231__ap_start;
  wire PE_wrapper_231__ap_ready;
  wire PE_wrapper_231__ap_done;
  wire PE_wrapper_231__ap_idle;
  wire PE_wrapper_232__ap_start;
  wire PE_wrapper_232__ap_ready;
  wire PE_wrapper_232__ap_done;
  wire PE_wrapper_232__ap_idle;
  wire PE_wrapper_233__ap_start;
  wire PE_wrapper_233__ap_ready;
  wire PE_wrapper_233__ap_done;
  wire PE_wrapper_233__ap_idle;
  wire PE_wrapper_234__ap_start;
  wire PE_wrapper_234__ap_ready;
  wire PE_wrapper_234__ap_done;
  wire PE_wrapper_234__ap_idle;
  wire PE_wrapper_235__ap_start;
  wire PE_wrapper_235__ap_ready;
  wire PE_wrapper_235__ap_done;
  wire PE_wrapper_235__ap_idle;
  wire PE_wrapper_236__ap_start;
  wire PE_wrapper_236__ap_ready;
  wire PE_wrapper_236__ap_done;
  wire PE_wrapper_236__ap_idle;
  wire PE_wrapper_237__ap_start;
  wire PE_wrapper_237__ap_ready;
  wire PE_wrapper_237__ap_done;
  wire PE_wrapper_237__ap_idle;
  wire PE_wrapper_238__ap_start;
  wire PE_wrapper_238__ap_ready;
  wire PE_wrapper_238__ap_done;
  wire PE_wrapper_238__ap_idle;
  wire PE_wrapper_239__ap_start;
  wire PE_wrapper_239__ap_ready;
  wire PE_wrapper_239__ap_done;
  wire PE_wrapper_239__ap_idle;
  wire PE_wrapper_240__ap_start;
  wire PE_wrapper_240__ap_ready;
  wire PE_wrapper_240__ap_done;
  wire PE_wrapper_240__ap_idle;
  wire PE_wrapper_241__ap_start;
  wire PE_wrapper_241__ap_ready;
  wire PE_wrapper_241__ap_done;
  wire PE_wrapper_241__ap_idle;
  wire PE_wrapper_242__ap_start;
  wire PE_wrapper_242__ap_ready;
  wire PE_wrapper_242__ap_done;
  wire PE_wrapper_242__ap_idle;
  wire PE_wrapper_243__ap_start;
  wire PE_wrapper_243__ap_ready;
  wire PE_wrapper_243__ap_done;
  wire PE_wrapper_243__ap_idle;
  wire PE_wrapper_244__ap_start;
  wire PE_wrapper_244__ap_ready;
  wire PE_wrapper_244__ap_done;
  wire PE_wrapper_244__ap_idle;
  wire PE_wrapper_245__ap_start;
  wire PE_wrapper_245__ap_ready;
  wire PE_wrapper_245__ap_done;
  wire PE_wrapper_245__ap_idle;
  wire PE_wrapper_246__ap_start;
  wire PE_wrapper_246__ap_ready;
  wire PE_wrapper_246__ap_done;
  wire PE_wrapper_246__ap_idle;
  wire PE_wrapper_247__ap_start;
  wire PE_wrapper_247__ap_ready;
  wire PE_wrapper_247__ap_done;
  wire PE_wrapper_247__ap_idle;
  wire PE_wrapper_248__ap_start;
  wire PE_wrapper_248__ap_ready;
  wire PE_wrapper_248__ap_done;
  wire PE_wrapper_248__ap_idle;
  wire PE_wrapper_249__ap_start;
  wire PE_wrapper_249__ap_ready;
  wire PE_wrapper_249__ap_done;
  wire PE_wrapper_249__ap_idle;
  wire PE_wrapper_250__ap_start;
  wire PE_wrapper_250__ap_ready;
  wire PE_wrapper_250__ap_done;
  wire PE_wrapper_250__ap_idle;
  wire PE_wrapper_251__ap_start;
  wire PE_wrapper_251__ap_ready;
  wire PE_wrapper_251__ap_done;
  wire PE_wrapper_251__ap_idle;
  wire PE_wrapper_252__ap_start;
  wire PE_wrapper_252__ap_ready;
  wire PE_wrapper_252__ap_done;
  wire PE_wrapper_252__ap_idle;
  wire PE_wrapper_253__ap_start;
  wire PE_wrapper_253__ap_ready;
  wire PE_wrapper_253__ap_done;
  wire PE_wrapper_253__ap_idle;
  wire PE_wrapper_254__ap_start;
  wire PE_wrapper_254__ap_ready;
  wire PE_wrapper_254__ap_done;
  wire PE_wrapper_254__ap_idle;
  wire PE_wrapper_255__ap_start;
  wire PE_wrapper_255__ap_ready;
  wire PE_wrapper_255__ap_done;
  wire PE_wrapper_255__ap_idle;
  wire PE_wrapper_256__ap_start;
  wire PE_wrapper_256__ap_ready;
  wire PE_wrapper_256__ap_done;
  wire PE_wrapper_256__ap_idle;
  wire PE_wrapper_257__ap_start;
  wire PE_wrapper_257__ap_ready;
  wire PE_wrapper_257__ap_done;
  wire PE_wrapper_257__ap_idle;
  wire PE_wrapper_258__ap_start;
  wire PE_wrapper_258__ap_ready;
  wire PE_wrapper_258__ap_done;
  wire PE_wrapper_258__ap_idle;
  wire PE_wrapper_259__ap_start;
  wire PE_wrapper_259__ap_ready;
  wire PE_wrapper_259__ap_done;
  wire PE_wrapper_259__ap_idle;
  wire PE_wrapper_260__ap_start;
  wire PE_wrapper_260__ap_ready;
  wire PE_wrapper_260__ap_done;
  wire PE_wrapper_260__ap_idle;
  wire PE_wrapper_261__ap_start;
  wire PE_wrapper_261__ap_ready;
  wire PE_wrapper_261__ap_done;
  wire PE_wrapper_261__ap_idle;
  wire PE_wrapper_262__ap_start;
  wire PE_wrapper_262__ap_ready;
  wire PE_wrapper_262__ap_done;
  wire PE_wrapper_262__ap_idle;
  wire PE_wrapper_263__ap_start;
  wire PE_wrapper_263__ap_ready;
  wire PE_wrapper_263__ap_done;
  wire PE_wrapper_263__ap_idle;
  wire PE_wrapper_264__ap_start;
  wire PE_wrapper_264__ap_ready;
  wire PE_wrapper_264__ap_done;
  wire PE_wrapper_264__ap_idle;
  wire PE_wrapper_265__ap_start;
  wire PE_wrapper_265__ap_ready;
  wire PE_wrapper_265__ap_done;
  wire PE_wrapper_265__ap_idle;
  wire PE_wrapper_266__ap_start;
  wire PE_wrapper_266__ap_ready;
  wire PE_wrapper_266__ap_done;
  wire PE_wrapper_266__ap_idle;
  wire PE_wrapper_267__ap_start;
  wire PE_wrapper_267__ap_ready;
  wire PE_wrapper_267__ap_done;
  wire PE_wrapper_267__ap_idle;
  wire PE_wrapper_268__ap_start;
  wire PE_wrapper_268__ap_ready;
  wire PE_wrapper_268__ap_done;
  wire PE_wrapper_268__ap_idle;
  wire PE_wrapper_269__ap_start;
  wire PE_wrapper_269__ap_ready;
  wire PE_wrapper_269__ap_done;
  wire PE_wrapper_269__ap_idle;
  wire PE_wrapper_270__ap_start;
  wire PE_wrapper_270__ap_ready;
  wire PE_wrapper_270__ap_done;
  wire PE_wrapper_270__ap_idle;
  wire PE_wrapper_271__ap_start;
  wire PE_wrapper_271__ap_ready;
  wire PE_wrapper_271__ap_done;
  wire PE_wrapper_271__ap_idle;
  wire PE_wrapper_272__ap_start;
  wire PE_wrapper_272__ap_ready;
  wire PE_wrapper_272__ap_done;
  wire PE_wrapper_272__ap_idle;
  wire PE_wrapper_273__ap_start;
  wire PE_wrapper_273__ap_ready;
  wire PE_wrapper_273__ap_done;
  wire PE_wrapper_273__ap_idle;
  wire PE_wrapper_274__ap_start;
  wire PE_wrapper_274__ap_ready;
  wire PE_wrapper_274__ap_done;
  wire PE_wrapper_274__ap_idle;
  wire PE_wrapper_275__ap_start;
  wire PE_wrapper_275__ap_ready;
  wire PE_wrapper_275__ap_done;
  wire PE_wrapper_275__ap_idle;
  wire PE_wrapper_276__ap_start;
  wire PE_wrapper_276__ap_ready;
  wire PE_wrapper_276__ap_done;
  wire PE_wrapper_276__ap_idle;
  wire PE_wrapper_277__ap_start;
  wire PE_wrapper_277__ap_ready;
  wire PE_wrapper_277__ap_done;
  wire PE_wrapper_277__ap_idle;
  wire PE_wrapper_278__ap_start;
  wire PE_wrapper_278__ap_ready;
  wire PE_wrapper_278__ap_done;
  wire PE_wrapper_278__ap_idle;
  wire PE_wrapper_279__ap_start;
  wire PE_wrapper_279__ap_ready;
  wire PE_wrapper_279__ap_done;
  wire PE_wrapper_279__ap_idle;
  wire PE_wrapper_280__ap_start;
  wire PE_wrapper_280__ap_ready;
  wire PE_wrapper_280__ap_done;
  wire PE_wrapper_280__ap_idle;
  wire PE_wrapper_281__ap_start;
  wire PE_wrapper_281__ap_ready;
  wire PE_wrapper_281__ap_done;
  wire PE_wrapper_281__ap_idle;
  wire PE_wrapper_282__ap_start;
  wire PE_wrapper_282__ap_ready;
  wire PE_wrapper_282__ap_done;
  wire PE_wrapper_282__ap_idle;
  wire PE_wrapper_283__ap_start;
  wire PE_wrapper_283__ap_ready;
  wire PE_wrapper_283__ap_done;
  wire PE_wrapper_283__ap_idle;
  wire PE_wrapper_284__ap_start;
  wire PE_wrapper_284__ap_ready;
  wire PE_wrapper_284__ap_done;
  wire PE_wrapper_284__ap_idle;
  wire PE_wrapper_285__ap_start;
  wire PE_wrapper_285__ap_ready;
  wire PE_wrapper_285__ap_done;
  wire PE_wrapper_285__ap_idle;
  wire PE_wrapper_286__ap_start;
  wire PE_wrapper_286__ap_ready;
  wire PE_wrapper_286__ap_done;
  wire PE_wrapper_286__ap_idle;
  wire PE_wrapper_287__ap_start;
  wire PE_wrapper_287__ap_ready;
  wire PE_wrapper_287__ap_done;
  wire PE_wrapper_287__ap_idle;
  wire PE_wrapper_288__ap_start;
  wire PE_wrapper_288__ap_ready;
  wire PE_wrapper_288__ap_done;
  wire PE_wrapper_288__ap_idle;
  wire PE_wrapper_289__ap_start;
  wire PE_wrapper_289__ap_ready;
  wire PE_wrapper_289__ap_done;
  wire PE_wrapper_289__ap_idle;
  wire PE_wrapper_290__ap_start;
  wire PE_wrapper_290__ap_ready;
  wire PE_wrapper_290__ap_done;
  wire PE_wrapper_290__ap_idle;
  wire PE_wrapper_291__ap_start;
  wire PE_wrapper_291__ap_ready;
  wire PE_wrapper_291__ap_done;
  wire PE_wrapper_291__ap_idle;
  wire PE_wrapper_292__ap_start;
  wire PE_wrapper_292__ap_ready;
  wire PE_wrapper_292__ap_done;
  wire PE_wrapper_292__ap_idle;
  wire PE_wrapper_293__ap_start;
  wire PE_wrapper_293__ap_ready;
  wire PE_wrapper_293__ap_done;
  wire PE_wrapper_293__ap_idle;
  wire PE_wrapper_294__ap_start;
  wire PE_wrapper_294__ap_ready;
  wire PE_wrapper_294__ap_done;
  wire PE_wrapper_294__ap_idle;
  wire PE_wrapper_295__ap_start;
  wire PE_wrapper_295__ap_ready;
  wire PE_wrapper_295__ap_done;
  wire PE_wrapper_295__ap_idle;
  wire PE_wrapper_296__ap_start;
  wire PE_wrapper_296__ap_ready;
  wire PE_wrapper_296__ap_done;
  wire PE_wrapper_296__ap_idle;
  wire PE_wrapper_297__ap_start;
  wire PE_wrapper_297__ap_ready;
  wire PE_wrapper_297__ap_done;
  wire PE_wrapper_297__ap_idle;
  wire PE_wrapper_298__ap_start;
  wire PE_wrapper_298__ap_ready;
  wire PE_wrapper_298__ap_done;
  wire PE_wrapper_298__ap_idle;
  wire PE_wrapper_299__ap_start;
  wire PE_wrapper_299__ap_ready;
  wire PE_wrapper_299__ap_done;
  wire PE_wrapper_299__ap_idle;
  wire PE_wrapper_300__ap_start;
  wire PE_wrapper_300__ap_ready;
  wire PE_wrapper_300__ap_done;
  wire PE_wrapper_300__ap_idle;
  wire PE_wrapper_301__ap_start;
  wire PE_wrapper_301__ap_ready;
  wire PE_wrapper_301__ap_done;
  wire PE_wrapper_301__ap_idle;
  wire PE_wrapper_302__ap_start;
  wire PE_wrapper_302__ap_ready;
  wire PE_wrapper_302__ap_done;
  wire PE_wrapper_302__ap_idle;
  wire PE_wrapper_303__ap_start;
  wire PE_wrapper_303__ap_ready;
  wire PE_wrapper_303__ap_done;
  wire PE_wrapper_303__ap_idle;
  wire PE_wrapper_304__ap_start;
  wire PE_wrapper_304__ap_ready;
  wire PE_wrapper_304__ap_done;
  wire PE_wrapper_304__ap_idle;
  wire PE_wrapper_305__ap_start;
  wire PE_wrapper_305__ap_ready;
  wire PE_wrapper_305__ap_done;
  wire PE_wrapper_305__ap_idle;
  wire ap_rst_n_inv;
  wire ap_done;
  wire ap_idle;
  wire ap_ready;

  kernel0_control_s_axi
  #(
    .C_S_AXI_ADDR_WIDTH(C_S_AXI_CONTROL_ADDR_WIDTH),
    .C_S_AXI_DATA_WIDTH(C_S_AXI_CONTROL_DATA_WIDTH)
  )
  control_s_axi_U
  (
    .AWVALID(s_axi_control_AWVALID),
    .AWREADY(s_axi_control_AWREADY),
    .AWADDR(s_axi_control_AWADDR),
    .WVALID(s_axi_control_WVALID),
    .WREADY(s_axi_control_WREADY),
    .WDATA(s_axi_control_WDATA),
    .WSTRB(s_axi_control_WSTRB),
    .ARVALID(s_axi_control_ARVALID),
    .ARREADY(s_axi_control_ARREADY),
    .ARADDR(s_axi_control_ARADDR),
    .RVALID(s_axi_control_RVALID),
    .RREADY(s_axi_control_RREADY),
    .RDATA(s_axi_control_RDATA),
    .RRESP(s_axi_control_RRESP),
    .BVALID(s_axi_control_BVALID),
    .BREADY(s_axi_control_BREADY),
    .BRESP(s_axi_control_BRESP),
    .ACLK(ap_clk),
    .ARESET(ap_rst_n_inv),
    .ACLK_EN(1'b1),
    .A(A),
    .B(B),
    .C(C),
    .ap_start(ap_start),
    .interrupt(interrupt),
    .ap_ready(ap_ready),
    .ap_done(ap_done),
    .ap_idle(ap_idle)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_A_IO_L2_in_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_A_IO_L2_in_0__dout),
    .if_empty_n(fifo_A_A_IO_L2_in_0__empty_n),
    .if_read(fifo_A_A_IO_L2_in_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_A_IO_L2_in_0__din),
    .if_full_n(fifo_A_A_IO_L2_in_0__full_n),
    .if_write(fifo_A_A_IO_L2_in_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_A_IO_L2_in_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_A_IO_L2_in_1__dout),
    .if_empty_n(fifo_A_A_IO_L2_in_1__empty_n),
    .if_read(fifo_A_A_IO_L2_in_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_A_IO_L2_in_1__din),
    .if_full_n(fifo_A_A_IO_L2_in_1__full_n),
    .if_write(fifo_A_A_IO_L2_in_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_A_IO_L2_in_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_A_IO_L2_in_10__dout),
    .if_empty_n(fifo_A_A_IO_L2_in_10__empty_n),
    .if_read(fifo_A_A_IO_L2_in_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_A_IO_L2_in_10__din),
    .if_full_n(fifo_A_A_IO_L2_in_10__full_n),
    .if_write(fifo_A_A_IO_L2_in_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_A_IO_L2_in_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_A_IO_L2_in_11__dout),
    .if_empty_n(fifo_A_A_IO_L2_in_11__empty_n),
    .if_read(fifo_A_A_IO_L2_in_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_A_IO_L2_in_11__din),
    .if_full_n(fifo_A_A_IO_L2_in_11__full_n),
    .if_write(fifo_A_A_IO_L2_in_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_A_IO_L2_in_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_A_IO_L2_in_12__dout),
    .if_empty_n(fifo_A_A_IO_L2_in_12__empty_n),
    .if_read(fifo_A_A_IO_L2_in_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_A_IO_L2_in_12__din),
    .if_full_n(fifo_A_A_IO_L2_in_12__full_n),
    .if_write(fifo_A_A_IO_L2_in_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_A_IO_L2_in_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_A_IO_L2_in_13__dout),
    .if_empty_n(fifo_A_A_IO_L2_in_13__empty_n),
    .if_read(fifo_A_A_IO_L2_in_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_A_IO_L2_in_13__din),
    .if_full_n(fifo_A_A_IO_L2_in_13__full_n),
    .if_write(fifo_A_A_IO_L2_in_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_A_IO_L2_in_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_A_IO_L2_in_14__dout),
    .if_empty_n(fifo_A_A_IO_L2_in_14__empty_n),
    .if_read(fifo_A_A_IO_L2_in_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_A_IO_L2_in_14__din),
    .if_full_n(fifo_A_A_IO_L2_in_14__full_n),
    .if_write(fifo_A_A_IO_L2_in_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_A_IO_L2_in_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_A_IO_L2_in_15__dout),
    .if_empty_n(fifo_A_A_IO_L2_in_15__empty_n),
    .if_read(fifo_A_A_IO_L2_in_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_A_IO_L2_in_15__din),
    .if_full_n(fifo_A_A_IO_L2_in_15__full_n),
    .if_write(fifo_A_A_IO_L2_in_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_A_IO_L2_in_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_A_IO_L2_in_16__dout),
    .if_empty_n(fifo_A_A_IO_L2_in_16__empty_n),
    .if_read(fifo_A_A_IO_L2_in_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_A_IO_L2_in_16__din),
    .if_full_n(fifo_A_A_IO_L2_in_16__full_n),
    .if_write(fifo_A_A_IO_L2_in_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_A_IO_L2_in_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_A_IO_L2_in_17__dout),
    .if_empty_n(fifo_A_A_IO_L2_in_17__empty_n),
    .if_read(fifo_A_A_IO_L2_in_17__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_A_IO_L2_in_17__din),
    .if_full_n(fifo_A_A_IO_L2_in_17__full_n),
    .if_write(fifo_A_A_IO_L2_in_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_A_IO_L2_in_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_A_IO_L2_in_2__dout),
    .if_empty_n(fifo_A_A_IO_L2_in_2__empty_n),
    .if_read(fifo_A_A_IO_L2_in_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_A_IO_L2_in_2__din),
    .if_full_n(fifo_A_A_IO_L2_in_2__full_n),
    .if_write(fifo_A_A_IO_L2_in_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_A_IO_L2_in_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_A_IO_L2_in_3__dout),
    .if_empty_n(fifo_A_A_IO_L2_in_3__empty_n),
    .if_read(fifo_A_A_IO_L2_in_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_A_IO_L2_in_3__din),
    .if_full_n(fifo_A_A_IO_L2_in_3__full_n),
    .if_write(fifo_A_A_IO_L2_in_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_A_IO_L2_in_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_A_IO_L2_in_4__dout),
    .if_empty_n(fifo_A_A_IO_L2_in_4__empty_n),
    .if_read(fifo_A_A_IO_L2_in_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_A_IO_L2_in_4__din),
    .if_full_n(fifo_A_A_IO_L2_in_4__full_n),
    .if_write(fifo_A_A_IO_L2_in_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_A_IO_L2_in_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_A_IO_L2_in_5__dout),
    .if_empty_n(fifo_A_A_IO_L2_in_5__empty_n),
    .if_read(fifo_A_A_IO_L2_in_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_A_IO_L2_in_5__din),
    .if_full_n(fifo_A_A_IO_L2_in_5__full_n),
    .if_write(fifo_A_A_IO_L2_in_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_A_IO_L2_in_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_A_IO_L2_in_6__dout),
    .if_empty_n(fifo_A_A_IO_L2_in_6__empty_n),
    .if_read(fifo_A_A_IO_L2_in_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_A_IO_L2_in_6__din),
    .if_full_n(fifo_A_A_IO_L2_in_6__full_n),
    .if_write(fifo_A_A_IO_L2_in_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_A_IO_L2_in_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_A_IO_L2_in_7__dout),
    .if_empty_n(fifo_A_A_IO_L2_in_7__empty_n),
    .if_read(fifo_A_A_IO_L2_in_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_A_IO_L2_in_7__din),
    .if_full_n(fifo_A_A_IO_L2_in_7__full_n),
    .if_write(fifo_A_A_IO_L2_in_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_A_IO_L2_in_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_A_IO_L2_in_8__dout),
    .if_empty_n(fifo_A_A_IO_L2_in_8__empty_n),
    .if_read(fifo_A_A_IO_L2_in_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_A_IO_L2_in_8__din),
    .if_full_n(fifo_A_A_IO_L2_in_8__full_n),
    .if_write(fifo_A_A_IO_L2_in_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_A_IO_L2_in_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_A_IO_L2_in_9__dout),
    .if_empty_n(fifo_A_A_IO_L2_in_9__empty_n),
    .if_read(fifo_A_A_IO_L2_in_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_A_IO_L2_in_9__din),
    .if_full_n(fifo_A_A_IO_L2_in_9__full_n),
    .if_write(fifo_A_A_IO_L2_in_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_A_IO_L3_in_serialize
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_A_IO_L3_in_serialize__dout),
    .if_empty_n(fifo_A_A_IO_L3_in_serialize__empty_n),
    .if_read(fifo_A_A_IO_L3_in_serialize__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_A_IO_L3_in_serialize__din),
    .if_full_n(fifo_A_A_IO_L3_in_serialize__full_n),
    .if_write(fifo_A_A_IO_L3_in_serialize__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_0_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_0_0__dout),
    .if_empty_n(fifo_A_PE_0_0__empty_n),
    .if_read(fifo_A_PE_0_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_0_0__din),
    .if_full_n(fifo_A_PE_0_0__full_n),
    .if_write(fifo_A_PE_0_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_0_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_0_1__dout),
    .if_empty_n(fifo_A_PE_0_1__empty_n),
    .if_read(fifo_A_PE_0_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_0_1__din),
    .if_full_n(fifo_A_PE_0_1__full_n),
    .if_write(fifo_A_PE_0_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_0_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_0_10__dout),
    .if_empty_n(fifo_A_PE_0_10__empty_n),
    .if_read(fifo_A_PE_0_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_0_10__din),
    .if_full_n(fifo_A_PE_0_10__full_n),
    .if_write(fifo_A_PE_0_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_0_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_0_11__dout),
    .if_empty_n(fifo_A_PE_0_11__empty_n),
    .if_read(fifo_A_PE_0_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_0_11__din),
    .if_full_n(fifo_A_PE_0_11__full_n),
    .if_write(fifo_A_PE_0_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_0_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_0_12__dout),
    .if_empty_n(fifo_A_PE_0_12__empty_n),
    .if_read(fifo_A_PE_0_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_0_12__din),
    .if_full_n(fifo_A_PE_0_12__full_n),
    .if_write(fifo_A_PE_0_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_0_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_0_13__dout),
    .if_empty_n(fifo_A_PE_0_13__empty_n),
    .if_read(fifo_A_PE_0_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_0_13__din),
    .if_full_n(fifo_A_PE_0_13__full_n),
    .if_write(fifo_A_PE_0_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_0_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_0_14__dout),
    .if_empty_n(fifo_A_PE_0_14__empty_n),
    .if_read(fifo_A_PE_0_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_0_14__din),
    .if_full_n(fifo_A_PE_0_14__full_n),
    .if_write(fifo_A_PE_0_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_0_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_0_15__dout),
    .if_empty_n(fifo_A_PE_0_15__empty_n),
    .if_read(fifo_A_PE_0_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_0_15__din),
    .if_full_n(fifo_A_PE_0_15__full_n),
    .if_write(fifo_A_PE_0_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_0_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_0_16__dout),
    .if_empty_n(fifo_A_PE_0_16__empty_n),
    .if_read(fifo_A_PE_0_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_0_16__din),
    .if_full_n(fifo_A_PE_0_16__full_n),
    .if_write(fifo_A_PE_0_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_0_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_0_17__dout),
    .if_empty_n(fifo_A_PE_0_17__empty_n),
    .if_read(fifo_A_PE_0_17__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_0_17__din),
    .if_full_n(fifo_A_PE_0_17__full_n),
    .if_write(fifo_A_PE_0_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_0_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_0_2__dout),
    .if_empty_n(fifo_A_PE_0_2__empty_n),
    .if_read(fifo_A_PE_0_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_0_2__din),
    .if_full_n(fifo_A_PE_0_2__full_n),
    .if_write(fifo_A_PE_0_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_0_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_0_3__dout),
    .if_empty_n(fifo_A_PE_0_3__empty_n),
    .if_read(fifo_A_PE_0_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_0_3__din),
    .if_full_n(fifo_A_PE_0_3__full_n),
    .if_write(fifo_A_PE_0_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_0_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_0_4__dout),
    .if_empty_n(fifo_A_PE_0_4__empty_n),
    .if_read(fifo_A_PE_0_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_0_4__din),
    .if_full_n(fifo_A_PE_0_4__full_n),
    .if_write(fifo_A_PE_0_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_0_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_0_5__dout),
    .if_empty_n(fifo_A_PE_0_5__empty_n),
    .if_read(fifo_A_PE_0_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_0_5__din),
    .if_full_n(fifo_A_PE_0_5__full_n),
    .if_write(fifo_A_PE_0_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_0_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_0_6__dout),
    .if_empty_n(fifo_A_PE_0_6__empty_n),
    .if_read(fifo_A_PE_0_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_0_6__din),
    .if_full_n(fifo_A_PE_0_6__full_n),
    .if_write(fifo_A_PE_0_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_0_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_0_7__dout),
    .if_empty_n(fifo_A_PE_0_7__empty_n),
    .if_read(fifo_A_PE_0_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_0_7__din),
    .if_full_n(fifo_A_PE_0_7__full_n),
    .if_write(fifo_A_PE_0_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_0_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_0_8__dout),
    .if_empty_n(fifo_A_PE_0_8__empty_n),
    .if_read(fifo_A_PE_0_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_0_8__din),
    .if_full_n(fifo_A_PE_0_8__full_n),
    .if_write(fifo_A_PE_0_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_0_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_0_9__dout),
    .if_empty_n(fifo_A_PE_0_9__empty_n),
    .if_read(fifo_A_PE_0_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_0_9__din),
    .if_full_n(fifo_A_PE_0_9__full_n),
    .if_write(fifo_A_PE_0_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_10_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_10_0__dout),
    .if_empty_n(fifo_A_PE_10_0__empty_n),
    .if_read(fifo_A_PE_10_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_10_0__din),
    .if_full_n(fifo_A_PE_10_0__full_n),
    .if_write(fifo_A_PE_10_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_10_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_10_1__dout),
    .if_empty_n(fifo_A_PE_10_1__empty_n),
    .if_read(fifo_A_PE_10_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_10_1__din),
    .if_full_n(fifo_A_PE_10_1__full_n),
    .if_write(fifo_A_PE_10_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_10_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_10_10__dout),
    .if_empty_n(fifo_A_PE_10_10__empty_n),
    .if_read(fifo_A_PE_10_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_10_10__din),
    .if_full_n(fifo_A_PE_10_10__full_n),
    .if_write(fifo_A_PE_10_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_10_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_10_11__dout),
    .if_empty_n(fifo_A_PE_10_11__empty_n),
    .if_read(fifo_A_PE_10_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_10_11__din),
    .if_full_n(fifo_A_PE_10_11__full_n),
    .if_write(fifo_A_PE_10_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_10_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_10_12__dout),
    .if_empty_n(fifo_A_PE_10_12__empty_n),
    .if_read(fifo_A_PE_10_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_10_12__din),
    .if_full_n(fifo_A_PE_10_12__full_n),
    .if_write(fifo_A_PE_10_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_10_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_10_13__dout),
    .if_empty_n(fifo_A_PE_10_13__empty_n),
    .if_read(fifo_A_PE_10_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_10_13__din),
    .if_full_n(fifo_A_PE_10_13__full_n),
    .if_write(fifo_A_PE_10_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_10_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_10_14__dout),
    .if_empty_n(fifo_A_PE_10_14__empty_n),
    .if_read(fifo_A_PE_10_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_10_14__din),
    .if_full_n(fifo_A_PE_10_14__full_n),
    .if_write(fifo_A_PE_10_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_10_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_10_15__dout),
    .if_empty_n(fifo_A_PE_10_15__empty_n),
    .if_read(fifo_A_PE_10_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_10_15__din),
    .if_full_n(fifo_A_PE_10_15__full_n),
    .if_write(fifo_A_PE_10_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_10_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_10_16__dout),
    .if_empty_n(fifo_A_PE_10_16__empty_n),
    .if_read(fifo_A_PE_10_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_10_16__din),
    .if_full_n(fifo_A_PE_10_16__full_n),
    .if_write(fifo_A_PE_10_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_10_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_10_17__dout),
    .if_empty_n(fifo_A_PE_10_17__empty_n),
    .if_read(fifo_A_PE_10_17__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_10_17__din),
    .if_full_n(fifo_A_PE_10_17__full_n),
    .if_write(fifo_A_PE_10_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_10_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_10_2__dout),
    .if_empty_n(fifo_A_PE_10_2__empty_n),
    .if_read(fifo_A_PE_10_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_10_2__din),
    .if_full_n(fifo_A_PE_10_2__full_n),
    .if_write(fifo_A_PE_10_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_10_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_10_3__dout),
    .if_empty_n(fifo_A_PE_10_3__empty_n),
    .if_read(fifo_A_PE_10_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_10_3__din),
    .if_full_n(fifo_A_PE_10_3__full_n),
    .if_write(fifo_A_PE_10_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_10_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_10_4__dout),
    .if_empty_n(fifo_A_PE_10_4__empty_n),
    .if_read(fifo_A_PE_10_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_10_4__din),
    .if_full_n(fifo_A_PE_10_4__full_n),
    .if_write(fifo_A_PE_10_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_10_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_10_5__dout),
    .if_empty_n(fifo_A_PE_10_5__empty_n),
    .if_read(fifo_A_PE_10_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_10_5__din),
    .if_full_n(fifo_A_PE_10_5__full_n),
    .if_write(fifo_A_PE_10_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_10_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_10_6__dout),
    .if_empty_n(fifo_A_PE_10_6__empty_n),
    .if_read(fifo_A_PE_10_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_10_6__din),
    .if_full_n(fifo_A_PE_10_6__full_n),
    .if_write(fifo_A_PE_10_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_10_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_10_7__dout),
    .if_empty_n(fifo_A_PE_10_7__empty_n),
    .if_read(fifo_A_PE_10_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_10_7__din),
    .if_full_n(fifo_A_PE_10_7__full_n),
    .if_write(fifo_A_PE_10_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_10_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_10_8__dout),
    .if_empty_n(fifo_A_PE_10_8__empty_n),
    .if_read(fifo_A_PE_10_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_10_8__din),
    .if_full_n(fifo_A_PE_10_8__full_n),
    .if_write(fifo_A_PE_10_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_10_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_10_9__dout),
    .if_empty_n(fifo_A_PE_10_9__empty_n),
    .if_read(fifo_A_PE_10_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_10_9__din),
    .if_full_n(fifo_A_PE_10_9__full_n),
    .if_write(fifo_A_PE_10_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_11_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_11_0__dout),
    .if_empty_n(fifo_A_PE_11_0__empty_n),
    .if_read(fifo_A_PE_11_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_11_0__din),
    .if_full_n(fifo_A_PE_11_0__full_n),
    .if_write(fifo_A_PE_11_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_11_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_11_1__dout),
    .if_empty_n(fifo_A_PE_11_1__empty_n),
    .if_read(fifo_A_PE_11_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_11_1__din),
    .if_full_n(fifo_A_PE_11_1__full_n),
    .if_write(fifo_A_PE_11_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_11_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_11_10__dout),
    .if_empty_n(fifo_A_PE_11_10__empty_n),
    .if_read(fifo_A_PE_11_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_11_10__din),
    .if_full_n(fifo_A_PE_11_10__full_n),
    .if_write(fifo_A_PE_11_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_11_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_11_11__dout),
    .if_empty_n(fifo_A_PE_11_11__empty_n),
    .if_read(fifo_A_PE_11_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_11_11__din),
    .if_full_n(fifo_A_PE_11_11__full_n),
    .if_write(fifo_A_PE_11_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_11_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_11_12__dout),
    .if_empty_n(fifo_A_PE_11_12__empty_n),
    .if_read(fifo_A_PE_11_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_11_12__din),
    .if_full_n(fifo_A_PE_11_12__full_n),
    .if_write(fifo_A_PE_11_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_11_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_11_13__dout),
    .if_empty_n(fifo_A_PE_11_13__empty_n),
    .if_read(fifo_A_PE_11_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_11_13__din),
    .if_full_n(fifo_A_PE_11_13__full_n),
    .if_write(fifo_A_PE_11_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_11_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_11_14__dout),
    .if_empty_n(fifo_A_PE_11_14__empty_n),
    .if_read(fifo_A_PE_11_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_11_14__din),
    .if_full_n(fifo_A_PE_11_14__full_n),
    .if_write(fifo_A_PE_11_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_11_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_11_15__dout),
    .if_empty_n(fifo_A_PE_11_15__empty_n),
    .if_read(fifo_A_PE_11_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_11_15__din),
    .if_full_n(fifo_A_PE_11_15__full_n),
    .if_write(fifo_A_PE_11_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_11_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_11_16__dout),
    .if_empty_n(fifo_A_PE_11_16__empty_n),
    .if_read(fifo_A_PE_11_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_11_16__din),
    .if_full_n(fifo_A_PE_11_16__full_n),
    .if_write(fifo_A_PE_11_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_11_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_11_17__dout),
    .if_empty_n(fifo_A_PE_11_17__empty_n),
    .if_read(fifo_A_PE_11_17__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_11_17__din),
    .if_full_n(fifo_A_PE_11_17__full_n),
    .if_write(fifo_A_PE_11_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_11_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_11_2__dout),
    .if_empty_n(fifo_A_PE_11_2__empty_n),
    .if_read(fifo_A_PE_11_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_11_2__din),
    .if_full_n(fifo_A_PE_11_2__full_n),
    .if_write(fifo_A_PE_11_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_11_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_11_3__dout),
    .if_empty_n(fifo_A_PE_11_3__empty_n),
    .if_read(fifo_A_PE_11_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_11_3__din),
    .if_full_n(fifo_A_PE_11_3__full_n),
    .if_write(fifo_A_PE_11_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_11_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_11_4__dout),
    .if_empty_n(fifo_A_PE_11_4__empty_n),
    .if_read(fifo_A_PE_11_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_11_4__din),
    .if_full_n(fifo_A_PE_11_4__full_n),
    .if_write(fifo_A_PE_11_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_11_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_11_5__dout),
    .if_empty_n(fifo_A_PE_11_5__empty_n),
    .if_read(fifo_A_PE_11_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_11_5__din),
    .if_full_n(fifo_A_PE_11_5__full_n),
    .if_write(fifo_A_PE_11_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_11_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_11_6__dout),
    .if_empty_n(fifo_A_PE_11_6__empty_n),
    .if_read(fifo_A_PE_11_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_11_6__din),
    .if_full_n(fifo_A_PE_11_6__full_n),
    .if_write(fifo_A_PE_11_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_11_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_11_7__dout),
    .if_empty_n(fifo_A_PE_11_7__empty_n),
    .if_read(fifo_A_PE_11_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_11_7__din),
    .if_full_n(fifo_A_PE_11_7__full_n),
    .if_write(fifo_A_PE_11_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_11_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_11_8__dout),
    .if_empty_n(fifo_A_PE_11_8__empty_n),
    .if_read(fifo_A_PE_11_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_11_8__din),
    .if_full_n(fifo_A_PE_11_8__full_n),
    .if_write(fifo_A_PE_11_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_11_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_11_9__dout),
    .if_empty_n(fifo_A_PE_11_9__empty_n),
    .if_read(fifo_A_PE_11_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_11_9__din),
    .if_full_n(fifo_A_PE_11_9__full_n),
    .if_write(fifo_A_PE_11_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_12_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_12_0__dout),
    .if_empty_n(fifo_A_PE_12_0__empty_n),
    .if_read(fifo_A_PE_12_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_12_0__din),
    .if_full_n(fifo_A_PE_12_0__full_n),
    .if_write(fifo_A_PE_12_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_12_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_12_1__dout),
    .if_empty_n(fifo_A_PE_12_1__empty_n),
    .if_read(fifo_A_PE_12_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_12_1__din),
    .if_full_n(fifo_A_PE_12_1__full_n),
    .if_write(fifo_A_PE_12_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_12_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_12_10__dout),
    .if_empty_n(fifo_A_PE_12_10__empty_n),
    .if_read(fifo_A_PE_12_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_12_10__din),
    .if_full_n(fifo_A_PE_12_10__full_n),
    .if_write(fifo_A_PE_12_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_12_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_12_11__dout),
    .if_empty_n(fifo_A_PE_12_11__empty_n),
    .if_read(fifo_A_PE_12_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_12_11__din),
    .if_full_n(fifo_A_PE_12_11__full_n),
    .if_write(fifo_A_PE_12_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_12_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_12_12__dout),
    .if_empty_n(fifo_A_PE_12_12__empty_n),
    .if_read(fifo_A_PE_12_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_12_12__din),
    .if_full_n(fifo_A_PE_12_12__full_n),
    .if_write(fifo_A_PE_12_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_12_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_12_13__dout),
    .if_empty_n(fifo_A_PE_12_13__empty_n),
    .if_read(fifo_A_PE_12_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_12_13__din),
    .if_full_n(fifo_A_PE_12_13__full_n),
    .if_write(fifo_A_PE_12_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_12_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_12_14__dout),
    .if_empty_n(fifo_A_PE_12_14__empty_n),
    .if_read(fifo_A_PE_12_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_12_14__din),
    .if_full_n(fifo_A_PE_12_14__full_n),
    .if_write(fifo_A_PE_12_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_12_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_12_15__dout),
    .if_empty_n(fifo_A_PE_12_15__empty_n),
    .if_read(fifo_A_PE_12_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_12_15__din),
    .if_full_n(fifo_A_PE_12_15__full_n),
    .if_write(fifo_A_PE_12_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_12_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_12_16__dout),
    .if_empty_n(fifo_A_PE_12_16__empty_n),
    .if_read(fifo_A_PE_12_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_12_16__din),
    .if_full_n(fifo_A_PE_12_16__full_n),
    .if_write(fifo_A_PE_12_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_12_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_12_17__dout),
    .if_empty_n(fifo_A_PE_12_17__empty_n),
    .if_read(fifo_A_PE_12_17__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_12_17__din),
    .if_full_n(fifo_A_PE_12_17__full_n),
    .if_write(fifo_A_PE_12_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_12_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_12_2__dout),
    .if_empty_n(fifo_A_PE_12_2__empty_n),
    .if_read(fifo_A_PE_12_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_12_2__din),
    .if_full_n(fifo_A_PE_12_2__full_n),
    .if_write(fifo_A_PE_12_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_12_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_12_3__dout),
    .if_empty_n(fifo_A_PE_12_3__empty_n),
    .if_read(fifo_A_PE_12_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_12_3__din),
    .if_full_n(fifo_A_PE_12_3__full_n),
    .if_write(fifo_A_PE_12_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_12_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_12_4__dout),
    .if_empty_n(fifo_A_PE_12_4__empty_n),
    .if_read(fifo_A_PE_12_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_12_4__din),
    .if_full_n(fifo_A_PE_12_4__full_n),
    .if_write(fifo_A_PE_12_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_12_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_12_5__dout),
    .if_empty_n(fifo_A_PE_12_5__empty_n),
    .if_read(fifo_A_PE_12_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_12_5__din),
    .if_full_n(fifo_A_PE_12_5__full_n),
    .if_write(fifo_A_PE_12_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_12_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_12_6__dout),
    .if_empty_n(fifo_A_PE_12_6__empty_n),
    .if_read(fifo_A_PE_12_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_12_6__din),
    .if_full_n(fifo_A_PE_12_6__full_n),
    .if_write(fifo_A_PE_12_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_12_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_12_7__dout),
    .if_empty_n(fifo_A_PE_12_7__empty_n),
    .if_read(fifo_A_PE_12_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_12_7__din),
    .if_full_n(fifo_A_PE_12_7__full_n),
    .if_write(fifo_A_PE_12_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_12_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_12_8__dout),
    .if_empty_n(fifo_A_PE_12_8__empty_n),
    .if_read(fifo_A_PE_12_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_12_8__din),
    .if_full_n(fifo_A_PE_12_8__full_n),
    .if_write(fifo_A_PE_12_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_12_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_12_9__dout),
    .if_empty_n(fifo_A_PE_12_9__empty_n),
    .if_read(fifo_A_PE_12_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_12_9__din),
    .if_full_n(fifo_A_PE_12_9__full_n),
    .if_write(fifo_A_PE_12_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_13_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_13_0__dout),
    .if_empty_n(fifo_A_PE_13_0__empty_n),
    .if_read(fifo_A_PE_13_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_13_0__din),
    .if_full_n(fifo_A_PE_13_0__full_n),
    .if_write(fifo_A_PE_13_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_13_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_13_1__dout),
    .if_empty_n(fifo_A_PE_13_1__empty_n),
    .if_read(fifo_A_PE_13_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_13_1__din),
    .if_full_n(fifo_A_PE_13_1__full_n),
    .if_write(fifo_A_PE_13_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_13_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_13_10__dout),
    .if_empty_n(fifo_A_PE_13_10__empty_n),
    .if_read(fifo_A_PE_13_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_13_10__din),
    .if_full_n(fifo_A_PE_13_10__full_n),
    .if_write(fifo_A_PE_13_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_13_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_13_11__dout),
    .if_empty_n(fifo_A_PE_13_11__empty_n),
    .if_read(fifo_A_PE_13_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_13_11__din),
    .if_full_n(fifo_A_PE_13_11__full_n),
    .if_write(fifo_A_PE_13_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_13_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_13_12__dout),
    .if_empty_n(fifo_A_PE_13_12__empty_n),
    .if_read(fifo_A_PE_13_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_13_12__din),
    .if_full_n(fifo_A_PE_13_12__full_n),
    .if_write(fifo_A_PE_13_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_13_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_13_13__dout),
    .if_empty_n(fifo_A_PE_13_13__empty_n),
    .if_read(fifo_A_PE_13_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_13_13__din),
    .if_full_n(fifo_A_PE_13_13__full_n),
    .if_write(fifo_A_PE_13_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_13_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_13_14__dout),
    .if_empty_n(fifo_A_PE_13_14__empty_n),
    .if_read(fifo_A_PE_13_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_13_14__din),
    .if_full_n(fifo_A_PE_13_14__full_n),
    .if_write(fifo_A_PE_13_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_13_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_13_15__dout),
    .if_empty_n(fifo_A_PE_13_15__empty_n),
    .if_read(fifo_A_PE_13_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_13_15__din),
    .if_full_n(fifo_A_PE_13_15__full_n),
    .if_write(fifo_A_PE_13_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_13_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_13_16__dout),
    .if_empty_n(fifo_A_PE_13_16__empty_n),
    .if_read(fifo_A_PE_13_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_13_16__din),
    .if_full_n(fifo_A_PE_13_16__full_n),
    .if_write(fifo_A_PE_13_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_13_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_13_17__dout),
    .if_empty_n(fifo_A_PE_13_17__empty_n),
    .if_read(fifo_A_PE_13_17__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_13_17__din),
    .if_full_n(fifo_A_PE_13_17__full_n),
    .if_write(fifo_A_PE_13_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_13_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_13_2__dout),
    .if_empty_n(fifo_A_PE_13_2__empty_n),
    .if_read(fifo_A_PE_13_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_13_2__din),
    .if_full_n(fifo_A_PE_13_2__full_n),
    .if_write(fifo_A_PE_13_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_13_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_13_3__dout),
    .if_empty_n(fifo_A_PE_13_3__empty_n),
    .if_read(fifo_A_PE_13_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_13_3__din),
    .if_full_n(fifo_A_PE_13_3__full_n),
    .if_write(fifo_A_PE_13_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_13_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_13_4__dout),
    .if_empty_n(fifo_A_PE_13_4__empty_n),
    .if_read(fifo_A_PE_13_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_13_4__din),
    .if_full_n(fifo_A_PE_13_4__full_n),
    .if_write(fifo_A_PE_13_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_13_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_13_5__dout),
    .if_empty_n(fifo_A_PE_13_5__empty_n),
    .if_read(fifo_A_PE_13_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_13_5__din),
    .if_full_n(fifo_A_PE_13_5__full_n),
    .if_write(fifo_A_PE_13_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_13_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_13_6__dout),
    .if_empty_n(fifo_A_PE_13_6__empty_n),
    .if_read(fifo_A_PE_13_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_13_6__din),
    .if_full_n(fifo_A_PE_13_6__full_n),
    .if_write(fifo_A_PE_13_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_13_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_13_7__dout),
    .if_empty_n(fifo_A_PE_13_7__empty_n),
    .if_read(fifo_A_PE_13_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_13_7__din),
    .if_full_n(fifo_A_PE_13_7__full_n),
    .if_write(fifo_A_PE_13_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_13_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_13_8__dout),
    .if_empty_n(fifo_A_PE_13_8__empty_n),
    .if_read(fifo_A_PE_13_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_13_8__din),
    .if_full_n(fifo_A_PE_13_8__full_n),
    .if_write(fifo_A_PE_13_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_13_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_13_9__dout),
    .if_empty_n(fifo_A_PE_13_9__empty_n),
    .if_read(fifo_A_PE_13_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_13_9__din),
    .if_full_n(fifo_A_PE_13_9__full_n),
    .if_write(fifo_A_PE_13_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_14_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_14_0__dout),
    .if_empty_n(fifo_A_PE_14_0__empty_n),
    .if_read(fifo_A_PE_14_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_14_0__din),
    .if_full_n(fifo_A_PE_14_0__full_n),
    .if_write(fifo_A_PE_14_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_14_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_14_1__dout),
    .if_empty_n(fifo_A_PE_14_1__empty_n),
    .if_read(fifo_A_PE_14_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_14_1__din),
    .if_full_n(fifo_A_PE_14_1__full_n),
    .if_write(fifo_A_PE_14_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_14_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_14_10__dout),
    .if_empty_n(fifo_A_PE_14_10__empty_n),
    .if_read(fifo_A_PE_14_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_14_10__din),
    .if_full_n(fifo_A_PE_14_10__full_n),
    .if_write(fifo_A_PE_14_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_14_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_14_11__dout),
    .if_empty_n(fifo_A_PE_14_11__empty_n),
    .if_read(fifo_A_PE_14_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_14_11__din),
    .if_full_n(fifo_A_PE_14_11__full_n),
    .if_write(fifo_A_PE_14_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_14_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_14_12__dout),
    .if_empty_n(fifo_A_PE_14_12__empty_n),
    .if_read(fifo_A_PE_14_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_14_12__din),
    .if_full_n(fifo_A_PE_14_12__full_n),
    .if_write(fifo_A_PE_14_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_14_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_14_13__dout),
    .if_empty_n(fifo_A_PE_14_13__empty_n),
    .if_read(fifo_A_PE_14_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_14_13__din),
    .if_full_n(fifo_A_PE_14_13__full_n),
    .if_write(fifo_A_PE_14_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_14_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_14_14__dout),
    .if_empty_n(fifo_A_PE_14_14__empty_n),
    .if_read(fifo_A_PE_14_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_14_14__din),
    .if_full_n(fifo_A_PE_14_14__full_n),
    .if_write(fifo_A_PE_14_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_14_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_14_15__dout),
    .if_empty_n(fifo_A_PE_14_15__empty_n),
    .if_read(fifo_A_PE_14_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_14_15__din),
    .if_full_n(fifo_A_PE_14_15__full_n),
    .if_write(fifo_A_PE_14_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_14_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_14_16__dout),
    .if_empty_n(fifo_A_PE_14_16__empty_n),
    .if_read(fifo_A_PE_14_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_14_16__din),
    .if_full_n(fifo_A_PE_14_16__full_n),
    .if_write(fifo_A_PE_14_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_14_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_14_17__dout),
    .if_empty_n(fifo_A_PE_14_17__empty_n),
    .if_read(fifo_A_PE_14_17__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_14_17__din),
    .if_full_n(fifo_A_PE_14_17__full_n),
    .if_write(fifo_A_PE_14_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_14_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_14_2__dout),
    .if_empty_n(fifo_A_PE_14_2__empty_n),
    .if_read(fifo_A_PE_14_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_14_2__din),
    .if_full_n(fifo_A_PE_14_2__full_n),
    .if_write(fifo_A_PE_14_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_14_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_14_3__dout),
    .if_empty_n(fifo_A_PE_14_3__empty_n),
    .if_read(fifo_A_PE_14_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_14_3__din),
    .if_full_n(fifo_A_PE_14_3__full_n),
    .if_write(fifo_A_PE_14_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_14_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_14_4__dout),
    .if_empty_n(fifo_A_PE_14_4__empty_n),
    .if_read(fifo_A_PE_14_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_14_4__din),
    .if_full_n(fifo_A_PE_14_4__full_n),
    .if_write(fifo_A_PE_14_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_14_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_14_5__dout),
    .if_empty_n(fifo_A_PE_14_5__empty_n),
    .if_read(fifo_A_PE_14_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_14_5__din),
    .if_full_n(fifo_A_PE_14_5__full_n),
    .if_write(fifo_A_PE_14_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_14_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_14_6__dout),
    .if_empty_n(fifo_A_PE_14_6__empty_n),
    .if_read(fifo_A_PE_14_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_14_6__din),
    .if_full_n(fifo_A_PE_14_6__full_n),
    .if_write(fifo_A_PE_14_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_14_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_14_7__dout),
    .if_empty_n(fifo_A_PE_14_7__empty_n),
    .if_read(fifo_A_PE_14_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_14_7__din),
    .if_full_n(fifo_A_PE_14_7__full_n),
    .if_write(fifo_A_PE_14_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_14_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_14_8__dout),
    .if_empty_n(fifo_A_PE_14_8__empty_n),
    .if_read(fifo_A_PE_14_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_14_8__din),
    .if_full_n(fifo_A_PE_14_8__full_n),
    .if_write(fifo_A_PE_14_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_14_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_14_9__dout),
    .if_empty_n(fifo_A_PE_14_9__empty_n),
    .if_read(fifo_A_PE_14_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_14_9__din),
    .if_full_n(fifo_A_PE_14_9__full_n),
    .if_write(fifo_A_PE_14_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_15_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_15_0__dout),
    .if_empty_n(fifo_A_PE_15_0__empty_n),
    .if_read(fifo_A_PE_15_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_15_0__din),
    .if_full_n(fifo_A_PE_15_0__full_n),
    .if_write(fifo_A_PE_15_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_15_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_15_1__dout),
    .if_empty_n(fifo_A_PE_15_1__empty_n),
    .if_read(fifo_A_PE_15_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_15_1__din),
    .if_full_n(fifo_A_PE_15_1__full_n),
    .if_write(fifo_A_PE_15_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_15_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_15_10__dout),
    .if_empty_n(fifo_A_PE_15_10__empty_n),
    .if_read(fifo_A_PE_15_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_15_10__din),
    .if_full_n(fifo_A_PE_15_10__full_n),
    .if_write(fifo_A_PE_15_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_15_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_15_11__dout),
    .if_empty_n(fifo_A_PE_15_11__empty_n),
    .if_read(fifo_A_PE_15_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_15_11__din),
    .if_full_n(fifo_A_PE_15_11__full_n),
    .if_write(fifo_A_PE_15_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_15_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_15_12__dout),
    .if_empty_n(fifo_A_PE_15_12__empty_n),
    .if_read(fifo_A_PE_15_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_15_12__din),
    .if_full_n(fifo_A_PE_15_12__full_n),
    .if_write(fifo_A_PE_15_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_15_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_15_13__dout),
    .if_empty_n(fifo_A_PE_15_13__empty_n),
    .if_read(fifo_A_PE_15_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_15_13__din),
    .if_full_n(fifo_A_PE_15_13__full_n),
    .if_write(fifo_A_PE_15_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_15_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_15_14__dout),
    .if_empty_n(fifo_A_PE_15_14__empty_n),
    .if_read(fifo_A_PE_15_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_15_14__din),
    .if_full_n(fifo_A_PE_15_14__full_n),
    .if_write(fifo_A_PE_15_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_15_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_15_15__dout),
    .if_empty_n(fifo_A_PE_15_15__empty_n),
    .if_read(fifo_A_PE_15_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_15_15__din),
    .if_full_n(fifo_A_PE_15_15__full_n),
    .if_write(fifo_A_PE_15_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_15_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_15_16__dout),
    .if_empty_n(fifo_A_PE_15_16__empty_n),
    .if_read(fifo_A_PE_15_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_15_16__din),
    .if_full_n(fifo_A_PE_15_16__full_n),
    .if_write(fifo_A_PE_15_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_15_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_15_17__dout),
    .if_empty_n(fifo_A_PE_15_17__empty_n),
    .if_read(fifo_A_PE_15_17__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_15_17__din),
    .if_full_n(fifo_A_PE_15_17__full_n),
    .if_write(fifo_A_PE_15_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_15_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_15_2__dout),
    .if_empty_n(fifo_A_PE_15_2__empty_n),
    .if_read(fifo_A_PE_15_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_15_2__din),
    .if_full_n(fifo_A_PE_15_2__full_n),
    .if_write(fifo_A_PE_15_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_15_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_15_3__dout),
    .if_empty_n(fifo_A_PE_15_3__empty_n),
    .if_read(fifo_A_PE_15_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_15_3__din),
    .if_full_n(fifo_A_PE_15_3__full_n),
    .if_write(fifo_A_PE_15_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_15_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_15_4__dout),
    .if_empty_n(fifo_A_PE_15_4__empty_n),
    .if_read(fifo_A_PE_15_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_15_4__din),
    .if_full_n(fifo_A_PE_15_4__full_n),
    .if_write(fifo_A_PE_15_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_15_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_15_5__dout),
    .if_empty_n(fifo_A_PE_15_5__empty_n),
    .if_read(fifo_A_PE_15_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_15_5__din),
    .if_full_n(fifo_A_PE_15_5__full_n),
    .if_write(fifo_A_PE_15_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_15_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_15_6__dout),
    .if_empty_n(fifo_A_PE_15_6__empty_n),
    .if_read(fifo_A_PE_15_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_15_6__din),
    .if_full_n(fifo_A_PE_15_6__full_n),
    .if_write(fifo_A_PE_15_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_15_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_15_7__dout),
    .if_empty_n(fifo_A_PE_15_7__empty_n),
    .if_read(fifo_A_PE_15_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_15_7__din),
    .if_full_n(fifo_A_PE_15_7__full_n),
    .if_write(fifo_A_PE_15_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_15_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_15_8__dout),
    .if_empty_n(fifo_A_PE_15_8__empty_n),
    .if_read(fifo_A_PE_15_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_15_8__din),
    .if_full_n(fifo_A_PE_15_8__full_n),
    .if_write(fifo_A_PE_15_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_15_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_15_9__dout),
    .if_empty_n(fifo_A_PE_15_9__empty_n),
    .if_read(fifo_A_PE_15_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_15_9__din),
    .if_full_n(fifo_A_PE_15_9__full_n),
    .if_write(fifo_A_PE_15_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_16_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_16_0__dout),
    .if_empty_n(fifo_A_PE_16_0__empty_n),
    .if_read(fifo_A_PE_16_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_16_0__din),
    .if_full_n(fifo_A_PE_16_0__full_n),
    .if_write(fifo_A_PE_16_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_16_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_16_1__dout),
    .if_empty_n(fifo_A_PE_16_1__empty_n),
    .if_read(fifo_A_PE_16_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_16_1__din),
    .if_full_n(fifo_A_PE_16_1__full_n),
    .if_write(fifo_A_PE_16_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_16_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_16_10__dout),
    .if_empty_n(fifo_A_PE_16_10__empty_n),
    .if_read(fifo_A_PE_16_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_16_10__din),
    .if_full_n(fifo_A_PE_16_10__full_n),
    .if_write(fifo_A_PE_16_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_16_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_16_11__dout),
    .if_empty_n(fifo_A_PE_16_11__empty_n),
    .if_read(fifo_A_PE_16_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_16_11__din),
    .if_full_n(fifo_A_PE_16_11__full_n),
    .if_write(fifo_A_PE_16_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_16_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_16_12__dout),
    .if_empty_n(fifo_A_PE_16_12__empty_n),
    .if_read(fifo_A_PE_16_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_16_12__din),
    .if_full_n(fifo_A_PE_16_12__full_n),
    .if_write(fifo_A_PE_16_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_16_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_16_13__dout),
    .if_empty_n(fifo_A_PE_16_13__empty_n),
    .if_read(fifo_A_PE_16_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_16_13__din),
    .if_full_n(fifo_A_PE_16_13__full_n),
    .if_write(fifo_A_PE_16_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_16_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_16_14__dout),
    .if_empty_n(fifo_A_PE_16_14__empty_n),
    .if_read(fifo_A_PE_16_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_16_14__din),
    .if_full_n(fifo_A_PE_16_14__full_n),
    .if_write(fifo_A_PE_16_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_16_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_16_15__dout),
    .if_empty_n(fifo_A_PE_16_15__empty_n),
    .if_read(fifo_A_PE_16_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_16_15__din),
    .if_full_n(fifo_A_PE_16_15__full_n),
    .if_write(fifo_A_PE_16_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_16_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_16_16__dout),
    .if_empty_n(fifo_A_PE_16_16__empty_n),
    .if_read(fifo_A_PE_16_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_16_16__din),
    .if_full_n(fifo_A_PE_16_16__full_n),
    .if_write(fifo_A_PE_16_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_16_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_16_17__dout),
    .if_empty_n(fifo_A_PE_16_17__empty_n),
    .if_read(fifo_A_PE_16_17__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_16_17__din),
    .if_full_n(fifo_A_PE_16_17__full_n),
    .if_write(fifo_A_PE_16_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_16_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_16_2__dout),
    .if_empty_n(fifo_A_PE_16_2__empty_n),
    .if_read(fifo_A_PE_16_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_16_2__din),
    .if_full_n(fifo_A_PE_16_2__full_n),
    .if_write(fifo_A_PE_16_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_16_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_16_3__dout),
    .if_empty_n(fifo_A_PE_16_3__empty_n),
    .if_read(fifo_A_PE_16_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_16_3__din),
    .if_full_n(fifo_A_PE_16_3__full_n),
    .if_write(fifo_A_PE_16_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_16_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_16_4__dout),
    .if_empty_n(fifo_A_PE_16_4__empty_n),
    .if_read(fifo_A_PE_16_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_16_4__din),
    .if_full_n(fifo_A_PE_16_4__full_n),
    .if_write(fifo_A_PE_16_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_16_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_16_5__dout),
    .if_empty_n(fifo_A_PE_16_5__empty_n),
    .if_read(fifo_A_PE_16_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_16_5__din),
    .if_full_n(fifo_A_PE_16_5__full_n),
    .if_write(fifo_A_PE_16_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_16_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_16_6__dout),
    .if_empty_n(fifo_A_PE_16_6__empty_n),
    .if_read(fifo_A_PE_16_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_16_6__din),
    .if_full_n(fifo_A_PE_16_6__full_n),
    .if_write(fifo_A_PE_16_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_16_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_16_7__dout),
    .if_empty_n(fifo_A_PE_16_7__empty_n),
    .if_read(fifo_A_PE_16_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_16_7__din),
    .if_full_n(fifo_A_PE_16_7__full_n),
    .if_write(fifo_A_PE_16_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_16_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_16_8__dout),
    .if_empty_n(fifo_A_PE_16_8__empty_n),
    .if_read(fifo_A_PE_16_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_16_8__din),
    .if_full_n(fifo_A_PE_16_8__full_n),
    .if_write(fifo_A_PE_16_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_16_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_16_9__dout),
    .if_empty_n(fifo_A_PE_16_9__empty_n),
    .if_read(fifo_A_PE_16_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_16_9__din),
    .if_full_n(fifo_A_PE_16_9__full_n),
    .if_write(fifo_A_PE_16_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_17_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_17_0__dout),
    .if_empty_n(fifo_A_PE_17_0__empty_n),
    .if_read(fifo_A_PE_17_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_17_0__din),
    .if_full_n(fifo_A_PE_17_0__full_n),
    .if_write(fifo_A_PE_17_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_17_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_17_1__dout),
    .if_empty_n(fifo_A_PE_17_1__empty_n),
    .if_read(fifo_A_PE_17_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_17_1__din),
    .if_full_n(fifo_A_PE_17_1__full_n),
    .if_write(fifo_A_PE_17_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_17_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_17_10__dout),
    .if_empty_n(fifo_A_PE_17_10__empty_n),
    .if_read(fifo_A_PE_17_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_17_10__din),
    .if_full_n(fifo_A_PE_17_10__full_n),
    .if_write(fifo_A_PE_17_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_17_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_17_11__dout),
    .if_empty_n(fifo_A_PE_17_11__empty_n),
    .if_read(fifo_A_PE_17_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_17_11__din),
    .if_full_n(fifo_A_PE_17_11__full_n),
    .if_write(fifo_A_PE_17_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_17_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_17_12__dout),
    .if_empty_n(fifo_A_PE_17_12__empty_n),
    .if_read(fifo_A_PE_17_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_17_12__din),
    .if_full_n(fifo_A_PE_17_12__full_n),
    .if_write(fifo_A_PE_17_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_17_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_17_13__dout),
    .if_empty_n(fifo_A_PE_17_13__empty_n),
    .if_read(fifo_A_PE_17_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_17_13__din),
    .if_full_n(fifo_A_PE_17_13__full_n),
    .if_write(fifo_A_PE_17_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_17_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_17_14__dout),
    .if_empty_n(fifo_A_PE_17_14__empty_n),
    .if_read(fifo_A_PE_17_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_17_14__din),
    .if_full_n(fifo_A_PE_17_14__full_n),
    .if_write(fifo_A_PE_17_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_17_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_17_15__dout),
    .if_empty_n(fifo_A_PE_17_15__empty_n),
    .if_read(fifo_A_PE_17_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_17_15__din),
    .if_full_n(fifo_A_PE_17_15__full_n),
    .if_write(fifo_A_PE_17_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_17_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_17_16__dout),
    .if_empty_n(fifo_A_PE_17_16__empty_n),
    .if_read(fifo_A_PE_17_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_17_16__din),
    .if_full_n(fifo_A_PE_17_16__full_n),
    .if_write(fifo_A_PE_17_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_17_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_17_17__dout),
    .if_empty_n(fifo_A_PE_17_17__empty_n),
    .if_read(fifo_A_PE_17_17__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_17_17__din),
    .if_full_n(fifo_A_PE_17_17__full_n),
    .if_write(fifo_A_PE_17_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_17_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_17_2__dout),
    .if_empty_n(fifo_A_PE_17_2__empty_n),
    .if_read(fifo_A_PE_17_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_17_2__din),
    .if_full_n(fifo_A_PE_17_2__full_n),
    .if_write(fifo_A_PE_17_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_17_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_17_3__dout),
    .if_empty_n(fifo_A_PE_17_3__empty_n),
    .if_read(fifo_A_PE_17_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_17_3__din),
    .if_full_n(fifo_A_PE_17_3__full_n),
    .if_write(fifo_A_PE_17_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_17_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_17_4__dout),
    .if_empty_n(fifo_A_PE_17_4__empty_n),
    .if_read(fifo_A_PE_17_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_17_4__din),
    .if_full_n(fifo_A_PE_17_4__full_n),
    .if_write(fifo_A_PE_17_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_17_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_17_5__dout),
    .if_empty_n(fifo_A_PE_17_5__empty_n),
    .if_read(fifo_A_PE_17_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_17_5__din),
    .if_full_n(fifo_A_PE_17_5__full_n),
    .if_write(fifo_A_PE_17_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_17_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_17_6__dout),
    .if_empty_n(fifo_A_PE_17_6__empty_n),
    .if_read(fifo_A_PE_17_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_17_6__din),
    .if_full_n(fifo_A_PE_17_6__full_n),
    .if_write(fifo_A_PE_17_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_17_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_17_7__dout),
    .if_empty_n(fifo_A_PE_17_7__empty_n),
    .if_read(fifo_A_PE_17_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_17_7__din),
    .if_full_n(fifo_A_PE_17_7__full_n),
    .if_write(fifo_A_PE_17_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_17_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_17_8__dout),
    .if_empty_n(fifo_A_PE_17_8__empty_n),
    .if_read(fifo_A_PE_17_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_17_8__din),
    .if_full_n(fifo_A_PE_17_8__full_n),
    .if_write(fifo_A_PE_17_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_17_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_17_9__dout),
    .if_empty_n(fifo_A_PE_17_9__empty_n),
    .if_read(fifo_A_PE_17_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_17_9__din),
    .if_full_n(fifo_A_PE_17_9__full_n),
    .if_write(fifo_A_PE_17_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_1_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_1_0__dout),
    .if_empty_n(fifo_A_PE_1_0__empty_n),
    .if_read(fifo_A_PE_1_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_1_0__din),
    .if_full_n(fifo_A_PE_1_0__full_n),
    .if_write(fifo_A_PE_1_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_1_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_1_1__dout),
    .if_empty_n(fifo_A_PE_1_1__empty_n),
    .if_read(fifo_A_PE_1_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_1_1__din),
    .if_full_n(fifo_A_PE_1_1__full_n),
    .if_write(fifo_A_PE_1_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_1_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_1_10__dout),
    .if_empty_n(fifo_A_PE_1_10__empty_n),
    .if_read(fifo_A_PE_1_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_1_10__din),
    .if_full_n(fifo_A_PE_1_10__full_n),
    .if_write(fifo_A_PE_1_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_1_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_1_11__dout),
    .if_empty_n(fifo_A_PE_1_11__empty_n),
    .if_read(fifo_A_PE_1_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_1_11__din),
    .if_full_n(fifo_A_PE_1_11__full_n),
    .if_write(fifo_A_PE_1_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_1_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_1_12__dout),
    .if_empty_n(fifo_A_PE_1_12__empty_n),
    .if_read(fifo_A_PE_1_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_1_12__din),
    .if_full_n(fifo_A_PE_1_12__full_n),
    .if_write(fifo_A_PE_1_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_1_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_1_13__dout),
    .if_empty_n(fifo_A_PE_1_13__empty_n),
    .if_read(fifo_A_PE_1_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_1_13__din),
    .if_full_n(fifo_A_PE_1_13__full_n),
    .if_write(fifo_A_PE_1_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_1_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_1_14__dout),
    .if_empty_n(fifo_A_PE_1_14__empty_n),
    .if_read(fifo_A_PE_1_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_1_14__din),
    .if_full_n(fifo_A_PE_1_14__full_n),
    .if_write(fifo_A_PE_1_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_1_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_1_15__dout),
    .if_empty_n(fifo_A_PE_1_15__empty_n),
    .if_read(fifo_A_PE_1_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_1_15__din),
    .if_full_n(fifo_A_PE_1_15__full_n),
    .if_write(fifo_A_PE_1_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_1_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_1_16__dout),
    .if_empty_n(fifo_A_PE_1_16__empty_n),
    .if_read(fifo_A_PE_1_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_1_16__din),
    .if_full_n(fifo_A_PE_1_16__full_n),
    .if_write(fifo_A_PE_1_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_1_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_1_17__dout),
    .if_empty_n(fifo_A_PE_1_17__empty_n),
    .if_read(fifo_A_PE_1_17__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_1_17__din),
    .if_full_n(fifo_A_PE_1_17__full_n),
    .if_write(fifo_A_PE_1_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_1_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_1_2__dout),
    .if_empty_n(fifo_A_PE_1_2__empty_n),
    .if_read(fifo_A_PE_1_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_1_2__din),
    .if_full_n(fifo_A_PE_1_2__full_n),
    .if_write(fifo_A_PE_1_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_1_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_1_3__dout),
    .if_empty_n(fifo_A_PE_1_3__empty_n),
    .if_read(fifo_A_PE_1_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_1_3__din),
    .if_full_n(fifo_A_PE_1_3__full_n),
    .if_write(fifo_A_PE_1_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_1_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_1_4__dout),
    .if_empty_n(fifo_A_PE_1_4__empty_n),
    .if_read(fifo_A_PE_1_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_1_4__din),
    .if_full_n(fifo_A_PE_1_4__full_n),
    .if_write(fifo_A_PE_1_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_1_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_1_5__dout),
    .if_empty_n(fifo_A_PE_1_5__empty_n),
    .if_read(fifo_A_PE_1_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_1_5__din),
    .if_full_n(fifo_A_PE_1_5__full_n),
    .if_write(fifo_A_PE_1_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_1_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_1_6__dout),
    .if_empty_n(fifo_A_PE_1_6__empty_n),
    .if_read(fifo_A_PE_1_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_1_6__din),
    .if_full_n(fifo_A_PE_1_6__full_n),
    .if_write(fifo_A_PE_1_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_1_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_1_7__dout),
    .if_empty_n(fifo_A_PE_1_7__empty_n),
    .if_read(fifo_A_PE_1_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_1_7__din),
    .if_full_n(fifo_A_PE_1_7__full_n),
    .if_write(fifo_A_PE_1_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_1_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_1_8__dout),
    .if_empty_n(fifo_A_PE_1_8__empty_n),
    .if_read(fifo_A_PE_1_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_1_8__din),
    .if_full_n(fifo_A_PE_1_8__full_n),
    .if_write(fifo_A_PE_1_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_1_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_1_9__dout),
    .if_empty_n(fifo_A_PE_1_9__empty_n),
    .if_read(fifo_A_PE_1_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_1_9__din),
    .if_full_n(fifo_A_PE_1_9__full_n),
    .if_write(fifo_A_PE_1_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_2_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_2_0__dout),
    .if_empty_n(fifo_A_PE_2_0__empty_n),
    .if_read(fifo_A_PE_2_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_2_0__din),
    .if_full_n(fifo_A_PE_2_0__full_n),
    .if_write(fifo_A_PE_2_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_2_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_2_1__dout),
    .if_empty_n(fifo_A_PE_2_1__empty_n),
    .if_read(fifo_A_PE_2_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_2_1__din),
    .if_full_n(fifo_A_PE_2_1__full_n),
    .if_write(fifo_A_PE_2_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_2_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_2_10__dout),
    .if_empty_n(fifo_A_PE_2_10__empty_n),
    .if_read(fifo_A_PE_2_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_2_10__din),
    .if_full_n(fifo_A_PE_2_10__full_n),
    .if_write(fifo_A_PE_2_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_2_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_2_11__dout),
    .if_empty_n(fifo_A_PE_2_11__empty_n),
    .if_read(fifo_A_PE_2_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_2_11__din),
    .if_full_n(fifo_A_PE_2_11__full_n),
    .if_write(fifo_A_PE_2_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_2_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_2_12__dout),
    .if_empty_n(fifo_A_PE_2_12__empty_n),
    .if_read(fifo_A_PE_2_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_2_12__din),
    .if_full_n(fifo_A_PE_2_12__full_n),
    .if_write(fifo_A_PE_2_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_2_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_2_13__dout),
    .if_empty_n(fifo_A_PE_2_13__empty_n),
    .if_read(fifo_A_PE_2_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_2_13__din),
    .if_full_n(fifo_A_PE_2_13__full_n),
    .if_write(fifo_A_PE_2_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_2_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_2_14__dout),
    .if_empty_n(fifo_A_PE_2_14__empty_n),
    .if_read(fifo_A_PE_2_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_2_14__din),
    .if_full_n(fifo_A_PE_2_14__full_n),
    .if_write(fifo_A_PE_2_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_2_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_2_15__dout),
    .if_empty_n(fifo_A_PE_2_15__empty_n),
    .if_read(fifo_A_PE_2_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_2_15__din),
    .if_full_n(fifo_A_PE_2_15__full_n),
    .if_write(fifo_A_PE_2_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_2_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_2_16__dout),
    .if_empty_n(fifo_A_PE_2_16__empty_n),
    .if_read(fifo_A_PE_2_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_2_16__din),
    .if_full_n(fifo_A_PE_2_16__full_n),
    .if_write(fifo_A_PE_2_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_2_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_2_17__dout),
    .if_empty_n(fifo_A_PE_2_17__empty_n),
    .if_read(fifo_A_PE_2_17__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_2_17__din),
    .if_full_n(fifo_A_PE_2_17__full_n),
    .if_write(fifo_A_PE_2_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_2_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_2_2__dout),
    .if_empty_n(fifo_A_PE_2_2__empty_n),
    .if_read(fifo_A_PE_2_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_2_2__din),
    .if_full_n(fifo_A_PE_2_2__full_n),
    .if_write(fifo_A_PE_2_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_2_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_2_3__dout),
    .if_empty_n(fifo_A_PE_2_3__empty_n),
    .if_read(fifo_A_PE_2_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_2_3__din),
    .if_full_n(fifo_A_PE_2_3__full_n),
    .if_write(fifo_A_PE_2_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_2_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_2_4__dout),
    .if_empty_n(fifo_A_PE_2_4__empty_n),
    .if_read(fifo_A_PE_2_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_2_4__din),
    .if_full_n(fifo_A_PE_2_4__full_n),
    .if_write(fifo_A_PE_2_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_2_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_2_5__dout),
    .if_empty_n(fifo_A_PE_2_5__empty_n),
    .if_read(fifo_A_PE_2_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_2_5__din),
    .if_full_n(fifo_A_PE_2_5__full_n),
    .if_write(fifo_A_PE_2_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_2_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_2_6__dout),
    .if_empty_n(fifo_A_PE_2_6__empty_n),
    .if_read(fifo_A_PE_2_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_2_6__din),
    .if_full_n(fifo_A_PE_2_6__full_n),
    .if_write(fifo_A_PE_2_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_2_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_2_7__dout),
    .if_empty_n(fifo_A_PE_2_7__empty_n),
    .if_read(fifo_A_PE_2_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_2_7__din),
    .if_full_n(fifo_A_PE_2_7__full_n),
    .if_write(fifo_A_PE_2_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_2_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_2_8__dout),
    .if_empty_n(fifo_A_PE_2_8__empty_n),
    .if_read(fifo_A_PE_2_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_2_8__din),
    .if_full_n(fifo_A_PE_2_8__full_n),
    .if_write(fifo_A_PE_2_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_2_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_2_9__dout),
    .if_empty_n(fifo_A_PE_2_9__empty_n),
    .if_read(fifo_A_PE_2_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_2_9__din),
    .if_full_n(fifo_A_PE_2_9__full_n),
    .if_write(fifo_A_PE_2_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_3_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_3_0__dout),
    .if_empty_n(fifo_A_PE_3_0__empty_n),
    .if_read(fifo_A_PE_3_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_3_0__din),
    .if_full_n(fifo_A_PE_3_0__full_n),
    .if_write(fifo_A_PE_3_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_3_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_3_1__dout),
    .if_empty_n(fifo_A_PE_3_1__empty_n),
    .if_read(fifo_A_PE_3_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_3_1__din),
    .if_full_n(fifo_A_PE_3_1__full_n),
    .if_write(fifo_A_PE_3_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_3_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_3_10__dout),
    .if_empty_n(fifo_A_PE_3_10__empty_n),
    .if_read(fifo_A_PE_3_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_3_10__din),
    .if_full_n(fifo_A_PE_3_10__full_n),
    .if_write(fifo_A_PE_3_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_3_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_3_11__dout),
    .if_empty_n(fifo_A_PE_3_11__empty_n),
    .if_read(fifo_A_PE_3_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_3_11__din),
    .if_full_n(fifo_A_PE_3_11__full_n),
    .if_write(fifo_A_PE_3_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_3_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_3_12__dout),
    .if_empty_n(fifo_A_PE_3_12__empty_n),
    .if_read(fifo_A_PE_3_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_3_12__din),
    .if_full_n(fifo_A_PE_3_12__full_n),
    .if_write(fifo_A_PE_3_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_3_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_3_13__dout),
    .if_empty_n(fifo_A_PE_3_13__empty_n),
    .if_read(fifo_A_PE_3_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_3_13__din),
    .if_full_n(fifo_A_PE_3_13__full_n),
    .if_write(fifo_A_PE_3_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_3_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_3_14__dout),
    .if_empty_n(fifo_A_PE_3_14__empty_n),
    .if_read(fifo_A_PE_3_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_3_14__din),
    .if_full_n(fifo_A_PE_3_14__full_n),
    .if_write(fifo_A_PE_3_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_3_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_3_15__dout),
    .if_empty_n(fifo_A_PE_3_15__empty_n),
    .if_read(fifo_A_PE_3_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_3_15__din),
    .if_full_n(fifo_A_PE_3_15__full_n),
    .if_write(fifo_A_PE_3_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_3_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_3_16__dout),
    .if_empty_n(fifo_A_PE_3_16__empty_n),
    .if_read(fifo_A_PE_3_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_3_16__din),
    .if_full_n(fifo_A_PE_3_16__full_n),
    .if_write(fifo_A_PE_3_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_3_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_3_17__dout),
    .if_empty_n(fifo_A_PE_3_17__empty_n),
    .if_read(fifo_A_PE_3_17__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_3_17__din),
    .if_full_n(fifo_A_PE_3_17__full_n),
    .if_write(fifo_A_PE_3_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_3_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_3_2__dout),
    .if_empty_n(fifo_A_PE_3_2__empty_n),
    .if_read(fifo_A_PE_3_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_3_2__din),
    .if_full_n(fifo_A_PE_3_2__full_n),
    .if_write(fifo_A_PE_3_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_3_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_3_3__dout),
    .if_empty_n(fifo_A_PE_3_3__empty_n),
    .if_read(fifo_A_PE_3_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_3_3__din),
    .if_full_n(fifo_A_PE_3_3__full_n),
    .if_write(fifo_A_PE_3_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_3_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_3_4__dout),
    .if_empty_n(fifo_A_PE_3_4__empty_n),
    .if_read(fifo_A_PE_3_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_3_4__din),
    .if_full_n(fifo_A_PE_3_4__full_n),
    .if_write(fifo_A_PE_3_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_3_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_3_5__dout),
    .if_empty_n(fifo_A_PE_3_5__empty_n),
    .if_read(fifo_A_PE_3_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_3_5__din),
    .if_full_n(fifo_A_PE_3_5__full_n),
    .if_write(fifo_A_PE_3_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_3_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_3_6__dout),
    .if_empty_n(fifo_A_PE_3_6__empty_n),
    .if_read(fifo_A_PE_3_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_3_6__din),
    .if_full_n(fifo_A_PE_3_6__full_n),
    .if_write(fifo_A_PE_3_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_3_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_3_7__dout),
    .if_empty_n(fifo_A_PE_3_7__empty_n),
    .if_read(fifo_A_PE_3_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_3_7__din),
    .if_full_n(fifo_A_PE_3_7__full_n),
    .if_write(fifo_A_PE_3_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_3_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_3_8__dout),
    .if_empty_n(fifo_A_PE_3_8__empty_n),
    .if_read(fifo_A_PE_3_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_3_8__din),
    .if_full_n(fifo_A_PE_3_8__full_n),
    .if_write(fifo_A_PE_3_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_3_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_3_9__dout),
    .if_empty_n(fifo_A_PE_3_9__empty_n),
    .if_read(fifo_A_PE_3_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_3_9__din),
    .if_full_n(fifo_A_PE_3_9__full_n),
    .if_write(fifo_A_PE_3_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_4_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_4_0__dout),
    .if_empty_n(fifo_A_PE_4_0__empty_n),
    .if_read(fifo_A_PE_4_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_4_0__din),
    .if_full_n(fifo_A_PE_4_0__full_n),
    .if_write(fifo_A_PE_4_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_4_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_4_1__dout),
    .if_empty_n(fifo_A_PE_4_1__empty_n),
    .if_read(fifo_A_PE_4_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_4_1__din),
    .if_full_n(fifo_A_PE_4_1__full_n),
    .if_write(fifo_A_PE_4_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_4_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_4_10__dout),
    .if_empty_n(fifo_A_PE_4_10__empty_n),
    .if_read(fifo_A_PE_4_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_4_10__din),
    .if_full_n(fifo_A_PE_4_10__full_n),
    .if_write(fifo_A_PE_4_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_4_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_4_11__dout),
    .if_empty_n(fifo_A_PE_4_11__empty_n),
    .if_read(fifo_A_PE_4_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_4_11__din),
    .if_full_n(fifo_A_PE_4_11__full_n),
    .if_write(fifo_A_PE_4_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_4_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_4_12__dout),
    .if_empty_n(fifo_A_PE_4_12__empty_n),
    .if_read(fifo_A_PE_4_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_4_12__din),
    .if_full_n(fifo_A_PE_4_12__full_n),
    .if_write(fifo_A_PE_4_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_4_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_4_13__dout),
    .if_empty_n(fifo_A_PE_4_13__empty_n),
    .if_read(fifo_A_PE_4_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_4_13__din),
    .if_full_n(fifo_A_PE_4_13__full_n),
    .if_write(fifo_A_PE_4_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_4_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_4_14__dout),
    .if_empty_n(fifo_A_PE_4_14__empty_n),
    .if_read(fifo_A_PE_4_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_4_14__din),
    .if_full_n(fifo_A_PE_4_14__full_n),
    .if_write(fifo_A_PE_4_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_4_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_4_15__dout),
    .if_empty_n(fifo_A_PE_4_15__empty_n),
    .if_read(fifo_A_PE_4_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_4_15__din),
    .if_full_n(fifo_A_PE_4_15__full_n),
    .if_write(fifo_A_PE_4_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_4_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_4_16__dout),
    .if_empty_n(fifo_A_PE_4_16__empty_n),
    .if_read(fifo_A_PE_4_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_4_16__din),
    .if_full_n(fifo_A_PE_4_16__full_n),
    .if_write(fifo_A_PE_4_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_4_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_4_17__dout),
    .if_empty_n(fifo_A_PE_4_17__empty_n),
    .if_read(fifo_A_PE_4_17__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_4_17__din),
    .if_full_n(fifo_A_PE_4_17__full_n),
    .if_write(fifo_A_PE_4_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_4_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_4_2__dout),
    .if_empty_n(fifo_A_PE_4_2__empty_n),
    .if_read(fifo_A_PE_4_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_4_2__din),
    .if_full_n(fifo_A_PE_4_2__full_n),
    .if_write(fifo_A_PE_4_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_4_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_4_3__dout),
    .if_empty_n(fifo_A_PE_4_3__empty_n),
    .if_read(fifo_A_PE_4_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_4_3__din),
    .if_full_n(fifo_A_PE_4_3__full_n),
    .if_write(fifo_A_PE_4_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_4_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_4_4__dout),
    .if_empty_n(fifo_A_PE_4_4__empty_n),
    .if_read(fifo_A_PE_4_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_4_4__din),
    .if_full_n(fifo_A_PE_4_4__full_n),
    .if_write(fifo_A_PE_4_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_4_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_4_5__dout),
    .if_empty_n(fifo_A_PE_4_5__empty_n),
    .if_read(fifo_A_PE_4_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_4_5__din),
    .if_full_n(fifo_A_PE_4_5__full_n),
    .if_write(fifo_A_PE_4_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_4_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_4_6__dout),
    .if_empty_n(fifo_A_PE_4_6__empty_n),
    .if_read(fifo_A_PE_4_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_4_6__din),
    .if_full_n(fifo_A_PE_4_6__full_n),
    .if_write(fifo_A_PE_4_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_4_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_4_7__dout),
    .if_empty_n(fifo_A_PE_4_7__empty_n),
    .if_read(fifo_A_PE_4_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_4_7__din),
    .if_full_n(fifo_A_PE_4_7__full_n),
    .if_write(fifo_A_PE_4_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_4_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_4_8__dout),
    .if_empty_n(fifo_A_PE_4_8__empty_n),
    .if_read(fifo_A_PE_4_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_4_8__din),
    .if_full_n(fifo_A_PE_4_8__full_n),
    .if_write(fifo_A_PE_4_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_4_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_4_9__dout),
    .if_empty_n(fifo_A_PE_4_9__empty_n),
    .if_read(fifo_A_PE_4_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_4_9__din),
    .if_full_n(fifo_A_PE_4_9__full_n),
    .if_write(fifo_A_PE_4_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_5_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_5_0__dout),
    .if_empty_n(fifo_A_PE_5_0__empty_n),
    .if_read(fifo_A_PE_5_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_5_0__din),
    .if_full_n(fifo_A_PE_5_0__full_n),
    .if_write(fifo_A_PE_5_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_5_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_5_1__dout),
    .if_empty_n(fifo_A_PE_5_1__empty_n),
    .if_read(fifo_A_PE_5_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_5_1__din),
    .if_full_n(fifo_A_PE_5_1__full_n),
    .if_write(fifo_A_PE_5_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_5_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_5_10__dout),
    .if_empty_n(fifo_A_PE_5_10__empty_n),
    .if_read(fifo_A_PE_5_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_5_10__din),
    .if_full_n(fifo_A_PE_5_10__full_n),
    .if_write(fifo_A_PE_5_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_5_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_5_11__dout),
    .if_empty_n(fifo_A_PE_5_11__empty_n),
    .if_read(fifo_A_PE_5_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_5_11__din),
    .if_full_n(fifo_A_PE_5_11__full_n),
    .if_write(fifo_A_PE_5_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_5_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_5_12__dout),
    .if_empty_n(fifo_A_PE_5_12__empty_n),
    .if_read(fifo_A_PE_5_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_5_12__din),
    .if_full_n(fifo_A_PE_5_12__full_n),
    .if_write(fifo_A_PE_5_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_5_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_5_13__dout),
    .if_empty_n(fifo_A_PE_5_13__empty_n),
    .if_read(fifo_A_PE_5_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_5_13__din),
    .if_full_n(fifo_A_PE_5_13__full_n),
    .if_write(fifo_A_PE_5_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_5_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_5_14__dout),
    .if_empty_n(fifo_A_PE_5_14__empty_n),
    .if_read(fifo_A_PE_5_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_5_14__din),
    .if_full_n(fifo_A_PE_5_14__full_n),
    .if_write(fifo_A_PE_5_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_5_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_5_15__dout),
    .if_empty_n(fifo_A_PE_5_15__empty_n),
    .if_read(fifo_A_PE_5_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_5_15__din),
    .if_full_n(fifo_A_PE_5_15__full_n),
    .if_write(fifo_A_PE_5_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_5_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_5_16__dout),
    .if_empty_n(fifo_A_PE_5_16__empty_n),
    .if_read(fifo_A_PE_5_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_5_16__din),
    .if_full_n(fifo_A_PE_5_16__full_n),
    .if_write(fifo_A_PE_5_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_5_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_5_17__dout),
    .if_empty_n(fifo_A_PE_5_17__empty_n),
    .if_read(fifo_A_PE_5_17__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_5_17__din),
    .if_full_n(fifo_A_PE_5_17__full_n),
    .if_write(fifo_A_PE_5_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_5_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_5_2__dout),
    .if_empty_n(fifo_A_PE_5_2__empty_n),
    .if_read(fifo_A_PE_5_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_5_2__din),
    .if_full_n(fifo_A_PE_5_2__full_n),
    .if_write(fifo_A_PE_5_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_5_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_5_3__dout),
    .if_empty_n(fifo_A_PE_5_3__empty_n),
    .if_read(fifo_A_PE_5_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_5_3__din),
    .if_full_n(fifo_A_PE_5_3__full_n),
    .if_write(fifo_A_PE_5_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_5_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_5_4__dout),
    .if_empty_n(fifo_A_PE_5_4__empty_n),
    .if_read(fifo_A_PE_5_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_5_4__din),
    .if_full_n(fifo_A_PE_5_4__full_n),
    .if_write(fifo_A_PE_5_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_5_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_5_5__dout),
    .if_empty_n(fifo_A_PE_5_5__empty_n),
    .if_read(fifo_A_PE_5_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_5_5__din),
    .if_full_n(fifo_A_PE_5_5__full_n),
    .if_write(fifo_A_PE_5_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_5_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_5_6__dout),
    .if_empty_n(fifo_A_PE_5_6__empty_n),
    .if_read(fifo_A_PE_5_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_5_6__din),
    .if_full_n(fifo_A_PE_5_6__full_n),
    .if_write(fifo_A_PE_5_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_5_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_5_7__dout),
    .if_empty_n(fifo_A_PE_5_7__empty_n),
    .if_read(fifo_A_PE_5_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_5_7__din),
    .if_full_n(fifo_A_PE_5_7__full_n),
    .if_write(fifo_A_PE_5_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_5_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_5_8__dout),
    .if_empty_n(fifo_A_PE_5_8__empty_n),
    .if_read(fifo_A_PE_5_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_5_8__din),
    .if_full_n(fifo_A_PE_5_8__full_n),
    .if_write(fifo_A_PE_5_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_5_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_5_9__dout),
    .if_empty_n(fifo_A_PE_5_9__empty_n),
    .if_read(fifo_A_PE_5_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_5_9__din),
    .if_full_n(fifo_A_PE_5_9__full_n),
    .if_write(fifo_A_PE_5_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_6_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_6_0__dout),
    .if_empty_n(fifo_A_PE_6_0__empty_n),
    .if_read(fifo_A_PE_6_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_6_0__din),
    .if_full_n(fifo_A_PE_6_0__full_n),
    .if_write(fifo_A_PE_6_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_6_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_6_1__dout),
    .if_empty_n(fifo_A_PE_6_1__empty_n),
    .if_read(fifo_A_PE_6_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_6_1__din),
    .if_full_n(fifo_A_PE_6_1__full_n),
    .if_write(fifo_A_PE_6_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_6_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_6_10__dout),
    .if_empty_n(fifo_A_PE_6_10__empty_n),
    .if_read(fifo_A_PE_6_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_6_10__din),
    .if_full_n(fifo_A_PE_6_10__full_n),
    .if_write(fifo_A_PE_6_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_6_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_6_11__dout),
    .if_empty_n(fifo_A_PE_6_11__empty_n),
    .if_read(fifo_A_PE_6_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_6_11__din),
    .if_full_n(fifo_A_PE_6_11__full_n),
    .if_write(fifo_A_PE_6_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_6_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_6_12__dout),
    .if_empty_n(fifo_A_PE_6_12__empty_n),
    .if_read(fifo_A_PE_6_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_6_12__din),
    .if_full_n(fifo_A_PE_6_12__full_n),
    .if_write(fifo_A_PE_6_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_6_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_6_13__dout),
    .if_empty_n(fifo_A_PE_6_13__empty_n),
    .if_read(fifo_A_PE_6_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_6_13__din),
    .if_full_n(fifo_A_PE_6_13__full_n),
    .if_write(fifo_A_PE_6_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_6_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_6_14__dout),
    .if_empty_n(fifo_A_PE_6_14__empty_n),
    .if_read(fifo_A_PE_6_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_6_14__din),
    .if_full_n(fifo_A_PE_6_14__full_n),
    .if_write(fifo_A_PE_6_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_6_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_6_15__dout),
    .if_empty_n(fifo_A_PE_6_15__empty_n),
    .if_read(fifo_A_PE_6_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_6_15__din),
    .if_full_n(fifo_A_PE_6_15__full_n),
    .if_write(fifo_A_PE_6_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_6_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_6_16__dout),
    .if_empty_n(fifo_A_PE_6_16__empty_n),
    .if_read(fifo_A_PE_6_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_6_16__din),
    .if_full_n(fifo_A_PE_6_16__full_n),
    .if_write(fifo_A_PE_6_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_6_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_6_17__dout),
    .if_empty_n(fifo_A_PE_6_17__empty_n),
    .if_read(fifo_A_PE_6_17__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_6_17__din),
    .if_full_n(fifo_A_PE_6_17__full_n),
    .if_write(fifo_A_PE_6_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_6_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_6_2__dout),
    .if_empty_n(fifo_A_PE_6_2__empty_n),
    .if_read(fifo_A_PE_6_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_6_2__din),
    .if_full_n(fifo_A_PE_6_2__full_n),
    .if_write(fifo_A_PE_6_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_6_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_6_3__dout),
    .if_empty_n(fifo_A_PE_6_3__empty_n),
    .if_read(fifo_A_PE_6_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_6_3__din),
    .if_full_n(fifo_A_PE_6_3__full_n),
    .if_write(fifo_A_PE_6_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_6_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_6_4__dout),
    .if_empty_n(fifo_A_PE_6_4__empty_n),
    .if_read(fifo_A_PE_6_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_6_4__din),
    .if_full_n(fifo_A_PE_6_4__full_n),
    .if_write(fifo_A_PE_6_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_6_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_6_5__dout),
    .if_empty_n(fifo_A_PE_6_5__empty_n),
    .if_read(fifo_A_PE_6_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_6_5__din),
    .if_full_n(fifo_A_PE_6_5__full_n),
    .if_write(fifo_A_PE_6_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_6_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_6_6__dout),
    .if_empty_n(fifo_A_PE_6_6__empty_n),
    .if_read(fifo_A_PE_6_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_6_6__din),
    .if_full_n(fifo_A_PE_6_6__full_n),
    .if_write(fifo_A_PE_6_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_6_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_6_7__dout),
    .if_empty_n(fifo_A_PE_6_7__empty_n),
    .if_read(fifo_A_PE_6_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_6_7__din),
    .if_full_n(fifo_A_PE_6_7__full_n),
    .if_write(fifo_A_PE_6_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_6_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_6_8__dout),
    .if_empty_n(fifo_A_PE_6_8__empty_n),
    .if_read(fifo_A_PE_6_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_6_8__din),
    .if_full_n(fifo_A_PE_6_8__full_n),
    .if_write(fifo_A_PE_6_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_6_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_6_9__dout),
    .if_empty_n(fifo_A_PE_6_9__empty_n),
    .if_read(fifo_A_PE_6_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_6_9__din),
    .if_full_n(fifo_A_PE_6_9__full_n),
    .if_write(fifo_A_PE_6_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_7_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_7_0__dout),
    .if_empty_n(fifo_A_PE_7_0__empty_n),
    .if_read(fifo_A_PE_7_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_7_0__din),
    .if_full_n(fifo_A_PE_7_0__full_n),
    .if_write(fifo_A_PE_7_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_7_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_7_1__dout),
    .if_empty_n(fifo_A_PE_7_1__empty_n),
    .if_read(fifo_A_PE_7_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_7_1__din),
    .if_full_n(fifo_A_PE_7_1__full_n),
    .if_write(fifo_A_PE_7_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_7_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_7_10__dout),
    .if_empty_n(fifo_A_PE_7_10__empty_n),
    .if_read(fifo_A_PE_7_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_7_10__din),
    .if_full_n(fifo_A_PE_7_10__full_n),
    .if_write(fifo_A_PE_7_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_7_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_7_11__dout),
    .if_empty_n(fifo_A_PE_7_11__empty_n),
    .if_read(fifo_A_PE_7_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_7_11__din),
    .if_full_n(fifo_A_PE_7_11__full_n),
    .if_write(fifo_A_PE_7_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_7_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_7_12__dout),
    .if_empty_n(fifo_A_PE_7_12__empty_n),
    .if_read(fifo_A_PE_7_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_7_12__din),
    .if_full_n(fifo_A_PE_7_12__full_n),
    .if_write(fifo_A_PE_7_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_7_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_7_13__dout),
    .if_empty_n(fifo_A_PE_7_13__empty_n),
    .if_read(fifo_A_PE_7_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_7_13__din),
    .if_full_n(fifo_A_PE_7_13__full_n),
    .if_write(fifo_A_PE_7_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_7_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_7_14__dout),
    .if_empty_n(fifo_A_PE_7_14__empty_n),
    .if_read(fifo_A_PE_7_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_7_14__din),
    .if_full_n(fifo_A_PE_7_14__full_n),
    .if_write(fifo_A_PE_7_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_7_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_7_15__dout),
    .if_empty_n(fifo_A_PE_7_15__empty_n),
    .if_read(fifo_A_PE_7_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_7_15__din),
    .if_full_n(fifo_A_PE_7_15__full_n),
    .if_write(fifo_A_PE_7_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_7_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_7_16__dout),
    .if_empty_n(fifo_A_PE_7_16__empty_n),
    .if_read(fifo_A_PE_7_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_7_16__din),
    .if_full_n(fifo_A_PE_7_16__full_n),
    .if_write(fifo_A_PE_7_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_7_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_7_17__dout),
    .if_empty_n(fifo_A_PE_7_17__empty_n),
    .if_read(fifo_A_PE_7_17__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_7_17__din),
    .if_full_n(fifo_A_PE_7_17__full_n),
    .if_write(fifo_A_PE_7_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_7_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_7_2__dout),
    .if_empty_n(fifo_A_PE_7_2__empty_n),
    .if_read(fifo_A_PE_7_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_7_2__din),
    .if_full_n(fifo_A_PE_7_2__full_n),
    .if_write(fifo_A_PE_7_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_7_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_7_3__dout),
    .if_empty_n(fifo_A_PE_7_3__empty_n),
    .if_read(fifo_A_PE_7_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_7_3__din),
    .if_full_n(fifo_A_PE_7_3__full_n),
    .if_write(fifo_A_PE_7_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_7_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_7_4__dout),
    .if_empty_n(fifo_A_PE_7_4__empty_n),
    .if_read(fifo_A_PE_7_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_7_4__din),
    .if_full_n(fifo_A_PE_7_4__full_n),
    .if_write(fifo_A_PE_7_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_7_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_7_5__dout),
    .if_empty_n(fifo_A_PE_7_5__empty_n),
    .if_read(fifo_A_PE_7_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_7_5__din),
    .if_full_n(fifo_A_PE_7_5__full_n),
    .if_write(fifo_A_PE_7_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_7_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_7_6__dout),
    .if_empty_n(fifo_A_PE_7_6__empty_n),
    .if_read(fifo_A_PE_7_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_7_6__din),
    .if_full_n(fifo_A_PE_7_6__full_n),
    .if_write(fifo_A_PE_7_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_7_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_7_7__dout),
    .if_empty_n(fifo_A_PE_7_7__empty_n),
    .if_read(fifo_A_PE_7_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_7_7__din),
    .if_full_n(fifo_A_PE_7_7__full_n),
    .if_write(fifo_A_PE_7_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_7_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_7_8__dout),
    .if_empty_n(fifo_A_PE_7_8__empty_n),
    .if_read(fifo_A_PE_7_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_7_8__din),
    .if_full_n(fifo_A_PE_7_8__full_n),
    .if_write(fifo_A_PE_7_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_7_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_7_9__dout),
    .if_empty_n(fifo_A_PE_7_9__empty_n),
    .if_read(fifo_A_PE_7_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_7_9__din),
    .if_full_n(fifo_A_PE_7_9__full_n),
    .if_write(fifo_A_PE_7_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_8_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_8_0__dout),
    .if_empty_n(fifo_A_PE_8_0__empty_n),
    .if_read(fifo_A_PE_8_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_8_0__din),
    .if_full_n(fifo_A_PE_8_0__full_n),
    .if_write(fifo_A_PE_8_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_8_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_8_1__dout),
    .if_empty_n(fifo_A_PE_8_1__empty_n),
    .if_read(fifo_A_PE_8_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_8_1__din),
    .if_full_n(fifo_A_PE_8_1__full_n),
    .if_write(fifo_A_PE_8_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_8_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_8_10__dout),
    .if_empty_n(fifo_A_PE_8_10__empty_n),
    .if_read(fifo_A_PE_8_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_8_10__din),
    .if_full_n(fifo_A_PE_8_10__full_n),
    .if_write(fifo_A_PE_8_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_8_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_8_11__dout),
    .if_empty_n(fifo_A_PE_8_11__empty_n),
    .if_read(fifo_A_PE_8_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_8_11__din),
    .if_full_n(fifo_A_PE_8_11__full_n),
    .if_write(fifo_A_PE_8_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_8_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_8_12__dout),
    .if_empty_n(fifo_A_PE_8_12__empty_n),
    .if_read(fifo_A_PE_8_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_8_12__din),
    .if_full_n(fifo_A_PE_8_12__full_n),
    .if_write(fifo_A_PE_8_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_8_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_8_13__dout),
    .if_empty_n(fifo_A_PE_8_13__empty_n),
    .if_read(fifo_A_PE_8_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_8_13__din),
    .if_full_n(fifo_A_PE_8_13__full_n),
    .if_write(fifo_A_PE_8_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_8_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_8_14__dout),
    .if_empty_n(fifo_A_PE_8_14__empty_n),
    .if_read(fifo_A_PE_8_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_8_14__din),
    .if_full_n(fifo_A_PE_8_14__full_n),
    .if_write(fifo_A_PE_8_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_8_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_8_15__dout),
    .if_empty_n(fifo_A_PE_8_15__empty_n),
    .if_read(fifo_A_PE_8_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_8_15__din),
    .if_full_n(fifo_A_PE_8_15__full_n),
    .if_write(fifo_A_PE_8_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_8_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_8_16__dout),
    .if_empty_n(fifo_A_PE_8_16__empty_n),
    .if_read(fifo_A_PE_8_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_8_16__din),
    .if_full_n(fifo_A_PE_8_16__full_n),
    .if_write(fifo_A_PE_8_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_8_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_8_17__dout),
    .if_empty_n(fifo_A_PE_8_17__empty_n),
    .if_read(fifo_A_PE_8_17__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_8_17__din),
    .if_full_n(fifo_A_PE_8_17__full_n),
    .if_write(fifo_A_PE_8_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_8_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_8_2__dout),
    .if_empty_n(fifo_A_PE_8_2__empty_n),
    .if_read(fifo_A_PE_8_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_8_2__din),
    .if_full_n(fifo_A_PE_8_2__full_n),
    .if_write(fifo_A_PE_8_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_8_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_8_3__dout),
    .if_empty_n(fifo_A_PE_8_3__empty_n),
    .if_read(fifo_A_PE_8_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_8_3__din),
    .if_full_n(fifo_A_PE_8_3__full_n),
    .if_write(fifo_A_PE_8_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_8_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_8_4__dout),
    .if_empty_n(fifo_A_PE_8_4__empty_n),
    .if_read(fifo_A_PE_8_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_8_4__din),
    .if_full_n(fifo_A_PE_8_4__full_n),
    .if_write(fifo_A_PE_8_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_8_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_8_5__dout),
    .if_empty_n(fifo_A_PE_8_5__empty_n),
    .if_read(fifo_A_PE_8_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_8_5__din),
    .if_full_n(fifo_A_PE_8_5__full_n),
    .if_write(fifo_A_PE_8_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_8_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_8_6__dout),
    .if_empty_n(fifo_A_PE_8_6__empty_n),
    .if_read(fifo_A_PE_8_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_8_6__din),
    .if_full_n(fifo_A_PE_8_6__full_n),
    .if_write(fifo_A_PE_8_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_8_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_8_7__dout),
    .if_empty_n(fifo_A_PE_8_7__empty_n),
    .if_read(fifo_A_PE_8_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_8_7__din),
    .if_full_n(fifo_A_PE_8_7__full_n),
    .if_write(fifo_A_PE_8_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_8_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_8_8__dout),
    .if_empty_n(fifo_A_PE_8_8__empty_n),
    .if_read(fifo_A_PE_8_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_8_8__din),
    .if_full_n(fifo_A_PE_8_8__full_n),
    .if_write(fifo_A_PE_8_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_8_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_8_9__dout),
    .if_empty_n(fifo_A_PE_8_9__empty_n),
    .if_read(fifo_A_PE_8_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_8_9__din),
    .if_full_n(fifo_A_PE_8_9__full_n),
    .if_write(fifo_A_PE_8_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_9_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_9_0__dout),
    .if_empty_n(fifo_A_PE_9_0__empty_n),
    .if_read(fifo_A_PE_9_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_9_0__din),
    .if_full_n(fifo_A_PE_9_0__full_n),
    .if_write(fifo_A_PE_9_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_9_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_9_1__dout),
    .if_empty_n(fifo_A_PE_9_1__empty_n),
    .if_read(fifo_A_PE_9_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_9_1__din),
    .if_full_n(fifo_A_PE_9_1__full_n),
    .if_write(fifo_A_PE_9_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_9_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_9_10__dout),
    .if_empty_n(fifo_A_PE_9_10__empty_n),
    .if_read(fifo_A_PE_9_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_9_10__din),
    .if_full_n(fifo_A_PE_9_10__full_n),
    .if_write(fifo_A_PE_9_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_9_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_9_11__dout),
    .if_empty_n(fifo_A_PE_9_11__empty_n),
    .if_read(fifo_A_PE_9_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_9_11__din),
    .if_full_n(fifo_A_PE_9_11__full_n),
    .if_write(fifo_A_PE_9_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_9_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_9_12__dout),
    .if_empty_n(fifo_A_PE_9_12__empty_n),
    .if_read(fifo_A_PE_9_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_9_12__din),
    .if_full_n(fifo_A_PE_9_12__full_n),
    .if_write(fifo_A_PE_9_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_9_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_9_13__dout),
    .if_empty_n(fifo_A_PE_9_13__empty_n),
    .if_read(fifo_A_PE_9_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_9_13__din),
    .if_full_n(fifo_A_PE_9_13__full_n),
    .if_write(fifo_A_PE_9_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_9_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_9_14__dout),
    .if_empty_n(fifo_A_PE_9_14__empty_n),
    .if_read(fifo_A_PE_9_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_9_14__din),
    .if_full_n(fifo_A_PE_9_14__full_n),
    .if_write(fifo_A_PE_9_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_9_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_9_15__dout),
    .if_empty_n(fifo_A_PE_9_15__empty_n),
    .if_read(fifo_A_PE_9_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_9_15__din),
    .if_full_n(fifo_A_PE_9_15__full_n),
    .if_write(fifo_A_PE_9_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_9_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_9_16__dout),
    .if_empty_n(fifo_A_PE_9_16__empty_n),
    .if_read(fifo_A_PE_9_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_9_16__din),
    .if_full_n(fifo_A_PE_9_16__full_n),
    .if_write(fifo_A_PE_9_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_9_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_9_17__dout),
    .if_empty_n(fifo_A_PE_9_17__empty_n),
    .if_read(fifo_A_PE_9_17__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_9_17__din),
    .if_full_n(fifo_A_PE_9_17__full_n),
    .if_write(fifo_A_PE_9_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_9_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_9_2__dout),
    .if_empty_n(fifo_A_PE_9_2__empty_n),
    .if_read(fifo_A_PE_9_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_9_2__din),
    .if_full_n(fifo_A_PE_9_2__full_n),
    .if_write(fifo_A_PE_9_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_9_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_9_3__dout),
    .if_empty_n(fifo_A_PE_9_3__empty_n),
    .if_read(fifo_A_PE_9_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_9_3__din),
    .if_full_n(fifo_A_PE_9_3__full_n),
    .if_write(fifo_A_PE_9_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_9_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_9_4__dout),
    .if_empty_n(fifo_A_PE_9_4__empty_n),
    .if_read(fifo_A_PE_9_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_9_4__din),
    .if_full_n(fifo_A_PE_9_4__full_n),
    .if_write(fifo_A_PE_9_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_9_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_9_5__dout),
    .if_empty_n(fifo_A_PE_9_5__empty_n),
    .if_read(fifo_A_PE_9_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_9_5__din),
    .if_full_n(fifo_A_PE_9_5__full_n),
    .if_write(fifo_A_PE_9_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_9_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_9_6__dout),
    .if_empty_n(fifo_A_PE_9_6__empty_n),
    .if_read(fifo_A_PE_9_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_9_6__din),
    .if_full_n(fifo_A_PE_9_6__full_n),
    .if_write(fifo_A_PE_9_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_9_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_9_7__dout),
    .if_empty_n(fifo_A_PE_9_7__empty_n),
    .if_read(fifo_A_PE_9_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_9_7__din),
    .if_full_n(fifo_A_PE_9_7__full_n),
    .if_write(fifo_A_PE_9_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_9_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_9_8__dout),
    .if_empty_n(fifo_A_PE_9_8__empty_n),
    .if_read(fifo_A_PE_9_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_9_8__din),
    .if_full_n(fifo_A_PE_9_8__full_n),
    .if_write(fifo_A_PE_9_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_A_PE_9_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_A_PE_9_9__dout),
    .if_empty_n(fifo_A_PE_9_9__empty_n),
    .if_read(fifo_A_PE_9_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_A_PE_9_9__din),
    .if_full_n(fifo_A_PE_9_9__full_n),
    .if_write(fifo_A_PE_9_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_B_IO_L2_in_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_B_IO_L2_in_0__dout),
    .if_empty_n(fifo_B_B_IO_L2_in_0__empty_n),
    .if_read(fifo_B_B_IO_L2_in_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_B_IO_L2_in_0__din),
    .if_full_n(fifo_B_B_IO_L2_in_0__full_n),
    .if_write(fifo_B_B_IO_L2_in_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_B_IO_L2_in_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_B_IO_L2_in_1__dout),
    .if_empty_n(fifo_B_B_IO_L2_in_1__empty_n),
    .if_read(fifo_B_B_IO_L2_in_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_B_IO_L2_in_1__din),
    .if_full_n(fifo_B_B_IO_L2_in_1__full_n),
    .if_write(fifo_B_B_IO_L2_in_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_B_IO_L2_in_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_B_IO_L2_in_10__dout),
    .if_empty_n(fifo_B_B_IO_L2_in_10__empty_n),
    .if_read(fifo_B_B_IO_L2_in_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_B_IO_L2_in_10__din),
    .if_full_n(fifo_B_B_IO_L2_in_10__full_n),
    .if_write(fifo_B_B_IO_L2_in_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_B_IO_L2_in_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_B_IO_L2_in_11__dout),
    .if_empty_n(fifo_B_B_IO_L2_in_11__empty_n),
    .if_read(fifo_B_B_IO_L2_in_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_B_IO_L2_in_11__din),
    .if_full_n(fifo_B_B_IO_L2_in_11__full_n),
    .if_write(fifo_B_B_IO_L2_in_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_B_IO_L2_in_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_B_IO_L2_in_12__dout),
    .if_empty_n(fifo_B_B_IO_L2_in_12__empty_n),
    .if_read(fifo_B_B_IO_L2_in_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_B_IO_L2_in_12__din),
    .if_full_n(fifo_B_B_IO_L2_in_12__full_n),
    .if_write(fifo_B_B_IO_L2_in_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_B_IO_L2_in_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_B_IO_L2_in_13__dout),
    .if_empty_n(fifo_B_B_IO_L2_in_13__empty_n),
    .if_read(fifo_B_B_IO_L2_in_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_B_IO_L2_in_13__din),
    .if_full_n(fifo_B_B_IO_L2_in_13__full_n),
    .if_write(fifo_B_B_IO_L2_in_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_B_IO_L2_in_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_B_IO_L2_in_14__dout),
    .if_empty_n(fifo_B_B_IO_L2_in_14__empty_n),
    .if_read(fifo_B_B_IO_L2_in_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_B_IO_L2_in_14__din),
    .if_full_n(fifo_B_B_IO_L2_in_14__full_n),
    .if_write(fifo_B_B_IO_L2_in_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_B_IO_L2_in_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_B_IO_L2_in_15__dout),
    .if_empty_n(fifo_B_B_IO_L2_in_15__empty_n),
    .if_read(fifo_B_B_IO_L2_in_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_B_IO_L2_in_15__din),
    .if_full_n(fifo_B_B_IO_L2_in_15__full_n),
    .if_write(fifo_B_B_IO_L2_in_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_B_IO_L2_in_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_B_IO_L2_in_16__dout),
    .if_empty_n(fifo_B_B_IO_L2_in_16__empty_n),
    .if_read(fifo_B_B_IO_L2_in_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_B_IO_L2_in_16__din),
    .if_full_n(fifo_B_B_IO_L2_in_16__full_n),
    .if_write(fifo_B_B_IO_L2_in_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_B_IO_L2_in_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_B_IO_L2_in_2__dout),
    .if_empty_n(fifo_B_B_IO_L2_in_2__empty_n),
    .if_read(fifo_B_B_IO_L2_in_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_B_IO_L2_in_2__din),
    .if_full_n(fifo_B_B_IO_L2_in_2__full_n),
    .if_write(fifo_B_B_IO_L2_in_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_B_IO_L2_in_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_B_IO_L2_in_3__dout),
    .if_empty_n(fifo_B_B_IO_L2_in_3__empty_n),
    .if_read(fifo_B_B_IO_L2_in_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_B_IO_L2_in_3__din),
    .if_full_n(fifo_B_B_IO_L2_in_3__full_n),
    .if_write(fifo_B_B_IO_L2_in_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_B_IO_L2_in_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_B_IO_L2_in_4__dout),
    .if_empty_n(fifo_B_B_IO_L2_in_4__empty_n),
    .if_read(fifo_B_B_IO_L2_in_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_B_IO_L2_in_4__din),
    .if_full_n(fifo_B_B_IO_L2_in_4__full_n),
    .if_write(fifo_B_B_IO_L2_in_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_B_IO_L2_in_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_B_IO_L2_in_5__dout),
    .if_empty_n(fifo_B_B_IO_L2_in_5__empty_n),
    .if_read(fifo_B_B_IO_L2_in_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_B_IO_L2_in_5__din),
    .if_full_n(fifo_B_B_IO_L2_in_5__full_n),
    .if_write(fifo_B_B_IO_L2_in_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_B_IO_L2_in_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_B_IO_L2_in_6__dout),
    .if_empty_n(fifo_B_B_IO_L2_in_6__empty_n),
    .if_read(fifo_B_B_IO_L2_in_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_B_IO_L2_in_6__din),
    .if_full_n(fifo_B_B_IO_L2_in_6__full_n),
    .if_write(fifo_B_B_IO_L2_in_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_B_IO_L2_in_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_B_IO_L2_in_7__dout),
    .if_empty_n(fifo_B_B_IO_L2_in_7__empty_n),
    .if_read(fifo_B_B_IO_L2_in_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_B_IO_L2_in_7__din),
    .if_full_n(fifo_B_B_IO_L2_in_7__full_n),
    .if_write(fifo_B_B_IO_L2_in_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_B_IO_L2_in_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_B_IO_L2_in_8__dout),
    .if_empty_n(fifo_B_B_IO_L2_in_8__empty_n),
    .if_read(fifo_B_B_IO_L2_in_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_B_IO_L2_in_8__din),
    .if_full_n(fifo_B_B_IO_L2_in_8__full_n),
    .if_write(fifo_B_B_IO_L2_in_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_B_IO_L2_in_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_B_IO_L2_in_9__dout),
    .if_empty_n(fifo_B_B_IO_L2_in_9__empty_n),
    .if_read(fifo_B_B_IO_L2_in_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_B_IO_L2_in_9__din),
    .if_full_n(fifo_B_B_IO_L2_in_9__full_n),
    .if_write(fifo_B_B_IO_L2_in_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_B_IO_L3_in_serialize
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_B_IO_L3_in_serialize__dout),
    .if_empty_n(fifo_B_B_IO_L3_in_serialize__empty_n),
    .if_read(fifo_B_B_IO_L3_in_serialize__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_B_IO_L3_in_serialize__din),
    .if_full_n(fifo_B_B_IO_L3_in_serialize__full_n),
    .if_write(fifo_B_B_IO_L3_in_serialize__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_0_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_0_0__dout),
    .if_empty_n(fifo_B_PE_0_0__empty_n),
    .if_read(fifo_B_PE_0_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_0_0__din),
    .if_full_n(fifo_B_PE_0_0__full_n),
    .if_write(fifo_B_PE_0_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_0_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_0_1__dout),
    .if_empty_n(fifo_B_PE_0_1__empty_n),
    .if_read(fifo_B_PE_0_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_0_1__din),
    .if_full_n(fifo_B_PE_0_1__full_n),
    .if_write(fifo_B_PE_0_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_0_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_0_10__dout),
    .if_empty_n(fifo_B_PE_0_10__empty_n),
    .if_read(fifo_B_PE_0_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_0_10__din),
    .if_full_n(fifo_B_PE_0_10__full_n),
    .if_write(fifo_B_PE_0_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_0_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_0_11__dout),
    .if_empty_n(fifo_B_PE_0_11__empty_n),
    .if_read(fifo_B_PE_0_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_0_11__din),
    .if_full_n(fifo_B_PE_0_11__full_n),
    .if_write(fifo_B_PE_0_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_0_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_0_12__dout),
    .if_empty_n(fifo_B_PE_0_12__empty_n),
    .if_read(fifo_B_PE_0_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_0_12__din),
    .if_full_n(fifo_B_PE_0_12__full_n),
    .if_write(fifo_B_PE_0_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_0_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_0_13__dout),
    .if_empty_n(fifo_B_PE_0_13__empty_n),
    .if_read(fifo_B_PE_0_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_0_13__din),
    .if_full_n(fifo_B_PE_0_13__full_n),
    .if_write(fifo_B_PE_0_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_0_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_0_14__dout),
    .if_empty_n(fifo_B_PE_0_14__empty_n),
    .if_read(fifo_B_PE_0_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_0_14__din),
    .if_full_n(fifo_B_PE_0_14__full_n),
    .if_write(fifo_B_PE_0_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_0_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_0_15__dout),
    .if_empty_n(fifo_B_PE_0_15__empty_n),
    .if_read(fifo_B_PE_0_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_0_15__din),
    .if_full_n(fifo_B_PE_0_15__full_n),
    .if_write(fifo_B_PE_0_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_0_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_0_16__dout),
    .if_empty_n(fifo_B_PE_0_16__empty_n),
    .if_read(fifo_B_PE_0_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_0_16__din),
    .if_full_n(fifo_B_PE_0_16__full_n),
    .if_write(fifo_B_PE_0_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_0_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_0_2__dout),
    .if_empty_n(fifo_B_PE_0_2__empty_n),
    .if_read(fifo_B_PE_0_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_0_2__din),
    .if_full_n(fifo_B_PE_0_2__full_n),
    .if_write(fifo_B_PE_0_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_0_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_0_3__dout),
    .if_empty_n(fifo_B_PE_0_3__empty_n),
    .if_read(fifo_B_PE_0_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_0_3__din),
    .if_full_n(fifo_B_PE_0_3__full_n),
    .if_write(fifo_B_PE_0_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_0_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_0_4__dout),
    .if_empty_n(fifo_B_PE_0_4__empty_n),
    .if_read(fifo_B_PE_0_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_0_4__din),
    .if_full_n(fifo_B_PE_0_4__full_n),
    .if_write(fifo_B_PE_0_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_0_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_0_5__dout),
    .if_empty_n(fifo_B_PE_0_5__empty_n),
    .if_read(fifo_B_PE_0_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_0_5__din),
    .if_full_n(fifo_B_PE_0_5__full_n),
    .if_write(fifo_B_PE_0_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_0_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_0_6__dout),
    .if_empty_n(fifo_B_PE_0_6__empty_n),
    .if_read(fifo_B_PE_0_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_0_6__din),
    .if_full_n(fifo_B_PE_0_6__full_n),
    .if_write(fifo_B_PE_0_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_0_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_0_7__dout),
    .if_empty_n(fifo_B_PE_0_7__empty_n),
    .if_read(fifo_B_PE_0_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_0_7__din),
    .if_full_n(fifo_B_PE_0_7__full_n),
    .if_write(fifo_B_PE_0_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_0_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_0_8__dout),
    .if_empty_n(fifo_B_PE_0_8__empty_n),
    .if_read(fifo_B_PE_0_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_0_8__din),
    .if_full_n(fifo_B_PE_0_8__full_n),
    .if_write(fifo_B_PE_0_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_0_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_0_9__dout),
    .if_empty_n(fifo_B_PE_0_9__empty_n),
    .if_read(fifo_B_PE_0_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_0_9__din),
    .if_full_n(fifo_B_PE_0_9__full_n),
    .if_write(fifo_B_PE_0_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_10_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_10_0__dout),
    .if_empty_n(fifo_B_PE_10_0__empty_n),
    .if_read(fifo_B_PE_10_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_10_0__din),
    .if_full_n(fifo_B_PE_10_0__full_n),
    .if_write(fifo_B_PE_10_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_10_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_10_1__dout),
    .if_empty_n(fifo_B_PE_10_1__empty_n),
    .if_read(fifo_B_PE_10_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_10_1__din),
    .if_full_n(fifo_B_PE_10_1__full_n),
    .if_write(fifo_B_PE_10_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_10_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_10_10__dout),
    .if_empty_n(fifo_B_PE_10_10__empty_n),
    .if_read(fifo_B_PE_10_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_10_10__din),
    .if_full_n(fifo_B_PE_10_10__full_n),
    .if_write(fifo_B_PE_10_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_10_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_10_11__dout),
    .if_empty_n(fifo_B_PE_10_11__empty_n),
    .if_read(fifo_B_PE_10_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_10_11__din),
    .if_full_n(fifo_B_PE_10_11__full_n),
    .if_write(fifo_B_PE_10_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_10_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_10_12__dout),
    .if_empty_n(fifo_B_PE_10_12__empty_n),
    .if_read(fifo_B_PE_10_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_10_12__din),
    .if_full_n(fifo_B_PE_10_12__full_n),
    .if_write(fifo_B_PE_10_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_10_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_10_13__dout),
    .if_empty_n(fifo_B_PE_10_13__empty_n),
    .if_read(fifo_B_PE_10_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_10_13__din),
    .if_full_n(fifo_B_PE_10_13__full_n),
    .if_write(fifo_B_PE_10_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_10_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_10_14__dout),
    .if_empty_n(fifo_B_PE_10_14__empty_n),
    .if_read(fifo_B_PE_10_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_10_14__din),
    .if_full_n(fifo_B_PE_10_14__full_n),
    .if_write(fifo_B_PE_10_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_10_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_10_15__dout),
    .if_empty_n(fifo_B_PE_10_15__empty_n),
    .if_read(fifo_B_PE_10_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_10_15__din),
    .if_full_n(fifo_B_PE_10_15__full_n),
    .if_write(fifo_B_PE_10_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_10_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_10_16__dout),
    .if_empty_n(fifo_B_PE_10_16__empty_n),
    .if_read(fifo_B_PE_10_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_10_16__din),
    .if_full_n(fifo_B_PE_10_16__full_n),
    .if_write(fifo_B_PE_10_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_10_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_10_2__dout),
    .if_empty_n(fifo_B_PE_10_2__empty_n),
    .if_read(fifo_B_PE_10_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_10_2__din),
    .if_full_n(fifo_B_PE_10_2__full_n),
    .if_write(fifo_B_PE_10_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_10_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_10_3__dout),
    .if_empty_n(fifo_B_PE_10_3__empty_n),
    .if_read(fifo_B_PE_10_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_10_3__din),
    .if_full_n(fifo_B_PE_10_3__full_n),
    .if_write(fifo_B_PE_10_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_10_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_10_4__dout),
    .if_empty_n(fifo_B_PE_10_4__empty_n),
    .if_read(fifo_B_PE_10_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_10_4__din),
    .if_full_n(fifo_B_PE_10_4__full_n),
    .if_write(fifo_B_PE_10_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_10_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_10_5__dout),
    .if_empty_n(fifo_B_PE_10_5__empty_n),
    .if_read(fifo_B_PE_10_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_10_5__din),
    .if_full_n(fifo_B_PE_10_5__full_n),
    .if_write(fifo_B_PE_10_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_10_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_10_6__dout),
    .if_empty_n(fifo_B_PE_10_6__empty_n),
    .if_read(fifo_B_PE_10_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_10_6__din),
    .if_full_n(fifo_B_PE_10_6__full_n),
    .if_write(fifo_B_PE_10_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_10_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_10_7__dout),
    .if_empty_n(fifo_B_PE_10_7__empty_n),
    .if_read(fifo_B_PE_10_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_10_7__din),
    .if_full_n(fifo_B_PE_10_7__full_n),
    .if_write(fifo_B_PE_10_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_10_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_10_8__dout),
    .if_empty_n(fifo_B_PE_10_8__empty_n),
    .if_read(fifo_B_PE_10_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_10_8__din),
    .if_full_n(fifo_B_PE_10_8__full_n),
    .if_write(fifo_B_PE_10_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_10_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_10_9__dout),
    .if_empty_n(fifo_B_PE_10_9__empty_n),
    .if_read(fifo_B_PE_10_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_10_9__din),
    .if_full_n(fifo_B_PE_10_9__full_n),
    .if_write(fifo_B_PE_10_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_11_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_11_0__dout),
    .if_empty_n(fifo_B_PE_11_0__empty_n),
    .if_read(fifo_B_PE_11_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_11_0__din),
    .if_full_n(fifo_B_PE_11_0__full_n),
    .if_write(fifo_B_PE_11_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_11_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_11_1__dout),
    .if_empty_n(fifo_B_PE_11_1__empty_n),
    .if_read(fifo_B_PE_11_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_11_1__din),
    .if_full_n(fifo_B_PE_11_1__full_n),
    .if_write(fifo_B_PE_11_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_11_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_11_10__dout),
    .if_empty_n(fifo_B_PE_11_10__empty_n),
    .if_read(fifo_B_PE_11_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_11_10__din),
    .if_full_n(fifo_B_PE_11_10__full_n),
    .if_write(fifo_B_PE_11_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_11_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_11_11__dout),
    .if_empty_n(fifo_B_PE_11_11__empty_n),
    .if_read(fifo_B_PE_11_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_11_11__din),
    .if_full_n(fifo_B_PE_11_11__full_n),
    .if_write(fifo_B_PE_11_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_11_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_11_12__dout),
    .if_empty_n(fifo_B_PE_11_12__empty_n),
    .if_read(fifo_B_PE_11_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_11_12__din),
    .if_full_n(fifo_B_PE_11_12__full_n),
    .if_write(fifo_B_PE_11_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_11_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_11_13__dout),
    .if_empty_n(fifo_B_PE_11_13__empty_n),
    .if_read(fifo_B_PE_11_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_11_13__din),
    .if_full_n(fifo_B_PE_11_13__full_n),
    .if_write(fifo_B_PE_11_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_11_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_11_14__dout),
    .if_empty_n(fifo_B_PE_11_14__empty_n),
    .if_read(fifo_B_PE_11_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_11_14__din),
    .if_full_n(fifo_B_PE_11_14__full_n),
    .if_write(fifo_B_PE_11_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_11_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_11_15__dout),
    .if_empty_n(fifo_B_PE_11_15__empty_n),
    .if_read(fifo_B_PE_11_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_11_15__din),
    .if_full_n(fifo_B_PE_11_15__full_n),
    .if_write(fifo_B_PE_11_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_11_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_11_16__dout),
    .if_empty_n(fifo_B_PE_11_16__empty_n),
    .if_read(fifo_B_PE_11_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_11_16__din),
    .if_full_n(fifo_B_PE_11_16__full_n),
    .if_write(fifo_B_PE_11_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_11_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_11_2__dout),
    .if_empty_n(fifo_B_PE_11_2__empty_n),
    .if_read(fifo_B_PE_11_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_11_2__din),
    .if_full_n(fifo_B_PE_11_2__full_n),
    .if_write(fifo_B_PE_11_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_11_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_11_3__dout),
    .if_empty_n(fifo_B_PE_11_3__empty_n),
    .if_read(fifo_B_PE_11_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_11_3__din),
    .if_full_n(fifo_B_PE_11_3__full_n),
    .if_write(fifo_B_PE_11_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_11_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_11_4__dout),
    .if_empty_n(fifo_B_PE_11_4__empty_n),
    .if_read(fifo_B_PE_11_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_11_4__din),
    .if_full_n(fifo_B_PE_11_4__full_n),
    .if_write(fifo_B_PE_11_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_11_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_11_5__dout),
    .if_empty_n(fifo_B_PE_11_5__empty_n),
    .if_read(fifo_B_PE_11_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_11_5__din),
    .if_full_n(fifo_B_PE_11_5__full_n),
    .if_write(fifo_B_PE_11_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_11_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_11_6__dout),
    .if_empty_n(fifo_B_PE_11_6__empty_n),
    .if_read(fifo_B_PE_11_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_11_6__din),
    .if_full_n(fifo_B_PE_11_6__full_n),
    .if_write(fifo_B_PE_11_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_11_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_11_7__dout),
    .if_empty_n(fifo_B_PE_11_7__empty_n),
    .if_read(fifo_B_PE_11_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_11_7__din),
    .if_full_n(fifo_B_PE_11_7__full_n),
    .if_write(fifo_B_PE_11_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_11_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_11_8__dout),
    .if_empty_n(fifo_B_PE_11_8__empty_n),
    .if_read(fifo_B_PE_11_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_11_8__din),
    .if_full_n(fifo_B_PE_11_8__full_n),
    .if_write(fifo_B_PE_11_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_11_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_11_9__dout),
    .if_empty_n(fifo_B_PE_11_9__empty_n),
    .if_read(fifo_B_PE_11_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_11_9__din),
    .if_full_n(fifo_B_PE_11_9__full_n),
    .if_write(fifo_B_PE_11_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_12_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_12_0__dout),
    .if_empty_n(fifo_B_PE_12_0__empty_n),
    .if_read(fifo_B_PE_12_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_12_0__din),
    .if_full_n(fifo_B_PE_12_0__full_n),
    .if_write(fifo_B_PE_12_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_12_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_12_1__dout),
    .if_empty_n(fifo_B_PE_12_1__empty_n),
    .if_read(fifo_B_PE_12_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_12_1__din),
    .if_full_n(fifo_B_PE_12_1__full_n),
    .if_write(fifo_B_PE_12_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_12_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_12_10__dout),
    .if_empty_n(fifo_B_PE_12_10__empty_n),
    .if_read(fifo_B_PE_12_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_12_10__din),
    .if_full_n(fifo_B_PE_12_10__full_n),
    .if_write(fifo_B_PE_12_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_12_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_12_11__dout),
    .if_empty_n(fifo_B_PE_12_11__empty_n),
    .if_read(fifo_B_PE_12_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_12_11__din),
    .if_full_n(fifo_B_PE_12_11__full_n),
    .if_write(fifo_B_PE_12_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_12_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_12_12__dout),
    .if_empty_n(fifo_B_PE_12_12__empty_n),
    .if_read(fifo_B_PE_12_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_12_12__din),
    .if_full_n(fifo_B_PE_12_12__full_n),
    .if_write(fifo_B_PE_12_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_12_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_12_13__dout),
    .if_empty_n(fifo_B_PE_12_13__empty_n),
    .if_read(fifo_B_PE_12_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_12_13__din),
    .if_full_n(fifo_B_PE_12_13__full_n),
    .if_write(fifo_B_PE_12_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_12_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_12_14__dout),
    .if_empty_n(fifo_B_PE_12_14__empty_n),
    .if_read(fifo_B_PE_12_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_12_14__din),
    .if_full_n(fifo_B_PE_12_14__full_n),
    .if_write(fifo_B_PE_12_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_12_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_12_15__dout),
    .if_empty_n(fifo_B_PE_12_15__empty_n),
    .if_read(fifo_B_PE_12_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_12_15__din),
    .if_full_n(fifo_B_PE_12_15__full_n),
    .if_write(fifo_B_PE_12_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_12_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_12_16__dout),
    .if_empty_n(fifo_B_PE_12_16__empty_n),
    .if_read(fifo_B_PE_12_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_12_16__din),
    .if_full_n(fifo_B_PE_12_16__full_n),
    .if_write(fifo_B_PE_12_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_12_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_12_2__dout),
    .if_empty_n(fifo_B_PE_12_2__empty_n),
    .if_read(fifo_B_PE_12_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_12_2__din),
    .if_full_n(fifo_B_PE_12_2__full_n),
    .if_write(fifo_B_PE_12_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_12_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_12_3__dout),
    .if_empty_n(fifo_B_PE_12_3__empty_n),
    .if_read(fifo_B_PE_12_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_12_3__din),
    .if_full_n(fifo_B_PE_12_3__full_n),
    .if_write(fifo_B_PE_12_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_12_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_12_4__dout),
    .if_empty_n(fifo_B_PE_12_4__empty_n),
    .if_read(fifo_B_PE_12_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_12_4__din),
    .if_full_n(fifo_B_PE_12_4__full_n),
    .if_write(fifo_B_PE_12_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_12_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_12_5__dout),
    .if_empty_n(fifo_B_PE_12_5__empty_n),
    .if_read(fifo_B_PE_12_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_12_5__din),
    .if_full_n(fifo_B_PE_12_5__full_n),
    .if_write(fifo_B_PE_12_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_12_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_12_6__dout),
    .if_empty_n(fifo_B_PE_12_6__empty_n),
    .if_read(fifo_B_PE_12_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_12_6__din),
    .if_full_n(fifo_B_PE_12_6__full_n),
    .if_write(fifo_B_PE_12_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_12_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_12_7__dout),
    .if_empty_n(fifo_B_PE_12_7__empty_n),
    .if_read(fifo_B_PE_12_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_12_7__din),
    .if_full_n(fifo_B_PE_12_7__full_n),
    .if_write(fifo_B_PE_12_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_12_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_12_8__dout),
    .if_empty_n(fifo_B_PE_12_8__empty_n),
    .if_read(fifo_B_PE_12_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_12_8__din),
    .if_full_n(fifo_B_PE_12_8__full_n),
    .if_write(fifo_B_PE_12_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_12_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_12_9__dout),
    .if_empty_n(fifo_B_PE_12_9__empty_n),
    .if_read(fifo_B_PE_12_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_12_9__din),
    .if_full_n(fifo_B_PE_12_9__full_n),
    .if_write(fifo_B_PE_12_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_13_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_13_0__dout),
    .if_empty_n(fifo_B_PE_13_0__empty_n),
    .if_read(fifo_B_PE_13_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_13_0__din),
    .if_full_n(fifo_B_PE_13_0__full_n),
    .if_write(fifo_B_PE_13_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_13_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_13_1__dout),
    .if_empty_n(fifo_B_PE_13_1__empty_n),
    .if_read(fifo_B_PE_13_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_13_1__din),
    .if_full_n(fifo_B_PE_13_1__full_n),
    .if_write(fifo_B_PE_13_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_13_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_13_10__dout),
    .if_empty_n(fifo_B_PE_13_10__empty_n),
    .if_read(fifo_B_PE_13_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_13_10__din),
    .if_full_n(fifo_B_PE_13_10__full_n),
    .if_write(fifo_B_PE_13_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_13_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_13_11__dout),
    .if_empty_n(fifo_B_PE_13_11__empty_n),
    .if_read(fifo_B_PE_13_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_13_11__din),
    .if_full_n(fifo_B_PE_13_11__full_n),
    .if_write(fifo_B_PE_13_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_13_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_13_12__dout),
    .if_empty_n(fifo_B_PE_13_12__empty_n),
    .if_read(fifo_B_PE_13_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_13_12__din),
    .if_full_n(fifo_B_PE_13_12__full_n),
    .if_write(fifo_B_PE_13_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_13_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_13_13__dout),
    .if_empty_n(fifo_B_PE_13_13__empty_n),
    .if_read(fifo_B_PE_13_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_13_13__din),
    .if_full_n(fifo_B_PE_13_13__full_n),
    .if_write(fifo_B_PE_13_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_13_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_13_14__dout),
    .if_empty_n(fifo_B_PE_13_14__empty_n),
    .if_read(fifo_B_PE_13_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_13_14__din),
    .if_full_n(fifo_B_PE_13_14__full_n),
    .if_write(fifo_B_PE_13_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_13_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_13_15__dout),
    .if_empty_n(fifo_B_PE_13_15__empty_n),
    .if_read(fifo_B_PE_13_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_13_15__din),
    .if_full_n(fifo_B_PE_13_15__full_n),
    .if_write(fifo_B_PE_13_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_13_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_13_16__dout),
    .if_empty_n(fifo_B_PE_13_16__empty_n),
    .if_read(fifo_B_PE_13_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_13_16__din),
    .if_full_n(fifo_B_PE_13_16__full_n),
    .if_write(fifo_B_PE_13_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_13_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_13_2__dout),
    .if_empty_n(fifo_B_PE_13_2__empty_n),
    .if_read(fifo_B_PE_13_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_13_2__din),
    .if_full_n(fifo_B_PE_13_2__full_n),
    .if_write(fifo_B_PE_13_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_13_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_13_3__dout),
    .if_empty_n(fifo_B_PE_13_3__empty_n),
    .if_read(fifo_B_PE_13_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_13_3__din),
    .if_full_n(fifo_B_PE_13_3__full_n),
    .if_write(fifo_B_PE_13_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_13_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_13_4__dout),
    .if_empty_n(fifo_B_PE_13_4__empty_n),
    .if_read(fifo_B_PE_13_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_13_4__din),
    .if_full_n(fifo_B_PE_13_4__full_n),
    .if_write(fifo_B_PE_13_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_13_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_13_5__dout),
    .if_empty_n(fifo_B_PE_13_5__empty_n),
    .if_read(fifo_B_PE_13_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_13_5__din),
    .if_full_n(fifo_B_PE_13_5__full_n),
    .if_write(fifo_B_PE_13_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_13_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_13_6__dout),
    .if_empty_n(fifo_B_PE_13_6__empty_n),
    .if_read(fifo_B_PE_13_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_13_6__din),
    .if_full_n(fifo_B_PE_13_6__full_n),
    .if_write(fifo_B_PE_13_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_13_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_13_7__dout),
    .if_empty_n(fifo_B_PE_13_7__empty_n),
    .if_read(fifo_B_PE_13_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_13_7__din),
    .if_full_n(fifo_B_PE_13_7__full_n),
    .if_write(fifo_B_PE_13_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_13_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_13_8__dout),
    .if_empty_n(fifo_B_PE_13_8__empty_n),
    .if_read(fifo_B_PE_13_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_13_8__din),
    .if_full_n(fifo_B_PE_13_8__full_n),
    .if_write(fifo_B_PE_13_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_13_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_13_9__dout),
    .if_empty_n(fifo_B_PE_13_9__empty_n),
    .if_read(fifo_B_PE_13_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_13_9__din),
    .if_full_n(fifo_B_PE_13_9__full_n),
    .if_write(fifo_B_PE_13_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_14_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_14_0__dout),
    .if_empty_n(fifo_B_PE_14_0__empty_n),
    .if_read(fifo_B_PE_14_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_14_0__din),
    .if_full_n(fifo_B_PE_14_0__full_n),
    .if_write(fifo_B_PE_14_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_14_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_14_1__dout),
    .if_empty_n(fifo_B_PE_14_1__empty_n),
    .if_read(fifo_B_PE_14_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_14_1__din),
    .if_full_n(fifo_B_PE_14_1__full_n),
    .if_write(fifo_B_PE_14_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_14_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_14_10__dout),
    .if_empty_n(fifo_B_PE_14_10__empty_n),
    .if_read(fifo_B_PE_14_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_14_10__din),
    .if_full_n(fifo_B_PE_14_10__full_n),
    .if_write(fifo_B_PE_14_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_14_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_14_11__dout),
    .if_empty_n(fifo_B_PE_14_11__empty_n),
    .if_read(fifo_B_PE_14_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_14_11__din),
    .if_full_n(fifo_B_PE_14_11__full_n),
    .if_write(fifo_B_PE_14_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_14_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_14_12__dout),
    .if_empty_n(fifo_B_PE_14_12__empty_n),
    .if_read(fifo_B_PE_14_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_14_12__din),
    .if_full_n(fifo_B_PE_14_12__full_n),
    .if_write(fifo_B_PE_14_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_14_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_14_13__dout),
    .if_empty_n(fifo_B_PE_14_13__empty_n),
    .if_read(fifo_B_PE_14_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_14_13__din),
    .if_full_n(fifo_B_PE_14_13__full_n),
    .if_write(fifo_B_PE_14_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_14_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_14_14__dout),
    .if_empty_n(fifo_B_PE_14_14__empty_n),
    .if_read(fifo_B_PE_14_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_14_14__din),
    .if_full_n(fifo_B_PE_14_14__full_n),
    .if_write(fifo_B_PE_14_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_14_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_14_15__dout),
    .if_empty_n(fifo_B_PE_14_15__empty_n),
    .if_read(fifo_B_PE_14_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_14_15__din),
    .if_full_n(fifo_B_PE_14_15__full_n),
    .if_write(fifo_B_PE_14_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_14_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_14_16__dout),
    .if_empty_n(fifo_B_PE_14_16__empty_n),
    .if_read(fifo_B_PE_14_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_14_16__din),
    .if_full_n(fifo_B_PE_14_16__full_n),
    .if_write(fifo_B_PE_14_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_14_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_14_2__dout),
    .if_empty_n(fifo_B_PE_14_2__empty_n),
    .if_read(fifo_B_PE_14_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_14_2__din),
    .if_full_n(fifo_B_PE_14_2__full_n),
    .if_write(fifo_B_PE_14_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_14_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_14_3__dout),
    .if_empty_n(fifo_B_PE_14_3__empty_n),
    .if_read(fifo_B_PE_14_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_14_3__din),
    .if_full_n(fifo_B_PE_14_3__full_n),
    .if_write(fifo_B_PE_14_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_14_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_14_4__dout),
    .if_empty_n(fifo_B_PE_14_4__empty_n),
    .if_read(fifo_B_PE_14_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_14_4__din),
    .if_full_n(fifo_B_PE_14_4__full_n),
    .if_write(fifo_B_PE_14_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_14_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_14_5__dout),
    .if_empty_n(fifo_B_PE_14_5__empty_n),
    .if_read(fifo_B_PE_14_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_14_5__din),
    .if_full_n(fifo_B_PE_14_5__full_n),
    .if_write(fifo_B_PE_14_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_14_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_14_6__dout),
    .if_empty_n(fifo_B_PE_14_6__empty_n),
    .if_read(fifo_B_PE_14_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_14_6__din),
    .if_full_n(fifo_B_PE_14_6__full_n),
    .if_write(fifo_B_PE_14_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_14_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_14_7__dout),
    .if_empty_n(fifo_B_PE_14_7__empty_n),
    .if_read(fifo_B_PE_14_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_14_7__din),
    .if_full_n(fifo_B_PE_14_7__full_n),
    .if_write(fifo_B_PE_14_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_14_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_14_8__dout),
    .if_empty_n(fifo_B_PE_14_8__empty_n),
    .if_read(fifo_B_PE_14_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_14_8__din),
    .if_full_n(fifo_B_PE_14_8__full_n),
    .if_write(fifo_B_PE_14_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_14_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_14_9__dout),
    .if_empty_n(fifo_B_PE_14_9__empty_n),
    .if_read(fifo_B_PE_14_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_14_9__din),
    .if_full_n(fifo_B_PE_14_9__full_n),
    .if_write(fifo_B_PE_14_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_15_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_15_0__dout),
    .if_empty_n(fifo_B_PE_15_0__empty_n),
    .if_read(fifo_B_PE_15_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_15_0__din),
    .if_full_n(fifo_B_PE_15_0__full_n),
    .if_write(fifo_B_PE_15_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_15_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_15_1__dout),
    .if_empty_n(fifo_B_PE_15_1__empty_n),
    .if_read(fifo_B_PE_15_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_15_1__din),
    .if_full_n(fifo_B_PE_15_1__full_n),
    .if_write(fifo_B_PE_15_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_15_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_15_10__dout),
    .if_empty_n(fifo_B_PE_15_10__empty_n),
    .if_read(fifo_B_PE_15_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_15_10__din),
    .if_full_n(fifo_B_PE_15_10__full_n),
    .if_write(fifo_B_PE_15_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_15_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_15_11__dout),
    .if_empty_n(fifo_B_PE_15_11__empty_n),
    .if_read(fifo_B_PE_15_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_15_11__din),
    .if_full_n(fifo_B_PE_15_11__full_n),
    .if_write(fifo_B_PE_15_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_15_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_15_12__dout),
    .if_empty_n(fifo_B_PE_15_12__empty_n),
    .if_read(fifo_B_PE_15_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_15_12__din),
    .if_full_n(fifo_B_PE_15_12__full_n),
    .if_write(fifo_B_PE_15_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_15_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_15_13__dout),
    .if_empty_n(fifo_B_PE_15_13__empty_n),
    .if_read(fifo_B_PE_15_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_15_13__din),
    .if_full_n(fifo_B_PE_15_13__full_n),
    .if_write(fifo_B_PE_15_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_15_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_15_14__dout),
    .if_empty_n(fifo_B_PE_15_14__empty_n),
    .if_read(fifo_B_PE_15_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_15_14__din),
    .if_full_n(fifo_B_PE_15_14__full_n),
    .if_write(fifo_B_PE_15_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_15_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_15_15__dout),
    .if_empty_n(fifo_B_PE_15_15__empty_n),
    .if_read(fifo_B_PE_15_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_15_15__din),
    .if_full_n(fifo_B_PE_15_15__full_n),
    .if_write(fifo_B_PE_15_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_15_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_15_16__dout),
    .if_empty_n(fifo_B_PE_15_16__empty_n),
    .if_read(fifo_B_PE_15_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_15_16__din),
    .if_full_n(fifo_B_PE_15_16__full_n),
    .if_write(fifo_B_PE_15_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_15_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_15_2__dout),
    .if_empty_n(fifo_B_PE_15_2__empty_n),
    .if_read(fifo_B_PE_15_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_15_2__din),
    .if_full_n(fifo_B_PE_15_2__full_n),
    .if_write(fifo_B_PE_15_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_15_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_15_3__dout),
    .if_empty_n(fifo_B_PE_15_3__empty_n),
    .if_read(fifo_B_PE_15_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_15_3__din),
    .if_full_n(fifo_B_PE_15_3__full_n),
    .if_write(fifo_B_PE_15_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_15_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_15_4__dout),
    .if_empty_n(fifo_B_PE_15_4__empty_n),
    .if_read(fifo_B_PE_15_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_15_4__din),
    .if_full_n(fifo_B_PE_15_4__full_n),
    .if_write(fifo_B_PE_15_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_15_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_15_5__dout),
    .if_empty_n(fifo_B_PE_15_5__empty_n),
    .if_read(fifo_B_PE_15_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_15_5__din),
    .if_full_n(fifo_B_PE_15_5__full_n),
    .if_write(fifo_B_PE_15_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_15_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_15_6__dout),
    .if_empty_n(fifo_B_PE_15_6__empty_n),
    .if_read(fifo_B_PE_15_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_15_6__din),
    .if_full_n(fifo_B_PE_15_6__full_n),
    .if_write(fifo_B_PE_15_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_15_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_15_7__dout),
    .if_empty_n(fifo_B_PE_15_7__empty_n),
    .if_read(fifo_B_PE_15_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_15_7__din),
    .if_full_n(fifo_B_PE_15_7__full_n),
    .if_write(fifo_B_PE_15_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_15_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_15_8__dout),
    .if_empty_n(fifo_B_PE_15_8__empty_n),
    .if_read(fifo_B_PE_15_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_15_8__din),
    .if_full_n(fifo_B_PE_15_8__full_n),
    .if_write(fifo_B_PE_15_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_15_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_15_9__dout),
    .if_empty_n(fifo_B_PE_15_9__empty_n),
    .if_read(fifo_B_PE_15_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_15_9__din),
    .if_full_n(fifo_B_PE_15_9__full_n),
    .if_write(fifo_B_PE_15_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_16_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_16_0__dout),
    .if_empty_n(fifo_B_PE_16_0__empty_n),
    .if_read(fifo_B_PE_16_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_16_0__din),
    .if_full_n(fifo_B_PE_16_0__full_n),
    .if_write(fifo_B_PE_16_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_16_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_16_1__dout),
    .if_empty_n(fifo_B_PE_16_1__empty_n),
    .if_read(fifo_B_PE_16_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_16_1__din),
    .if_full_n(fifo_B_PE_16_1__full_n),
    .if_write(fifo_B_PE_16_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_16_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_16_10__dout),
    .if_empty_n(fifo_B_PE_16_10__empty_n),
    .if_read(fifo_B_PE_16_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_16_10__din),
    .if_full_n(fifo_B_PE_16_10__full_n),
    .if_write(fifo_B_PE_16_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_16_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_16_11__dout),
    .if_empty_n(fifo_B_PE_16_11__empty_n),
    .if_read(fifo_B_PE_16_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_16_11__din),
    .if_full_n(fifo_B_PE_16_11__full_n),
    .if_write(fifo_B_PE_16_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_16_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_16_12__dout),
    .if_empty_n(fifo_B_PE_16_12__empty_n),
    .if_read(fifo_B_PE_16_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_16_12__din),
    .if_full_n(fifo_B_PE_16_12__full_n),
    .if_write(fifo_B_PE_16_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_16_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_16_13__dout),
    .if_empty_n(fifo_B_PE_16_13__empty_n),
    .if_read(fifo_B_PE_16_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_16_13__din),
    .if_full_n(fifo_B_PE_16_13__full_n),
    .if_write(fifo_B_PE_16_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_16_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_16_14__dout),
    .if_empty_n(fifo_B_PE_16_14__empty_n),
    .if_read(fifo_B_PE_16_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_16_14__din),
    .if_full_n(fifo_B_PE_16_14__full_n),
    .if_write(fifo_B_PE_16_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_16_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_16_15__dout),
    .if_empty_n(fifo_B_PE_16_15__empty_n),
    .if_read(fifo_B_PE_16_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_16_15__din),
    .if_full_n(fifo_B_PE_16_15__full_n),
    .if_write(fifo_B_PE_16_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_16_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_16_16__dout),
    .if_empty_n(fifo_B_PE_16_16__empty_n),
    .if_read(fifo_B_PE_16_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_16_16__din),
    .if_full_n(fifo_B_PE_16_16__full_n),
    .if_write(fifo_B_PE_16_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_16_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_16_2__dout),
    .if_empty_n(fifo_B_PE_16_2__empty_n),
    .if_read(fifo_B_PE_16_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_16_2__din),
    .if_full_n(fifo_B_PE_16_2__full_n),
    .if_write(fifo_B_PE_16_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_16_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_16_3__dout),
    .if_empty_n(fifo_B_PE_16_3__empty_n),
    .if_read(fifo_B_PE_16_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_16_3__din),
    .if_full_n(fifo_B_PE_16_3__full_n),
    .if_write(fifo_B_PE_16_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_16_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_16_4__dout),
    .if_empty_n(fifo_B_PE_16_4__empty_n),
    .if_read(fifo_B_PE_16_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_16_4__din),
    .if_full_n(fifo_B_PE_16_4__full_n),
    .if_write(fifo_B_PE_16_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_16_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_16_5__dout),
    .if_empty_n(fifo_B_PE_16_5__empty_n),
    .if_read(fifo_B_PE_16_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_16_5__din),
    .if_full_n(fifo_B_PE_16_5__full_n),
    .if_write(fifo_B_PE_16_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_16_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_16_6__dout),
    .if_empty_n(fifo_B_PE_16_6__empty_n),
    .if_read(fifo_B_PE_16_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_16_6__din),
    .if_full_n(fifo_B_PE_16_6__full_n),
    .if_write(fifo_B_PE_16_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_16_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_16_7__dout),
    .if_empty_n(fifo_B_PE_16_7__empty_n),
    .if_read(fifo_B_PE_16_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_16_7__din),
    .if_full_n(fifo_B_PE_16_7__full_n),
    .if_write(fifo_B_PE_16_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_16_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_16_8__dout),
    .if_empty_n(fifo_B_PE_16_8__empty_n),
    .if_read(fifo_B_PE_16_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_16_8__din),
    .if_full_n(fifo_B_PE_16_8__full_n),
    .if_write(fifo_B_PE_16_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_16_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_16_9__dout),
    .if_empty_n(fifo_B_PE_16_9__empty_n),
    .if_read(fifo_B_PE_16_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_16_9__din),
    .if_full_n(fifo_B_PE_16_9__full_n),
    .if_write(fifo_B_PE_16_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_17_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_17_0__dout),
    .if_empty_n(fifo_B_PE_17_0__empty_n),
    .if_read(fifo_B_PE_17_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_17_0__din),
    .if_full_n(fifo_B_PE_17_0__full_n),
    .if_write(fifo_B_PE_17_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_17_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_17_1__dout),
    .if_empty_n(fifo_B_PE_17_1__empty_n),
    .if_read(fifo_B_PE_17_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_17_1__din),
    .if_full_n(fifo_B_PE_17_1__full_n),
    .if_write(fifo_B_PE_17_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_17_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_17_10__dout),
    .if_empty_n(fifo_B_PE_17_10__empty_n),
    .if_read(fifo_B_PE_17_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_17_10__din),
    .if_full_n(fifo_B_PE_17_10__full_n),
    .if_write(fifo_B_PE_17_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_17_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_17_11__dout),
    .if_empty_n(fifo_B_PE_17_11__empty_n),
    .if_read(fifo_B_PE_17_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_17_11__din),
    .if_full_n(fifo_B_PE_17_11__full_n),
    .if_write(fifo_B_PE_17_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_17_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_17_12__dout),
    .if_empty_n(fifo_B_PE_17_12__empty_n),
    .if_read(fifo_B_PE_17_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_17_12__din),
    .if_full_n(fifo_B_PE_17_12__full_n),
    .if_write(fifo_B_PE_17_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_17_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_17_13__dout),
    .if_empty_n(fifo_B_PE_17_13__empty_n),
    .if_read(fifo_B_PE_17_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_17_13__din),
    .if_full_n(fifo_B_PE_17_13__full_n),
    .if_write(fifo_B_PE_17_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_17_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_17_14__dout),
    .if_empty_n(fifo_B_PE_17_14__empty_n),
    .if_read(fifo_B_PE_17_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_17_14__din),
    .if_full_n(fifo_B_PE_17_14__full_n),
    .if_write(fifo_B_PE_17_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_17_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_17_15__dout),
    .if_empty_n(fifo_B_PE_17_15__empty_n),
    .if_read(fifo_B_PE_17_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_17_15__din),
    .if_full_n(fifo_B_PE_17_15__full_n),
    .if_write(fifo_B_PE_17_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_17_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_17_16__dout),
    .if_empty_n(fifo_B_PE_17_16__empty_n),
    .if_read(fifo_B_PE_17_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_17_16__din),
    .if_full_n(fifo_B_PE_17_16__full_n),
    .if_write(fifo_B_PE_17_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_17_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_17_2__dout),
    .if_empty_n(fifo_B_PE_17_2__empty_n),
    .if_read(fifo_B_PE_17_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_17_2__din),
    .if_full_n(fifo_B_PE_17_2__full_n),
    .if_write(fifo_B_PE_17_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_17_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_17_3__dout),
    .if_empty_n(fifo_B_PE_17_3__empty_n),
    .if_read(fifo_B_PE_17_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_17_3__din),
    .if_full_n(fifo_B_PE_17_3__full_n),
    .if_write(fifo_B_PE_17_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_17_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_17_4__dout),
    .if_empty_n(fifo_B_PE_17_4__empty_n),
    .if_read(fifo_B_PE_17_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_17_4__din),
    .if_full_n(fifo_B_PE_17_4__full_n),
    .if_write(fifo_B_PE_17_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_17_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_17_5__dout),
    .if_empty_n(fifo_B_PE_17_5__empty_n),
    .if_read(fifo_B_PE_17_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_17_5__din),
    .if_full_n(fifo_B_PE_17_5__full_n),
    .if_write(fifo_B_PE_17_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_17_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_17_6__dout),
    .if_empty_n(fifo_B_PE_17_6__empty_n),
    .if_read(fifo_B_PE_17_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_17_6__din),
    .if_full_n(fifo_B_PE_17_6__full_n),
    .if_write(fifo_B_PE_17_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_17_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_17_7__dout),
    .if_empty_n(fifo_B_PE_17_7__empty_n),
    .if_read(fifo_B_PE_17_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_17_7__din),
    .if_full_n(fifo_B_PE_17_7__full_n),
    .if_write(fifo_B_PE_17_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_17_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_17_8__dout),
    .if_empty_n(fifo_B_PE_17_8__empty_n),
    .if_read(fifo_B_PE_17_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_17_8__din),
    .if_full_n(fifo_B_PE_17_8__full_n),
    .if_write(fifo_B_PE_17_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_17_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_17_9__dout),
    .if_empty_n(fifo_B_PE_17_9__empty_n),
    .if_read(fifo_B_PE_17_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_17_9__din),
    .if_full_n(fifo_B_PE_17_9__full_n),
    .if_write(fifo_B_PE_17_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_18_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_18_0__dout),
    .if_empty_n(fifo_B_PE_18_0__empty_n),
    .if_read(fifo_B_PE_18_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_18_0__din),
    .if_full_n(fifo_B_PE_18_0__full_n),
    .if_write(fifo_B_PE_18_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_18_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_18_1__dout),
    .if_empty_n(fifo_B_PE_18_1__empty_n),
    .if_read(fifo_B_PE_18_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_18_1__din),
    .if_full_n(fifo_B_PE_18_1__full_n),
    .if_write(fifo_B_PE_18_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_18_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_18_10__dout),
    .if_empty_n(fifo_B_PE_18_10__empty_n),
    .if_read(fifo_B_PE_18_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_18_10__din),
    .if_full_n(fifo_B_PE_18_10__full_n),
    .if_write(fifo_B_PE_18_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_18_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_18_11__dout),
    .if_empty_n(fifo_B_PE_18_11__empty_n),
    .if_read(fifo_B_PE_18_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_18_11__din),
    .if_full_n(fifo_B_PE_18_11__full_n),
    .if_write(fifo_B_PE_18_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_18_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_18_12__dout),
    .if_empty_n(fifo_B_PE_18_12__empty_n),
    .if_read(fifo_B_PE_18_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_18_12__din),
    .if_full_n(fifo_B_PE_18_12__full_n),
    .if_write(fifo_B_PE_18_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_18_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_18_13__dout),
    .if_empty_n(fifo_B_PE_18_13__empty_n),
    .if_read(fifo_B_PE_18_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_18_13__din),
    .if_full_n(fifo_B_PE_18_13__full_n),
    .if_write(fifo_B_PE_18_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_18_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_18_14__dout),
    .if_empty_n(fifo_B_PE_18_14__empty_n),
    .if_read(fifo_B_PE_18_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_18_14__din),
    .if_full_n(fifo_B_PE_18_14__full_n),
    .if_write(fifo_B_PE_18_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_18_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_18_15__dout),
    .if_empty_n(fifo_B_PE_18_15__empty_n),
    .if_read(fifo_B_PE_18_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_18_15__din),
    .if_full_n(fifo_B_PE_18_15__full_n),
    .if_write(fifo_B_PE_18_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_18_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_18_16__dout),
    .if_empty_n(fifo_B_PE_18_16__empty_n),
    .if_read(fifo_B_PE_18_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_18_16__din),
    .if_full_n(fifo_B_PE_18_16__full_n),
    .if_write(fifo_B_PE_18_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_18_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_18_2__dout),
    .if_empty_n(fifo_B_PE_18_2__empty_n),
    .if_read(fifo_B_PE_18_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_18_2__din),
    .if_full_n(fifo_B_PE_18_2__full_n),
    .if_write(fifo_B_PE_18_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_18_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_18_3__dout),
    .if_empty_n(fifo_B_PE_18_3__empty_n),
    .if_read(fifo_B_PE_18_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_18_3__din),
    .if_full_n(fifo_B_PE_18_3__full_n),
    .if_write(fifo_B_PE_18_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_18_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_18_4__dout),
    .if_empty_n(fifo_B_PE_18_4__empty_n),
    .if_read(fifo_B_PE_18_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_18_4__din),
    .if_full_n(fifo_B_PE_18_4__full_n),
    .if_write(fifo_B_PE_18_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_18_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_18_5__dout),
    .if_empty_n(fifo_B_PE_18_5__empty_n),
    .if_read(fifo_B_PE_18_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_18_5__din),
    .if_full_n(fifo_B_PE_18_5__full_n),
    .if_write(fifo_B_PE_18_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_18_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_18_6__dout),
    .if_empty_n(fifo_B_PE_18_6__empty_n),
    .if_read(fifo_B_PE_18_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_18_6__din),
    .if_full_n(fifo_B_PE_18_6__full_n),
    .if_write(fifo_B_PE_18_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_18_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_18_7__dout),
    .if_empty_n(fifo_B_PE_18_7__empty_n),
    .if_read(fifo_B_PE_18_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_18_7__din),
    .if_full_n(fifo_B_PE_18_7__full_n),
    .if_write(fifo_B_PE_18_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_18_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_18_8__dout),
    .if_empty_n(fifo_B_PE_18_8__empty_n),
    .if_read(fifo_B_PE_18_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_18_8__din),
    .if_full_n(fifo_B_PE_18_8__full_n),
    .if_write(fifo_B_PE_18_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_18_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_18_9__dout),
    .if_empty_n(fifo_B_PE_18_9__empty_n),
    .if_read(fifo_B_PE_18_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_18_9__din),
    .if_full_n(fifo_B_PE_18_9__full_n),
    .if_write(fifo_B_PE_18_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_1_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_1_0__dout),
    .if_empty_n(fifo_B_PE_1_0__empty_n),
    .if_read(fifo_B_PE_1_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_1_0__din),
    .if_full_n(fifo_B_PE_1_0__full_n),
    .if_write(fifo_B_PE_1_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_1_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_1_1__dout),
    .if_empty_n(fifo_B_PE_1_1__empty_n),
    .if_read(fifo_B_PE_1_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_1_1__din),
    .if_full_n(fifo_B_PE_1_1__full_n),
    .if_write(fifo_B_PE_1_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_1_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_1_10__dout),
    .if_empty_n(fifo_B_PE_1_10__empty_n),
    .if_read(fifo_B_PE_1_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_1_10__din),
    .if_full_n(fifo_B_PE_1_10__full_n),
    .if_write(fifo_B_PE_1_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_1_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_1_11__dout),
    .if_empty_n(fifo_B_PE_1_11__empty_n),
    .if_read(fifo_B_PE_1_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_1_11__din),
    .if_full_n(fifo_B_PE_1_11__full_n),
    .if_write(fifo_B_PE_1_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_1_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_1_12__dout),
    .if_empty_n(fifo_B_PE_1_12__empty_n),
    .if_read(fifo_B_PE_1_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_1_12__din),
    .if_full_n(fifo_B_PE_1_12__full_n),
    .if_write(fifo_B_PE_1_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_1_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_1_13__dout),
    .if_empty_n(fifo_B_PE_1_13__empty_n),
    .if_read(fifo_B_PE_1_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_1_13__din),
    .if_full_n(fifo_B_PE_1_13__full_n),
    .if_write(fifo_B_PE_1_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_1_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_1_14__dout),
    .if_empty_n(fifo_B_PE_1_14__empty_n),
    .if_read(fifo_B_PE_1_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_1_14__din),
    .if_full_n(fifo_B_PE_1_14__full_n),
    .if_write(fifo_B_PE_1_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_1_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_1_15__dout),
    .if_empty_n(fifo_B_PE_1_15__empty_n),
    .if_read(fifo_B_PE_1_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_1_15__din),
    .if_full_n(fifo_B_PE_1_15__full_n),
    .if_write(fifo_B_PE_1_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_1_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_1_16__dout),
    .if_empty_n(fifo_B_PE_1_16__empty_n),
    .if_read(fifo_B_PE_1_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_1_16__din),
    .if_full_n(fifo_B_PE_1_16__full_n),
    .if_write(fifo_B_PE_1_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_1_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_1_2__dout),
    .if_empty_n(fifo_B_PE_1_2__empty_n),
    .if_read(fifo_B_PE_1_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_1_2__din),
    .if_full_n(fifo_B_PE_1_2__full_n),
    .if_write(fifo_B_PE_1_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_1_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_1_3__dout),
    .if_empty_n(fifo_B_PE_1_3__empty_n),
    .if_read(fifo_B_PE_1_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_1_3__din),
    .if_full_n(fifo_B_PE_1_3__full_n),
    .if_write(fifo_B_PE_1_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_1_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_1_4__dout),
    .if_empty_n(fifo_B_PE_1_4__empty_n),
    .if_read(fifo_B_PE_1_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_1_4__din),
    .if_full_n(fifo_B_PE_1_4__full_n),
    .if_write(fifo_B_PE_1_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_1_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_1_5__dout),
    .if_empty_n(fifo_B_PE_1_5__empty_n),
    .if_read(fifo_B_PE_1_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_1_5__din),
    .if_full_n(fifo_B_PE_1_5__full_n),
    .if_write(fifo_B_PE_1_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_1_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_1_6__dout),
    .if_empty_n(fifo_B_PE_1_6__empty_n),
    .if_read(fifo_B_PE_1_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_1_6__din),
    .if_full_n(fifo_B_PE_1_6__full_n),
    .if_write(fifo_B_PE_1_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_1_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_1_7__dout),
    .if_empty_n(fifo_B_PE_1_7__empty_n),
    .if_read(fifo_B_PE_1_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_1_7__din),
    .if_full_n(fifo_B_PE_1_7__full_n),
    .if_write(fifo_B_PE_1_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_1_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_1_8__dout),
    .if_empty_n(fifo_B_PE_1_8__empty_n),
    .if_read(fifo_B_PE_1_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_1_8__din),
    .if_full_n(fifo_B_PE_1_8__full_n),
    .if_write(fifo_B_PE_1_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_1_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_1_9__dout),
    .if_empty_n(fifo_B_PE_1_9__empty_n),
    .if_read(fifo_B_PE_1_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_1_9__din),
    .if_full_n(fifo_B_PE_1_9__full_n),
    .if_write(fifo_B_PE_1_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_2_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_2_0__dout),
    .if_empty_n(fifo_B_PE_2_0__empty_n),
    .if_read(fifo_B_PE_2_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_2_0__din),
    .if_full_n(fifo_B_PE_2_0__full_n),
    .if_write(fifo_B_PE_2_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_2_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_2_1__dout),
    .if_empty_n(fifo_B_PE_2_1__empty_n),
    .if_read(fifo_B_PE_2_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_2_1__din),
    .if_full_n(fifo_B_PE_2_1__full_n),
    .if_write(fifo_B_PE_2_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_2_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_2_10__dout),
    .if_empty_n(fifo_B_PE_2_10__empty_n),
    .if_read(fifo_B_PE_2_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_2_10__din),
    .if_full_n(fifo_B_PE_2_10__full_n),
    .if_write(fifo_B_PE_2_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_2_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_2_11__dout),
    .if_empty_n(fifo_B_PE_2_11__empty_n),
    .if_read(fifo_B_PE_2_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_2_11__din),
    .if_full_n(fifo_B_PE_2_11__full_n),
    .if_write(fifo_B_PE_2_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_2_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_2_12__dout),
    .if_empty_n(fifo_B_PE_2_12__empty_n),
    .if_read(fifo_B_PE_2_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_2_12__din),
    .if_full_n(fifo_B_PE_2_12__full_n),
    .if_write(fifo_B_PE_2_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_2_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_2_13__dout),
    .if_empty_n(fifo_B_PE_2_13__empty_n),
    .if_read(fifo_B_PE_2_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_2_13__din),
    .if_full_n(fifo_B_PE_2_13__full_n),
    .if_write(fifo_B_PE_2_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_2_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_2_14__dout),
    .if_empty_n(fifo_B_PE_2_14__empty_n),
    .if_read(fifo_B_PE_2_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_2_14__din),
    .if_full_n(fifo_B_PE_2_14__full_n),
    .if_write(fifo_B_PE_2_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_2_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_2_15__dout),
    .if_empty_n(fifo_B_PE_2_15__empty_n),
    .if_read(fifo_B_PE_2_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_2_15__din),
    .if_full_n(fifo_B_PE_2_15__full_n),
    .if_write(fifo_B_PE_2_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_2_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_2_16__dout),
    .if_empty_n(fifo_B_PE_2_16__empty_n),
    .if_read(fifo_B_PE_2_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_2_16__din),
    .if_full_n(fifo_B_PE_2_16__full_n),
    .if_write(fifo_B_PE_2_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_2_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_2_2__dout),
    .if_empty_n(fifo_B_PE_2_2__empty_n),
    .if_read(fifo_B_PE_2_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_2_2__din),
    .if_full_n(fifo_B_PE_2_2__full_n),
    .if_write(fifo_B_PE_2_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_2_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_2_3__dout),
    .if_empty_n(fifo_B_PE_2_3__empty_n),
    .if_read(fifo_B_PE_2_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_2_3__din),
    .if_full_n(fifo_B_PE_2_3__full_n),
    .if_write(fifo_B_PE_2_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_2_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_2_4__dout),
    .if_empty_n(fifo_B_PE_2_4__empty_n),
    .if_read(fifo_B_PE_2_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_2_4__din),
    .if_full_n(fifo_B_PE_2_4__full_n),
    .if_write(fifo_B_PE_2_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_2_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_2_5__dout),
    .if_empty_n(fifo_B_PE_2_5__empty_n),
    .if_read(fifo_B_PE_2_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_2_5__din),
    .if_full_n(fifo_B_PE_2_5__full_n),
    .if_write(fifo_B_PE_2_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_2_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_2_6__dout),
    .if_empty_n(fifo_B_PE_2_6__empty_n),
    .if_read(fifo_B_PE_2_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_2_6__din),
    .if_full_n(fifo_B_PE_2_6__full_n),
    .if_write(fifo_B_PE_2_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_2_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_2_7__dout),
    .if_empty_n(fifo_B_PE_2_7__empty_n),
    .if_read(fifo_B_PE_2_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_2_7__din),
    .if_full_n(fifo_B_PE_2_7__full_n),
    .if_write(fifo_B_PE_2_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_2_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_2_8__dout),
    .if_empty_n(fifo_B_PE_2_8__empty_n),
    .if_read(fifo_B_PE_2_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_2_8__din),
    .if_full_n(fifo_B_PE_2_8__full_n),
    .if_write(fifo_B_PE_2_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_2_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_2_9__dout),
    .if_empty_n(fifo_B_PE_2_9__empty_n),
    .if_read(fifo_B_PE_2_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_2_9__din),
    .if_full_n(fifo_B_PE_2_9__full_n),
    .if_write(fifo_B_PE_2_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_3_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_3_0__dout),
    .if_empty_n(fifo_B_PE_3_0__empty_n),
    .if_read(fifo_B_PE_3_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_3_0__din),
    .if_full_n(fifo_B_PE_3_0__full_n),
    .if_write(fifo_B_PE_3_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_3_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_3_1__dout),
    .if_empty_n(fifo_B_PE_3_1__empty_n),
    .if_read(fifo_B_PE_3_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_3_1__din),
    .if_full_n(fifo_B_PE_3_1__full_n),
    .if_write(fifo_B_PE_3_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_3_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_3_10__dout),
    .if_empty_n(fifo_B_PE_3_10__empty_n),
    .if_read(fifo_B_PE_3_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_3_10__din),
    .if_full_n(fifo_B_PE_3_10__full_n),
    .if_write(fifo_B_PE_3_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_3_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_3_11__dout),
    .if_empty_n(fifo_B_PE_3_11__empty_n),
    .if_read(fifo_B_PE_3_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_3_11__din),
    .if_full_n(fifo_B_PE_3_11__full_n),
    .if_write(fifo_B_PE_3_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_3_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_3_12__dout),
    .if_empty_n(fifo_B_PE_3_12__empty_n),
    .if_read(fifo_B_PE_3_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_3_12__din),
    .if_full_n(fifo_B_PE_3_12__full_n),
    .if_write(fifo_B_PE_3_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_3_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_3_13__dout),
    .if_empty_n(fifo_B_PE_3_13__empty_n),
    .if_read(fifo_B_PE_3_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_3_13__din),
    .if_full_n(fifo_B_PE_3_13__full_n),
    .if_write(fifo_B_PE_3_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_3_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_3_14__dout),
    .if_empty_n(fifo_B_PE_3_14__empty_n),
    .if_read(fifo_B_PE_3_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_3_14__din),
    .if_full_n(fifo_B_PE_3_14__full_n),
    .if_write(fifo_B_PE_3_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_3_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_3_15__dout),
    .if_empty_n(fifo_B_PE_3_15__empty_n),
    .if_read(fifo_B_PE_3_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_3_15__din),
    .if_full_n(fifo_B_PE_3_15__full_n),
    .if_write(fifo_B_PE_3_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_3_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_3_16__dout),
    .if_empty_n(fifo_B_PE_3_16__empty_n),
    .if_read(fifo_B_PE_3_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_3_16__din),
    .if_full_n(fifo_B_PE_3_16__full_n),
    .if_write(fifo_B_PE_3_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_3_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_3_2__dout),
    .if_empty_n(fifo_B_PE_3_2__empty_n),
    .if_read(fifo_B_PE_3_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_3_2__din),
    .if_full_n(fifo_B_PE_3_2__full_n),
    .if_write(fifo_B_PE_3_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_3_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_3_3__dout),
    .if_empty_n(fifo_B_PE_3_3__empty_n),
    .if_read(fifo_B_PE_3_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_3_3__din),
    .if_full_n(fifo_B_PE_3_3__full_n),
    .if_write(fifo_B_PE_3_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_3_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_3_4__dout),
    .if_empty_n(fifo_B_PE_3_4__empty_n),
    .if_read(fifo_B_PE_3_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_3_4__din),
    .if_full_n(fifo_B_PE_3_4__full_n),
    .if_write(fifo_B_PE_3_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_3_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_3_5__dout),
    .if_empty_n(fifo_B_PE_3_5__empty_n),
    .if_read(fifo_B_PE_3_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_3_5__din),
    .if_full_n(fifo_B_PE_3_5__full_n),
    .if_write(fifo_B_PE_3_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_3_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_3_6__dout),
    .if_empty_n(fifo_B_PE_3_6__empty_n),
    .if_read(fifo_B_PE_3_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_3_6__din),
    .if_full_n(fifo_B_PE_3_6__full_n),
    .if_write(fifo_B_PE_3_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_3_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_3_7__dout),
    .if_empty_n(fifo_B_PE_3_7__empty_n),
    .if_read(fifo_B_PE_3_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_3_7__din),
    .if_full_n(fifo_B_PE_3_7__full_n),
    .if_write(fifo_B_PE_3_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_3_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_3_8__dout),
    .if_empty_n(fifo_B_PE_3_8__empty_n),
    .if_read(fifo_B_PE_3_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_3_8__din),
    .if_full_n(fifo_B_PE_3_8__full_n),
    .if_write(fifo_B_PE_3_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_3_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_3_9__dout),
    .if_empty_n(fifo_B_PE_3_9__empty_n),
    .if_read(fifo_B_PE_3_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_3_9__din),
    .if_full_n(fifo_B_PE_3_9__full_n),
    .if_write(fifo_B_PE_3_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_4_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_4_0__dout),
    .if_empty_n(fifo_B_PE_4_0__empty_n),
    .if_read(fifo_B_PE_4_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_4_0__din),
    .if_full_n(fifo_B_PE_4_0__full_n),
    .if_write(fifo_B_PE_4_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_4_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_4_1__dout),
    .if_empty_n(fifo_B_PE_4_1__empty_n),
    .if_read(fifo_B_PE_4_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_4_1__din),
    .if_full_n(fifo_B_PE_4_1__full_n),
    .if_write(fifo_B_PE_4_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_4_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_4_10__dout),
    .if_empty_n(fifo_B_PE_4_10__empty_n),
    .if_read(fifo_B_PE_4_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_4_10__din),
    .if_full_n(fifo_B_PE_4_10__full_n),
    .if_write(fifo_B_PE_4_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_4_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_4_11__dout),
    .if_empty_n(fifo_B_PE_4_11__empty_n),
    .if_read(fifo_B_PE_4_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_4_11__din),
    .if_full_n(fifo_B_PE_4_11__full_n),
    .if_write(fifo_B_PE_4_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_4_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_4_12__dout),
    .if_empty_n(fifo_B_PE_4_12__empty_n),
    .if_read(fifo_B_PE_4_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_4_12__din),
    .if_full_n(fifo_B_PE_4_12__full_n),
    .if_write(fifo_B_PE_4_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_4_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_4_13__dout),
    .if_empty_n(fifo_B_PE_4_13__empty_n),
    .if_read(fifo_B_PE_4_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_4_13__din),
    .if_full_n(fifo_B_PE_4_13__full_n),
    .if_write(fifo_B_PE_4_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_4_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_4_14__dout),
    .if_empty_n(fifo_B_PE_4_14__empty_n),
    .if_read(fifo_B_PE_4_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_4_14__din),
    .if_full_n(fifo_B_PE_4_14__full_n),
    .if_write(fifo_B_PE_4_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_4_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_4_15__dout),
    .if_empty_n(fifo_B_PE_4_15__empty_n),
    .if_read(fifo_B_PE_4_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_4_15__din),
    .if_full_n(fifo_B_PE_4_15__full_n),
    .if_write(fifo_B_PE_4_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_4_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_4_16__dout),
    .if_empty_n(fifo_B_PE_4_16__empty_n),
    .if_read(fifo_B_PE_4_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_4_16__din),
    .if_full_n(fifo_B_PE_4_16__full_n),
    .if_write(fifo_B_PE_4_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_4_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_4_2__dout),
    .if_empty_n(fifo_B_PE_4_2__empty_n),
    .if_read(fifo_B_PE_4_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_4_2__din),
    .if_full_n(fifo_B_PE_4_2__full_n),
    .if_write(fifo_B_PE_4_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_4_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_4_3__dout),
    .if_empty_n(fifo_B_PE_4_3__empty_n),
    .if_read(fifo_B_PE_4_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_4_3__din),
    .if_full_n(fifo_B_PE_4_3__full_n),
    .if_write(fifo_B_PE_4_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_4_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_4_4__dout),
    .if_empty_n(fifo_B_PE_4_4__empty_n),
    .if_read(fifo_B_PE_4_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_4_4__din),
    .if_full_n(fifo_B_PE_4_4__full_n),
    .if_write(fifo_B_PE_4_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_4_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_4_5__dout),
    .if_empty_n(fifo_B_PE_4_5__empty_n),
    .if_read(fifo_B_PE_4_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_4_5__din),
    .if_full_n(fifo_B_PE_4_5__full_n),
    .if_write(fifo_B_PE_4_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_4_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_4_6__dout),
    .if_empty_n(fifo_B_PE_4_6__empty_n),
    .if_read(fifo_B_PE_4_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_4_6__din),
    .if_full_n(fifo_B_PE_4_6__full_n),
    .if_write(fifo_B_PE_4_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_4_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_4_7__dout),
    .if_empty_n(fifo_B_PE_4_7__empty_n),
    .if_read(fifo_B_PE_4_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_4_7__din),
    .if_full_n(fifo_B_PE_4_7__full_n),
    .if_write(fifo_B_PE_4_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_4_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_4_8__dout),
    .if_empty_n(fifo_B_PE_4_8__empty_n),
    .if_read(fifo_B_PE_4_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_4_8__din),
    .if_full_n(fifo_B_PE_4_8__full_n),
    .if_write(fifo_B_PE_4_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_4_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_4_9__dout),
    .if_empty_n(fifo_B_PE_4_9__empty_n),
    .if_read(fifo_B_PE_4_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_4_9__din),
    .if_full_n(fifo_B_PE_4_9__full_n),
    .if_write(fifo_B_PE_4_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_5_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_5_0__dout),
    .if_empty_n(fifo_B_PE_5_0__empty_n),
    .if_read(fifo_B_PE_5_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_5_0__din),
    .if_full_n(fifo_B_PE_5_0__full_n),
    .if_write(fifo_B_PE_5_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_5_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_5_1__dout),
    .if_empty_n(fifo_B_PE_5_1__empty_n),
    .if_read(fifo_B_PE_5_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_5_1__din),
    .if_full_n(fifo_B_PE_5_1__full_n),
    .if_write(fifo_B_PE_5_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_5_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_5_10__dout),
    .if_empty_n(fifo_B_PE_5_10__empty_n),
    .if_read(fifo_B_PE_5_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_5_10__din),
    .if_full_n(fifo_B_PE_5_10__full_n),
    .if_write(fifo_B_PE_5_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_5_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_5_11__dout),
    .if_empty_n(fifo_B_PE_5_11__empty_n),
    .if_read(fifo_B_PE_5_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_5_11__din),
    .if_full_n(fifo_B_PE_5_11__full_n),
    .if_write(fifo_B_PE_5_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_5_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_5_12__dout),
    .if_empty_n(fifo_B_PE_5_12__empty_n),
    .if_read(fifo_B_PE_5_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_5_12__din),
    .if_full_n(fifo_B_PE_5_12__full_n),
    .if_write(fifo_B_PE_5_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_5_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_5_13__dout),
    .if_empty_n(fifo_B_PE_5_13__empty_n),
    .if_read(fifo_B_PE_5_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_5_13__din),
    .if_full_n(fifo_B_PE_5_13__full_n),
    .if_write(fifo_B_PE_5_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_5_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_5_14__dout),
    .if_empty_n(fifo_B_PE_5_14__empty_n),
    .if_read(fifo_B_PE_5_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_5_14__din),
    .if_full_n(fifo_B_PE_5_14__full_n),
    .if_write(fifo_B_PE_5_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_5_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_5_15__dout),
    .if_empty_n(fifo_B_PE_5_15__empty_n),
    .if_read(fifo_B_PE_5_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_5_15__din),
    .if_full_n(fifo_B_PE_5_15__full_n),
    .if_write(fifo_B_PE_5_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_5_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_5_16__dout),
    .if_empty_n(fifo_B_PE_5_16__empty_n),
    .if_read(fifo_B_PE_5_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_5_16__din),
    .if_full_n(fifo_B_PE_5_16__full_n),
    .if_write(fifo_B_PE_5_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_5_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_5_2__dout),
    .if_empty_n(fifo_B_PE_5_2__empty_n),
    .if_read(fifo_B_PE_5_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_5_2__din),
    .if_full_n(fifo_B_PE_5_2__full_n),
    .if_write(fifo_B_PE_5_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_5_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_5_3__dout),
    .if_empty_n(fifo_B_PE_5_3__empty_n),
    .if_read(fifo_B_PE_5_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_5_3__din),
    .if_full_n(fifo_B_PE_5_3__full_n),
    .if_write(fifo_B_PE_5_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_5_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_5_4__dout),
    .if_empty_n(fifo_B_PE_5_4__empty_n),
    .if_read(fifo_B_PE_5_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_5_4__din),
    .if_full_n(fifo_B_PE_5_4__full_n),
    .if_write(fifo_B_PE_5_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_5_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_5_5__dout),
    .if_empty_n(fifo_B_PE_5_5__empty_n),
    .if_read(fifo_B_PE_5_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_5_5__din),
    .if_full_n(fifo_B_PE_5_5__full_n),
    .if_write(fifo_B_PE_5_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_5_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_5_6__dout),
    .if_empty_n(fifo_B_PE_5_6__empty_n),
    .if_read(fifo_B_PE_5_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_5_6__din),
    .if_full_n(fifo_B_PE_5_6__full_n),
    .if_write(fifo_B_PE_5_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_5_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_5_7__dout),
    .if_empty_n(fifo_B_PE_5_7__empty_n),
    .if_read(fifo_B_PE_5_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_5_7__din),
    .if_full_n(fifo_B_PE_5_7__full_n),
    .if_write(fifo_B_PE_5_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_5_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_5_8__dout),
    .if_empty_n(fifo_B_PE_5_8__empty_n),
    .if_read(fifo_B_PE_5_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_5_8__din),
    .if_full_n(fifo_B_PE_5_8__full_n),
    .if_write(fifo_B_PE_5_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_5_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_5_9__dout),
    .if_empty_n(fifo_B_PE_5_9__empty_n),
    .if_read(fifo_B_PE_5_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_5_9__din),
    .if_full_n(fifo_B_PE_5_9__full_n),
    .if_write(fifo_B_PE_5_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_6_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_6_0__dout),
    .if_empty_n(fifo_B_PE_6_0__empty_n),
    .if_read(fifo_B_PE_6_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_6_0__din),
    .if_full_n(fifo_B_PE_6_0__full_n),
    .if_write(fifo_B_PE_6_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_6_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_6_1__dout),
    .if_empty_n(fifo_B_PE_6_1__empty_n),
    .if_read(fifo_B_PE_6_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_6_1__din),
    .if_full_n(fifo_B_PE_6_1__full_n),
    .if_write(fifo_B_PE_6_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_6_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_6_10__dout),
    .if_empty_n(fifo_B_PE_6_10__empty_n),
    .if_read(fifo_B_PE_6_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_6_10__din),
    .if_full_n(fifo_B_PE_6_10__full_n),
    .if_write(fifo_B_PE_6_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_6_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_6_11__dout),
    .if_empty_n(fifo_B_PE_6_11__empty_n),
    .if_read(fifo_B_PE_6_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_6_11__din),
    .if_full_n(fifo_B_PE_6_11__full_n),
    .if_write(fifo_B_PE_6_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_6_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_6_12__dout),
    .if_empty_n(fifo_B_PE_6_12__empty_n),
    .if_read(fifo_B_PE_6_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_6_12__din),
    .if_full_n(fifo_B_PE_6_12__full_n),
    .if_write(fifo_B_PE_6_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_6_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_6_13__dout),
    .if_empty_n(fifo_B_PE_6_13__empty_n),
    .if_read(fifo_B_PE_6_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_6_13__din),
    .if_full_n(fifo_B_PE_6_13__full_n),
    .if_write(fifo_B_PE_6_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_6_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_6_14__dout),
    .if_empty_n(fifo_B_PE_6_14__empty_n),
    .if_read(fifo_B_PE_6_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_6_14__din),
    .if_full_n(fifo_B_PE_6_14__full_n),
    .if_write(fifo_B_PE_6_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_6_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_6_15__dout),
    .if_empty_n(fifo_B_PE_6_15__empty_n),
    .if_read(fifo_B_PE_6_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_6_15__din),
    .if_full_n(fifo_B_PE_6_15__full_n),
    .if_write(fifo_B_PE_6_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_6_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_6_16__dout),
    .if_empty_n(fifo_B_PE_6_16__empty_n),
    .if_read(fifo_B_PE_6_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_6_16__din),
    .if_full_n(fifo_B_PE_6_16__full_n),
    .if_write(fifo_B_PE_6_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_6_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_6_2__dout),
    .if_empty_n(fifo_B_PE_6_2__empty_n),
    .if_read(fifo_B_PE_6_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_6_2__din),
    .if_full_n(fifo_B_PE_6_2__full_n),
    .if_write(fifo_B_PE_6_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_6_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_6_3__dout),
    .if_empty_n(fifo_B_PE_6_3__empty_n),
    .if_read(fifo_B_PE_6_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_6_3__din),
    .if_full_n(fifo_B_PE_6_3__full_n),
    .if_write(fifo_B_PE_6_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_6_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_6_4__dout),
    .if_empty_n(fifo_B_PE_6_4__empty_n),
    .if_read(fifo_B_PE_6_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_6_4__din),
    .if_full_n(fifo_B_PE_6_4__full_n),
    .if_write(fifo_B_PE_6_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_6_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_6_5__dout),
    .if_empty_n(fifo_B_PE_6_5__empty_n),
    .if_read(fifo_B_PE_6_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_6_5__din),
    .if_full_n(fifo_B_PE_6_5__full_n),
    .if_write(fifo_B_PE_6_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_6_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_6_6__dout),
    .if_empty_n(fifo_B_PE_6_6__empty_n),
    .if_read(fifo_B_PE_6_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_6_6__din),
    .if_full_n(fifo_B_PE_6_6__full_n),
    .if_write(fifo_B_PE_6_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_6_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_6_7__dout),
    .if_empty_n(fifo_B_PE_6_7__empty_n),
    .if_read(fifo_B_PE_6_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_6_7__din),
    .if_full_n(fifo_B_PE_6_7__full_n),
    .if_write(fifo_B_PE_6_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_6_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_6_8__dout),
    .if_empty_n(fifo_B_PE_6_8__empty_n),
    .if_read(fifo_B_PE_6_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_6_8__din),
    .if_full_n(fifo_B_PE_6_8__full_n),
    .if_write(fifo_B_PE_6_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_6_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_6_9__dout),
    .if_empty_n(fifo_B_PE_6_9__empty_n),
    .if_read(fifo_B_PE_6_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_6_9__din),
    .if_full_n(fifo_B_PE_6_9__full_n),
    .if_write(fifo_B_PE_6_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_7_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_7_0__dout),
    .if_empty_n(fifo_B_PE_7_0__empty_n),
    .if_read(fifo_B_PE_7_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_7_0__din),
    .if_full_n(fifo_B_PE_7_0__full_n),
    .if_write(fifo_B_PE_7_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_7_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_7_1__dout),
    .if_empty_n(fifo_B_PE_7_1__empty_n),
    .if_read(fifo_B_PE_7_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_7_1__din),
    .if_full_n(fifo_B_PE_7_1__full_n),
    .if_write(fifo_B_PE_7_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_7_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_7_10__dout),
    .if_empty_n(fifo_B_PE_7_10__empty_n),
    .if_read(fifo_B_PE_7_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_7_10__din),
    .if_full_n(fifo_B_PE_7_10__full_n),
    .if_write(fifo_B_PE_7_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_7_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_7_11__dout),
    .if_empty_n(fifo_B_PE_7_11__empty_n),
    .if_read(fifo_B_PE_7_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_7_11__din),
    .if_full_n(fifo_B_PE_7_11__full_n),
    .if_write(fifo_B_PE_7_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_7_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_7_12__dout),
    .if_empty_n(fifo_B_PE_7_12__empty_n),
    .if_read(fifo_B_PE_7_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_7_12__din),
    .if_full_n(fifo_B_PE_7_12__full_n),
    .if_write(fifo_B_PE_7_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_7_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_7_13__dout),
    .if_empty_n(fifo_B_PE_7_13__empty_n),
    .if_read(fifo_B_PE_7_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_7_13__din),
    .if_full_n(fifo_B_PE_7_13__full_n),
    .if_write(fifo_B_PE_7_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_7_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_7_14__dout),
    .if_empty_n(fifo_B_PE_7_14__empty_n),
    .if_read(fifo_B_PE_7_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_7_14__din),
    .if_full_n(fifo_B_PE_7_14__full_n),
    .if_write(fifo_B_PE_7_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_7_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_7_15__dout),
    .if_empty_n(fifo_B_PE_7_15__empty_n),
    .if_read(fifo_B_PE_7_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_7_15__din),
    .if_full_n(fifo_B_PE_7_15__full_n),
    .if_write(fifo_B_PE_7_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_7_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_7_16__dout),
    .if_empty_n(fifo_B_PE_7_16__empty_n),
    .if_read(fifo_B_PE_7_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_7_16__din),
    .if_full_n(fifo_B_PE_7_16__full_n),
    .if_write(fifo_B_PE_7_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_7_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_7_2__dout),
    .if_empty_n(fifo_B_PE_7_2__empty_n),
    .if_read(fifo_B_PE_7_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_7_2__din),
    .if_full_n(fifo_B_PE_7_2__full_n),
    .if_write(fifo_B_PE_7_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_7_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_7_3__dout),
    .if_empty_n(fifo_B_PE_7_3__empty_n),
    .if_read(fifo_B_PE_7_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_7_3__din),
    .if_full_n(fifo_B_PE_7_3__full_n),
    .if_write(fifo_B_PE_7_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_7_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_7_4__dout),
    .if_empty_n(fifo_B_PE_7_4__empty_n),
    .if_read(fifo_B_PE_7_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_7_4__din),
    .if_full_n(fifo_B_PE_7_4__full_n),
    .if_write(fifo_B_PE_7_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_7_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_7_5__dout),
    .if_empty_n(fifo_B_PE_7_5__empty_n),
    .if_read(fifo_B_PE_7_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_7_5__din),
    .if_full_n(fifo_B_PE_7_5__full_n),
    .if_write(fifo_B_PE_7_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_7_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_7_6__dout),
    .if_empty_n(fifo_B_PE_7_6__empty_n),
    .if_read(fifo_B_PE_7_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_7_6__din),
    .if_full_n(fifo_B_PE_7_6__full_n),
    .if_write(fifo_B_PE_7_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_7_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_7_7__dout),
    .if_empty_n(fifo_B_PE_7_7__empty_n),
    .if_read(fifo_B_PE_7_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_7_7__din),
    .if_full_n(fifo_B_PE_7_7__full_n),
    .if_write(fifo_B_PE_7_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_7_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_7_8__dout),
    .if_empty_n(fifo_B_PE_7_8__empty_n),
    .if_read(fifo_B_PE_7_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_7_8__din),
    .if_full_n(fifo_B_PE_7_8__full_n),
    .if_write(fifo_B_PE_7_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_7_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_7_9__dout),
    .if_empty_n(fifo_B_PE_7_9__empty_n),
    .if_read(fifo_B_PE_7_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_7_9__din),
    .if_full_n(fifo_B_PE_7_9__full_n),
    .if_write(fifo_B_PE_7_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_8_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_8_0__dout),
    .if_empty_n(fifo_B_PE_8_0__empty_n),
    .if_read(fifo_B_PE_8_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_8_0__din),
    .if_full_n(fifo_B_PE_8_0__full_n),
    .if_write(fifo_B_PE_8_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_8_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_8_1__dout),
    .if_empty_n(fifo_B_PE_8_1__empty_n),
    .if_read(fifo_B_PE_8_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_8_1__din),
    .if_full_n(fifo_B_PE_8_1__full_n),
    .if_write(fifo_B_PE_8_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_8_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_8_10__dout),
    .if_empty_n(fifo_B_PE_8_10__empty_n),
    .if_read(fifo_B_PE_8_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_8_10__din),
    .if_full_n(fifo_B_PE_8_10__full_n),
    .if_write(fifo_B_PE_8_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_8_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_8_11__dout),
    .if_empty_n(fifo_B_PE_8_11__empty_n),
    .if_read(fifo_B_PE_8_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_8_11__din),
    .if_full_n(fifo_B_PE_8_11__full_n),
    .if_write(fifo_B_PE_8_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_8_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_8_12__dout),
    .if_empty_n(fifo_B_PE_8_12__empty_n),
    .if_read(fifo_B_PE_8_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_8_12__din),
    .if_full_n(fifo_B_PE_8_12__full_n),
    .if_write(fifo_B_PE_8_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_8_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_8_13__dout),
    .if_empty_n(fifo_B_PE_8_13__empty_n),
    .if_read(fifo_B_PE_8_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_8_13__din),
    .if_full_n(fifo_B_PE_8_13__full_n),
    .if_write(fifo_B_PE_8_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_8_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_8_14__dout),
    .if_empty_n(fifo_B_PE_8_14__empty_n),
    .if_read(fifo_B_PE_8_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_8_14__din),
    .if_full_n(fifo_B_PE_8_14__full_n),
    .if_write(fifo_B_PE_8_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_8_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_8_15__dout),
    .if_empty_n(fifo_B_PE_8_15__empty_n),
    .if_read(fifo_B_PE_8_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_8_15__din),
    .if_full_n(fifo_B_PE_8_15__full_n),
    .if_write(fifo_B_PE_8_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_8_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_8_16__dout),
    .if_empty_n(fifo_B_PE_8_16__empty_n),
    .if_read(fifo_B_PE_8_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_8_16__din),
    .if_full_n(fifo_B_PE_8_16__full_n),
    .if_write(fifo_B_PE_8_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_8_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_8_2__dout),
    .if_empty_n(fifo_B_PE_8_2__empty_n),
    .if_read(fifo_B_PE_8_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_8_2__din),
    .if_full_n(fifo_B_PE_8_2__full_n),
    .if_write(fifo_B_PE_8_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_8_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_8_3__dout),
    .if_empty_n(fifo_B_PE_8_3__empty_n),
    .if_read(fifo_B_PE_8_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_8_3__din),
    .if_full_n(fifo_B_PE_8_3__full_n),
    .if_write(fifo_B_PE_8_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_8_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_8_4__dout),
    .if_empty_n(fifo_B_PE_8_4__empty_n),
    .if_read(fifo_B_PE_8_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_8_4__din),
    .if_full_n(fifo_B_PE_8_4__full_n),
    .if_write(fifo_B_PE_8_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_8_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_8_5__dout),
    .if_empty_n(fifo_B_PE_8_5__empty_n),
    .if_read(fifo_B_PE_8_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_8_5__din),
    .if_full_n(fifo_B_PE_8_5__full_n),
    .if_write(fifo_B_PE_8_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_8_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_8_6__dout),
    .if_empty_n(fifo_B_PE_8_6__empty_n),
    .if_read(fifo_B_PE_8_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_8_6__din),
    .if_full_n(fifo_B_PE_8_6__full_n),
    .if_write(fifo_B_PE_8_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_8_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_8_7__dout),
    .if_empty_n(fifo_B_PE_8_7__empty_n),
    .if_read(fifo_B_PE_8_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_8_7__din),
    .if_full_n(fifo_B_PE_8_7__full_n),
    .if_write(fifo_B_PE_8_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_8_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_8_8__dout),
    .if_empty_n(fifo_B_PE_8_8__empty_n),
    .if_read(fifo_B_PE_8_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_8_8__din),
    .if_full_n(fifo_B_PE_8_8__full_n),
    .if_write(fifo_B_PE_8_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_8_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_8_9__dout),
    .if_empty_n(fifo_B_PE_8_9__empty_n),
    .if_read(fifo_B_PE_8_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_8_9__din),
    .if_full_n(fifo_B_PE_8_9__full_n),
    .if_write(fifo_B_PE_8_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_9_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_9_0__dout),
    .if_empty_n(fifo_B_PE_9_0__empty_n),
    .if_read(fifo_B_PE_9_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_9_0__din),
    .if_full_n(fifo_B_PE_9_0__full_n),
    .if_write(fifo_B_PE_9_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_9_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_9_1__dout),
    .if_empty_n(fifo_B_PE_9_1__empty_n),
    .if_read(fifo_B_PE_9_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_9_1__din),
    .if_full_n(fifo_B_PE_9_1__full_n),
    .if_write(fifo_B_PE_9_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_9_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_9_10__dout),
    .if_empty_n(fifo_B_PE_9_10__empty_n),
    .if_read(fifo_B_PE_9_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_9_10__din),
    .if_full_n(fifo_B_PE_9_10__full_n),
    .if_write(fifo_B_PE_9_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_9_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_9_11__dout),
    .if_empty_n(fifo_B_PE_9_11__empty_n),
    .if_read(fifo_B_PE_9_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_9_11__din),
    .if_full_n(fifo_B_PE_9_11__full_n),
    .if_write(fifo_B_PE_9_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_9_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_9_12__dout),
    .if_empty_n(fifo_B_PE_9_12__empty_n),
    .if_read(fifo_B_PE_9_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_9_12__din),
    .if_full_n(fifo_B_PE_9_12__full_n),
    .if_write(fifo_B_PE_9_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_9_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_9_13__dout),
    .if_empty_n(fifo_B_PE_9_13__empty_n),
    .if_read(fifo_B_PE_9_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_9_13__din),
    .if_full_n(fifo_B_PE_9_13__full_n),
    .if_write(fifo_B_PE_9_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_9_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_9_14__dout),
    .if_empty_n(fifo_B_PE_9_14__empty_n),
    .if_read(fifo_B_PE_9_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_9_14__din),
    .if_full_n(fifo_B_PE_9_14__full_n),
    .if_write(fifo_B_PE_9_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_9_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_9_15__dout),
    .if_empty_n(fifo_B_PE_9_15__empty_n),
    .if_read(fifo_B_PE_9_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_9_15__din),
    .if_full_n(fifo_B_PE_9_15__full_n),
    .if_write(fifo_B_PE_9_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_9_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_9_16__dout),
    .if_empty_n(fifo_B_PE_9_16__empty_n),
    .if_read(fifo_B_PE_9_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_9_16__din),
    .if_full_n(fifo_B_PE_9_16__full_n),
    .if_write(fifo_B_PE_9_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_9_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_9_2__dout),
    .if_empty_n(fifo_B_PE_9_2__empty_n),
    .if_read(fifo_B_PE_9_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_9_2__din),
    .if_full_n(fifo_B_PE_9_2__full_n),
    .if_write(fifo_B_PE_9_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_9_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_9_3__dout),
    .if_empty_n(fifo_B_PE_9_3__empty_n),
    .if_read(fifo_B_PE_9_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_9_3__din),
    .if_full_n(fifo_B_PE_9_3__full_n),
    .if_write(fifo_B_PE_9_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_9_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_9_4__dout),
    .if_empty_n(fifo_B_PE_9_4__empty_n),
    .if_read(fifo_B_PE_9_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_9_4__din),
    .if_full_n(fifo_B_PE_9_4__full_n),
    .if_write(fifo_B_PE_9_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_9_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_9_5__dout),
    .if_empty_n(fifo_B_PE_9_5__empty_n),
    .if_read(fifo_B_PE_9_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_9_5__din),
    .if_full_n(fifo_B_PE_9_5__full_n),
    .if_write(fifo_B_PE_9_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_9_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_9_6__dout),
    .if_empty_n(fifo_B_PE_9_6__empty_n),
    .if_read(fifo_B_PE_9_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_9_6__din),
    .if_full_n(fifo_B_PE_9_6__full_n),
    .if_write(fifo_B_PE_9_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_9_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_9_7__dout),
    .if_empty_n(fifo_B_PE_9_7__empty_n),
    .if_read(fifo_B_PE_9_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_9_7__din),
    .if_full_n(fifo_B_PE_9_7__full_n),
    .if_write(fifo_B_PE_9_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_9_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_9_8__dout),
    .if_empty_n(fifo_B_PE_9_8__empty_n),
    .if_read(fifo_B_PE_9_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_9_8__din),
    .if_full_n(fifo_B_PE_9_8__full_n),
    .if_write(fifo_B_PE_9_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(513),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_B_PE_9_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_B_PE_9_9__dout),
    .if_empty_n(fifo_B_PE_9_9__empty_n),
    .if_read(fifo_B_PE_9_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_B_PE_9_9__din),
    .if_full_n(fifo_B_PE_9_9__full_n),
    .if_write(fifo_B_PE_9_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_0_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_0_0__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_0__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_0_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_0_0__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_0_0__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_0_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_0_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_0_1__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_1__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_0_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_0_1__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_0_1__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_0_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_0_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_0_10__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_10__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_0_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_0_10__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_0_10__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_0_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_0_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_0_11__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_11__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_0_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_0_11__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_0_11__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_0_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_0_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_0_12__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_12__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_0_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_0_12__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_0_12__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_0_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_0_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_0_13__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_13__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_0_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_0_13__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_0_13__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_0_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_0_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_0_14__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_14__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_0_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_0_14__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_0_14__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_0_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_0_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_0_15__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_15__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_0_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_0_15__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_0_15__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_0_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_0_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_0_16__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_16__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_0_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_0_16__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_0_16__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_0_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_0_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_0_17__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_17__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_0_17__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_0_17__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_0_17__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_0_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_0_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_0_2__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_2__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_0_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_0_2__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_0_2__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_0_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_0_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_0_3__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_3__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_0_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_0_3__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_0_3__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_0_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_0_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_0_4__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_4__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_0_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_0_4__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_0_4__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_0_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_0_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_0_5__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_5__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_0_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_0_5__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_0_5__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_0_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_0_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_0_6__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_6__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_0_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_0_6__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_0_6__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_0_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_0_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_0_7__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_7__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_0_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_0_7__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_0_7__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_0_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_0_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_0_8__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_8__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_0_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_0_8__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_0_8__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_0_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_0_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_0_9__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_9__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_0_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_0_9__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_0_9__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_0_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_10_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_10_0__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_0__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_10_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_10_0__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_10_0__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_10_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_10_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_10_1__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_1__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_10_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_10_1__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_10_1__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_10_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_10_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_10_10__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_10__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_10_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_10_10__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_10_10__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_10_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_10_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_10_11__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_11__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_10_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_10_11__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_10_11__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_10_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_10_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_10_12__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_12__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_10_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_10_12__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_10_12__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_10_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_10_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_10_13__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_13__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_10_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_10_13__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_10_13__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_10_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_10_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_10_14__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_14__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_10_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_10_14__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_10_14__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_10_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_10_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_10_15__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_15__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_10_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_10_15__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_10_15__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_10_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_10_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_10_16__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_16__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_10_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_10_16__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_10_16__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_10_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_10_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_10_17__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_17__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_10_17__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_10_17__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_10_17__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_10_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_10_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_10_2__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_2__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_10_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_10_2__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_10_2__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_10_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_10_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_10_3__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_3__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_10_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_10_3__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_10_3__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_10_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_10_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_10_4__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_4__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_10_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_10_4__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_10_4__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_10_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_10_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_10_5__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_5__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_10_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_10_5__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_10_5__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_10_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_10_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_10_6__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_6__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_10_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_10_6__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_10_6__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_10_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_10_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_10_7__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_7__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_10_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_10_7__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_10_7__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_10_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_10_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_10_8__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_8__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_10_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_10_8__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_10_8__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_10_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_10_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_10_9__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_9__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_10_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_10_9__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_10_9__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_10_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_11_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_11_0__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_0__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_11_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_11_0__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_11_0__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_11_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_11_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_11_1__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_1__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_11_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_11_1__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_11_1__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_11_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_11_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_11_10__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_10__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_11_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_11_10__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_11_10__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_11_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_11_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_11_11__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_11__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_11_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_11_11__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_11_11__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_11_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_11_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_11_12__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_12__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_11_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_11_12__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_11_12__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_11_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_11_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_11_13__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_13__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_11_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_11_13__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_11_13__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_11_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_11_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_11_14__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_14__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_11_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_11_14__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_11_14__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_11_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_11_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_11_15__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_15__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_11_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_11_15__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_11_15__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_11_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_11_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_11_16__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_16__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_11_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_11_16__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_11_16__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_11_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_11_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_11_17__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_17__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_11_17__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_11_17__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_11_17__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_11_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_11_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_11_2__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_2__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_11_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_11_2__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_11_2__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_11_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_11_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_11_3__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_3__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_11_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_11_3__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_11_3__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_11_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_11_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_11_4__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_4__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_11_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_11_4__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_11_4__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_11_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_11_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_11_5__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_5__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_11_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_11_5__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_11_5__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_11_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_11_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_11_6__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_6__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_11_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_11_6__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_11_6__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_11_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_11_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_11_7__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_7__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_11_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_11_7__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_11_7__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_11_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_11_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_11_8__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_8__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_11_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_11_8__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_11_8__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_11_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_11_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_11_9__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_9__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_11_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_11_9__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_11_9__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_11_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_12_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_12_0__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_0__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_12_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_12_0__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_12_0__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_12_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_12_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_12_1__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_1__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_12_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_12_1__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_12_1__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_12_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_12_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_12_10__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_10__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_12_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_12_10__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_12_10__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_12_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_12_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_12_11__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_11__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_12_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_12_11__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_12_11__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_12_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_12_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_12_12__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_12__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_12_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_12_12__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_12_12__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_12_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_12_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_12_13__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_13__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_12_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_12_13__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_12_13__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_12_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_12_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_12_14__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_14__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_12_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_12_14__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_12_14__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_12_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_12_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_12_15__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_15__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_12_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_12_15__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_12_15__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_12_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_12_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_12_16__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_16__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_12_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_12_16__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_12_16__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_12_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_12_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_12_17__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_17__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_12_17__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_12_17__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_12_17__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_12_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_12_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_12_2__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_2__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_12_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_12_2__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_12_2__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_12_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_12_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_12_3__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_3__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_12_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_12_3__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_12_3__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_12_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_12_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_12_4__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_4__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_12_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_12_4__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_12_4__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_12_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_12_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_12_5__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_5__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_12_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_12_5__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_12_5__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_12_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_12_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_12_6__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_6__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_12_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_12_6__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_12_6__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_12_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_12_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_12_7__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_7__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_12_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_12_7__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_12_7__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_12_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_12_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_12_8__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_8__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_12_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_12_8__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_12_8__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_12_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_12_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_12_9__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_9__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_12_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_12_9__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_12_9__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_12_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_13_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_13_0__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_0__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_13_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_13_0__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_13_0__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_13_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_13_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_13_1__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_1__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_13_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_13_1__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_13_1__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_13_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_13_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_13_10__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_10__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_13_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_13_10__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_13_10__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_13_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_13_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_13_11__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_11__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_13_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_13_11__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_13_11__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_13_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_13_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_13_12__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_12__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_13_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_13_12__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_13_12__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_13_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_13_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_13_13__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_13__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_13_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_13_13__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_13_13__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_13_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_13_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_13_14__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_14__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_13_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_13_14__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_13_14__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_13_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_13_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_13_15__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_15__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_13_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_13_15__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_13_15__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_13_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_13_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_13_16__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_16__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_13_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_13_16__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_13_16__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_13_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_13_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_13_17__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_17__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_13_17__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_13_17__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_13_17__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_13_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_13_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_13_2__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_2__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_13_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_13_2__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_13_2__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_13_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_13_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_13_3__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_3__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_13_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_13_3__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_13_3__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_13_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_13_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_13_4__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_4__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_13_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_13_4__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_13_4__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_13_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_13_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_13_5__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_5__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_13_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_13_5__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_13_5__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_13_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_13_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_13_6__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_6__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_13_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_13_6__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_13_6__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_13_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_13_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_13_7__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_7__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_13_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_13_7__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_13_7__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_13_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_13_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_13_8__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_8__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_13_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_13_8__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_13_8__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_13_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_13_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_13_9__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_9__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_13_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_13_9__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_13_9__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_13_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_14_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_14_0__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_0__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_14_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_14_0__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_14_0__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_14_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_14_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_14_1__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_1__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_14_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_14_1__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_14_1__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_14_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_14_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_14_10__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_10__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_14_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_14_10__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_14_10__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_14_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_14_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_14_11__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_11__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_14_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_14_11__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_14_11__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_14_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_14_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_14_12__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_12__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_14_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_14_12__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_14_12__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_14_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_14_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_14_13__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_13__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_14_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_14_13__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_14_13__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_14_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_14_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_14_14__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_14__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_14_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_14_14__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_14_14__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_14_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_14_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_14_15__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_15__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_14_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_14_15__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_14_15__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_14_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_14_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_14_16__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_16__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_14_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_14_16__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_14_16__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_14_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_14_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_14_17__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_17__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_14_17__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_14_17__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_14_17__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_14_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_14_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_14_2__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_2__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_14_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_14_2__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_14_2__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_14_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_14_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_14_3__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_3__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_14_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_14_3__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_14_3__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_14_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_14_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_14_4__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_4__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_14_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_14_4__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_14_4__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_14_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_14_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_14_5__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_5__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_14_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_14_5__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_14_5__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_14_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_14_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_14_6__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_6__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_14_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_14_6__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_14_6__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_14_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_14_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_14_7__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_7__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_14_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_14_7__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_14_7__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_14_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_14_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_14_8__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_8__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_14_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_14_8__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_14_8__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_14_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_14_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_14_9__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_9__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_14_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_14_9__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_14_9__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_14_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_15_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_15_0__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_0__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_15_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_15_0__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_15_0__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_15_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_15_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_15_1__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_1__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_15_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_15_1__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_15_1__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_15_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_15_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_15_10__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_10__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_15_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_15_10__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_15_10__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_15_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_15_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_15_11__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_11__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_15_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_15_11__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_15_11__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_15_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_15_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_15_12__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_12__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_15_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_15_12__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_15_12__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_15_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_15_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_15_13__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_13__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_15_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_15_13__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_15_13__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_15_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_15_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_15_14__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_14__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_15_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_15_14__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_15_14__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_15_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_15_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_15_15__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_15__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_15_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_15_15__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_15_15__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_15_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_15_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_15_16__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_16__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_15_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_15_16__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_15_16__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_15_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_15_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_15_17__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_17__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_15_17__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_15_17__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_15_17__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_15_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_15_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_15_2__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_2__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_15_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_15_2__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_15_2__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_15_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_15_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_15_3__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_3__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_15_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_15_3__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_15_3__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_15_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_15_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_15_4__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_4__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_15_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_15_4__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_15_4__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_15_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_15_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_15_5__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_5__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_15_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_15_5__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_15_5__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_15_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_15_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_15_6__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_6__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_15_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_15_6__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_15_6__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_15_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_15_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_15_7__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_7__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_15_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_15_7__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_15_7__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_15_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_15_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_15_8__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_8__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_15_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_15_8__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_15_8__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_15_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_15_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_15_9__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_9__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_15_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_15_9__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_15_9__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_15_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_16_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_16_0__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_0__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_16_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_16_0__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_16_0__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_16_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_16_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_16_1__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_1__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_16_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_16_1__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_16_1__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_16_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_16_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_16_10__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_10__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_16_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_16_10__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_16_10__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_16_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_16_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_16_11__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_11__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_16_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_16_11__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_16_11__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_16_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_16_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_16_12__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_12__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_16_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_16_12__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_16_12__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_16_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_16_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_16_13__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_13__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_16_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_16_13__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_16_13__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_16_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_16_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_16_14__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_14__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_16_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_16_14__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_16_14__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_16_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_16_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_16_15__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_15__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_16_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_16_15__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_16_15__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_16_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_16_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_16_16__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_16__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_16_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_16_16__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_16_16__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_16_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_16_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_16_17__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_17__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_16_17__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_16_17__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_16_17__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_16_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_16_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_16_2__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_2__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_16_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_16_2__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_16_2__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_16_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_16_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_16_3__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_3__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_16_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_16_3__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_16_3__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_16_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_16_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_16_4__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_4__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_16_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_16_4__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_16_4__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_16_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_16_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_16_5__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_5__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_16_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_16_5__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_16_5__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_16_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_16_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_16_6__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_6__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_16_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_16_6__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_16_6__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_16_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_16_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_16_7__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_7__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_16_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_16_7__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_16_7__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_16_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_16_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_16_8__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_8__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_16_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_16_8__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_16_8__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_16_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_16_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_16_9__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_9__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_16_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_16_9__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_16_9__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_16_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_1_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_1_0__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_0__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_1_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_1_0__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_1_0__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_1_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_1_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_1_1__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_1__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_1_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_1_1__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_1_1__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_1_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_1_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_1_10__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_10__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_1_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_1_10__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_1_10__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_1_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_1_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_1_11__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_11__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_1_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_1_11__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_1_11__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_1_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_1_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_1_12__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_12__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_1_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_1_12__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_1_12__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_1_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_1_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_1_13__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_13__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_1_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_1_13__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_1_13__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_1_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_1_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_1_14__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_14__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_1_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_1_14__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_1_14__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_1_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_1_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_1_15__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_15__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_1_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_1_15__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_1_15__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_1_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_1_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_1_16__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_16__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_1_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_1_16__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_1_16__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_1_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_1_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_1_17__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_17__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_1_17__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_1_17__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_1_17__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_1_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_1_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_1_2__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_2__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_1_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_1_2__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_1_2__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_1_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_1_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_1_3__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_3__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_1_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_1_3__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_1_3__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_1_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_1_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_1_4__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_4__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_1_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_1_4__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_1_4__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_1_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_1_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_1_5__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_5__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_1_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_1_5__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_1_5__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_1_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_1_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_1_6__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_6__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_1_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_1_6__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_1_6__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_1_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_1_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_1_7__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_7__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_1_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_1_7__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_1_7__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_1_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_1_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_1_8__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_8__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_1_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_1_8__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_1_8__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_1_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_1_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_1_9__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_9__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_1_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_1_9__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_1_9__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_1_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_2_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_2_0__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_0__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_2_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_2_0__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_2_0__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_2_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_2_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_2_1__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_1__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_2_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_2_1__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_2_1__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_2_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_2_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_2_10__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_10__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_2_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_2_10__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_2_10__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_2_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_2_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_2_11__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_11__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_2_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_2_11__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_2_11__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_2_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_2_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_2_12__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_12__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_2_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_2_12__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_2_12__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_2_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_2_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_2_13__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_13__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_2_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_2_13__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_2_13__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_2_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_2_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_2_14__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_14__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_2_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_2_14__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_2_14__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_2_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_2_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_2_15__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_15__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_2_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_2_15__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_2_15__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_2_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_2_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_2_16__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_16__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_2_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_2_16__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_2_16__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_2_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_2_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_2_17__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_17__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_2_17__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_2_17__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_2_17__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_2_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_2_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_2_2__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_2__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_2_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_2_2__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_2_2__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_2_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_2_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_2_3__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_3__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_2_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_2_3__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_2_3__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_2_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_2_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_2_4__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_4__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_2_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_2_4__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_2_4__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_2_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_2_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_2_5__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_5__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_2_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_2_5__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_2_5__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_2_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_2_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_2_6__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_6__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_2_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_2_6__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_2_6__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_2_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_2_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_2_7__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_7__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_2_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_2_7__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_2_7__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_2_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_2_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_2_8__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_8__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_2_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_2_8__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_2_8__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_2_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_2_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_2_9__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_9__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_2_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_2_9__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_2_9__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_2_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_3_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_3_0__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_0__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_3_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_3_0__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_3_0__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_3_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_3_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_3_1__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_1__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_3_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_3_1__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_3_1__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_3_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_3_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_3_10__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_10__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_3_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_3_10__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_3_10__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_3_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_3_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_3_11__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_11__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_3_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_3_11__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_3_11__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_3_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_3_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_3_12__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_12__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_3_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_3_12__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_3_12__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_3_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_3_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_3_13__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_13__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_3_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_3_13__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_3_13__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_3_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_3_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_3_14__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_14__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_3_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_3_14__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_3_14__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_3_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_3_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_3_15__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_15__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_3_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_3_15__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_3_15__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_3_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_3_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_3_16__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_16__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_3_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_3_16__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_3_16__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_3_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_3_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_3_17__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_17__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_3_17__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_3_17__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_3_17__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_3_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_3_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_3_2__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_2__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_3_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_3_2__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_3_2__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_3_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_3_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_3_3__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_3__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_3_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_3_3__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_3_3__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_3_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_3_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_3_4__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_4__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_3_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_3_4__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_3_4__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_3_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_3_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_3_5__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_5__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_3_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_3_5__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_3_5__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_3_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_3_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_3_6__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_6__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_3_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_3_6__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_3_6__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_3_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_3_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_3_7__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_7__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_3_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_3_7__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_3_7__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_3_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_3_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_3_8__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_8__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_3_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_3_8__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_3_8__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_3_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_3_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_3_9__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_9__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_3_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_3_9__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_3_9__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_3_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_4_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_4_0__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_0__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_4_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_4_0__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_4_0__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_4_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_4_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_4_1__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_1__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_4_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_4_1__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_4_1__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_4_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_4_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_4_10__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_10__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_4_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_4_10__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_4_10__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_4_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_4_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_4_11__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_11__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_4_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_4_11__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_4_11__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_4_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_4_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_4_12__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_12__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_4_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_4_12__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_4_12__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_4_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_4_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_4_13__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_13__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_4_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_4_13__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_4_13__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_4_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_4_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_4_14__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_14__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_4_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_4_14__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_4_14__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_4_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_4_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_4_15__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_15__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_4_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_4_15__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_4_15__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_4_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_4_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_4_16__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_16__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_4_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_4_16__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_4_16__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_4_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_4_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_4_17__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_17__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_4_17__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_4_17__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_4_17__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_4_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_4_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_4_2__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_2__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_4_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_4_2__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_4_2__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_4_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_4_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_4_3__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_3__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_4_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_4_3__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_4_3__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_4_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_4_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_4_4__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_4__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_4_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_4_4__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_4_4__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_4_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_4_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_4_5__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_5__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_4_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_4_5__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_4_5__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_4_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_4_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_4_6__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_6__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_4_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_4_6__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_4_6__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_4_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_4_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_4_7__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_7__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_4_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_4_7__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_4_7__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_4_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_4_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_4_8__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_8__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_4_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_4_8__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_4_8__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_4_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_4_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_4_9__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_9__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_4_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_4_9__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_4_9__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_4_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_5_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_5_0__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_0__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_5_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_5_0__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_5_0__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_5_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_5_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_5_1__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_1__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_5_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_5_1__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_5_1__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_5_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_5_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_5_10__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_10__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_5_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_5_10__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_5_10__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_5_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_5_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_5_11__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_11__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_5_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_5_11__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_5_11__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_5_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_5_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_5_12__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_12__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_5_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_5_12__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_5_12__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_5_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_5_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_5_13__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_13__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_5_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_5_13__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_5_13__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_5_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_5_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_5_14__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_14__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_5_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_5_14__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_5_14__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_5_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_5_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_5_15__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_15__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_5_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_5_15__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_5_15__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_5_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_5_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_5_16__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_16__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_5_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_5_16__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_5_16__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_5_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_5_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_5_17__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_17__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_5_17__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_5_17__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_5_17__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_5_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_5_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_5_2__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_2__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_5_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_5_2__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_5_2__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_5_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_5_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_5_3__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_3__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_5_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_5_3__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_5_3__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_5_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_5_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_5_4__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_4__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_5_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_5_4__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_5_4__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_5_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_5_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_5_5__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_5__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_5_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_5_5__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_5_5__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_5_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_5_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_5_6__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_6__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_5_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_5_6__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_5_6__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_5_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_5_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_5_7__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_7__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_5_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_5_7__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_5_7__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_5_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_5_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_5_8__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_8__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_5_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_5_8__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_5_8__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_5_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_5_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_5_9__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_9__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_5_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_5_9__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_5_9__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_5_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_6_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_6_0__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_0__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_6_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_6_0__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_6_0__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_6_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_6_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_6_1__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_1__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_6_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_6_1__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_6_1__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_6_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_6_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_6_10__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_10__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_6_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_6_10__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_6_10__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_6_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_6_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_6_11__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_11__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_6_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_6_11__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_6_11__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_6_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_6_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_6_12__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_12__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_6_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_6_12__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_6_12__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_6_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_6_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_6_13__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_13__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_6_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_6_13__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_6_13__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_6_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_6_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_6_14__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_14__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_6_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_6_14__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_6_14__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_6_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_6_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_6_15__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_15__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_6_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_6_15__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_6_15__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_6_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_6_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_6_16__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_16__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_6_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_6_16__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_6_16__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_6_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_6_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_6_17__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_17__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_6_17__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_6_17__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_6_17__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_6_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_6_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_6_2__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_2__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_6_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_6_2__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_6_2__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_6_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_6_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_6_3__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_3__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_6_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_6_3__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_6_3__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_6_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_6_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_6_4__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_4__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_6_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_6_4__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_6_4__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_6_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_6_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_6_5__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_5__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_6_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_6_5__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_6_5__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_6_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_6_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_6_6__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_6__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_6_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_6_6__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_6_6__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_6_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_6_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_6_7__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_7__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_6_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_6_7__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_6_7__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_6_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_6_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_6_8__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_8__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_6_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_6_8__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_6_8__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_6_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_6_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_6_9__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_9__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_6_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_6_9__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_6_9__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_6_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_7_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_7_0__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_0__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_7_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_7_0__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_7_0__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_7_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_7_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_7_1__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_1__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_7_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_7_1__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_7_1__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_7_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_7_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_7_10__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_10__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_7_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_7_10__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_7_10__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_7_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_7_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_7_11__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_11__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_7_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_7_11__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_7_11__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_7_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_7_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_7_12__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_12__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_7_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_7_12__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_7_12__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_7_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_7_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_7_13__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_13__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_7_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_7_13__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_7_13__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_7_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_7_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_7_14__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_14__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_7_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_7_14__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_7_14__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_7_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_7_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_7_15__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_15__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_7_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_7_15__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_7_15__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_7_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_7_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_7_16__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_16__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_7_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_7_16__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_7_16__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_7_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_7_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_7_17__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_17__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_7_17__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_7_17__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_7_17__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_7_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_7_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_7_2__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_2__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_7_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_7_2__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_7_2__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_7_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_7_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_7_3__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_3__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_7_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_7_3__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_7_3__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_7_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_7_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_7_4__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_4__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_7_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_7_4__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_7_4__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_7_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_7_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_7_5__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_5__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_7_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_7_5__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_7_5__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_7_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_7_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_7_6__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_6__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_7_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_7_6__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_7_6__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_7_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_7_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_7_7__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_7__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_7_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_7_7__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_7_7__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_7_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_7_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_7_8__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_8__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_7_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_7_8__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_7_8__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_7_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_7_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_7_9__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_9__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_7_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_7_9__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_7_9__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_7_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_8_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_8_0__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_0__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_8_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_8_0__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_8_0__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_8_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_8_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_8_1__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_1__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_8_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_8_1__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_8_1__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_8_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_8_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_8_10__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_10__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_8_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_8_10__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_8_10__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_8_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_8_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_8_11__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_11__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_8_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_8_11__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_8_11__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_8_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_8_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_8_12__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_12__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_8_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_8_12__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_8_12__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_8_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_8_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_8_13__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_13__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_8_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_8_13__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_8_13__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_8_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_8_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_8_14__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_14__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_8_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_8_14__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_8_14__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_8_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_8_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_8_15__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_15__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_8_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_8_15__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_8_15__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_8_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_8_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_8_16__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_16__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_8_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_8_16__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_8_16__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_8_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_8_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_8_17__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_17__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_8_17__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_8_17__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_8_17__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_8_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_8_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_8_2__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_2__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_8_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_8_2__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_8_2__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_8_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_8_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_8_3__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_3__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_8_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_8_3__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_8_3__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_8_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_8_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_8_4__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_4__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_8_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_8_4__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_8_4__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_8_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_8_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_8_5__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_5__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_8_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_8_5__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_8_5__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_8_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_8_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_8_6__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_6__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_8_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_8_6__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_8_6__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_8_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_8_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_8_7__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_7__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_8_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_8_7__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_8_7__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_8_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_8_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_8_8__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_8__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_8_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_8_8__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_8_8__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_8_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_8_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_8_9__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_9__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_8_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_8_9__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_8_9__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_8_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_9_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_9_0__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_0__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_9_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_9_0__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_9_0__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_9_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_9_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_9_1__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_1__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_9_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_9_1__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_9_1__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_9_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_9_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_9_10__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_10__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_9_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_9_10__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_9_10__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_9_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_9_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_9_11__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_11__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_9_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_9_11__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_9_11__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_9_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_9_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_9_12__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_12__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_9_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_9_12__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_9_12__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_9_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_9_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_9_13__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_13__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_9_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_9_13__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_9_13__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_9_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_9_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_9_14__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_14__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_9_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_9_14__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_9_14__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_9_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_9_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_9_15__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_15__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_9_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_9_15__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_9_15__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_9_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_9_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_9_16__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_16__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_9_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_9_16__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_9_16__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_9_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_9_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_9_17__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_17__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_9_17__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_9_17__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_9_17__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_9_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_9_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_9_2__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_2__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_9_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_9_2__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_9_2__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_9_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_9_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_9_3__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_3__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_9_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_9_3__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_9_3__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_9_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_9_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_9_4__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_4__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_9_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_9_4__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_9_4__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_9_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_9_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_9_5__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_5__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_9_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_9_5__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_9_5__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_9_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_9_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_9_6__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_6__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_9_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_9_6__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_9_6__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_9_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_9_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_9_7__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_7__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_9_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_9_7__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_9_7__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_9_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_9_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_9_8__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_8__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_9_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_9_8__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_9_8__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_9_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L1_out_9_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L1_out_9_9__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_9__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L1_out_9_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L1_out_9_9__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L1_out_9_9__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L1_out_9_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L2_out_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L2_out_0__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L2_out_0__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L2_out_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L2_out_0__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L2_out_0__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L2_out_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L2_out_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L2_out_1__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L2_out_1__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L2_out_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L2_out_1__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L2_out_1__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L2_out_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L2_out_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L2_out_10__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L2_out_10__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L2_out_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L2_out_10__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L2_out_10__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L2_out_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L2_out_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L2_out_11__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L2_out_11__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L2_out_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L2_out_11__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L2_out_11__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L2_out_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L2_out_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L2_out_12__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L2_out_12__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L2_out_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L2_out_12__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L2_out_12__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L2_out_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L2_out_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L2_out_13__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L2_out_13__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L2_out_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L2_out_13__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L2_out_13__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L2_out_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L2_out_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L2_out_14__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L2_out_14__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L2_out_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L2_out_14__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L2_out_14__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L2_out_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L2_out_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L2_out_15__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L2_out_15__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L2_out_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L2_out_15__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L2_out_15__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L2_out_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L2_out_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L2_out_16__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L2_out_16__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L2_out_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L2_out_16__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L2_out_16__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L2_out_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L2_out_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L2_out_2__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L2_out_2__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L2_out_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L2_out_2__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L2_out_2__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L2_out_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L2_out_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L2_out_3__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L2_out_3__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L2_out_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L2_out_3__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L2_out_3__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L2_out_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L2_out_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L2_out_4__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L2_out_4__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L2_out_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L2_out_4__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L2_out_4__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L2_out_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L2_out_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L2_out_5__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L2_out_5__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L2_out_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L2_out_5__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L2_out_5__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L2_out_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L2_out_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L2_out_6__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L2_out_6__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L2_out_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L2_out_6__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L2_out_6__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L2_out_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L2_out_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L2_out_7__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L2_out_7__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L2_out_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L2_out_7__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L2_out_7__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L2_out_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L2_out_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L2_out_8__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L2_out_8__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L2_out_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L2_out_8__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L2_out_8__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L2_out_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L2_out_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L2_out_9__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L2_out_9__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L2_out_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L2_out_9__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L2_out_9__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L2_out_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(129),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_C_drain_IO_L3_out_serialize
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_C_drain_IO_L3_out_serialize__dout),
    .if_empty_n(fifo_C_drain_C_drain_IO_L3_out_serialize__empty_n),
    .if_read(fifo_C_drain_C_drain_IO_L3_out_serialize__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_C_drain_IO_L3_out_serialize__din),
    .if_full_n(fifo_C_drain_C_drain_IO_L3_out_serialize__full_n),
    .if_write(fifo_C_drain_C_drain_IO_L3_out_serialize__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_0_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_0_0__dout),
    .if_empty_n(fifo_C_drain_PE_0_0__empty_n),
    .if_read(fifo_C_drain_PE_0_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_0_0__din),
    .if_full_n(fifo_C_drain_PE_0_0__full_n),
    .if_write(fifo_C_drain_PE_0_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_0_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_0_1__dout),
    .if_empty_n(fifo_C_drain_PE_0_1__empty_n),
    .if_read(fifo_C_drain_PE_0_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_0_1__din),
    .if_full_n(fifo_C_drain_PE_0_1__full_n),
    .if_write(fifo_C_drain_PE_0_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_0_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_0_10__dout),
    .if_empty_n(fifo_C_drain_PE_0_10__empty_n),
    .if_read(fifo_C_drain_PE_0_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_0_10__din),
    .if_full_n(fifo_C_drain_PE_0_10__full_n),
    .if_write(fifo_C_drain_PE_0_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_0_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_0_11__dout),
    .if_empty_n(fifo_C_drain_PE_0_11__empty_n),
    .if_read(fifo_C_drain_PE_0_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_0_11__din),
    .if_full_n(fifo_C_drain_PE_0_11__full_n),
    .if_write(fifo_C_drain_PE_0_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_0_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_0_12__dout),
    .if_empty_n(fifo_C_drain_PE_0_12__empty_n),
    .if_read(fifo_C_drain_PE_0_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_0_12__din),
    .if_full_n(fifo_C_drain_PE_0_12__full_n),
    .if_write(fifo_C_drain_PE_0_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_0_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_0_13__dout),
    .if_empty_n(fifo_C_drain_PE_0_13__empty_n),
    .if_read(fifo_C_drain_PE_0_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_0_13__din),
    .if_full_n(fifo_C_drain_PE_0_13__full_n),
    .if_write(fifo_C_drain_PE_0_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_0_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_0_14__dout),
    .if_empty_n(fifo_C_drain_PE_0_14__empty_n),
    .if_read(fifo_C_drain_PE_0_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_0_14__din),
    .if_full_n(fifo_C_drain_PE_0_14__full_n),
    .if_write(fifo_C_drain_PE_0_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_0_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_0_15__dout),
    .if_empty_n(fifo_C_drain_PE_0_15__empty_n),
    .if_read(fifo_C_drain_PE_0_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_0_15__din),
    .if_full_n(fifo_C_drain_PE_0_15__full_n),
    .if_write(fifo_C_drain_PE_0_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_0_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_0_16__dout),
    .if_empty_n(fifo_C_drain_PE_0_16__empty_n),
    .if_read(fifo_C_drain_PE_0_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_0_16__din),
    .if_full_n(fifo_C_drain_PE_0_16__full_n),
    .if_write(fifo_C_drain_PE_0_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_0_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_0_2__dout),
    .if_empty_n(fifo_C_drain_PE_0_2__empty_n),
    .if_read(fifo_C_drain_PE_0_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_0_2__din),
    .if_full_n(fifo_C_drain_PE_0_2__full_n),
    .if_write(fifo_C_drain_PE_0_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_0_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_0_3__dout),
    .if_empty_n(fifo_C_drain_PE_0_3__empty_n),
    .if_read(fifo_C_drain_PE_0_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_0_3__din),
    .if_full_n(fifo_C_drain_PE_0_3__full_n),
    .if_write(fifo_C_drain_PE_0_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_0_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_0_4__dout),
    .if_empty_n(fifo_C_drain_PE_0_4__empty_n),
    .if_read(fifo_C_drain_PE_0_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_0_4__din),
    .if_full_n(fifo_C_drain_PE_0_4__full_n),
    .if_write(fifo_C_drain_PE_0_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_0_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_0_5__dout),
    .if_empty_n(fifo_C_drain_PE_0_5__empty_n),
    .if_read(fifo_C_drain_PE_0_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_0_5__din),
    .if_full_n(fifo_C_drain_PE_0_5__full_n),
    .if_write(fifo_C_drain_PE_0_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_0_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_0_6__dout),
    .if_empty_n(fifo_C_drain_PE_0_6__empty_n),
    .if_read(fifo_C_drain_PE_0_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_0_6__din),
    .if_full_n(fifo_C_drain_PE_0_6__full_n),
    .if_write(fifo_C_drain_PE_0_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_0_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_0_7__dout),
    .if_empty_n(fifo_C_drain_PE_0_7__empty_n),
    .if_read(fifo_C_drain_PE_0_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_0_7__din),
    .if_full_n(fifo_C_drain_PE_0_7__full_n),
    .if_write(fifo_C_drain_PE_0_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_0_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_0_8__dout),
    .if_empty_n(fifo_C_drain_PE_0_8__empty_n),
    .if_read(fifo_C_drain_PE_0_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_0_8__din),
    .if_full_n(fifo_C_drain_PE_0_8__full_n),
    .if_write(fifo_C_drain_PE_0_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_0_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_0_9__dout),
    .if_empty_n(fifo_C_drain_PE_0_9__empty_n),
    .if_read(fifo_C_drain_PE_0_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_0_9__din),
    .if_full_n(fifo_C_drain_PE_0_9__full_n),
    .if_write(fifo_C_drain_PE_0_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_10_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_10_0__dout),
    .if_empty_n(fifo_C_drain_PE_10_0__empty_n),
    .if_read(fifo_C_drain_PE_10_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_10_0__din),
    .if_full_n(fifo_C_drain_PE_10_0__full_n),
    .if_write(fifo_C_drain_PE_10_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_10_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_10_1__dout),
    .if_empty_n(fifo_C_drain_PE_10_1__empty_n),
    .if_read(fifo_C_drain_PE_10_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_10_1__din),
    .if_full_n(fifo_C_drain_PE_10_1__full_n),
    .if_write(fifo_C_drain_PE_10_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_10_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_10_10__dout),
    .if_empty_n(fifo_C_drain_PE_10_10__empty_n),
    .if_read(fifo_C_drain_PE_10_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_10_10__din),
    .if_full_n(fifo_C_drain_PE_10_10__full_n),
    .if_write(fifo_C_drain_PE_10_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_10_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_10_11__dout),
    .if_empty_n(fifo_C_drain_PE_10_11__empty_n),
    .if_read(fifo_C_drain_PE_10_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_10_11__din),
    .if_full_n(fifo_C_drain_PE_10_11__full_n),
    .if_write(fifo_C_drain_PE_10_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_10_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_10_12__dout),
    .if_empty_n(fifo_C_drain_PE_10_12__empty_n),
    .if_read(fifo_C_drain_PE_10_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_10_12__din),
    .if_full_n(fifo_C_drain_PE_10_12__full_n),
    .if_write(fifo_C_drain_PE_10_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_10_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_10_13__dout),
    .if_empty_n(fifo_C_drain_PE_10_13__empty_n),
    .if_read(fifo_C_drain_PE_10_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_10_13__din),
    .if_full_n(fifo_C_drain_PE_10_13__full_n),
    .if_write(fifo_C_drain_PE_10_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_10_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_10_14__dout),
    .if_empty_n(fifo_C_drain_PE_10_14__empty_n),
    .if_read(fifo_C_drain_PE_10_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_10_14__din),
    .if_full_n(fifo_C_drain_PE_10_14__full_n),
    .if_write(fifo_C_drain_PE_10_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_10_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_10_15__dout),
    .if_empty_n(fifo_C_drain_PE_10_15__empty_n),
    .if_read(fifo_C_drain_PE_10_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_10_15__din),
    .if_full_n(fifo_C_drain_PE_10_15__full_n),
    .if_write(fifo_C_drain_PE_10_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_10_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_10_16__dout),
    .if_empty_n(fifo_C_drain_PE_10_16__empty_n),
    .if_read(fifo_C_drain_PE_10_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_10_16__din),
    .if_full_n(fifo_C_drain_PE_10_16__full_n),
    .if_write(fifo_C_drain_PE_10_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_10_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_10_2__dout),
    .if_empty_n(fifo_C_drain_PE_10_2__empty_n),
    .if_read(fifo_C_drain_PE_10_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_10_2__din),
    .if_full_n(fifo_C_drain_PE_10_2__full_n),
    .if_write(fifo_C_drain_PE_10_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_10_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_10_3__dout),
    .if_empty_n(fifo_C_drain_PE_10_3__empty_n),
    .if_read(fifo_C_drain_PE_10_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_10_3__din),
    .if_full_n(fifo_C_drain_PE_10_3__full_n),
    .if_write(fifo_C_drain_PE_10_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_10_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_10_4__dout),
    .if_empty_n(fifo_C_drain_PE_10_4__empty_n),
    .if_read(fifo_C_drain_PE_10_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_10_4__din),
    .if_full_n(fifo_C_drain_PE_10_4__full_n),
    .if_write(fifo_C_drain_PE_10_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_10_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_10_5__dout),
    .if_empty_n(fifo_C_drain_PE_10_5__empty_n),
    .if_read(fifo_C_drain_PE_10_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_10_5__din),
    .if_full_n(fifo_C_drain_PE_10_5__full_n),
    .if_write(fifo_C_drain_PE_10_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_10_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_10_6__dout),
    .if_empty_n(fifo_C_drain_PE_10_6__empty_n),
    .if_read(fifo_C_drain_PE_10_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_10_6__din),
    .if_full_n(fifo_C_drain_PE_10_6__full_n),
    .if_write(fifo_C_drain_PE_10_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_10_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_10_7__dout),
    .if_empty_n(fifo_C_drain_PE_10_7__empty_n),
    .if_read(fifo_C_drain_PE_10_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_10_7__din),
    .if_full_n(fifo_C_drain_PE_10_7__full_n),
    .if_write(fifo_C_drain_PE_10_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_10_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_10_8__dout),
    .if_empty_n(fifo_C_drain_PE_10_8__empty_n),
    .if_read(fifo_C_drain_PE_10_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_10_8__din),
    .if_full_n(fifo_C_drain_PE_10_8__full_n),
    .if_write(fifo_C_drain_PE_10_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_10_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_10_9__dout),
    .if_empty_n(fifo_C_drain_PE_10_9__empty_n),
    .if_read(fifo_C_drain_PE_10_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_10_9__din),
    .if_full_n(fifo_C_drain_PE_10_9__full_n),
    .if_write(fifo_C_drain_PE_10_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_11_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_11_0__dout),
    .if_empty_n(fifo_C_drain_PE_11_0__empty_n),
    .if_read(fifo_C_drain_PE_11_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_11_0__din),
    .if_full_n(fifo_C_drain_PE_11_0__full_n),
    .if_write(fifo_C_drain_PE_11_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_11_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_11_1__dout),
    .if_empty_n(fifo_C_drain_PE_11_1__empty_n),
    .if_read(fifo_C_drain_PE_11_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_11_1__din),
    .if_full_n(fifo_C_drain_PE_11_1__full_n),
    .if_write(fifo_C_drain_PE_11_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_11_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_11_10__dout),
    .if_empty_n(fifo_C_drain_PE_11_10__empty_n),
    .if_read(fifo_C_drain_PE_11_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_11_10__din),
    .if_full_n(fifo_C_drain_PE_11_10__full_n),
    .if_write(fifo_C_drain_PE_11_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_11_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_11_11__dout),
    .if_empty_n(fifo_C_drain_PE_11_11__empty_n),
    .if_read(fifo_C_drain_PE_11_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_11_11__din),
    .if_full_n(fifo_C_drain_PE_11_11__full_n),
    .if_write(fifo_C_drain_PE_11_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_11_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_11_12__dout),
    .if_empty_n(fifo_C_drain_PE_11_12__empty_n),
    .if_read(fifo_C_drain_PE_11_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_11_12__din),
    .if_full_n(fifo_C_drain_PE_11_12__full_n),
    .if_write(fifo_C_drain_PE_11_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_11_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_11_13__dout),
    .if_empty_n(fifo_C_drain_PE_11_13__empty_n),
    .if_read(fifo_C_drain_PE_11_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_11_13__din),
    .if_full_n(fifo_C_drain_PE_11_13__full_n),
    .if_write(fifo_C_drain_PE_11_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_11_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_11_14__dout),
    .if_empty_n(fifo_C_drain_PE_11_14__empty_n),
    .if_read(fifo_C_drain_PE_11_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_11_14__din),
    .if_full_n(fifo_C_drain_PE_11_14__full_n),
    .if_write(fifo_C_drain_PE_11_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_11_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_11_15__dout),
    .if_empty_n(fifo_C_drain_PE_11_15__empty_n),
    .if_read(fifo_C_drain_PE_11_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_11_15__din),
    .if_full_n(fifo_C_drain_PE_11_15__full_n),
    .if_write(fifo_C_drain_PE_11_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_11_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_11_16__dout),
    .if_empty_n(fifo_C_drain_PE_11_16__empty_n),
    .if_read(fifo_C_drain_PE_11_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_11_16__din),
    .if_full_n(fifo_C_drain_PE_11_16__full_n),
    .if_write(fifo_C_drain_PE_11_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_11_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_11_2__dout),
    .if_empty_n(fifo_C_drain_PE_11_2__empty_n),
    .if_read(fifo_C_drain_PE_11_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_11_2__din),
    .if_full_n(fifo_C_drain_PE_11_2__full_n),
    .if_write(fifo_C_drain_PE_11_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_11_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_11_3__dout),
    .if_empty_n(fifo_C_drain_PE_11_3__empty_n),
    .if_read(fifo_C_drain_PE_11_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_11_3__din),
    .if_full_n(fifo_C_drain_PE_11_3__full_n),
    .if_write(fifo_C_drain_PE_11_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_11_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_11_4__dout),
    .if_empty_n(fifo_C_drain_PE_11_4__empty_n),
    .if_read(fifo_C_drain_PE_11_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_11_4__din),
    .if_full_n(fifo_C_drain_PE_11_4__full_n),
    .if_write(fifo_C_drain_PE_11_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_11_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_11_5__dout),
    .if_empty_n(fifo_C_drain_PE_11_5__empty_n),
    .if_read(fifo_C_drain_PE_11_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_11_5__din),
    .if_full_n(fifo_C_drain_PE_11_5__full_n),
    .if_write(fifo_C_drain_PE_11_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_11_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_11_6__dout),
    .if_empty_n(fifo_C_drain_PE_11_6__empty_n),
    .if_read(fifo_C_drain_PE_11_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_11_6__din),
    .if_full_n(fifo_C_drain_PE_11_6__full_n),
    .if_write(fifo_C_drain_PE_11_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_11_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_11_7__dout),
    .if_empty_n(fifo_C_drain_PE_11_7__empty_n),
    .if_read(fifo_C_drain_PE_11_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_11_7__din),
    .if_full_n(fifo_C_drain_PE_11_7__full_n),
    .if_write(fifo_C_drain_PE_11_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_11_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_11_8__dout),
    .if_empty_n(fifo_C_drain_PE_11_8__empty_n),
    .if_read(fifo_C_drain_PE_11_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_11_8__din),
    .if_full_n(fifo_C_drain_PE_11_8__full_n),
    .if_write(fifo_C_drain_PE_11_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_11_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_11_9__dout),
    .if_empty_n(fifo_C_drain_PE_11_9__empty_n),
    .if_read(fifo_C_drain_PE_11_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_11_9__din),
    .if_full_n(fifo_C_drain_PE_11_9__full_n),
    .if_write(fifo_C_drain_PE_11_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_12_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_12_0__dout),
    .if_empty_n(fifo_C_drain_PE_12_0__empty_n),
    .if_read(fifo_C_drain_PE_12_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_12_0__din),
    .if_full_n(fifo_C_drain_PE_12_0__full_n),
    .if_write(fifo_C_drain_PE_12_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_12_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_12_1__dout),
    .if_empty_n(fifo_C_drain_PE_12_1__empty_n),
    .if_read(fifo_C_drain_PE_12_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_12_1__din),
    .if_full_n(fifo_C_drain_PE_12_1__full_n),
    .if_write(fifo_C_drain_PE_12_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_12_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_12_10__dout),
    .if_empty_n(fifo_C_drain_PE_12_10__empty_n),
    .if_read(fifo_C_drain_PE_12_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_12_10__din),
    .if_full_n(fifo_C_drain_PE_12_10__full_n),
    .if_write(fifo_C_drain_PE_12_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_12_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_12_11__dout),
    .if_empty_n(fifo_C_drain_PE_12_11__empty_n),
    .if_read(fifo_C_drain_PE_12_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_12_11__din),
    .if_full_n(fifo_C_drain_PE_12_11__full_n),
    .if_write(fifo_C_drain_PE_12_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_12_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_12_12__dout),
    .if_empty_n(fifo_C_drain_PE_12_12__empty_n),
    .if_read(fifo_C_drain_PE_12_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_12_12__din),
    .if_full_n(fifo_C_drain_PE_12_12__full_n),
    .if_write(fifo_C_drain_PE_12_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_12_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_12_13__dout),
    .if_empty_n(fifo_C_drain_PE_12_13__empty_n),
    .if_read(fifo_C_drain_PE_12_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_12_13__din),
    .if_full_n(fifo_C_drain_PE_12_13__full_n),
    .if_write(fifo_C_drain_PE_12_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_12_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_12_14__dout),
    .if_empty_n(fifo_C_drain_PE_12_14__empty_n),
    .if_read(fifo_C_drain_PE_12_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_12_14__din),
    .if_full_n(fifo_C_drain_PE_12_14__full_n),
    .if_write(fifo_C_drain_PE_12_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_12_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_12_15__dout),
    .if_empty_n(fifo_C_drain_PE_12_15__empty_n),
    .if_read(fifo_C_drain_PE_12_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_12_15__din),
    .if_full_n(fifo_C_drain_PE_12_15__full_n),
    .if_write(fifo_C_drain_PE_12_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_12_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_12_16__dout),
    .if_empty_n(fifo_C_drain_PE_12_16__empty_n),
    .if_read(fifo_C_drain_PE_12_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_12_16__din),
    .if_full_n(fifo_C_drain_PE_12_16__full_n),
    .if_write(fifo_C_drain_PE_12_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_12_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_12_2__dout),
    .if_empty_n(fifo_C_drain_PE_12_2__empty_n),
    .if_read(fifo_C_drain_PE_12_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_12_2__din),
    .if_full_n(fifo_C_drain_PE_12_2__full_n),
    .if_write(fifo_C_drain_PE_12_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_12_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_12_3__dout),
    .if_empty_n(fifo_C_drain_PE_12_3__empty_n),
    .if_read(fifo_C_drain_PE_12_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_12_3__din),
    .if_full_n(fifo_C_drain_PE_12_3__full_n),
    .if_write(fifo_C_drain_PE_12_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_12_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_12_4__dout),
    .if_empty_n(fifo_C_drain_PE_12_4__empty_n),
    .if_read(fifo_C_drain_PE_12_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_12_4__din),
    .if_full_n(fifo_C_drain_PE_12_4__full_n),
    .if_write(fifo_C_drain_PE_12_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_12_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_12_5__dout),
    .if_empty_n(fifo_C_drain_PE_12_5__empty_n),
    .if_read(fifo_C_drain_PE_12_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_12_5__din),
    .if_full_n(fifo_C_drain_PE_12_5__full_n),
    .if_write(fifo_C_drain_PE_12_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_12_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_12_6__dout),
    .if_empty_n(fifo_C_drain_PE_12_6__empty_n),
    .if_read(fifo_C_drain_PE_12_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_12_6__din),
    .if_full_n(fifo_C_drain_PE_12_6__full_n),
    .if_write(fifo_C_drain_PE_12_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_12_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_12_7__dout),
    .if_empty_n(fifo_C_drain_PE_12_7__empty_n),
    .if_read(fifo_C_drain_PE_12_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_12_7__din),
    .if_full_n(fifo_C_drain_PE_12_7__full_n),
    .if_write(fifo_C_drain_PE_12_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_12_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_12_8__dout),
    .if_empty_n(fifo_C_drain_PE_12_8__empty_n),
    .if_read(fifo_C_drain_PE_12_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_12_8__din),
    .if_full_n(fifo_C_drain_PE_12_8__full_n),
    .if_write(fifo_C_drain_PE_12_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_12_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_12_9__dout),
    .if_empty_n(fifo_C_drain_PE_12_9__empty_n),
    .if_read(fifo_C_drain_PE_12_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_12_9__din),
    .if_full_n(fifo_C_drain_PE_12_9__full_n),
    .if_write(fifo_C_drain_PE_12_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_13_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_13_0__dout),
    .if_empty_n(fifo_C_drain_PE_13_0__empty_n),
    .if_read(fifo_C_drain_PE_13_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_13_0__din),
    .if_full_n(fifo_C_drain_PE_13_0__full_n),
    .if_write(fifo_C_drain_PE_13_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_13_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_13_1__dout),
    .if_empty_n(fifo_C_drain_PE_13_1__empty_n),
    .if_read(fifo_C_drain_PE_13_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_13_1__din),
    .if_full_n(fifo_C_drain_PE_13_1__full_n),
    .if_write(fifo_C_drain_PE_13_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_13_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_13_10__dout),
    .if_empty_n(fifo_C_drain_PE_13_10__empty_n),
    .if_read(fifo_C_drain_PE_13_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_13_10__din),
    .if_full_n(fifo_C_drain_PE_13_10__full_n),
    .if_write(fifo_C_drain_PE_13_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_13_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_13_11__dout),
    .if_empty_n(fifo_C_drain_PE_13_11__empty_n),
    .if_read(fifo_C_drain_PE_13_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_13_11__din),
    .if_full_n(fifo_C_drain_PE_13_11__full_n),
    .if_write(fifo_C_drain_PE_13_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_13_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_13_12__dout),
    .if_empty_n(fifo_C_drain_PE_13_12__empty_n),
    .if_read(fifo_C_drain_PE_13_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_13_12__din),
    .if_full_n(fifo_C_drain_PE_13_12__full_n),
    .if_write(fifo_C_drain_PE_13_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_13_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_13_13__dout),
    .if_empty_n(fifo_C_drain_PE_13_13__empty_n),
    .if_read(fifo_C_drain_PE_13_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_13_13__din),
    .if_full_n(fifo_C_drain_PE_13_13__full_n),
    .if_write(fifo_C_drain_PE_13_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_13_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_13_14__dout),
    .if_empty_n(fifo_C_drain_PE_13_14__empty_n),
    .if_read(fifo_C_drain_PE_13_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_13_14__din),
    .if_full_n(fifo_C_drain_PE_13_14__full_n),
    .if_write(fifo_C_drain_PE_13_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_13_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_13_15__dout),
    .if_empty_n(fifo_C_drain_PE_13_15__empty_n),
    .if_read(fifo_C_drain_PE_13_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_13_15__din),
    .if_full_n(fifo_C_drain_PE_13_15__full_n),
    .if_write(fifo_C_drain_PE_13_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_13_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_13_16__dout),
    .if_empty_n(fifo_C_drain_PE_13_16__empty_n),
    .if_read(fifo_C_drain_PE_13_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_13_16__din),
    .if_full_n(fifo_C_drain_PE_13_16__full_n),
    .if_write(fifo_C_drain_PE_13_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_13_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_13_2__dout),
    .if_empty_n(fifo_C_drain_PE_13_2__empty_n),
    .if_read(fifo_C_drain_PE_13_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_13_2__din),
    .if_full_n(fifo_C_drain_PE_13_2__full_n),
    .if_write(fifo_C_drain_PE_13_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_13_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_13_3__dout),
    .if_empty_n(fifo_C_drain_PE_13_3__empty_n),
    .if_read(fifo_C_drain_PE_13_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_13_3__din),
    .if_full_n(fifo_C_drain_PE_13_3__full_n),
    .if_write(fifo_C_drain_PE_13_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_13_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_13_4__dout),
    .if_empty_n(fifo_C_drain_PE_13_4__empty_n),
    .if_read(fifo_C_drain_PE_13_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_13_4__din),
    .if_full_n(fifo_C_drain_PE_13_4__full_n),
    .if_write(fifo_C_drain_PE_13_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_13_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_13_5__dout),
    .if_empty_n(fifo_C_drain_PE_13_5__empty_n),
    .if_read(fifo_C_drain_PE_13_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_13_5__din),
    .if_full_n(fifo_C_drain_PE_13_5__full_n),
    .if_write(fifo_C_drain_PE_13_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_13_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_13_6__dout),
    .if_empty_n(fifo_C_drain_PE_13_6__empty_n),
    .if_read(fifo_C_drain_PE_13_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_13_6__din),
    .if_full_n(fifo_C_drain_PE_13_6__full_n),
    .if_write(fifo_C_drain_PE_13_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_13_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_13_7__dout),
    .if_empty_n(fifo_C_drain_PE_13_7__empty_n),
    .if_read(fifo_C_drain_PE_13_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_13_7__din),
    .if_full_n(fifo_C_drain_PE_13_7__full_n),
    .if_write(fifo_C_drain_PE_13_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_13_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_13_8__dout),
    .if_empty_n(fifo_C_drain_PE_13_8__empty_n),
    .if_read(fifo_C_drain_PE_13_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_13_8__din),
    .if_full_n(fifo_C_drain_PE_13_8__full_n),
    .if_write(fifo_C_drain_PE_13_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_13_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_13_9__dout),
    .if_empty_n(fifo_C_drain_PE_13_9__empty_n),
    .if_read(fifo_C_drain_PE_13_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_13_9__din),
    .if_full_n(fifo_C_drain_PE_13_9__full_n),
    .if_write(fifo_C_drain_PE_13_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_14_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_14_0__dout),
    .if_empty_n(fifo_C_drain_PE_14_0__empty_n),
    .if_read(fifo_C_drain_PE_14_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_14_0__din),
    .if_full_n(fifo_C_drain_PE_14_0__full_n),
    .if_write(fifo_C_drain_PE_14_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_14_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_14_1__dout),
    .if_empty_n(fifo_C_drain_PE_14_1__empty_n),
    .if_read(fifo_C_drain_PE_14_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_14_1__din),
    .if_full_n(fifo_C_drain_PE_14_1__full_n),
    .if_write(fifo_C_drain_PE_14_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_14_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_14_10__dout),
    .if_empty_n(fifo_C_drain_PE_14_10__empty_n),
    .if_read(fifo_C_drain_PE_14_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_14_10__din),
    .if_full_n(fifo_C_drain_PE_14_10__full_n),
    .if_write(fifo_C_drain_PE_14_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_14_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_14_11__dout),
    .if_empty_n(fifo_C_drain_PE_14_11__empty_n),
    .if_read(fifo_C_drain_PE_14_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_14_11__din),
    .if_full_n(fifo_C_drain_PE_14_11__full_n),
    .if_write(fifo_C_drain_PE_14_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_14_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_14_12__dout),
    .if_empty_n(fifo_C_drain_PE_14_12__empty_n),
    .if_read(fifo_C_drain_PE_14_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_14_12__din),
    .if_full_n(fifo_C_drain_PE_14_12__full_n),
    .if_write(fifo_C_drain_PE_14_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_14_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_14_13__dout),
    .if_empty_n(fifo_C_drain_PE_14_13__empty_n),
    .if_read(fifo_C_drain_PE_14_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_14_13__din),
    .if_full_n(fifo_C_drain_PE_14_13__full_n),
    .if_write(fifo_C_drain_PE_14_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_14_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_14_14__dout),
    .if_empty_n(fifo_C_drain_PE_14_14__empty_n),
    .if_read(fifo_C_drain_PE_14_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_14_14__din),
    .if_full_n(fifo_C_drain_PE_14_14__full_n),
    .if_write(fifo_C_drain_PE_14_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_14_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_14_15__dout),
    .if_empty_n(fifo_C_drain_PE_14_15__empty_n),
    .if_read(fifo_C_drain_PE_14_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_14_15__din),
    .if_full_n(fifo_C_drain_PE_14_15__full_n),
    .if_write(fifo_C_drain_PE_14_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_14_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_14_16__dout),
    .if_empty_n(fifo_C_drain_PE_14_16__empty_n),
    .if_read(fifo_C_drain_PE_14_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_14_16__din),
    .if_full_n(fifo_C_drain_PE_14_16__full_n),
    .if_write(fifo_C_drain_PE_14_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_14_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_14_2__dout),
    .if_empty_n(fifo_C_drain_PE_14_2__empty_n),
    .if_read(fifo_C_drain_PE_14_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_14_2__din),
    .if_full_n(fifo_C_drain_PE_14_2__full_n),
    .if_write(fifo_C_drain_PE_14_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_14_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_14_3__dout),
    .if_empty_n(fifo_C_drain_PE_14_3__empty_n),
    .if_read(fifo_C_drain_PE_14_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_14_3__din),
    .if_full_n(fifo_C_drain_PE_14_3__full_n),
    .if_write(fifo_C_drain_PE_14_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_14_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_14_4__dout),
    .if_empty_n(fifo_C_drain_PE_14_4__empty_n),
    .if_read(fifo_C_drain_PE_14_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_14_4__din),
    .if_full_n(fifo_C_drain_PE_14_4__full_n),
    .if_write(fifo_C_drain_PE_14_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_14_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_14_5__dout),
    .if_empty_n(fifo_C_drain_PE_14_5__empty_n),
    .if_read(fifo_C_drain_PE_14_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_14_5__din),
    .if_full_n(fifo_C_drain_PE_14_5__full_n),
    .if_write(fifo_C_drain_PE_14_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_14_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_14_6__dout),
    .if_empty_n(fifo_C_drain_PE_14_6__empty_n),
    .if_read(fifo_C_drain_PE_14_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_14_6__din),
    .if_full_n(fifo_C_drain_PE_14_6__full_n),
    .if_write(fifo_C_drain_PE_14_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_14_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_14_7__dout),
    .if_empty_n(fifo_C_drain_PE_14_7__empty_n),
    .if_read(fifo_C_drain_PE_14_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_14_7__din),
    .if_full_n(fifo_C_drain_PE_14_7__full_n),
    .if_write(fifo_C_drain_PE_14_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_14_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_14_8__dout),
    .if_empty_n(fifo_C_drain_PE_14_8__empty_n),
    .if_read(fifo_C_drain_PE_14_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_14_8__din),
    .if_full_n(fifo_C_drain_PE_14_8__full_n),
    .if_write(fifo_C_drain_PE_14_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_14_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_14_9__dout),
    .if_empty_n(fifo_C_drain_PE_14_9__empty_n),
    .if_read(fifo_C_drain_PE_14_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_14_9__din),
    .if_full_n(fifo_C_drain_PE_14_9__full_n),
    .if_write(fifo_C_drain_PE_14_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_15_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_15_0__dout),
    .if_empty_n(fifo_C_drain_PE_15_0__empty_n),
    .if_read(fifo_C_drain_PE_15_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_15_0__din),
    .if_full_n(fifo_C_drain_PE_15_0__full_n),
    .if_write(fifo_C_drain_PE_15_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_15_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_15_1__dout),
    .if_empty_n(fifo_C_drain_PE_15_1__empty_n),
    .if_read(fifo_C_drain_PE_15_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_15_1__din),
    .if_full_n(fifo_C_drain_PE_15_1__full_n),
    .if_write(fifo_C_drain_PE_15_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_15_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_15_10__dout),
    .if_empty_n(fifo_C_drain_PE_15_10__empty_n),
    .if_read(fifo_C_drain_PE_15_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_15_10__din),
    .if_full_n(fifo_C_drain_PE_15_10__full_n),
    .if_write(fifo_C_drain_PE_15_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_15_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_15_11__dout),
    .if_empty_n(fifo_C_drain_PE_15_11__empty_n),
    .if_read(fifo_C_drain_PE_15_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_15_11__din),
    .if_full_n(fifo_C_drain_PE_15_11__full_n),
    .if_write(fifo_C_drain_PE_15_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_15_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_15_12__dout),
    .if_empty_n(fifo_C_drain_PE_15_12__empty_n),
    .if_read(fifo_C_drain_PE_15_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_15_12__din),
    .if_full_n(fifo_C_drain_PE_15_12__full_n),
    .if_write(fifo_C_drain_PE_15_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_15_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_15_13__dout),
    .if_empty_n(fifo_C_drain_PE_15_13__empty_n),
    .if_read(fifo_C_drain_PE_15_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_15_13__din),
    .if_full_n(fifo_C_drain_PE_15_13__full_n),
    .if_write(fifo_C_drain_PE_15_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_15_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_15_14__dout),
    .if_empty_n(fifo_C_drain_PE_15_14__empty_n),
    .if_read(fifo_C_drain_PE_15_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_15_14__din),
    .if_full_n(fifo_C_drain_PE_15_14__full_n),
    .if_write(fifo_C_drain_PE_15_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_15_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_15_15__dout),
    .if_empty_n(fifo_C_drain_PE_15_15__empty_n),
    .if_read(fifo_C_drain_PE_15_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_15_15__din),
    .if_full_n(fifo_C_drain_PE_15_15__full_n),
    .if_write(fifo_C_drain_PE_15_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_15_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_15_16__dout),
    .if_empty_n(fifo_C_drain_PE_15_16__empty_n),
    .if_read(fifo_C_drain_PE_15_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_15_16__din),
    .if_full_n(fifo_C_drain_PE_15_16__full_n),
    .if_write(fifo_C_drain_PE_15_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_15_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_15_2__dout),
    .if_empty_n(fifo_C_drain_PE_15_2__empty_n),
    .if_read(fifo_C_drain_PE_15_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_15_2__din),
    .if_full_n(fifo_C_drain_PE_15_2__full_n),
    .if_write(fifo_C_drain_PE_15_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_15_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_15_3__dout),
    .if_empty_n(fifo_C_drain_PE_15_3__empty_n),
    .if_read(fifo_C_drain_PE_15_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_15_3__din),
    .if_full_n(fifo_C_drain_PE_15_3__full_n),
    .if_write(fifo_C_drain_PE_15_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_15_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_15_4__dout),
    .if_empty_n(fifo_C_drain_PE_15_4__empty_n),
    .if_read(fifo_C_drain_PE_15_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_15_4__din),
    .if_full_n(fifo_C_drain_PE_15_4__full_n),
    .if_write(fifo_C_drain_PE_15_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_15_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_15_5__dout),
    .if_empty_n(fifo_C_drain_PE_15_5__empty_n),
    .if_read(fifo_C_drain_PE_15_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_15_5__din),
    .if_full_n(fifo_C_drain_PE_15_5__full_n),
    .if_write(fifo_C_drain_PE_15_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_15_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_15_6__dout),
    .if_empty_n(fifo_C_drain_PE_15_6__empty_n),
    .if_read(fifo_C_drain_PE_15_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_15_6__din),
    .if_full_n(fifo_C_drain_PE_15_6__full_n),
    .if_write(fifo_C_drain_PE_15_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_15_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_15_7__dout),
    .if_empty_n(fifo_C_drain_PE_15_7__empty_n),
    .if_read(fifo_C_drain_PE_15_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_15_7__din),
    .if_full_n(fifo_C_drain_PE_15_7__full_n),
    .if_write(fifo_C_drain_PE_15_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_15_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_15_8__dout),
    .if_empty_n(fifo_C_drain_PE_15_8__empty_n),
    .if_read(fifo_C_drain_PE_15_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_15_8__din),
    .if_full_n(fifo_C_drain_PE_15_8__full_n),
    .if_write(fifo_C_drain_PE_15_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_15_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_15_9__dout),
    .if_empty_n(fifo_C_drain_PE_15_9__empty_n),
    .if_read(fifo_C_drain_PE_15_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_15_9__din),
    .if_full_n(fifo_C_drain_PE_15_9__full_n),
    .if_write(fifo_C_drain_PE_15_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_16_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_16_0__dout),
    .if_empty_n(fifo_C_drain_PE_16_0__empty_n),
    .if_read(fifo_C_drain_PE_16_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_16_0__din),
    .if_full_n(fifo_C_drain_PE_16_0__full_n),
    .if_write(fifo_C_drain_PE_16_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_16_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_16_1__dout),
    .if_empty_n(fifo_C_drain_PE_16_1__empty_n),
    .if_read(fifo_C_drain_PE_16_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_16_1__din),
    .if_full_n(fifo_C_drain_PE_16_1__full_n),
    .if_write(fifo_C_drain_PE_16_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_16_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_16_10__dout),
    .if_empty_n(fifo_C_drain_PE_16_10__empty_n),
    .if_read(fifo_C_drain_PE_16_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_16_10__din),
    .if_full_n(fifo_C_drain_PE_16_10__full_n),
    .if_write(fifo_C_drain_PE_16_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_16_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_16_11__dout),
    .if_empty_n(fifo_C_drain_PE_16_11__empty_n),
    .if_read(fifo_C_drain_PE_16_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_16_11__din),
    .if_full_n(fifo_C_drain_PE_16_11__full_n),
    .if_write(fifo_C_drain_PE_16_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_16_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_16_12__dout),
    .if_empty_n(fifo_C_drain_PE_16_12__empty_n),
    .if_read(fifo_C_drain_PE_16_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_16_12__din),
    .if_full_n(fifo_C_drain_PE_16_12__full_n),
    .if_write(fifo_C_drain_PE_16_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_16_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_16_13__dout),
    .if_empty_n(fifo_C_drain_PE_16_13__empty_n),
    .if_read(fifo_C_drain_PE_16_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_16_13__din),
    .if_full_n(fifo_C_drain_PE_16_13__full_n),
    .if_write(fifo_C_drain_PE_16_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_16_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_16_14__dout),
    .if_empty_n(fifo_C_drain_PE_16_14__empty_n),
    .if_read(fifo_C_drain_PE_16_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_16_14__din),
    .if_full_n(fifo_C_drain_PE_16_14__full_n),
    .if_write(fifo_C_drain_PE_16_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_16_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_16_15__dout),
    .if_empty_n(fifo_C_drain_PE_16_15__empty_n),
    .if_read(fifo_C_drain_PE_16_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_16_15__din),
    .if_full_n(fifo_C_drain_PE_16_15__full_n),
    .if_write(fifo_C_drain_PE_16_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_16_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_16_16__dout),
    .if_empty_n(fifo_C_drain_PE_16_16__empty_n),
    .if_read(fifo_C_drain_PE_16_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_16_16__din),
    .if_full_n(fifo_C_drain_PE_16_16__full_n),
    .if_write(fifo_C_drain_PE_16_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_16_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_16_2__dout),
    .if_empty_n(fifo_C_drain_PE_16_2__empty_n),
    .if_read(fifo_C_drain_PE_16_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_16_2__din),
    .if_full_n(fifo_C_drain_PE_16_2__full_n),
    .if_write(fifo_C_drain_PE_16_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_16_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_16_3__dout),
    .if_empty_n(fifo_C_drain_PE_16_3__empty_n),
    .if_read(fifo_C_drain_PE_16_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_16_3__din),
    .if_full_n(fifo_C_drain_PE_16_3__full_n),
    .if_write(fifo_C_drain_PE_16_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_16_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_16_4__dout),
    .if_empty_n(fifo_C_drain_PE_16_4__empty_n),
    .if_read(fifo_C_drain_PE_16_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_16_4__din),
    .if_full_n(fifo_C_drain_PE_16_4__full_n),
    .if_write(fifo_C_drain_PE_16_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_16_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_16_5__dout),
    .if_empty_n(fifo_C_drain_PE_16_5__empty_n),
    .if_read(fifo_C_drain_PE_16_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_16_5__din),
    .if_full_n(fifo_C_drain_PE_16_5__full_n),
    .if_write(fifo_C_drain_PE_16_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_16_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_16_6__dout),
    .if_empty_n(fifo_C_drain_PE_16_6__empty_n),
    .if_read(fifo_C_drain_PE_16_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_16_6__din),
    .if_full_n(fifo_C_drain_PE_16_6__full_n),
    .if_write(fifo_C_drain_PE_16_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_16_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_16_7__dout),
    .if_empty_n(fifo_C_drain_PE_16_7__empty_n),
    .if_read(fifo_C_drain_PE_16_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_16_7__din),
    .if_full_n(fifo_C_drain_PE_16_7__full_n),
    .if_write(fifo_C_drain_PE_16_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_16_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_16_8__dout),
    .if_empty_n(fifo_C_drain_PE_16_8__empty_n),
    .if_read(fifo_C_drain_PE_16_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_16_8__din),
    .if_full_n(fifo_C_drain_PE_16_8__full_n),
    .if_write(fifo_C_drain_PE_16_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_16_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_16_9__dout),
    .if_empty_n(fifo_C_drain_PE_16_9__empty_n),
    .if_read(fifo_C_drain_PE_16_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_16_9__din),
    .if_full_n(fifo_C_drain_PE_16_9__full_n),
    .if_write(fifo_C_drain_PE_16_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_17_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_17_0__dout),
    .if_empty_n(fifo_C_drain_PE_17_0__empty_n),
    .if_read(fifo_C_drain_PE_17_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_17_0__din),
    .if_full_n(fifo_C_drain_PE_17_0__full_n),
    .if_write(fifo_C_drain_PE_17_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_17_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_17_1__dout),
    .if_empty_n(fifo_C_drain_PE_17_1__empty_n),
    .if_read(fifo_C_drain_PE_17_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_17_1__din),
    .if_full_n(fifo_C_drain_PE_17_1__full_n),
    .if_write(fifo_C_drain_PE_17_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_17_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_17_10__dout),
    .if_empty_n(fifo_C_drain_PE_17_10__empty_n),
    .if_read(fifo_C_drain_PE_17_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_17_10__din),
    .if_full_n(fifo_C_drain_PE_17_10__full_n),
    .if_write(fifo_C_drain_PE_17_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_17_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_17_11__dout),
    .if_empty_n(fifo_C_drain_PE_17_11__empty_n),
    .if_read(fifo_C_drain_PE_17_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_17_11__din),
    .if_full_n(fifo_C_drain_PE_17_11__full_n),
    .if_write(fifo_C_drain_PE_17_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_17_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_17_12__dout),
    .if_empty_n(fifo_C_drain_PE_17_12__empty_n),
    .if_read(fifo_C_drain_PE_17_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_17_12__din),
    .if_full_n(fifo_C_drain_PE_17_12__full_n),
    .if_write(fifo_C_drain_PE_17_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_17_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_17_13__dout),
    .if_empty_n(fifo_C_drain_PE_17_13__empty_n),
    .if_read(fifo_C_drain_PE_17_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_17_13__din),
    .if_full_n(fifo_C_drain_PE_17_13__full_n),
    .if_write(fifo_C_drain_PE_17_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_17_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_17_14__dout),
    .if_empty_n(fifo_C_drain_PE_17_14__empty_n),
    .if_read(fifo_C_drain_PE_17_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_17_14__din),
    .if_full_n(fifo_C_drain_PE_17_14__full_n),
    .if_write(fifo_C_drain_PE_17_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_17_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_17_15__dout),
    .if_empty_n(fifo_C_drain_PE_17_15__empty_n),
    .if_read(fifo_C_drain_PE_17_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_17_15__din),
    .if_full_n(fifo_C_drain_PE_17_15__full_n),
    .if_write(fifo_C_drain_PE_17_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_17_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_17_16__dout),
    .if_empty_n(fifo_C_drain_PE_17_16__empty_n),
    .if_read(fifo_C_drain_PE_17_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_17_16__din),
    .if_full_n(fifo_C_drain_PE_17_16__full_n),
    .if_write(fifo_C_drain_PE_17_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_17_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_17_2__dout),
    .if_empty_n(fifo_C_drain_PE_17_2__empty_n),
    .if_read(fifo_C_drain_PE_17_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_17_2__din),
    .if_full_n(fifo_C_drain_PE_17_2__full_n),
    .if_write(fifo_C_drain_PE_17_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_17_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_17_3__dout),
    .if_empty_n(fifo_C_drain_PE_17_3__empty_n),
    .if_read(fifo_C_drain_PE_17_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_17_3__din),
    .if_full_n(fifo_C_drain_PE_17_3__full_n),
    .if_write(fifo_C_drain_PE_17_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_17_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_17_4__dout),
    .if_empty_n(fifo_C_drain_PE_17_4__empty_n),
    .if_read(fifo_C_drain_PE_17_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_17_4__din),
    .if_full_n(fifo_C_drain_PE_17_4__full_n),
    .if_write(fifo_C_drain_PE_17_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_17_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_17_5__dout),
    .if_empty_n(fifo_C_drain_PE_17_5__empty_n),
    .if_read(fifo_C_drain_PE_17_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_17_5__din),
    .if_full_n(fifo_C_drain_PE_17_5__full_n),
    .if_write(fifo_C_drain_PE_17_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_17_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_17_6__dout),
    .if_empty_n(fifo_C_drain_PE_17_6__empty_n),
    .if_read(fifo_C_drain_PE_17_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_17_6__din),
    .if_full_n(fifo_C_drain_PE_17_6__full_n),
    .if_write(fifo_C_drain_PE_17_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_17_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_17_7__dout),
    .if_empty_n(fifo_C_drain_PE_17_7__empty_n),
    .if_read(fifo_C_drain_PE_17_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_17_7__din),
    .if_full_n(fifo_C_drain_PE_17_7__full_n),
    .if_write(fifo_C_drain_PE_17_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_17_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_17_8__dout),
    .if_empty_n(fifo_C_drain_PE_17_8__empty_n),
    .if_read(fifo_C_drain_PE_17_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_17_8__din),
    .if_full_n(fifo_C_drain_PE_17_8__full_n),
    .if_write(fifo_C_drain_PE_17_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_17_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_17_9__dout),
    .if_empty_n(fifo_C_drain_PE_17_9__empty_n),
    .if_read(fifo_C_drain_PE_17_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_17_9__din),
    .if_full_n(fifo_C_drain_PE_17_9__full_n),
    .if_write(fifo_C_drain_PE_17_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_1_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_1_0__dout),
    .if_empty_n(fifo_C_drain_PE_1_0__empty_n),
    .if_read(fifo_C_drain_PE_1_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_1_0__din),
    .if_full_n(fifo_C_drain_PE_1_0__full_n),
    .if_write(fifo_C_drain_PE_1_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_1_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_1_1__dout),
    .if_empty_n(fifo_C_drain_PE_1_1__empty_n),
    .if_read(fifo_C_drain_PE_1_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_1_1__din),
    .if_full_n(fifo_C_drain_PE_1_1__full_n),
    .if_write(fifo_C_drain_PE_1_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_1_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_1_10__dout),
    .if_empty_n(fifo_C_drain_PE_1_10__empty_n),
    .if_read(fifo_C_drain_PE_1_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_1_10__din),
    .if_full_n(fifo_C_drain_PE_1_10__full_n),
    .if_write(fifo_C_drain_PE_1_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_1_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_1_11__dout),
    .if_empty_n(fifo_C_drain_PE_1_11__empty_n),
    .if_read(fifo_C_drain_PE_1_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_1_11__din),
    .if_full_n(fifo_C_drain_PE_1_11__full_n),
    .if_write(fifo_C_drain_PE_1_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_1_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_1_12__dout),
    .if_empty_n(fifo_C_drain_PE_1_12__empty_n),
    .if_read(fifo_C_drain_PE_1_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_1_12__din),
    .if_full_n(fifo_C_drain_PE_1_12__full_n),
    .if_write(fifo_C_drain_PE_1_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_1_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_1_13__dout),
    .if_empty_n(fifo_C_drain_PE_1_13__empty_n),
    .if_read(fifo_C_drain_PE_1_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_1_13__din),
    .if_full_n(fifo_C_drain_PE_1_13__full_n),
    .if_write(fifo_C_drain_PE_1_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_1_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_1_14__dout),
    .if_empty_n(fifo_C_drain_PE_1_14__empty_n),
    .if_read(fifo_C_drain_PE_1_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_1_14__din),
    .if_full_n(fifo_C_drain_PE_1_14__full_n),
    .if_write(fifo_C_drain_PE_1_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_1_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_1_15__dout),
    .if_empty_n(fifo_C_drain_PE_1_15__empty_n),
    .if_read(fifo_C_drain_PE_1_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_1_15__din),
    .if_full_n(fifo_C_drain_PE_1_15__full_n),
    .if_write(fifo_C_drain_PE_1_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_1_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_1_16__dout),
    .if_empty_n(fifo_C_drain_PE_1_16__empty_n),
    .if_read(fifo_C_drain_PE_1_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_1_16__din),
    .if_full_n(fifo_C_drain_PE_1_16__full_n),
    .if_write(fifo_C_drain_PE_1_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_1_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_1_2__dout),
    .if_empty_n(fifo_C_drain_PE_1_2__empty_n),
    .if_read(fifo_C_drain_PE_1_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_1_2__din),
    .if_full_n(fifo_C_drain_PE_1_2__full_n),
    .if_write(fifo_C_drain_PE_1_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_1_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_1_3__dout),
    .if_empty_n(fifo_C_drain_PE_1_3__empty_n),
    .if_read(fifo_C_drain_PE_1_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_1_3__din),
    .if_full_n(fifo_C_drain_PE_1_3__full_n),
    .if_write(fifo_C_drain_PE_1_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_1_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_1_4__dout),
    .if_empty_n(fifo_C_drain_PE_1_4__empty_n),
    .if_read(fifo_C_drain_PE_1_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_1_4__din),
    .if_full_n(fifo_C_drain_PE_1_4__full_n),
    .if_write(fifo_C_drain_PE_1_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_1_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_1_5__dout),
    .if_empty_n(fifo_C_drain_PE_1_5__empty_n),
    .if_read(fifo_C_drain_PE_1_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_1_5__din),
    .if_full_n(fifo_C_drain_PE_1_5__full_n),
    .if_write(fifo_C_drain_PE_1_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_1_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_1_6__dout),
    .if_empty_n(fifo_C_drain_PE_1_6__empty_n),
    .if_read(fifo_C_drain_PE_1_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_1_6__din),
    .if_full_n(fifo_C_drain_PE_1_6__full_n),
    .if_write(fifo_C_drain_PE_1_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_1_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_1_7__dout),
    .if_empty_n(fifo_C_drain_PE_1_7__empty_n),
    .if_read(fifo_C_drain_PE_1_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_1_7__din),
    .if_full_n(fifo_C_drain_PE_1_7__full_n),
    .if_write(fifo_C_drain_PE_1_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_1_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_1_8__dout),
    .if_empty_n(fifo_C_drain_PE_1_8__empty_n),
    .if_read(fifo_C_drain_PE_1_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_1_8__din),
    .if_full_n(fifo_C_drain_PE_1_8__full_n),
    .if_write(fifo_C_drain_PE_1_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_1_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_1_9__dout),
    .if_empty_n(fifo_C_drain_PE_1_9__empty_n),
    .if_read(fifo_C_drain_PE_1_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_1_9__din),
    .if_full_n(fifo_C_drain_PE_1_9__full_n),
    .if_write(fifo_C_drain_PE_1_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_2_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_2_0__dout),
    .if_empty_n(fifo_C_drain_PE_2_0__empty_n),
    .if_read(fifo_C_drain_PE_2_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_2_0__din),
    .if_full_n(fifo_C_drain_PE_2_0__full_n),
    .if_write(fifo_C_drain_PE_2_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_2_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_2_1__dout),
    .if_empty_n(fifo_C_drain_PE_2_1__empty_n),
    .if_read(fifo_C_drain_PE_2_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_2_1__din),
    .if_full_n(fifo_C_drain_PE_2_1__full_n),
    .if_write(fifo_C_drain_PE_2_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_2_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_2_10__dout),
    .if_empty_n(fifo_C_drain_PE_2_10__empty_n),
    .if_read(fifo_C_drain_PE_2_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_2_10__din),
    .if_full_n(fifo_C_drain_PE_2_10__full_n),
    .if_write(fifo_C_drain_PE_2_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_2_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_2_11__dout),
    .if_empty_n(fifo_C_drain_PE_2_11__empty_n),
    .if_read(fifo_C_drain_PE_2_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_2_11__din),
    .if_full_n(fifo_C_drain_PE_2_11__full_n),
    .if_write(fifo_C_drain_PE_2_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_2_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_2_12__dout),
    .if_empty_n(fifo_C_drain_PE_2_12__empty_n),
    .if_read(fifo_C_drain_PE_2_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_2_12__din),
    .if_full_n(fifo_C_drain_PE_2_12__full_n),
    .if_write(fifo_C_drain_PE_2_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_2_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_2_13__dout),
    .if_empty_n(fifo_C_drain_PE_2_13__empty_n),
    .if_read(fifo_C_drain_PE_2_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_2_13__din),
    .if_full_n(fifo_C_drain_PE_2_13__full_n),
    .if_write(fifo_C_drain_PE_2_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_2_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_2_14__dout),
    .if_empty_n(fifo_C_drain_PE_2_14__empty_n),
    .if_read(fifo_C_drain_PE_2_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_2_14__din),
    .if_full_n(fifo_C_drain_PE_2_14__full_n),
    .if_write(fifo_C_drain_PE_2_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_2_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_2_15__dout),
    .if_empty_n(fifo_C_drain_PE_2_15__empty_n),
    .if_read(fifo_C_drain_PE_2_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_2_15__din),
    .if_full_n(fifo_C_drain_PE_2_15__full_n),
    .if_write(fifo_C_drain_PE_2_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_2_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_2_16__dout),
    .if_empty_n(fifo_C_drain_PE_2_16__empty_n),
    .if_read(fifo_C_drain_PE_2_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_2_16__din),
    .if_full_n(fifo_C_drain_PE_2_16__full_n),
    .if_write(fifo_C_drain_PE_2_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_2_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_2_2__dout),
    .if_empty_n(fifo_C_drain_PE_2_2__empty_n),
    .if_read(fifo_C_drain_PE_2_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_2_2__din),
    .if_full_n(fifo_C_drain_PE_2_2__full_n),
    .if_write(fifo_C_drain_PE_2_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_2_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_2_3__dout),
    .if_empty_n(fifo_C_drain_PE_2_3__empty_n),
    .if_read(fifo_C_drain_PE_2_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_2_3__din),
    .if_full_n(fifo_C_drain_PE_2_3__full_n),
    .if_write(fifo_C_drain_PE_2_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_2_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_2_4__dout),
    .if_empty_n(fifo_C_drain_PE_2_4__empty_n),
    .if_read(fifo_C_drain_PE_2_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_2_4__din),
    .if_full_n(fifo_C_drain_PE_2_4__full_n),
    .if_write(fifo_C_drain_PE_2_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_2_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_2_5__dout),
    .if_empty_n(fifo_C_drain_PE_2_5__empty_n),
    .if_read(fifo_C_drain_PE_2_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_2_5__din),
    .if_full_n(fifo_C_drain_PE_2_5__full_n),
    .if_write(fifo_C_drain_PE_2_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_2_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_2_6__dout),
    .if_empty_n(fifo_C_drain_PE_2_6__empty_n),
    .if_read(fifo_C_drain_PE_2_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_2_6__din),
    .if_full_n(fifo_C_drain_PE_2_6__full_n),
    .if_write(fifo_C_drain_PE_2_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_2_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_2_7__dout),
    .if_empty_n(fifo_C_drain_PE_2_7__empty_n),
    .if_read(fifo_C_drain_PE_2_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_2_7__din),
    .if_full_n(fifo_C_drain_PE_2_7__full_n),
    .if_write(fifo_C_drain_PE_2_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_2_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_2_8__dout),
    .if_empty_n(fifo_C_drain_PE_2_8__empty_n),
    .if_read(fifo_C_drain_PE_2_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_2_8__din),
    .if_full_n(fifo_C_drain_PE_2_8__full_n),
    .if_write(fifo_C_drain_PE_2_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_2_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_2_9__dout),
    .if_empty_n(fifo_C_drain_PE_2_9__empty_n),
    .if_read(fifo_C_drain_PE_2_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_2_9__din),
    .if_full_n(fifo_C_drain_PE_2_9__full_n),
    .if_write(fifo_C_drain_PE_2_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_3_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_3_0__dout),
    .if_empty_n(fifo_C_drain_PE_3_0__empty_n),
    .if_read(fifo_C_drain_PE_3_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_3_0__din),
    .if_full_n(fifo_C_drain_PE_3_0__full_n),
    .if_write(fifo_C_drain_PE_3_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_3_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_3_1__dout),
    .if_empty_n(fifo_C_drain_PE_3_1__empty_n),
    .if_read(fifo_C_drain_PE_3_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_3_1__din),
    .if_full_n(fifo_C_drain_PE_3_1__full_n),
    .if_write(fifo_C_drain_PE_3_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_3_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_3_10__dout),
    .if_empty_n(fifo_C_drain_PE_3_10__empty_n),
    .if_read(fifo_C_drain_PE_3_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_3_10__din),
    .if_full_n(fifo_C_drain_PE_3_10__full_n),
    .if_write(fifo_C_drain_PE_3_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_3_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_3_11__dout),
    .if_empty_n(fifo_C_drain_PE_3_11__empty_n),
    .if_read(fifo_C_drain_PE_3_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_3_11__din),
    .if_full_n(fifo_C_drain_PE_3_11__full_n),
    .if_write(fifo_C_drain_PE_3_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_3_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_3_12__dout),
    .if_empty_n(fifo_C_drain_PE_3_12__empty_n),
    .if_read(fifo_C_drain_PE_3_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_3_12__din),
    .if_full_n(fifo_C_drain_PE_3_12__full_n),
    .if_write(fifo_C_drain_PE_3_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_3_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_3_13__dout),
    .if_empty_n(fifo_C_drain_PE_3_13__empty_n),
    .if_read(fifo_C_drain_PE_3_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_3_13__din),
    .if_full_n(fifo_C_drain_PE_3_13__full_n),
    .if_write(fifo_C_drain_PE_3_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_3_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_3_14__dout),
    .if_empty_n(fifo_C_drain_PE_3_14__empty_n),
    .if_read(fifo_C_drain_PE_3_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_3_14__din),
    .if_full_n(fifo_C_drain_PE_3_14__full_n),
    .if_write(fifo_C_drain_PE_3_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_3_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_3_15__dout),
    .if_empty_n(fifo_C_drain_PE_3_15__empty_n),
    .if_read(fifo_C_drain_PE_3_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_3_15__din),
    .if_full_n(fifo_C_drain_PE_3_15__full_n),
    .if_write(fifo_C_drain_PE_3_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_3_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_3_16__dout),
    .if_empty_n(fifo_C_drain_PE_3_16__empty_n),
    .if_read(fifo_C_drain_PE_3_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_3_16__din),
    .if_full_n(fifo_C_drain_PE_3_16__full_n),
    .if_write(fifo_C_drain_PE_3_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_3_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_3_2__dout),
    .if_empty_n(fifo_C_drain_PE_3_2__empty_n),
    .if_read(fifo_C_drain_PE_3_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_3_2__din),
    .if_full_n(fifo_C_drain_PE_3_2__full_n),
    .if_write(fifo_C_drain_PE_3_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_3_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_3_3__dout),
    .if_empty_n(fifo_C_drain_PE_3_3__empty_n),
    .if_read(fifo_C_drain_PE_3_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_3_3__din),
    .if_full_n(fifo_C_drain_PE_3_3__full_n),
    .if_write(fifo_C_drain_PE_3_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_3_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_3_4__dout),
    .if_empty_n(fifo_C_drain_PE_3_4__empty_n),
    .if_read(fifo_C_drain_PE_3_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_3_4__din),
    .if_full_n(fifo_C_drain_PE_3_4__full_n),
    .if_write(fifo_C_drain_PE_3_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_3_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_3_5__dout),
    .if_empty_n(fifo_C_drain_PE_3_5__empty_n),
    .if_read(fifo_C_drain_PE_3_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_3_5__din),
    .if_full_n(fifo_C_drain_PE_3_5__full_n),
    .if_write(fifo_C_drain_PE_3_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_3_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_3_6__dout),
    .if_empty_n(fifo_C_drain_PE_3_6__empty_n),
    .if_read(fifo_C_drain_PE_3_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_3_6__din),
    .if_full_n(fifo_C_drain_PE_3_6__full_n),
    .if_write(fifo_C_drain_PE_3_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_3_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_3_7__dout),
    .if_empty_n(fifo_C_drain_PE_3_7__empty_n),
    .if_read(fifo_C_drain_PE_3_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_3_7__din),
    .if_full_n(fifo_C_drain_PE_3_7__full_n),
    .if_write(fifo_C_drain_PE_3_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_3_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_3_8__dout),
    .if_empty_n(fifo_C_drain_PE_3_8__empty_n),
    .if_read(fifo_C_drain_PE_3_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_3_8__din),
    .if_full_n(fifo_C_drain_PE_3_8__full_n),
    .if_write(fifo_C_drain_PE_3_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_3_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_3_9__dout),
    .if_empty_n(fifo_C_drain_PE_3_9__empty_n),
    .if_read(fifo_C_drain_PE_3_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_3_9__din),
    .if_full_n(fifo_C_drain_PE_3_9__full_n),
    .if_write(fifo_C_drain_PE_3_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_4_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_4_0__dout),
    .if_empty_n(fifo_C_drain_PE_4_0__empty_n),
    .if_read(fifo_C_drain_PE_4_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_4_0__din),
    .if_full_n(fifo_C_drain_PE_4_0__full_n),
    .if_write(fifo_C_drain_PE_4_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_4_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_4_1__dout),
    .if_empty_n(fifo_C_drain_PE_4_1__empty_n),
    .if_read(fifo_C_drain_PE_4_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_4_1__din),
    .if_full_n(fifo_C_drain_PE_4_1__full_n),
    .if_write(fifo_C_drain_PE_4_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_4_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_4_10__dout),
    .if_empty_n(fifo_C_drain_PE_4_10__empty_n),
    .if_read(fifo_C_drain_PE_4_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_4_10__din),
    .if_full_n(fifo_C_drain_PE_4_10__full_n),
    .if_write(fifo_C_drain_PE_4_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_4_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_4_11__dout),
    .if_empty_n(fifo_C_drain_PE_4_11__empty_n),
    .if_read(fifo_C_drain_PE_4_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_4_11__din),
    .if_full_n(fifo_C_drain_PE_4_11__full_n),
    .if_write(fifo_C_drain_PE_4_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_4_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_4_12__dout),
    .if_empty_n(fifo_C_drain_PE_4_12__empty_n),
    .if_read(fifo_C_drain_PE_4_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_4_12__din),
    .if_full_n(fifo_C_drain_PE_4_12__full_n),
    .if_write(fifo_C_drain_PE_4_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_4_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_4_13__dout),
    .if_empty_n(fifo_C_drain_PE_4_13__empty_n),
    .if_read(fifo_C_drain_PE_4_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_4_13__din),
    .if_full_n(fifo_C_drain_PE_4_13__full_n),
    .if_write(fifo_C_drain_PE_4_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_4_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_4_14__dout),
    .if_empty_n(fifo_C_drain_PE_4_14__empty_n),
    .if_read(fifo_C_drain_PE_4_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_4_14__din),
    .if_full_n(fifo_C_drain_PE_4_14__full_n),
    .if_write(fifo_C_drain_PE_4_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_4_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_4_15__dout),
    .if_empty_n(fifo_C_drain_PE_4_15__empty_n),
    .if_read(fifo_C_drain_PE_4_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_4_15__din),
    .if_full_n(fifo_C_drain_PE_4_15__full_n),
    .if_write(fifo_C_drain_PE_4_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_4_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_4_16__dout),
    .if_empty_n(fifo_C_drain_PE_4_16__empty_n),
    .if_read(fifo_C_drain_PE_4_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_4_16__din),
    .if_full_n(fifo_C_drain_PE_4_16__full_n),
    .if_write(fifo_C_drain_PE_4_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_4_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_4_2__dout),
    .if_empty_n(fifo_C_drain_PE_4_2__empty_n),
    .if_read(fifo_C_drain_PE_4_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_4_2__din),
    .if_full_n(fifo_C_drain_PE_4_2__full_n),
    .if_write(fifo_C_drain_PE_4_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_4_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_4_3__dout),
    .if_empty_n(fifo_C_drain_PE_4_3__empty_n),
    .if_read(fifo_C_drain_PE_4_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_4_3__din),
    .if_full_n(fifo_C_drain_PE_4_3__full_n),
    .if_write(fifo_C_drain_PE_4_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_4_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_4_4__dout),
    .if_empty_n(fifo_C_drain_PE_4_4__empty_n),
    .if_read(fifo_C_drain_PE_4_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_4_4__din),
    .if_full_n(fifo_C_drain_PE_4_4__full_n),
    .if_write(fifo_C_drain_PE_4_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_4_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_4_5__dout),
    .if_empty_n(fifo_C_drain_PE_4_5__empty_n),
    .if_read(fifo_C_drain_PE_4_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_4_5__din),
    .if_full_n(fifo_C_drain_PE_4_5__full_n),
    .if_write(fifo_C_drain_PE_4_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_4_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_4_6__dout),
    .if_empty_n(fifo_C_drain_PE_4_6__empty_n),
    .if_read(fifo_C_drain_PE_4_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_4_6__din),
    .if_full_n(fifo_C_drain_PE_4_6__full_n),
    .if_write(fifo_C_drain_PE_4_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_4_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_4_7__dout),
    .if_empty_n(fifo_C_drain_PE_4_7__empty_n),
    .if_read(fifo_C_drain_PE_4_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_4_7__din),
    .if_full_n(fifo_C_drain_PE_4_7__full_n),
    .if_write(fifo_C_drain_PE_4_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_4_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_4_8__dout),
    .if_empty_n(fifo_C_drain_PE_4_8__empty_n),
    .if_read(fifo_C_drain_PE_4_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_4_8__din),
    .if_full_n(fifo_C_drain_PE_4_8__full_n),
    .if_write(fifo_C_drain_PE_4_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_4_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_4_9__dout),
    .if_empty_n(fifo_C_drain_PE_4_9__empty_n),
    .if_read(fifo_C_drain_PE_4_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_4_9__din),
    .if_full_n(fifo_C_drain_PE_4_9__full_n),
    .if_write(fifo_C_drain_PE_4_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_5_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_5_0__dout),
    .if_empty_n(fifo_C_drain_PE_5_0__empty_n),
    .if_read(fifo_C_drain_PE_5_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_5_0__din),
    .if_full_n(fifo_C_drain_PE_5_0__full_n),
    .if_write(fifo_C_drain_PE_5_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_5_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_5_1__dout),
    .if_empty_n(fifo_C_drain_PE_5_1__empty_n),
    .if_read(fifo_C_drain_PE_5_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_5_1__din),
    .if_full_n(fifo_C_drain_PE_5_1__full_n),
    .if_write(fifo_C_drain_PE_5_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_5_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_5_10__dout),
    .if_empty_n(fifo_C_drain_PE_5_10__empty_n),
    .if_read(fifo_C_drain_PE_5_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_5_10__din),
    .if_full_n(fifo_C_drain_PE_5_10__full_n),
    .if_write(fifo_C_drain_PE_5_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_5_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_5_11__dout),
    .if_empty_n(fifo_C_drain_PE_5_11__empty_n),
    .if_read(fifo_C_drain_PE_5_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_5_11__din),
    .if_full_n(fifo_C_drain_PE_5_11__full_n),
    .if_write(fifo_C_drain_PE_5_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_5_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_5_12__dout),
    .if_empty_n(fifo_C_drain_PE_5_12__empty_n),
    .if_read(fifo_C_drain_PE_5_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_5_12__din),
    .if_full_n(fifo_C_drain_PE_5_12__full_n),
    .if_write(fifo_C_drain_PE_5_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_5_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_5_13__dout),
    .if_empty_n(fifo_C_drain_PE_5_13__empty_n),
    .if_read(fifo_C_drain_PE_5_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_5_13__din),
    .if_full_n(fifo_C_drain_PE_5_13__full_n),
    .if_write(fifo_C_drain_PE_5_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_5_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_5_14__dout),
    .if_empty_n(fifo_C_drain_PE_5_14__empty_n),
    .if_read(fifo_C_drain_PE_5_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_5_14__din),
    .if_full_n(fifo_C_drain_PE_5_14__full_n),
    .if_write(fifo_C_drain_PE_5_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_5_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_5_15__dout),
    .if_empty_n(fifo_C_drain_PE_5_15__empty_n),
    .if_read(fifo_C_drain_PE_5_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_5_15__din),
    .if_full_n(fifo_C_drain_PE_5_15__full_n),
    .if_write(fifo_C_drain_PE_5_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_5_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_5_16__dout),
    .if_empty_n(fifo_C_drain_PE_5_16__empty_n),
    .if_read(fifo_C_drain_PE_5_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_5_16__din),
    .if_full_n(fifo_C_drain_PE_5_16__full_n),
    .if_write(fifo_C_drain_PE_5_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_5_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_5_2__dout),
    .if_empty_n(fifo_C_drain_PE_5_2__empty_n),
    .if_read(fifo_C_drain_PE_5_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_5_2__din),
    .if_full_n(fifo_C_drain_PE_5_2__full_n),
    .if_write(fifo_C_drain_PE_5_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_5_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_5_3__dout),
    .if_empty_n(fifo_C_drain_PE_5_3__empty_n),
    .if_read(fifo_C_drain_PE_5_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_5_3__din),
    .if_full_n(fifo_C_drain_PE_5_3__full_n),
    .if_write(fifo_C_drain_PE_5_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_5_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_5_4__dout),
    .if_empty_n(fifo_C_drain_PE_5_4__empty_n),
    .if_read(fifo_C_drain_PE_5_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_5_4__din),
    .if_full_n(fifo_C_drain_PE_5_4__full_n),
    .if_write(fifo_C_drain_PE_5_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_5_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_5_5__dout),
    .if_empty_n(fifo_C_drain_PE_5_5__empty_n),
    .if_read(fifo_C_drain_PE_5_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_5_5__din),
    .if_full_n(fifo_C_drain_PE_5_5__full_n),
    .if_write(fifo_C_drain_PE_5_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_5_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_5_6__dout),
    .if_empty_n(fifo_C_drain_PE_5_6__empty_n),
    .if_read(fifo_C_drain_PE_5_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_5_6__din),
    .if_full_n(fifo_C_drain_PE_5_6__full_n),
    .if_write(fifo_C_drain_PE_5_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_5_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_5_7__dout),
    .if_empty_n(fifo_C_drain_PE_5_7__empty_n),
    .if_read(fifo_C_drain_PE_5_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_5_7__din),
    .if_full_n(fifo_C_drain_PE_5_7__full_n),
    .if_write(fifo_C_drain_PE_5_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_5_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_5_8__dout),
    .if_empty_n(fifo_C_drain_PE_5_8__empty_n),
    .if_read(fifo_C_drain_PE_5_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_5_8__din),
    .if_full_n(fifo_C_drain_PE_5_8__full_n),
    .if_write(fifo_C_drain_PE_5_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_5_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_5_9__dout),
    .if_empty_n(fifo_C_drain_PE_5_9__empty_n),
    .if_read(fifo_C_drain_PE_5_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_5_9__din),
    .if_full_n(fifo_C_drain_PE_5_9__full_n),
    .if_write(fifo_C_drain_PE_5_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_6_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_6_0__dout),
    .if_empty_n(fifo_C_drain_PE_6_0__empty_n),
    .if_read(fifo_C_drain_PE_6_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_6_0__din),
    .if_full_n(fifo_C_drain_PE_6_0__full_n),
    .if_write(fifo_C_drain_PE_6_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_6_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_6_1__dout),
    .if_empty_n(fifo_C_drain_PE_6_1__empty_n),
    .if_read(fifo_C_drain_PE_6_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_6_1__din),
    .if_full_n(fifo_C_drain_PE_6_1__full_n),
    .if_write(fifo_C_drain_PE_6_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_6_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_6_10__dout),
    .if_empty_n(fifo_C_drain_PE_6_10__empty_n),
    .if_read(fifo_C_drain_PE_6_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_6_10__din),
    .if_full_n(fifo_C_drain_PE_6_10__full_n),
    .if_write(fifo_C_drain_PE_6_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_6_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_6_11__dout),
    .if_empty_n(fifo_C_drain_PE_6_11__empty_n),
    .if_read(fifo_C_drain_PE_6_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_6_11__din),
    .if_full_n(fifo_C_drain_PE_6_11__full_n),
    .if_write(fifo_C_drain_PE_6_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_6_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_6_12__dout),
    .if_empty_n(fifo_C_drain_PE_6_12__empty_n),
    .if_read(fifo_C_drain_PE_6_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_6_12__din),
    .if_full_n(fifo_C_drain_PE_6_12__full_n),
    .if_write(fifo_C_drain_PE_6_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_6_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_6_13__dout),
    .if_empty_n(fifo_C_drain_PE_6_13__empty_n),
    .if_read(fifo_C_drain_PE_6_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_6_13__din),
    .if_full_n(fifo_C_drain_PE_6_13__full_n),
    .if_write(fifo_C_drain_PE_6_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_6_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_6_14__dout),
    .if_empty_n(fifo_C_drain_PE_6_14__empty_n),
    .if_read(fifo_C_drain_PE_6_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_6_14__din),
    .if_full_n(fifo_C_drain_PE_6_14__full_n),
    .if_write(fifo_C_drain_PE_6_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_6_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_6_15__dout),
    .if_empty_n(fifo_C_drain_PE_6_15__empty_n),
    .if_read(fifo_C_drain_PE_6_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_6_15__din),
    .if_full_n(fifo_C_drain_PE_6_15__full_n),
    .if_write(fifo_C_drain_PE_6_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_6_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_6_16__dout),
    .if_empty_n(fifo_C_drain_PE_6_16__empty_n),
    .if_read(fifo_C_drain_PE_6_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_6_16__din),
    .if_full_n(fifo_C_drain_PE_6_16__full_n),
    .if_write(fifo_C_drain_PE_6_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_6_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_6_2__dout),
    .if_empty_n(fifo_C_drain_PE_6_2__empty_n),
    .if_read(fifo_C_drain_PE_6_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_6_2__din),
    .if_full_n(fifo_C_drain_PE_6_2__full_n),
    .if_write(fifo_C_drain_PE_6_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_6_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_6_3__dout),
    .if_empty_n(fifo_C_drain_PE_6_3__empty_n),
    .if_read(fifo_C_drain_PE_6_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_6_3__din),
    .if_full_n(fifo_C_drain_PE_6_3__full_n),
    .if_write(fifo_C_drain_PE_6_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_6_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_6_4__dout),
    .if_empty_n(fifo_C_drain_PE_6_4__empty_n),
    .if_read(fifo_C_drain_PE_6_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_6_4__din),
    .if_full_n(fifo_C_drain_PE_6_4__full_n),
    .if_write(fifo_C_drain_PE_6_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_6_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_6_5__dout),
    .if_empty_n(fifo_C_drain_PE_6_5__empty_n),
    .if_read(fifo_C_drain_PE_6_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_6_5__din),
    .if_full_n(fifo_C_drain_PE_6_5__full_n),
    .if_write(fifo_C_drain_PE_6_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_6_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_6_6__dout),
    .if_empty_n(fifo_C_drain_PE_6_6__empty_n),
    .if_read(fifo_C_drain_PE_6_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_6_6__din),
    .if_full_n(fifo_C_drain_PE_6_6__full_n),
    .if_write(fifo_C_drain_PE_6_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_6_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_6_7__dout),
    .if_empty_n(fifo_C_drain_PE_6_7__empty_n),
    .if_read(fifo_C_drain_PE_6_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_6_7__din),
    .if_full_n(fifo_C_drain_PE_6_7__full_n),
    .if_write(fifo_C_drain_PE_6_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_6_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_6_8__dout),
    .if_empty_n(fifo_C_drain_PE_6_8__empty_n),
    .if_read(fifo_C_drain_PE_6_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_6_8__din),
    .if_full_n(fifo_C_drain_PE_6_8__full_n),
    .if_write(fifo_C_drain_PE_6_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_6_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_6_9__dout),
    .if_empty_n(fifo_C_drain_PE_6_9__empty_n),
    .if_read(fifo_C_drain_PE_6_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_6_9__din),
    .if_full_n(fifo_C_drain_PE_6_9__full_n),
    .if_write(fifo_C_drain_PE_6_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_7_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_7_0__dout),
    .if_empty_n(fifo_C_drain_PE_7_0__empty_n),
    .if_read(fifo_C_drain_PE_7_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_7_0__din),
    .if_full_n(fifo_C_drain_PE_7_0__full_n),
    .if_write(fifo_C_drain_PE_7_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_7_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_7_1__dout),
    .if_empty_n(fifo_C_drain_PE_7_1__empty_n),
    .if_read(fifo_C_drain_PE_7_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_7_1__din),
    .if_full_n(fifo_C_drain_PE_7_1__full_n),
    .if_write(fifo_C_drain_PE_7_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_7_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_7_10__dout),
    .if_empty_n(fifo_C_drain_PE_7_10__empty_n),
    .if_read(fifo_C_drain_PE_7_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_7_10__din),
    .if_full_n(fifo_C_drain_PE_7_10__full_n),
    .if_write(fifo_C_drain_PE_7_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_7_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_7_11__dout),
    .if_empty_n(fifo_C_drain_PE_7_11__empty_n),
    .if_read(fifo_C_drain_PE_7_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_7_11__din),
    .if_full_n(fifo_C_drain_PE_7_11__full_n),
    .if_write(fifo_C_drain_PE_7_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_7_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_7_12__dout),
    .if_empty_n(fifo_C_drain_PE_7_12__empty_n),
    .if_read(fifo_C_drain_PE_7_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_7_12__din),
    .if_full_n(fifo_C_drain_PE_7_12__full_n),
    .if_write(fifo_C_drain_PE_7_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_7_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_7_13__dout),
    .if_empty_n(fifo_C_drain_PE_7_13__empty_n),
    .if_read(fifo_C_drain_PE_7_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_7_13__din),
    .if_full_n(fifo_C_drain_PE_7_13__full_n),
    .if_write(fifo_C_drain_PE_7_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_7_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_7_14__dout),
    .if_empty_n(fifo_C_drain_PE_7_14__empty_n),
    .if_read(fifo_C_drain_PE_7_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_7_14__din),
    .if_full_n(fifo_C_drain_PE_7_14__full_n),
    .if_write(fifo_C_drain_PE_7_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_7_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_7_15__dout),
    .if_empty_n(fifo_C_drain_PE_7_15__empty_n),
    .if_read(fifo_C_drain_PE_7_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_7_15__din),
    .if_full_n(fifo_C_drain_PE_7_15__full_n),
    .if_write(fifo_C_drain_PE_7_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_7_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_7_16__dout),
    .if_empty_n(fifo_C_drain_PE_7_16__empty_n),
    .if_read(fifo_C_drain_PE_7_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_7_16__din),
    .if_full_n(fifo_C_drain_PE_7_16__full_n),
    .if_write(fifo_C_drain_PE_7_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_7_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_7_2__dout),
    .if_empty_n(fifo_C_drain_PE_7_2__empty_n),
    .if_read(fifo_C_drain_PE_7_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_7_2__din),
    .if_full_n(fifo_C_drain_PE_7_2__full_n),
    .if_write(fifo_C_drain_PE_7_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_7_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_7_3__dout),
    .if_empty_n(fifo_C_drain_PE_7_3__empty_n),
    .if_read(fifo_C_drain_PE_7_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_7_3__din),
    .if_full_n(fifo_C_drain_PE_7_3__full_n),
    .if_write(fifo_C_drain_PE_7_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_7_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_7_4__dout),
    .if_empty_n(fifo_C_drain_PE_7_4__empty_n),
    .if_read(fifo_C_drain_PE_7_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_7_4__din),
    .if_full_n(fifo_C_drain_PE_7_4__full_n),
    .if_write(fifo_C_drain_PE_7_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_7_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_7_5__dout),
    .if_empty_n(fifo_C_drain_PE_7_5__empty_n),
    .if_read(fifo_C_drain_PE_7_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_7_5__din),
    .if_full_n(fifo_C_drain_PE_7_5__full_n),
    .if_write(fifo_C_drain_PE_7_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_7_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_7_6__dout),
    .if_empty_n(fifo_C_drain_PE_7_6__empty_n),
    .if_read(fifo_C_drain_PE_7_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_7_6__din),
    .if_full_n(fifo_C_drain_PE_7_6__full_n),
    .if_write(fifo_C_drain_PE_7_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_7_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_7_7__dout),
    .if_empty_n(fifo_C_drain_PE_7_7__empty_n),
    .if_read(fifo_C_drain_PE_7_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_7_7__din),
    .if_full_n(fifo_C_drain_PE_7_7__full_n),
    .if_write(fifo_C_drain_PE_7_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_7_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_7_8__dout),
    .if_empty_n(fifo_C_drain_PE_7_8__empty_n),
    .if_read(fifo_C_drain_PE_7_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_7_8__din),
    .if_full_n(fifo_C_drain_PE_7_8__full_n),
    .if_write(fifo_C_drain_PE_7_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_7_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_7_9__dout),
    .if_empty_n(fifo_C_drain_PE_7_9__empty_n),
    .if_read(fifo_C_drain_PE_7_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_7_9__din),
    .if_full_n(fifo_C_drain_PE_7_9__full_n),
    .if_write(fifo_C_drain_PE_7_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_8_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_8_0__dout),
    .if_empty_n(fifo_C_drain_PE_8_0__empty_n),
    .if_read(fifo_C_drain_PE_8_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_8_0__din),
    .if_full_n(fifo_C_drain_PE_8_0__full_n),
    .if_write(fifo_C_drain_PE_8_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_8_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_8_1__dout),
    .if_empty_n(fifo_C_drain_PE_8_1__empty_n),
    .if_read(fifo_C_drain_PE_8_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_8_1__din),
    .if_full_n(fifo_C_drain_PE_8_1__full_n),
    .if_write(fifo_C_drain_PE_8_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_8_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_8_10__dout),
    .if_empty_n(fifo_C_drain_PE_8_10__empty_n),
    .if_read(fifo_C_drain_PE_8_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_8_10__din),
    .if_full_n(fifo_C_drain_PE_8_10__full_n),
    .if_write(fifo_C_drain_PE_8_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_8_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_8_11__dout),
    .if_empty_n(fifo_C_drain_PE_8_11__empty_n),
    .if_read(fifo_C_drain_PE_8_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_8_11__din),
    .if_full_n(fifo_C_drain_PE_8_11__full_n),
    .if_write(fifo_C_drain_PE_8_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_8_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_8_12__dout),
    .if_empty_n(fifo_C_drain_PE_8_12__empty_n),
    .if_read(fifo_C_drain_PE_8_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_8_12__din),
    .if_full_n(fifo_C_drain_PE_8_12__full_n),
    .if_write(fifo_C_drain_PE_8_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_8_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_8_13__dout),
    .if_empty_n(fifo_C_drain_PE_8_13__empty_n),
    .if_read(fifo_C_drain_PE_8_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_8_13__din),
    .if_full_n(fifo_C_drain_PE_8_13__full_n),
    .if_write(fifo_C_drain_PE_8_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_8_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_8_14__dout),
    .if_empty_n(fifo_C_drain_PE_8_14__empty_n),
    .if_read(fifo_C_drain_PE_8_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_8_14__din),
    .if_full_n(fifo_C_drain_PE_8_14__full_n),
    .if_write(fifo_C_drain_PE_8_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_8_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_8_15__dout),
    .if_empty_n(fifo_C_drain_PE_8_15__empty_n),
    .if_read(fifo_C_drain_PE_8_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_8_15__din),
    .if_full_n(fifo_C_drain_PE_8_15__full_n),
    .if_write(fifo_C_drain_PE_8_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_8_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_8_16__dout),
    .if_empty_n(fifo_C_drain_PE_8_16__empty_n),
    .if_read(fifo_C_drain_PE_8_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_8_16__din),
    .if_full_n(fifo_C_drain_PE_8_16__full_n),
    .if_write(fifo_C_drain_PE_8_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_8_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_8_2__dout),
    .if_empty_n(fifo_C_drain_PE_8_2__empty_n),
    .if_read(fifo_C_drain_PE_8_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_8_2__din),
    .if_full_n(fifo_C_drain_PE_8_2__full_n),
    .if_write(fifo_C_drain_PE_8_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_8_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_8_3__dout),
    .if_empty_n(fifo_C_drain_PE_8_3__empty_n),
    .if_read(fifo_C_drain_PE_8_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_8_3__din),
    .if_full_n(fifo_C_drain_PE_8_3__full_n),
    .if_write(fifo_C_drain_PE_8_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_8_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_8_4__dout),
    .if_empty_n(fifo_C_drain_PE_8_4__empty_n),
    .if_read(fifo_C_drain_PE_8_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_8_4__din),
    .if_full_n(fifo_C_drain_PE_8_4__full_n),
    .if_write(fifo_C_drain_PE_8_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_8_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_8_5__dout),
    .if_empty_n(fifo_C_drain_PE_8_5__empty_n),
    .if_read(fifo_C_drain_PE_8_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_8_5__din),
    .if_full_n(fifo_C_drain_PE_8_5__full_n),
    .if_write(fifo_C_drain_PE_8_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_8_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_8_6__dout),
    .if_empty_n(fifo_C_drain_PE_8_6__empty_n),
    .if_read(fifo_C_drain_PE_8_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_8_6__din),
    .if_full_n(fifo_C_drain_PE_8_6__full_n),
    .if_write(fifo_C_drain_PE_8_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_8_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_8_7__dout),
    .if_empty_n(fifo_C_drain_PE_8_7__empty_n),
    .if_read(fifo_C_drain_PE_8_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_8_7__din),
    .if_full_n(fifo_C_drain_PE_8_7__full_n),
    .if_write(fifo_C_drain_PE_8_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_8_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_8_8__dout),
    .if_empty_n(fifo_C_drain_PE_8_8__empty_n),
    .if_read(fifo_C_drain_PE_8_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_8_8__din),
    .if_full_n(fifo_C_drain_PE_8_8__full_n),
    .if_write(fifo_C_drain_PE_8_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_8_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_8_9__dout),
    .if_empty_n(fifo_C_drain_PE_8_9__empty_n),
    .if_read(fifo_C_drain_PE_8_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_8_9__din),
    .if_full_n(fifo_C_drain_PE_8_9__full_n),
    .if_write(fifo_C_drain_PE_8_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_9_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_9_0__dout),
    .if_empty_n(fifo_C_drain_PE_9_0__empty_n),
    .if_read(fifo_C_drain_PE_9_0__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_9_0__din),
    .if_full_n(fifo_C_drain_PE_9_0__full_n),
    .if_write(fifo_C_drain_PE_9_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_9_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_9_1__dout),
    .if_empty_n(fifo_C_drain_PE_9_1__empty_n),
    .if_read(fifo_C_drain_PE_9_1__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_9_1__din),
    .if_full_n(fifo_C_drain_PE_9_1__full_n),
    .if_write(fifo_C_drain_PE_9_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_9_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_9_10__dout),
    .if_empty_n(fifo_C_drain_PE_9_10__empty_n),
    .if_read(fifo_C_drain_PE_9_10__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_9_10__din),
    .if_full_n(fifo_C_drain_PE_9_10__full_n),
    .if_write(fifo_C_drain_PE_9_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_9_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_9_11__dout),
    .if_empty_n(fifo_C_drain_PE_9_11__empty_n),
    .if_read(fifo_C_drain_PE_9_11__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_9_11__din),
    .if_full_n(fifo_C_drain_PE_9_11__full_n),
    .if_write(fifo_C_drain_PE_9_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_9_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_9_12__dout),
    .if_empty_n(fifo_C_drain_PE_9_12__empty_n),
    .if_read(fifo_C_drain_PE_9_12__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_9_12__din),
    .if_full_n(fifo_C_drain_PE_9_12__full_n),
    .if_write(fifo_C_drain_PE_9_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_9_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_9_13__dout),
    .if_empty_n(fifo_C_drain_PE_9_13__empty_n),
    .if_read(fifo_C_drain_PE_9_13__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_9_13__din),
    .if_full_n(fifo_C_drain_PE_9_13__full_n),
    .if_write(fifo_C_drain_PE_9_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_9_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_9_14__dout),
    .if_empty_n(fifo_C_drain_PE_9_14__empty_n),
    .if_read(fifo_C_drain_PE_9_14__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_9_14__din),
    .if_full_n(fifo_C_drain_PE_9_14__full_n),
    .if_write(fifo_C_drain_PE_9_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_9_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_9_15__dout),
    .if_empty_n(fifo_C_drain_PE_9_15__empty_n),
    .if_read(fifo_C_drain_PE_9_15__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_9_15__din),
    .if_full_n(fifo_C_drain_PE_9_15__full_n),
    .if_write(fifo_C_drain_PE_9_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_9_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_9_16__dout),
    .if_empty_n(fifo_C_drain_PE_9_16__empty_n),
    .if_read(fifo_C_drain_PE_9_16__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_9_16__din),
    .if_full_n(fifo_C_drain_PE_9_16__full_n),
    .if_write(fifo_C_drain_PE_9_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_9_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_9_2__dout),
    .if_empty_n(fifo_C_drain_PE_9_2__empty_n),
    .if_read(fifo_C_drain_PE_9_2__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_9_2__din),
    .if_full_n(fifo_C_drain_PE_9_2__full_n),
    .if_write(fifo_C_drain_PE_9_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_9_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_9_3__dout),
    .if_empty_n(fifo_C_drain_PE_9_3__empty_n),
    .if_read(fifo_C_drain_PE_9_3__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_9_3__din),
    .if_full_n(fifo_C_drain_PE_9_3__full_n),
    .if_write(fifo_C_drain_PE_9_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_9_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_9_4__dout),
    .if_empty_n(fifo_C_drain_PE_9_4__empty_n),
    .if_read(fifo_C_drain_PE_9_4__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_9_4__din),
    .if_full_n(fifo_C_drain_PE_9_4__full_n),
    .if_write(fifo_C_drain_PE_9_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_9_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_9_5__dout),
    .if_empty_n(fifo_C_drain_PE_9_5__empty_n),
    .if_read(fifo_C_drain_PE_9_5__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_9_5__din),
    .if_full_n(fifo_C_drain_PE_9_5__full_n),
    .if_write(fifo_C_drain_PE_9_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_9_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_9_6__dout),
    .if_empty_n(fifo_C_drain_PE_9_6__empty_n),
    .if_read(fifo_C_drain_PE_9_6__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_9_6__din),
    .if_full_n(fifo_C_drain_PE_9_6__full_n),
    .if_write(fifo_C_drain_PE_9_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_9_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_9_7__dout),
    .if_empty_n(fifo_C_drain_PE_9_7__empty_n),
    .if_read(fifo_C_drain_PE_9_7__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_9_7__din),
    .if_full_n(fifo_C_drain_PE_9_7__full_n),
    .if_write(fifo_C_drain_PE_9_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_9_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_9_8__dout),
    .if_empty_n(fifo_C_drain_PE_9_8__empty_n),
    .if_read(fifo_C_drain_PE_9_8__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_9_8__din),
    .if_full_n(fifo_C_drain_PE_9_8__full_n),
    .if_write(fifo_C_drain_PE_9_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(17),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  fifo_C_drain_PE_9_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(fifo_C_drain_PE_9_9__dout),
    .if_empty_n(fifo_C_drain_PE_9_9__empty_n),
    .if_read(fifo_C_drain_PE_9_9__read),
    .if_read_ce(1'b1),
    .if_din(fifo_C_drain_PE_9_9__din),
    .if_full_n(fifo_C_drain_PE_9_9__full_n),
    .if_write(fifo_C_drain_PE_9_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) A_IO_L2_in
  A_IO_L2_in_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(A_IO_L2_in_0__ap_start),
    .ap_done(A_IO_L2_in_0__ap_done),
    .ap_idle(A_IO_L2_in_0__ap_idle),
    .ap_ready(A_IO_L2_in_0__ap_ready),
    .idx(64'd0),
    .fifo_A_in_s_dout(fifo_A_A_IO_L2_in_0__dout),
    .fifo_A_in_peek_dout(fifo_A_A_IO_L2_in_0__dout),
    .fifo_A_in_s_empty_n(fifo_A_A_IO_L2_in_0__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_A_IO_L2_in_0__empty_n),
    .fifo_A_in_s_read(fifo_A_A_IO_L2_in_0__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_A_IO_L2_in_1__din),
    .fifo_A_out_full_n(fifo_A_A_IO_L2_in_1__full_n),
    .fifo_A_out_write(fifo_A_A_IO_L2_in_1__write),
    .fifo_A_local_out_din(fifo_A_PE_0_0__din),
    .fifo_A_local_out_full_n(fifo_A_PE_0_0__full_n),
    .fifo_A_local_out_write(fifo_A_PE_0_0__write)
  );


  (* keep_hierarchy = "yes" *) A_IO_L2_in
  A_IO_L2_in_1
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(A_IO_L2_in_1__ap_start),
    .ap_done(A_IO_L2_in_1__ap_done),
    .ap_idle(A_IO_L2_in_1__ap_idle),
    .ap_ready(A_IO_L2_in_1__ap_ready),
    .idx(64'd1),
    .fifo_A_in_s_dout(fifo_A_A_IO_L2_in_1__dout),
    .fifo_A_in_peek_dout(fifo_A_A_IO_L2_in_1__dout),
    .fifo_A_in_s_empty_n(fifo_A_A_IO_L2_in_1__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_A_IO_L2_in_1__empty_n),
    .fifo_A_in_s_read(fifo_A_A_IO_L2_in_1__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_A_IO_L2_in_2__din),
    .fifo_A_out_full_n(fifo_A_A_IO_L2_in_2__full_n),
    .fifo_A_out_write(fifo_A_A_IO_L2_in_2__write),
    .fifo_A_local_out_din(fifo_A_PE_1_0__din),
    .fifo_A_local_out_full_n(fifo_A_PE_1_0__full_n),
    .fifo_A_local_out_write(fifo_A_PE_1_0__write)
  );


  (* keep_hierarchy = "yes" *) A_IO_L2_in
  A_IO_L2_in_2
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(A_IO_L2_in_2__ap_start),
    .ap_done(A_IO_L2_in_2__ap_done),
    .ap_idle(A_IO_L2_in_2__ap_idle),
    .ap_ready(A_IO_L2_in_2__ap_ready),
    .idx(64'd2),
    .fifo_A_in_s_dout(fifo_A_A_IO_L2_in_2__dout),
    .fifo_A_in_peek_dout(fifo_A_A_IO_L2_in_2__dout),
    .fifo_A_in_s_empty_n(fifo_A_A_IO_L2_in_2__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_A_IO_L2_in_2__empty_n),
    .fifo_A_in_s_read(fifo_A_A_IO_L2_in_2__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_A_IO_L2_in_3__din),
    .fifo_A_out_full_n(fifo_A_A_IO_L2_in_3__full_n),
    .fifo_A_out_write(fifo_A_A_IO_L2_in_3__write),
    .fifo_A_local_out_din(fifo_A_PE_2_0__din),
    .fifo_A_local_out_full_n(fifo_A_PE_2_0__full_n),
    .fifo_A_local_out_write(fifo_A_PE_2_0__write)
  );


  (* keep_hierarchy = "yes" *) A_IO_L2_in
  A_IO_L2_in_3
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(A_IO_L2_in_3__ap_start),
    .ap_done(A_IO_L2_in_3__ap_done),
    .ap_idle(A_IO_L2_in_3__ap_idle),
    .ap_ready(A_IO_L2_in_3__ap_ready),
    .idx(64'd3),
    .fifo_A_in_s_dout(fifo_A_A_IO_L2_in_3__dout),
    .fifo_A_in_peek_dout(fifo_A_A_IO_L2_in_3__dout),
    .fifo_A_in_s_empty_n(fifo_A_A_IO_L2_in_3__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_A_IO_L2_in_3__empty_n),
    .fifo_A_in_s_read(fifo_A_A_IO_L2_in_3__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_A_IO_L2_in_4__din),
    .fifo_A_out_full_n(fifo_A_A_IO_L2_in_4__full_n),
    .fifo_A_out_write(fifo_A_A_IO_L2_in_4__write),
    .fifo_A_local_out_din(fifo_A_PE_3_0__din),
    .fifo_A_local_out_full_n(fifo_A_PE_3_0__full_n),
    .fifo_A_local_out_write(fifo_A_PE_3_0__write)
  );


  (* keep_hierarchy = "yes" *) A_IO_L2_in
  A_IO_L2_in_4
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(A_IO_L2_in_4__ap_start),
    .ap_done(A_IO_L2_in_4__ap_done),
    .ap_idle(A_IO_L2_in_4__ap_idle),
    .ap_ready(A_IO_L2_in_4__ap_ready),
    .idx(64'd4),
    .fifo_A_in_s_dout(fifo_A_A_IO_L2_in_4__dout),
    .fifo_A_in_peek_dout(fifo_A_A_IO_L2_in_4__dout),
    .fifo_A_in_s_empty_n(fifo_A_A_IO_L2_in_4__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_A_IO_L2_in_4__empty_n),
    .fifo_A_in_s_read(fifo_A_A_IO_L2_in_4__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_A_IO_L2_in_5__din),
    .fifo_A_out_full_n(fifo_A_A_IO_L2_in_5__full_n),
    .fifo_A_out_write(fifo_A_A_IO_L2_in_5__write),
    .fifo_A_local_out_din(fifo_A_PE_4_0__din),
    .fifo_A_local_out_full_n(fifo_A_PE_4_0__full_n),
    .fifo_A_local_out_write(fifo_A_PE_4_0__write)
  );


  (* keep_hierarchy = "yes" *) A_IO_L2_in
  A_IO_L2_in_5
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(A_IO_L2_in_5__ap_start),
    .ap_done(A_IO_L2_in_5__ap_done),
    .ap_idle(A_IO_L2_in_5__ap_idle),
    .ap_ready(A_IO_L2_in_5__ap_ready),
    .idx(64'd5),
    .fifo_A_in_s_dout(fifo_A_A_IO_L2_in_5__dout),
    .fifo_A_in_peek_dout(fifo_A_A_IO_L2_in_5__dout),
    .fifo_A_in_s_empty_n(fifo_A_A_IO_L2_in_5__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_A_IO_L2_in_5__empty_n),
    .fifo_A_in_s_read(fifo_A_A_IO_L2_in_5__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_A_IO_L2_in_6__din),
    .fifo_A_out_full_n(fifo_A_A_IO_L2_in_6__full_n),
    .fifo_A_out_write(fifo_A_A_IO_L2_in_6__write),
    .fifo_A_local_out_din(fifo_A_PE_5_0__din),
    .fifo_A_local_out_full_n(fifo_A_PE_5_0__full_n),
    .fifo_A_local_out_write(fifo_A_PE_5_0__write)
  );


  (* keep_hierarchy = "yes" *) A_IO_L2_in
  A_IO_L2_in_6
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(A_IO_L2_in_6__ap_start),
    .ap_done(A_IO_L2_in_6__ap_done),
    .ap_idle(A_IO_L2_in_6__ap_idle),
    .ap_ready(A_IO_L2_in_6__ap_ready),
    .idx(64'd6),
    .fifo_A_in_s_dout(fifo_A_A_IO_L2_in_6__dout),
    .fifo_A_in_peek_dout(fifo_A_A_IO_L2_in_6__dout),
    .fifo_A_in_s_empty_n(fifo_A_A_IO_L2_in_6__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_A_IO_L2_in_6__empty_n),
    .fifo_A_in_s_read(fifo_A_A_IO_L2_in_6__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_A_IO_L2_in_7__din),
    .fifo_A_out_full_n(fifo_A_A_IO_L2_in_7__full_n),
    .fifo_A_out_write(fifo_A_A_IO_L2_in_7__write),
    .fifo_A_local_out_din(fifo_A_PE_6_0__din),
    .fifo_A_local_out_full_n(fifo_A_PE_6_0__full_n),
    .fifo_A_local_out_write(fifo_A_PE_6_0__write)
  );


  (* keep_hierarchy = "yes" *) A_IO_L2_in
  A_IO_L2_in_7
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(A_IO_L2_in_7__ap_start),
    .ap_done(A_IO_L2_in_7__ap_done),
    .ap_idle(A_IO_L2_in_7__ap_idle),
    .ap_ready(A_IO_L2_in_7__ap_ready),
    .idx(64'd7),
    .fifo_A_in_s_dout(fifo_A_A_IO_L2_in_7__dout),
    .fifo_A_in_peek_dout(fifo_A_A_IO_L2_in_7__dout),
    .fifo_A_in_s_empty_n(fifo_A_A_IO_L2_in_7__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_A_IO_L2_in_7__empty_n),
    .fifo_A_in_s_read(fifo_A_A_IO_L2_in_7__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_A_IO_L2_in_8__din),
    .fifo_A_out_full_n(fifo_A_A_IO_L2_in_8__full_n),
    .fifo_A_out_write(fifo_A_A_IO_L2_in_8__write),
    .fifo_A_local_out_din(fifo_A_PE_7_0__din),
    .fifo_A_local_out_full_n(fifo_A_PE_7_0__full_n),
    .fifo_A_local_out_write(fifo_A_PE_7_0__write)
  );


  (* keep_hierarchy = "yes" *) A_IO_L2_in
  A_IO_L2_in_8
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(A_IO_L2_in_8__ap_start),
    .ap_done(A_IO_L2_in_8__ap_done),
    .ap_idle(A_IO_L2_in_8__ap_idle),
    .ap_ready(A_IO_L2_in_8__ap_ready),
    .idx(64'd8),
    .fifo_A_in_s_dout(fifo_A_A_IO_L2_in_8__dout),
    .fifo_A_in_peek_dout(fifo_A_A_IO_L2_in_8__dout),
    .fifo_A_in_s_empty_n(fifo_A_A_IO_L2_in_8__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_A_IO_L2_in_8__empty_n),
    .fifo_A_in_s_read(fifo_A_A_IO_L2_in_8__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_A_IO_L2_in_9__din),
    .fifo_A_out_full_n(fifo_A_A_IO_L2_in_9__full_n),
    .fifo_A_out_write(fifo_A_A_IO_L2_in_9__write),
    .fifo_A_local_out_din(fifo_A_PE_8_0__din),
    .fifo_A_local_out_full_n(fifo_A_PE_8_0__full_n),
    .fifo_A_local_out_write(fifo_A_PE_8_0__write)
  );


  (* keep_hierarchy = "yes" *) A_IO_L2_in
  A_IO_L2_in_9
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(A_IO_L2_in_9__ap_start),
    .ap_done(A_IO_L2_in_9__ap_done),
    .ap_idle(A_IO_L2_in_9__ap_idle),
    .ap_ready(A_IO_L2_in_9__ap_ready),
    .idx(64'd9),
    .fifo_A_out_din(fifo_A_A_IO_L2_in_10__din),
    .fifo_A_out_full_n(fifo_A_A_IO_L2_in_10__full_n),
    .fifo_A_out_write(fifo_A_A_IO_L2_in_10__write),
    .fifo_A_in_s_dout(fifo_A_A_IO_L2_in_9__dout),
    .fifo_A_in_peek_dout(fifo_A_A_IO_L2_in_9__dout),
    .fifo_A_in_s_empty_n(fifo_A_A_IO_L2_in_9__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_A_IO_L2_in_9__empty_n),
    .fifo_A_in_s_read(fifo_A_A_IO_L2_in_9__read),
    .fifo_A_in_peek_read(),
    .fifo_A_local_out_din(fifo_A_PE_9_0__din),
    .fifo_A_local_out_full_n(fifo_A_PE_9_0__full_n),
    .fifo_A_local_out_write(fifo_A_PE_9_0__write)
  );


  (* keep_hierarchy = "yes" *) A_IO_L2_in
  A_IO_L2_in_10
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(A_IO_L2_in_10__ap_start),
    .ap_done(A_IO_L2_in_10__ap_done),
    .ap_idle(A_IO_L2_in_10__ap_idle),
    .ap_ready(A_IO_L2_in_10__ap_ready),
    .idx(64'd10),
    .fifo_A_in_s_dout(fifo_A_A_IO_L2_in_10__dout),
    .fifo_A_in_peek_dout(fifo_A_A_IO_L2_in_10__dout),
    .fifo_A_in_s_empty_n(fifo_A_A_IO_L2_in_10__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_A_IO_L2_in_10__empty_n),
    .fifo_A_in_s_read(fifo_A_A_IO_L2_in_10__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_A_IO_L2_in_11__din),
    .fifo_A_out_full_n(fifo_A_A_IO_L2_in_11__full_n),
    .fifo_A_out_write(fifo_A_A_IO_L2_in_11__write),
    .fifo_A_local_out_din(fifo_A_PE_10_0__din),
    .fifo_A_local_out_full_n(fifo_A_PE_10_0__full_n),
    .fifo_A_local_out_write(fifo_A_PE_10_0__write)
  );


  (* keep_hierarchy = "yes" *) A_IO_L2_in
  A_IO_L2_in_11
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(A_IO_L2_in_11__ap_start),
    .ap_done(A_IO_L2_in_11__ap_done),
    .ap_idle(A_IO_L2_in_11__ap_idle),
    .ap_ready(A_IO_L2_in_11__ap_ready),
    .idx(64'd11),
    .fifo_A_in_s_dout(fifo_A_A_IO_L2_in_11__dout),
    .fifo_A_in_peek_dout(fifo_A_A_IO_L2_in_11__dout),
    .fifo_A_in_s_empty_n(fifo_A_A_IO_L2_in_11__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_A_IO_L2_in_11__empty_n),
    .fifo_A_in_s_read(fifo_A_A_IO_L2_in_11__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_A_IO_L2_in_12__din),
    .fifo_A_out_full_n(fifo_A_A_IO_L2_in_12__full_n),
    .fifo_A_out_write(fifo_A_A_IO_L2_in_12__write),
    .fifo_A_local_out_din(fifo_A_PE_11_0__din),
    .fifo_A_local_out_full_n(fifo_A_PE_11_0__full_n),
    .fifo_A_local_out_write(fifo_A_PE_11_0__write)
  );


  (* keep_hierarchy = "yes" *) A_IO_L2_in
  A_IO_L2_in_12
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(A_IO_L2_in_12__ap_start),
    .ap_done(A_IO_L2_in_12__ap_done),
    .ap_idle(A_IO_L2_in_12__ap_idle),
    .ap_ready(A_IO_L2_in_12__ap_ready),
    .idx(64'd12),
    .fifo_A_in_s_dout(fifo_A_A_IO_L2_in_12__dout),
    .fifo_A_in_peek_dout(fifo_A_A_IO_L2_in_12__dout),
    .fifo_A_in_s_empty_n(fifo_A_A_IO_L2_in_12__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_A_IO_L2_in_12__empty_n),
    .fifo_A_in_s_read(fifo_A_A_IO_L2_in_12__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_A_IO_L2_in_13__din),
    .fifo_A_out_full_n(fifo_A_A_IO_L2_in_13__full_n),
    .fifo_A_out_write(fifo_A_A_IO_L2_in_13__write),
    .fifo_A_local_out_din(fifo_A_PE_12_0__din),
    .fifo_A_local_out_full_n(fifo_A_PE_12_0__full_n),
    .fifo_A_local_out_write(fifo_A_PE_12_0__write)
  );


  (* keep_hierarchy = "yes" *) A_IO_L2_in
  A_IO_L2_in_13
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(A_IO_L2_in_13__ap_start),
    .ap_done(A_IO_L2_in_13__ap_done),
    .ap_idle(A_IO_L2_in_13__ap_idle),
    .ap_ready(A_IO_L2_in_13__ap_ready),
    .idx(64'd13),
    .fifo_A_in_s_dout(fifo_A_A_IO_L2_in_13__dout),
    .fifo_A_in_peek_dout(fifo_A_A_IO_L2_in_13__dout),
    .fifo_A_in_s_empty_n(fifo_A_A_IO_L2_in_13__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_A_IO_L2_in_13__empty_n),
    .fifo_A_in_s_read(fifo_A_A_IO_L2_in_13__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_A_IO_L2_in_14__din),
    .fifo_A_out_full_n(fifo_A_A_IO_L2_in_14__full_n),
    .fifo_A_out_write(fifo_A_A_IO_L2_in_14__write),
    .fifo_A_local_out_din(fifo_A_PE_13_0__din),
    .fifo_A_local_out_full_n(fifo_A_PE_13_0__full_n),
    .fifo_A_local_out_write(fifo_A_PE_13_0__write)
  );


  (* keep_hierarchy = "yes" *) A_IO_L2_in
  A_IO_L2_in_14
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(A_IO_L2_in_14__ap_start),
    .ap_done(A_IO_L2_in_14__ap_done),
    .ap_idle(A_IO_L2_in_14__ap_idle),
    .ap_ready(A_IO_L2_in_14__ap_ready),
    .idx(64'd14),
    .fifo_A_in_s_dout(fifo_A_A_IO_L2_in_14__dout),
    .fifo_A_in_peek_dout(fifo_A_A_IO_L2_in_14__dout),
    .fifo_A_in_s_empty_n(fifo_A_A_IO_L2_in_14__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_A_IO_L2_in_14__empty_n),
    .fifo_A_in_s_read(fifo_A_A_IO_L2_in_14__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_A_IO_L2_in_15__din),
    .fifo_A_out_full_n(fifo_A_A_IO_L2_in_15__full_n),
    .fifo_A_out_write(fifo_A_A_IO_L2_in_15__write),
    .fifo_A_local_out_din(fifo_A_PE_14_0__din),
    .fifo_A_local_out_full_n(fifo_A_PE_14_0__full_n),
    .fifo_A_local_out_write(fifo_A_PE_14_0__write)
  );


  (* keep_hierarchy = "yes" *) A_IO_L2_in
  A_IO_L2_in_15
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(A_IO_L2_in_15__ap_start),
    .ap_done(A_IO_L2_in_15__ap_done),
    .ap_idle(A_IO_L2_in_15__ap_idle),
    .ap_ready(A_IO_L2_in_15__ap_ready),
    .idx(64'd15),
    .fifo_A_in_s_dout(fifo_A_A_IO_L2_in_15__dout),
    .fifo_A_in_peek_dout(fifo_A_A_IO_L2_in_15__dout),
    .fifo_A_in_s_empty_n(fifo_A_A_IO_L2_in_15__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_A_IO_L2_in_15__empty_n),
    .fifo_A_in_s_read(fifo_A_A_IO_L2_in_15__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_A_IO_L2_in_16__din),
    .fifo_A_out_full_n(fifo_A_A_IO_L2_in_16__full_n),
    .fifo_A_out_write(fifo_A_A_IO_L2_in_16__write),
    .fifo_A_local_out_din(fifo_A_PE_15_0__din),
    .fifo_A_local_out_full_n(fifo_A_PE_15_0__full_n),
    .fifo_A_local_out_write(fifo_A_PE_15_0__write)
  );


  (* keep_hierarchy = "yes" *) A_IO_L2_in
  A_IO_L2_in_16
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(A_IO_L2_in_16__ap_start),
    .ap_done(A_IO_L2_in_16__ap_done),
    .ap_idle(A_IO_L2_in_16__ap_idle),
    .ap_ready(A_IO_L2_in_16__ap_ready),
    .idx(64'd16),
    .fifo_A_in_s_dout(fifo_A_A_IO_L2_in_16__dout),
    .fifo_A_in_peek_dout(fifo_A_A_IO_L2_in_16__dout),
    .fifo_A_in_s_empty_n(fifo_A_A_IO_L2_in_16__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_A_IO_L2_in_16__empty_n),
    .fifo_A_in_s_read(fifo_A_A_IO_L2_in_16__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_A_IO_L2_in_17__din),
    .fifo_A_out_full_n(fifo_A_A_IO_L2_in_17__full_n),
    .fifo_A_out_write(fifo_A_A_IO_L2_in_17__write),
    .fifo_A_local_out_din(fifo_A_PE_16_0__din),
    .fifo_A_local_out_full_n(fifo_A_PE_16_0__full_n),
    .fifo_A_local_out_write(fifo_A_PE_16_0__write)
  );


  (* keep_hierarchy = "yes" *) A_IO_L2_in_boundary
  A_IO_L2_in_boundary_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(A_IO_L2_in_boundary_0__ap_start),
    .ap_done(A_IO_L2_in_boundary_0__ap_done),
    .ap_idle(A_IO_L2_in_boundary_0__ap_idle),
    .ap_ready(A_IO_L2_in_boundary_0__ap_ready),
    .idx(64'd17),
    .fifo_A_in_s_dout(fifo_A_A_IO_L2_in_17__dout),
    .fifo_A_in_peek_dout(fifo_A_A_IO_L2_in_17__dout),
    .fifo_A_in_s_empty_n(fifo_A_A_IO_L2_in_17__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_A_IO_L2_in_17__empty_n),
    .fifo_A_in_s_read(fifo_A_A_IO_L2_in_17__read),
    .fifo_A_in_peek_read(),
    .fifo_A_local_out_din(fifo_A_PE_17_0__din),
    .fifo_A_local_out_full_n(fifo_A_PE_17_0__full_n),
    .fifo_A_local_out_write(fifo_A_PE_17_0__write)
  );


  (* keep_hierarchy = "yes" *) A_IO_L3_in
  A_IO_L3_in_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(A_IO_L3_in_0__ap_start),
    .ap_done(A_IO_L3_in_0__ap_done),
    .ap_idle(A_IO_L3_in_0__ap_idle),
    .ap_ready(A_IO_L3_in_0__ap_ready),
    .fifo_A_local_out_din(fifo_A_A_IO_L2_in_0__din),
    .fifo_A_local_out_full_n(fifo_A_A_IO_L2_in_0__full_n),
    .fifo_A_local_out_write(fifo_A_A_IO_L2_in_0__write),
    .fifo_A_in_s_dout(fifo_A_A_IO_L3_in_serialize__dout),
    .fifo_A_in_peek_dout(fifo_A_A_IO_L3_in_serialize__dout),
    .fifo_A_in_s_empty_n(fifo_A_A_IO_L3_in_serialize__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_A_IO_L3_in_serialize__empty_n),
    .fifo_A_in_s_read(fifo_A_A_IO_L3_in_serialize__read),
    .fifo_A_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) A_IO_L3_in_serialize
  A_IO_L3_in_serialize_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(A_IO_L3_in_serialize_0__ap_start),
    .ap_done(A_IO_L3_in_serialize_0__ap_done),
    .ap_idle(A_IO_L3_in_serialize_0__ap_idle),
    .ap_ready(A_IO_L3_in_serialize_0__ap_ready),
    .m_axi_A_ARADDR(m_axi_A_ARADDR),
    .m_axi_A_ARBURST(m_axi_A_ARBURST),
    .m_axi_A_ARID(m_axi_A_ARID),
    .m_axi_A_ARLEN(m_axi_A_ARLEN),
    .m_axi_A_ARREADY(m_axi_A_ARREADY),
    .m_axi_A_ARSIZE(m_axi_A_ARSIZE),
    .m_axi_A_ARVALID(m_axi_A_ARVALID),
    .m_axi_A_AWADDR(m_axi_A_AWADDR),
    .m_axi_A_AWBURST(m_axi_A_AWBURST),
    .m_axi_A_AWID(m_axi_A_AWID),
    .m_axi_A_AWLEN(m_axi_A_AWLEN),
    .m_axi_A_AWREADY(m_axi_A_AWREADY),
    .m_axi_A_AWSIZE(m_axi_A_AWSIZE),
    .m_axi_A_AWVALID(m_axi_A_AWVALID),
    .m_axi_A_BID(m_axi_A_BID),
    .m_axi_A_BREADY(m_axi_A_BREADY),
    .m_axi_A_BRESP(m_axi_A_BRESP),
    .m_axi_A_BVALID(m_axi_A_BVALID),
    .m_axi_A_RDATA(m_axi_A_RDATA),
    .m_axi_A_RID(m_axi_A_RID),
    .m_axi_A_RLAST(m_axi_A_RLAST),
    .m_axi_A_RREADY(m_axi_A_RREADY),
    .m_axi_A_RRESP(m_axi_A_RRESP),
    .m_axi_A_RVALID(m_axi_A_RVALID),
    .m_axi_A_WDATA(m_axi_A_WDATA),
    .m_axi_A_WLAST(m_axi_A_WLAST),
    .m_axi_A_WREADY(m_axi_A_WREADY),
    .m_axi_A_WSTRB(m_axi_A_WSTRB),
    .m_axi_A_WVALID(m_axi_A_WVALID),
    .m_axi_A_ARLOCK(m_axi_A_ARLOCK),
    .m_axi_A_ARPROT(m_axi_A_ARPROT),
    .m_axi_A_ARQOS(m_axi_A_ARQOS),
    .m_axi_A_ARCACHE(m_axi_A_ARCACHE),
    .m_axi_A_AWCACHE(m_axi_A_AWCACHE),
    .m_axi_A_AWLOCK(m_axi_A_AWLOCK),
    .m_axi_A_AWPROT(m_axi_A_AWPROT),
    .m_axi_A_AWQOS(m_axi_A_AWQOS),
    .A_offset(A_IO_L3_in_serialize_0___A__q0),
    .fifo_A_local_out_din(fifo_A_A_IO_L3_in_serialize__din),
    .fifo_A_local_out_full_n(fifo_A_A_IO_L3_in_serialize__full_n),
    .fifo_A_local_out_write(fifo_A_A_IO_L3_in_serialize__write)
  );


  (* keep_hierarchy = "yes" *) A_PE_dummy_in
  A_PE_dummy_in_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(A_PE_dummy_in_0__ap_start),
    .ap_done(A_PE_dummy_in_0__ap_done),
    .ap_idle(A_PE_dummy_in_0__ap_idle),
    .ap_ready(A_PE_dummy_in_0__ap_ready),
    .idx(64'd0),
    .idy(64'd16),
    .fifo_A_in_s_dout(fifo_A_PE_0_17__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_0_17__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_0_17__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_0_17__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_0_17__read),
    .fifo_A_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) A_PE_dummy_in
  A_PE_dummy_in_1
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(A_PE_dummy_in_1__ap_start),
    .ap_done(A_PE_dummy_in_1__ap_done),
    .ap_idle(A_PE_dummy_in_1__ap_idle),
    .ap_ready(A_PE_dummy_in_1__ap_ready),
    .idx(64'd1),
    .idy(64'd16),
    .fifo_A_in_s_dout(fifo_A_PE_1_17__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_1_17__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_1_17__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_1_17__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_1_17__read),
    .fifo_A_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) A_PE_dummy_in
  A_PE_dummy_in_2
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(A_PE_dummy_in_2__ap_start),
    .ap_done(A_PE_dummy_in_2__ap_done),
    .ap_idle(A_PE_dummy_in_2__ap_idle),
    .ap_ready(A_PE_dummy_in_2__ap_ready),
    .idy(64'd16),
    .idx(64'd2),
    .fifo_A_in_s_dout(fifo_A_PE_2_17__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_2_17__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_2_17__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_2_17__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_2_17__read),
    .fifo_A_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) A_PE_dummy_in
  A_PE_dummy_in_3
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(A_PE_dummy_in_3__ap_start),
    .ap_done(A_PE_dummy_in_3__ap_done),
    .ap_idle(A_PE_dummy_in_3__ap_idle),
    .ap_ready(A_PE_dummy_in_3__ap_ready),
    .idy(64'd16),
    .idx(64'd3),
    .fifo_A_in_s_dout(fifo_A_PE_3_17__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_3_17__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_3_17__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_3_17__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_3_17__read),
    .fifo_A_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) A_PE_dummy_in
  A_PE_dummy_in_4
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(A_PE_dummy_in_4__ap_start),
    .ap_done(A_PE_dummy_in_4__ap_done),
    .ap_idle(A_PE_dummy_in_4__ap_idle),
    .ap_ready(A_PE_dummy_in_4__ap_ready),
    .idy(64'd16),
    .idx(64'd4),
    .fifo_A_in_s_dout(fifo_A_PE_4_17__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_4_17__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_4_17__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_4_17__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_4_17__read),
    .fifo_A_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) A_PE_dummy_in
  A_PE_dummy_in_5
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(A_PE_dummy_in_5__ap_start),
    .ap_done(A_PE_dummy_in_5__ap_done),
    .ap_idle(A_PE_dummy_in_5__ap_idle),
    .ap_ready(A_PE_dummy_in_5__ap_ready),
    .idy(64'd16),
    .idx(64'd5),
    .fifo_A_in_s_dout(fifo_A_PE_5_17__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_5_17__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_5_17__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_5_17__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_5_17__read),
    .fifo_A_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) A_PE_dummy_in
  A_PE_dummy_in_6
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(A_PE_dummy_in_6__ap_start),
    .ap_done(A_PE_dummy_in_6__ap_done),
    .ap_idle(A_PE_dummy_in_6__ap_idle),
    .ap_ready(A_PE_dummy_in_6__ap_ready),
    .idy(64'd16),
    .idx(64'd6),
    .fifo_A_in_s_dout(fifo_A_PE_6_17__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_6_17__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_6_17__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_6_17__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_6_17__read),
    .fifo_A_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) A_PE_dummy_in
  A_PE_dummy_in_7
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(A_PE_dummy_in_7__ap_start),
    .ap_done(A_PE_dummy_in_7__ap_done),
    .ap_idle(A_PE_dummy_in_7__ap_idle),
    .ap_ready(A_PE_dummy_in_7__ap_ready),
    .idy(64'd16),
    .idx(64'd7),
    .fifo_A_in_s_dout(fifo_A_PE_7_17__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_7_17__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_7_17__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_7_17__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_7_17__read),
    .fifo_A_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) A_PE_dummy_in
  A_PE_dummy_in_8
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(A_PE_dummy_in_8__ap_start),
    .ap_done(A_PE_dummy_in_8__ap_done),
    .ap_idle(A_PE_dummy_in_8__ap_idle),
    .ap_ready(A_PE_dummy_in_8__ap_ready),
    .idy(64'd16),
    .idx(64'd8),
    .fifo_A_in_s_dout(fifo_A_PE_8_17__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_8_17__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_8_17__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_8_17__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_8_17__read),
    .fifo_A_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) A_PE_dummy_in
  A_PE_dummy_in_9
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(A_PE_dummy_in_9__ap_start),
    .ap_done(A_PE_dummy_in_9__ap_done),
    .ap_idle(A_PE_dummy_in_9__ap_idle),
    .ap_ready(A_PE_dummy_in_9__ap_ready),
    .idy(64'd16),
    .idx(64'd9),
    .fifo_A_in_s_dout(fifo_A_PE_9_17__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_9_17__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_9_17__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_9_17__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_9_17__read),
    .fifo_A_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) A_PE_dummy_in
  A_PE_dummy_in_10
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(A_PE_dummy_in_10__ap_start),
    .ap_done(A_PE_dummy_in_10__ap_done),
    .ap_idle(A_PE_dummy_in_10__ap_idle),
    .ap_ready(A_PE_dummy_in_10__ap_ready),
    .idx(64'd10),
    .idy(64'd16),
    .fifo_A_in_s_dout(fifo_A_PE_10_17__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_10_17__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_10_17__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_10_17__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_10_17__read),
    .fifo_A_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) A_PE_dummy_in
  A_PE_dummy_in_11
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(A_PE_dummy_in_11__ap_start),
    .ap_done(A_PE_dummy_in_11__ap_done),
    .ap_idle(A_PE_dummy_in_11__ap_idle),
    .ap_ready(A_PE_dummy_in_11__ap_ready),
    .idx(64'd11),
    .idy(64'd16),
    .fifo_A_in_s_dout(fifo_A_PE_11_17__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_11_17__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_11_17__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_11_17__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_11_17__read),
    .fifo_A_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) A_PE_dummy_in
  A_PE_dummy_in_12
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(A_PE_dummy_in_12__ap_start),
    .ap_done(A_PE_dummy_in_12__ap_done),
    .ap_idle(A_PE_dummy_in_12__ap_idle),
    .ap_ready(A_PE_dummy_in_12__ap_ready),
    .idx(64'd12),
    .idy(64'd16),
    .fifo_A_in_s_dout(fifo_A_PE_12_17__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_12_17__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_12_17__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_12_17__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_12_17__read),
    .fifo_A_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) A_PE_dummy_in
  A_PE_dummy_in_13
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(A_PE_dummy_in_13__ap_start),
    .ap_done(A_PE_dummy_in_13__ap_done),
    .ap_idle(A_PE_dummy_in_13__ap_idle),
    .ap_ready(A_PE_dummy_in_13__ap_ready),
    .idx(64'd13),
    .idy(64'd16),
    .fifo_A_in_s_dout(fifo_A_PE_13_17__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_13_17__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_13_17__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_13_17__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_13_17__read),
    .fifo_A_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) A_PE_dummy_in
  A_PE_dummy_in_14
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(A_PE_dummy_in_14__ap_start),
    .ap_done(A_PE_dummy_in_14__ap_done),
    .ap_idle(A_PE_dummy_in_14__ap_idle),
    .ap_ready(A_PE_dummy_in_14__ap_ready),
    .idx(64'd14),
    .idy(64'd16),
    .fifo_A_in_s_dout(fifo_A_PE_14_17__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_14_17__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_14_17__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_14_17__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_14_17__read),
    .fifo_A_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) A_PE_dummy_in
  A_PE_dummy_in_15
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(A_PE_dummy_in_15__ap_start),
    .ap_done(A_PE_dummy_in_15__ap_done),
    .ap_idle(A_PE_dummy_in_15__ap_idle),
    .ap_ready(A_PE_dummy_in_15__ap_ready),
    .idx(64'd15),
    .idy(64'd16),
    .fifo_A_in_s_dout(fifo_A_PE_15_17__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_15_17__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_15_17__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_15_17__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_15_17__read),
    .fifo_A_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) A_PE_dummy_in
  A_PE_dummy_in_16
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(A_PE_dummy_in_16__ap_start),
    .ap_done(A_PE_dummy_in_16__ap_done),
    .ap_idle(A_PE_dummy_in_16__ap_idle),
    .ap_ready(A_PE_dummy_in_16__ap_ready),
    .idx(64'd16),
    .idy(64'd16),
    .fifo_A_in_s_dout(fifo_A_PE_16_17__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_16_17__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_16_17__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_16_17__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_16_17__read),
    .fifo_A_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) A_PE_dummy_in
  A_PE_dummy_in_17
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(A_PE_dummy_in_17__ap_start),
    .ap_done(A_PE_dummy_in_17__ap_done),
    .ap_idle(A_PE_dummy_in_17__ap_idle),
    .ap_ready(A_PE_dummy_in_17__ap_ready),
    .idy(64'd16),
    .idx(64'd17),
    .fifo_A_in_s_dout(fifo_A_PE_17_17__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_17_17__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_17_17__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_17_17__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_17_17__read),
    .fifo_A_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) B_IO_L2_in
  B_IO_L2_in_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(B_IO_L2_in_0__ap_start),
    .ap_done(B_IO_L2_in_0__ap_done),
    .ap_idle(B_IO_L2_in_0__ap_idle),
    .ap_ready(B_IO_L2_in_0__ap_ready),
    .idx(64'd0),
    .fifo_B_in_s_dout(fifo_B_B_IO_L2_in_0__dout),
    .fifo_B_in_peek_dout(fifo_B_B_IO_L2_in_0__dout),
    .fifo_B_in_s_empty_n(fifo_B_B_IO_L2_in_0__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_B_IO_L2_in_0__empty_n),
    .fifo_B_in_s_read(fifo_B_B_IO_L2_in_0__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_B_IO_L2_in_1__din),
    .fifo_B_out_full_n(fifo_B_B_IO_L2_in_1__full_n),
    .fifo_B_out_write(fifo_B_B_IO_L2_in_1__write),
    .fifo_B_local_out_din(fifo_B_PE_0_0__din),
    .fifo_B_local_out_full_n(fifo_B_PE_0_0__full_n),
    .fifo_B_local_out_write(fifo_B_PE_0_0__write)
  );


  (* keep_hierarchy = "yes" *) B_IO_L2_in
  B_IO_L2_in_1
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(B_IO_L2_in_1__ap_start),
    .ap_done(B_IO_L2_in_1__ap_done),
    .ap_idle(B_IO_L2_in_1__ap_idle),
    .ap_ready(B_IO_L2_in_1__ap_ready),
    .idx(64'd1),
    .fifo_B_in_s_dout(fifo_B_B_IO_L2_in_1__dout),
    .fifo_B_in_peek_dout(fifo_B_B_IO_L2_in_1__dout),
    .fifo_B_in_s_empty_n(fifo_B_B_IO_L2_in_1__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_B_IO_L2_in_1__empty_n),
    .fifo_B_in_s_read(fifo_B_B_IO_L2_in_1__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_B_IO_L2_in_2__din),
    .fifo_B_out_full_n(fifo_B_B_IO_L2_in_2__full_n),
    .fifo_B_out_write(fifo_B_B_IO_L2_in_2__write),
    .fifo_B_local_out_din(fifo_B_PE_0_1__din),
    .fifo_B_local_out_full_n(fifo_B_PE_0_1__full_n),
    .fifo_B_local_out_write(fifo_B_PE_0_1__write)
  );


  (* keep_hierarchy = "yes" *) B_IO_L2_in
  B_IO_L2_in_2
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(B_IO_L2_in_2__ap_start),
    .ap_done(B_IO_L2_in_2__ap_done),
    .ap_idle(B_IO_L2_in_2__ap_idle),
    .ap_ready(B_IO_L2_in_2__ap_ready),
    .idx(64'd2),
    .fifo_B_in_s_dout(fifo_B_B_IO_L2_in_2__dout),
    .fifo_B_in_peek_dout(fifo_B_B_IO_L2_in_2__dout),
    .fifo_B_in_s_empty_n(fifo_B_B_IO_L2_in_2__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_B_IO_L2_in_2__empty_n),
    .fifo_B_in_s_read(fifo_B_B_IO_L2_in_2__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_B_IO_L2_in_3__din),
    .fifo_B_out_full_n(fifo_B_B_IO_L2_in_3__full_n),
    .fifo_B_out_write(fifo_B_B_IO_L2_in_3__write),
    .fifo_B_local_out_din(fifo_B_PE_0_2__din),
    .fifo_B_local_out_full_n(fifo_B_PE_0_2__full_n),
    .fifo_B_local_out_write(fifo_B_PE_0_2__write)
  );


  (* keep_hierarchy = "yes" *) B_IO_L2_in
  B_IO_L2_in_3
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(B_IO_L2_in_3__ap_start),
    .ap_done(B_IO_L2_in_3__ap_done),
    .ap_idle(B_IO_L2_in_3__ap_idle),
    .ap_ready(B_IO_L2_in_3__ap_ready),
    .idx(64'd3),
    .fifo_B_in_s_dout(fifo_B_B_IO_L2_in_3__dout),
    .fifo_B_in_peek_dout(fifo_B_B_IO_L2_in_3__dout),
    .fifo_B_in_s_empty_n(fifo_B_B_IO_L2_in_3__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_B_IO_L2_in_3__empty_n),
    .fifo_B_in_s_read(fifo_B_B_IO_L2_in_3__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_B_IO_L2_in_4__din),
    .fifo_B_out_full_n(fifo_B_B_IO_L2_in_4__full_n),
    .fifo_B_out_write(fifo_B_B_IO_L2_in_4__write),
    .fifo_B_local_out_din(fifo_B_PE_0_3__din),
    .fifo_B_local_out_full_n(fifo_B_PE_0_3__full_n),
    .fifo_B_local_out_write(fifo_B_PE_0_3__write)
  );


  (* keep_hierarchy = "yes" *) B_IO_L2_in
  B_IO_L2_in_4
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(B_IO_L2_in_4__ap_start),
    .ap_done(B_IO_L2_in_4__ap_done),
    .ap_idle(B_IO_L2_in_4__ap_idle),
    .ap_ready(B_IO_L2_in_4__ap_ready),
    .idx(64'd4),
    .fifo_B_in_s_dout(fifo_B_B_IO_L2_in_4__dout),
    .fifo_B_in_peek_dout(fifo_B_B_IO_L2_in_4__dout),
    .fifo_B_in_s_empty_n(fifo_B_B_IO_L2_in_4__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_B_IO_L2_in_4__empty_n),
    .fifo_B_in_s_read(fifo_B_B_IO_L2_in_4__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_B_IO_L2_in_5__din),
    .fifo_B_out_full_n(fifo_B_B_IO_L2_in_5__full_n),
    .fifo_B_out_write(fifo_B_B_IO_L2_in_5__write),
    .fifo_B_local_out_din(fifo_B_PE_0_4__din),
    .fifo_B_local_out_full_n(fifo_B_PE_0_4__full_n),
    .fifo_B_local_out_write(fifo_B_PE_0_4__write)
  );


  (* keep_hierarchy = "yes" *) B_IO_L2_in
  B_IO_L2_in_5
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(B_IO_L2_in_5__ap_start),
    .ap_done(B_IO_L2_in_5__ap_done),
    .ap_idle(B_IO_L2_in_5__ap_idle),
    .ap_ready(B_IO_L2_in_5__ap_ready),
    .idx(64'd5),
    .fifo_B_in_s_dout(fifo_B_B_IO_L2_in_5__dout),
    .fifo_B_in_peek_dout(fifo_B_B_IO_L2_in_5__dout),
    .fifo_B_in_s_empty_n(fifo_B_B_IO_L2_in_5__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_B_IO_L2_in_5__empty_n),
    .fifo_B_in_s_read(fifo_B_B_IO_L2_in_5__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_B_IO_L2_in_6__din),
    .fifo_B_out_full_n(fifo_B_B_IO_L2_in_6__full_n),
    .fifo_B_out_write(fifo_B_B_IO_L2_in_6__write),
    .fifo_B_local_out_din(fifo_B_PE_0_5__din),
    .fifo_B_local_out_full_n(fifo_B_PE_0_5__full_n),
    .fifo_B_local_out_write(fifo_B_PE_0_5__write)
  );


  (* keep_hierarchy = "yes" *) B_IO_L2_in
  B_IO_L2_in_6
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(B_IO_L2_in_6__ap_start),
    .ap_done(B_IO_L2_in_6__ap_done),
    .ap_idle(B_IO_L2_in_6__ap_idle),
    .ap_ready(B_IO_L2_in_6__ap_ready),
    .idx(64'd6),
    .fifo_B_in_s_dout(fifo_B_B_IO_L2_in_6__dout),
    .fifo_B_in_peek_dout(fifo_B_B_IO_L2_in_6__dout),
    .fifo_B_in_s_empty_n(fifo_B_B_IO_L2_in_6__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_B_IO_L2_in_6__empty_n),
    .fifo_B_in_s_read(fifo_B_B_IO_L2_in_6__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_B_IO_L2_in_7__din),
    .fifo_B_out_full_n(fifo_B_B_IO_L2_in_7__full_n),
    .fifo_B_out_write(fifo_B_B_IO_L2_in_7__write),
    .fifo_B_local_out_din(fifo_B_PE_0_6__din),
    .fifo_B_local_out_full_n(fifo_B_PE_0_6__full_n),
    .fifo_B_local_out_write(fifo_B_PE_0_6__write)
  );


  (* keep_hierarchy = "yes" *) B_IO_L2_in
  B_IO_L2_in_7
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(B_IO_L2_in_7__ap_start),
    .ap_done(B_IO_L2_in_7__ap_done),
    .ap_idle(B_IO_L2_in_7__ap_idle),
    .ap_ready(B_IO_L2_in_7__ap_ready),
    .idx(64'd7),
    .fifo_B_in_s_dout(fifo_B_B_IO_L2_in_7__dout),
    .fifo_B_in_peek_dout(fifo_B_B_IO_L2_in_7__dout),
    .fifo_B_in_s_empty_n(fifo_B_B_IO_L2_in_7__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_B_IO_L2_in_7__empty_n),
    .fifo_B_in_s_read(fifo_B_B_IO_L2_in_7__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_B_IO_L2_in_8__din),
    .fifo_B_out_full_n(fifo_B_B_IO_L2_in_8__full_n),
    .fifo_B_out_write(fifo_B_B_IO_L2_in_8__write),
    .fifo_B_local_out_din(fifo_B_PE_0_7__din),
    .fifo_B_local_out_full_n(fifo_B_PE_0_7__full_n),
    .fifo_B_local_out_write(fifo_B_PE_0_7__write)
  );


  (* keep_hierarchy = "yes" *) B_IO_L2_in
  B_IO_L2_in_8
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(B_IO_L2_in_8__ap_start),
    .ap_done(B_IO_L2_in_8__ap_done),
    .ap_idle(B_IO_L2_in_8__ap_idle),
    .ap_ready(B_IO_L2_in_8__ap_ready),
    .idx(64'd8),
    .fifo_B_in_s_dout(fifo_B_B_IO_L2_in_8__dout),
    .fifo_B_in_peek_dout(fifo_B_B_IO_L2_in_8__dout),
    .fifo_B_in_s_empty_n(fifo_B_B_IO_L2_in_8__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_B_IO_L2_in_8__empty_n),
    .fifo_B_in_s_read(fifo_B_B_IO_L2_in_8__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_B_IO_L2_in_9__din),
    .fifo_B_out_full_n(fifo_B_B_IO_L2_in_9__full_n),
    .fifo_B_out_write(fifo_B_B_IO_L2_in_9__write),
    .fifo_B_local_out_din(fifo_B_PE_0_8__din),
    .fifo_B_local_out_full_n(fifo_B_PE_0_8__full_n),
    .fifo_B_local_out_write(fifo_B_PE_0_8__write)
  );


  (* keep_hierarchy = "yes" *) B_IO_L2_in
  B_IO_L2_in_9
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(B_IO_L2_in_9__ap_start),
    .ap_done(B_IO_L2_in_9__ap_done),
    .ap_idle(B_IO_L2_in_9__ap_idle),
    .ap_ready(B_IO_L2_in_9__ap_ready),
    .idx(64'd9),
    .fifo_B_out_din(fifo_B_B_IO_L2_in_10__din),
    .fifo_B_out_full_n(fifo_B_B_IO_L2_in_10__full_n),
    .fifo_B_out_write(fifo_B_B_IO_L2_in_10__write),
    .fifo_B_in_s_dout(fifo_B_B_IO_L2_in_9__dout),
    .fifo_B_in_peek_dout(fifo_B_B_IO_L2_in_9__dout),
    .fifo_B_in_s_empty_n(fifo_B_B_IO_L2_in_9__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_B_IO_L2_in_9__empty_n),
    .fifo_B_in_s_read(fifo_B_B_IO_L2_in_9__read),
    .fifo_B_in_peek_read(),
    .fifo_B_local_out_din(fifo_B_PE_0_9__din),
    .fifo_B_local_out_full_n(fifo_B_PE_0_9__full_n),
    .fifo_B_local_out_write(fifo_B_PE_0_9__write)
  );


  (* keep_hierarchy = "yes" *) B_IO_L2_in
  B_IO_L2_in_10
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(B_IO_L2_in_10__ap_start),
    .ap_done(B_IO_L2_in_10__ap_done),
    .ap_idle(B_IO_L2_in_10__ap_idle),
    .ap_ready(B_IO_L2_in_10__ap_ready),
    .idx(64'd10),
    .fifo_B_in_s_dout(fifo_B_B_IO_L2_in_10__dout),
    .fifo_B_in_peek_dout(fifo_B_B_IO_L2_in_10__dout),
    .fifo_B_in_s_empty_n(fifo_B_B_IO_L2_in_10__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_B_IO_L2_in_10__empty_n),
    .fifo_B_in_s_read(fifo_B_B_IO_L2_in_10__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_B_IO_L2_in_11__din),
    .fifo_B_out_full_n(fifo_B_B_IO_L2_in_11__full_n),
    .fifo_B_out_write(fifo_B_B_IO_L2_in_11__write),
    .fifo_B_local_out_din(fifo_B_PE_0_10__din),
    .fifo_B_local_out_full_n(fifo_B_PE_0_10__full_n),
    .fifo_B_local_out_write(fifo_B_PE_0_10__write)
  );


  (* keep_hierarchy = "yes" *) B_IO_L2_in
  B_IO_L2_in_11
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(B_IO_L2_in_11__ap_start),
    .ap_done(B_IO_L2_in_11__ap_done),
    .ap_idle(B_IO_L2_in_11__ap_idle),
    .ap_ready(B_IO_L2_in_11__ap_ready),
    .idx(64'd11),
    .fifo_B_in_s_dout(fifo_B_B_IO_L2_in_11__dout),
    .fifo_B_in_peek_dout(fifo_B_B_IO_L2_in_11__dout),
    .fifo_B_in_s_empty_n(fifo_B_B_IO_L2_in_11__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_B_IO_L2_in_11__empty_n),
    .fifo_B_in_s_read(fifo_B_B_IO_L2_in_11__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_B_IO_L2_in_12__din),
    .fifo_B_out_full_n(fifo_B_B_IO_L2_in_12__full_n),
    .fifo_B_out_write(fifo_B_B_IO_L2_in_12__write),
    .fifo_B_local_out_din(fifo_B_PE_0_11__din),
    .fifo_B_local_out_full_n(fifo_B_PE_0_11__full_n),
    .fifo_B_local_out_write(fifo_B_PE_0_11__write)
  );


  (* keep_hierarchy = "yes" *) B_IO_L2_in
  B_IO_L2_in_12
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(B_IO_L2_in_12__ap_start),
    .ap_done(B_IO_L2_in_12__ap_done),
    .ap_idle(B_IO_L2_in_12__ap_idle),
    .ap_ready(B_IO_L2_in_12__ap_ready),
    .idx(64'd12),
    .fifo_B_in_s_dout(fifo_B_B_IO_L2_in_12__dout),
    .fifo_B_in_peek_dout(fifo_B_B_IO_L2_in_12__dout),
    .fifo_B_in_s_empty_n(fifo_B_B_IO_L2_in_12__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_B_IO_L2_in_12__empty_n),
    .fifo_B_in_s_read(fifo_B_B_IO_L2_in_12__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_B_IO_L2_in_13__din),
    .fifo_B_out_full_n(fifo_B_B_IO_L2_in_13__full_n),
    .fifo_B_out_write(fifo_B_B_IO_L2_in_13__write),
    .fifo_B_local_out_din(fifo_B_PE_0_12__din),
    .fifo_B_local_out_full_n(fifo_B_PE_0_12__full_n),
    .fifo_B_local_out_write(fifo_B_PE_0_12__write)
  );


  (* keep_hierarchy = "yes" *) B_IO_L2_in
  B_IO_L2_in_13
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(B_IO_L2_in_13__ap_start),
    .ap_done(B_IO_L2_in_13__ap_done),
    .ap_idle(B_IO_L2_in_13__ap_idle),
    .ap_ready(B_IO_L2_in_13__ap_ready),
    .idx(64'd13),
    .fifo_B_in_s_dout(fifo_B_B_IO_L2_in_13__dout),
    .fifo_B_in_peek_dout(fifo_B_B_IO_L2_in_13__dout),
    .fifo_B_in_s_empty_n(fifo_B_B_IO_L2_in_13__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_B_IO_L2_in_13__empty_n),
    .fifo_B_in_s_read(fifo_B_B_IO_L2_in_13__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_B_IO_L2_in_14__din),
    .fifo_B_out_full_n(fifo_B_B_IO_L2_in_14__full_n),
    .fifo_B_out_write(fifo_B_B_IO_L2_in_14__write),
    .fifo_B_local_out_din(fifo_B_PE_0_13__din),
    .fifo_B_local_out_full_n(fifo_B_PE_0_13__full_n),
    .fifo_B_local_out_write(fifo_B_PE_0_13__write)
  );


  (* keep_hierarchy = "yes" *) B_IO_L2_in
  B_IO_L2_in_14
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(B_IO_L2_in_14__ap_start),
    .ap_done(B_IO_L2_in_14__ap_done),
    .ap_idle(B_IO_L2_in_14__ap_idle),
    .ap_ready(B_IO_L2_in_14__ap_ready),
    .idx(64'd14),
    .fifo_B_in_s_dout(fifo_B_B_IO_L2_in_14__dout),
    .fifo_B_in_peek_dout(fifo_B_B_IO_L2_in_14__dout),
    .fifo_B_in_s_empty_n(fifo_B_B_IO_L2_in_14__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_B_IO_L2_in_14__empty_n),
    .fifo_B_in_s_read(fifo_B_B_IO_L2_in_14__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_B_IO_L2_in_15__din),
    .fifo_B_out_full_n(fifo_B_B_IO_L2_in_15__full_n),
    .fifo_B_out_write(fifo_B_B_IO_L2_in_15__write),
    .fifo_B_local_out_din(fifo_B_PE_0_14__din),
    .fifo_B_local_out_full_n(fifo_B_PE_0_14__full_n),
    .fifo_B_local_out_write(fifo_B_PE_0_14__write)
  );


  (* keep_hierarchy = "yes" *) B_IO_L2_in
  B_IO_L2_in_15
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(B_IO_L2_in_15__ap_start),
    .ap_done(B_IO_L2_in_15__ap_done),
    .ap_idle(B_IO_L2_in_15__ap_idle),
    .ap_ready(B_IO_L2_in_15__ap_ready),
    .idx(64'd15),
    .fifo_B_in_s_dout(fifo_B_B_IO_L2_in_15__dout),
    .fifo_B_in_peek_dout(fifo_B_B_IO_L2_in_15__dout),
    .fifo_B_in_s_empty_n(fifo_B_B_IO_L2_in_15__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_B_IO_L2_in_15__empty_n),
    .fifo_B_in_s_read(fifo_B_B_IO_L2_in_15__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_B_IO_L2_in_16__din),
    .fifo_B_out_full_n(fifo_B_B_IO_L2_in_16__full_n),
    .fifo_B_out_write(fifo_B_B_IO_L2_in_16__write),
    .fifo_B_local_out_din(fifo_B_PE_0_15__din),
    .fifo_B_local_out_full_n(fifo_B_PE_0_15__full_n),
    .fifo_B_local_out_write(fifo_B_PE_0_15__write)
  );


  (* keep_hierarchy = "yes" *) B_IO_L2_in_boundary
  B_IO_L2_in_boundary_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(B_IO_L2_in_boundary_0__ap_start),
    .ap_done(B_IO_L2_in_boundary_0__ap_done),
    .ap_idle(B_IO_L2_in_boundary_0__ap_idle),
    .ap_ready(B_IO_L2_in_boundary_0__ap_ready),
    .idx(64'd16),
    .fifo_B_in_s_dout(fifo_B_B_IO_L2_in_16__dout),
    .fifo_B_in_peek_dout(fifo_B_B_IO_L2_in_16__dout),
    .fifo_B_in_s_empty_n(fifo_B_B_IO_L2_in_16__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_B_IO_L2_in_16__empty_n),
    .fifo_B_in_s_read(fifo_B_B_IO_L2_in_16__read),
    .fifo_B_in_peek_read(),
    .fifo_B_local_out_din(fifo_B_PE_0_16__din),
    .fifo_B_local_out_full_n(fifo_B_PE_0_16__full_n),
    .fifo_B_local_out_write(fifo_B_PE_0_16__write)
  );


  (* keep_hierarchy = "yes" *) B_IO_L3_in
  B_IO_L3_in_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(B_IO_L3_in_0__ap_start),
    .ap_done(B_IO_L3_in_0__ap_done),
    .ap_idle(B_IO_L3_in_0__ap_idle),
    .ap_ready(B_IO_L3_in_0__ap_ready),
    .fifo_B_local_out_din(fifo_B_B_IO_L2_in_0__din),
    .fifo_B_local_out_full_n(fifo_B_B_IO_L2_in_0__full_n),
    .fifo_B_local_out_write(fifo_B_B_IO_L2_in_0__write),
    .fifo_B_in_s_dout(fifo_B_B_IO_L3_in_serialize__dout),
    .fifo_B_in_peek_dout(fifo_B_B_IO_L3_in_serialize__dout),
    .fifo_B_in_s_empty_n(fifo_B_B_IO_L3_in_serialize__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_B_IO_L3_in_serialize__empty_n),
    .fifo_B_in_s_read(fifo_B_B_IO_L3_in_serialize__read),
    .fifo_B_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) B_IO_L3_in_serialize
  B_IO_L3_in_serialize_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(B_IO_L3_in_serialize_0__ap_start),
    .ap_done(B_IO_L3_in_serialize_0__ap_done),
    .ap_idle(B_IO_L3_in_serialize_0__ap_idle),
    .ap_ready(B_IO_L3_in_serialize_0__ap_ready),
    .m_axi_B_ARADDR(m_axi_B_ARADDR),
    .m_axi_B_ARBURST(m_axi_B_ARBURST),
    .m_axi_B_ARID(m_axi_B_ARID),
    .m_axi_B_ARLEN(m_axi_B_ARLEN),
    .m_axi_B_ARREADY(m_axi_B_ARREADY),
    .m_axi_B_ARSIZE(m_axi_B_ARSIZE),
    .m_axi_B_ARVALID(m_axi_B_ARVALID),
    .m_axi_B_AWADDR(m_axi_B_AWADDR),
    .m_axi_B_AWBURST(m_axi_B_AWBURST),
    .m_axi_B_AWID(m_axi_B_AWID),
    .m_axi_B_AWLEN(m_axi_B_AWLEN),
    .m_axi_B_AWREADY(m_axi_B_AWREADY),
    .m_axi_B_AWSIZE(m_axi_B_AWSIZE),
    .m_axi_B_AWVALID(m_axi_B_AWVALID),
    .m_axi_B_BID(m_axi_B_BID),
    .m_axi_B_BREADY(m_axi_B_BREADY),
    .m_axi_B_BRESP(m_axi_B_BRESP),
    .m_axi_B_BVALID(m_axi_B_BVALID),
    .m_axi_B_RDATA(m_axi_B_RDATA),
    .m_axi_B_RID(m_axi_B_RID),
    .m_axi_B_RLAST(m_axi_B_RLAST),
    .m_axi_B_RREADY(m_axi_B_RREADY),
    .m_axi_B_RRESP(m_axi_B_RRESP),
    .m_axi_B_RVALID(m_axi_B_RVALID),
    .m_axi_B_WDATA(m_axi_B_WDATA),
    .m_axi_B_WLAST(m_axi_B_WLAST),
    .m_axi_B_WREADY(m_axi_B_WREADY),
    .m_axi_B_WSTRB(m_axi_B_WSTRB),
    .m_axi_B_WVALID(m_axi_B_WVALID),
    .m_axi_B_ARLOCK(m_axi_B_ARLOCK),
    .m_axi_B_ARPROT(m_axi_B_ARPROT),
    .m_axi_B_ARQOS(m_axi_B_ARQOS),
    .m_axi_B_ARCACHE(m_axi_B_ARCACHE),
    .m_axi_B_AWCACHE(m_axi_B_AWCACHE),
    .m_axi_B_AWLOCK(m_axi_B_AWLOCK),
    .m_axi_B_AWPROT(m_axi_B_AWPROT),
    .m_axi_B_AWQOS(m_axi_B_AWQOS),
    .B_offset(B_IO_L3_in_serialize_0___B__q0),
    .fifo_B_local_out_din(fifo_B_B_IO_L3_in_serialize__din),
    .fifo_B_local_out_full_n(fifo_B_B_IO_L3_in_serialize__full_n),
    .fifo_B_local_out_write(fifo_B_B_IO_L3_in_serialize__write)
  );


  (* keep_hierarchy = "yes" *) B_PE_dummy_in
  B_PE_dummy_in_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(B_PE_dummy_in_0__ap_start),
    .ap_done(B_PE_dummy_in_0__ap_done),
    .ap_idle(B_PE_dummy_in_0__ap_idle),
    .ap_ready(B_PE_dummy_in_0__ap_ready),
    .idy(64'd0),
    .idx(64'd17),
    .fifo_B_in_s_dout(fifo_B_PE_18_0__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_18_0__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_18_0__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_18_0__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_18_0__read),
    .fifo_B_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) B_PE_dummy_in
  B_PE_dummy_in_1
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(B_PE_dummy_in_1__ap_start),
    .ap_done(B_PE_dummy_in_1__ap_done),
    .ap_idle(B_PE_dummy_in_1__ap_idle),
    .ap_ready(B_PE_dummy_in_1__ap_ready),
    .idy(64'd1),
    .idx(64'd17),
    .fifo_B_in_s_dout(fifo_B_PE_18_1__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_18_1__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_18_1__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_18_1__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_18_1__read),
    .fifo_B_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) B_PE_dummy_in
  B_PE_dummy_in_2
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(B_PE_dummy_in_2__ap_start),
    .ap_done(B_PE_dummy_in_2__ap_done),
    .ap_idle(B_PE_dummy_in_2__ap_idle),
    .ap_ready(B_PE_dummy_in_2__ap_ready),
    .idx(64'd17),
    .idy(64'd2),
    .fifo_B_in_s_dout(fifo_B_PE_18_2__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_18_2__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_18_2__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_18_2__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_18_2__read),
    .fifo_B_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) B_PE_dummy_in
  B_PE_dummy_in_3
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(B_PE_dummy_in_3__ap_start),
    .ap_done(B_PE_dummy_in_3__ap_done),
    .ap_idle(B_PE_dummy_in_3__ap_idle),
    .ap_ready(B_PE_dummy_in_3__ap_ready),
    .idx(64'd17),
    .idy(64'd3),
    .fifo_B_in_s_dout(fifo_B_PE_18_3__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_18_3__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_18_3__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_18_3__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_18_3__read),
    .fifo_B_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) B_PE_dummy_in
  B_PE_dummy_in_4
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(B_PE_dummy_in_4__ap_start),
    .ap_done(B_PE_dummy_in_4__ap_done),
    .ap_idle(B_PE_dummy_in_4__ap_idle),
    .ap_ready(B_PE_dummy_in_4__ap_ready),
    .idx(64'd17),
    .idy(64'd4),
    .fifo_B_in_s_dout(fifo_B_PE_18_4__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_18_4__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_18_4__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_18_4__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_18_4__read),
    .fifo_B_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) B_PE_dummy_in
  B_PE_dummy_in_5
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(B_PE_dummy_in_5__ap_start),
    .ap_done(B_PE_dummy_in_5__ap_done),
    .ap_idle(B_PE_dummy_in_5__ap_idle),
    .ap_ready(B_PE_dummy_in_5__ap_ready),
    .idx(64'd17),
    .idy(64'd5),
    .fifo_B_in_s_dout(fifo_B_PE_18_5__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_18_5__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_18_5__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_18_5__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_18_5__read),
    .fifo_B_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) B_PE_dummy_in
  B_PE_dummy_in_6
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(B_PE_dummy_in_6__ap_start),
    .ap_done(B_PE_dummy_in_6__ap_done),
    .ap_idle(B_PE_dummy_in_6__ap_idle),
    .ap_ready(B_PE_dummy_in_6__ap_ready),
    .idx(64'd17),
    .idy(64'd6),
    .fifo_B_in_s_dout(fifo_B_PE_18_6__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_18_6__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_18_6__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_18_6__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_18_6__read),
    .fifo_B_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) B_PE_dummy_in
  B_PE_dummy_in_7
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(B_PE_dummy_in_7__ap_start),
    .ap_done(B_PE_dummy_in_7__ap_done),
    .ap_idle(B_PE_dummy_in_7__ap_idle),
    .ap_ready(B_PE_dummy_in_7__ap_ready),
    .idx(64'd17),
    .idy(64'd7),
    .fifo_B_in_s_dout(fifo_B_PE_18_7__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_18_7__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_18_7__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_18_7__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_18_7__read),
    .fifo_B_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) B_PE_dummy_in
  B_PE_dummy_in_8
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(B_PE_dummy_in_8__ap_start),
    .ap_done(B_PE_dummy_in_8__ap_done),
    .ap_idle(B_PE_dummy_in_8__ap_idle),
    .ap_ready(B_PE_dummy_in_8__ap_ready),
    .idx(64'd17),
    .idy(64'd8),
    .fifo_B_in_s_dout(fifo_B_PE_18_8__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_18_8__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_18_8__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_18_8__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_18_8__read),
    .fifo_B_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) B_PE_dummy_in
  B_PE_dummy_in_9
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(B_PE_dummy_in_9__ap_start),
    .ap_done(B_PE_dummy_in_9__ap_done),
    .ap_idle(B_PE_dummy_in_9__ap_idle),
    .ap_ready(B_PE_dummy_in_9__ap_ready),
    .idx(64'd17),
    .idy(64'd9),
    .fifo_B_in_s_dout(fifo_B_PE_18_9__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_18_9__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_18_9__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_18_9__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_18_9__read),
    .fifo_B_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) B_PE_dummy_in
  B_PE_dummy_in_10
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(B_PE_dummy_in_10__ap_start),
    .ap_done(B_PE_dummy_in_10__ap_done),
    .ap_idle(B_PE_dummy_in_10__ap_idle),
    .ap_ready(B_PE_dummy_in_10__ap_ready),
    .idy(64'd10),
    .idx(64'd17),
    .fifo_B_in_s_dout(fifo_B_PE_18_10__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_18_10__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_18_10__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_18_10__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_18_10__read),
    .fifo_B_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) B_PE_dummy_in
  B_PE_dummy_in_11
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(B_PE_dummy_in_11__ap_start),
    .ap_done(B_PE_dummy_in_11__ap_done),
    .ap_idle(B_PE_dummy_in_11__ap_idle),
    .ap_ready(B_PE_dummy_in_11__ap_ready),
    .idy(64'd11),
    .idx(64'd17),
    .fifo_B_in_s_dout(fifo_B_PE_18_11__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_18_11__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_18_11__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_18_11__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_18_11__read),
    .fifo_B_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) B_PE_dummy_in
  B_PE_dummy_in_12
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(B_PE_dummy_in_12__ap_start),
    .ap_done(B_PE_dummy_in_12__ap_done),
    .ap_idle(B_PE_dummy_in_12__ap_idle),
    .ap_ready(B_PE_dummy_in_12__ap_ready),
    .idy(64'd12),
    .idx(64'd17),
    .fifo_B_in_s_dout(fifo_B_PE_18_12__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_18_12__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_18_12__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_18_12__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_18_12__read),
    .fifo_B_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) B_PE_dummy_in
  B_PE_dummy_in_13
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(B_PE_dummy_in_13__ap_start),
    .ap_done(B_PE_dummy_in_13__ap_done),
    .ap_idle(B_PE_dummy_in_13__ap_idle),
    .ap_ready(B_PE_dummy_in_13__ap_ready),
    .idy(64'd13),
    .idx(64'd17),
    .fifo_B_in_s_dout(fifo_B_PE_18_13__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_18_13__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_18_13__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_18_13__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_18_13__read),
    .fifo_B_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) B_PE_dummy_in
  B_PE_dummy_in_14
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(B_PE_dummy_in_14__ap_start),
    .ap_done(B_PE_dummy_in_14__ap_done),
    .ap_idle(B_PE_dummy_in_14__ap_idle),
    .ap_ready(B_PE_dummy_in_14__ap_ready),
    .idy(64'd14),
    .idx(64'd17),
    .fifo_B_in_s_dout(fifo_B_PE_18_14__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_18_14__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_18_14__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_18_14__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_18_14__read),
    .fifo_B_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) B_PE_dummy_in
  B_PE_dummy_in_15
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(B_PE_dummy_in_15__ap_start),
    .ap_done(B_PE_dummy_in_15__ap_done),
    .ap_idle(B_PE_dummy_in_15__ap_idle),
    .ap_ready(B_PE_dummy_in_15__ap_ready),
    .idy(64'd15),
    .idx(64'd17),
    .fifo_B_in_s_dout(fifo_B_PE_18_15__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_18_15__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_18_15__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_18_15__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_18_15__read),
    .fifo_B_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) B_PE_dummy_in
  B_PE_dummy_in_16
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(B_PE_dummy_in_16__ap_start),
    .ap_done(B_PE_dummy_in_16__ap_done),
    .ap_idle(B_PE_dummy_in_16__ap_idle),
    .ap_ready(B_PE_dummy_in_16__ap_ready),
    .idy(64'd16),
    .idx(64'd17),
    .fifo_B_in_s_dout(fifo_B_PE_18_16__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_18_16__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_18_16__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_18_16__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_18_16__read),
    .fifo_B_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_boundary_wrapper
  C_drain_IO_L1_out_boundary_wrapper_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_boundary_wrapper_0__ap_start),
    .ap_done(C_drain_IO_L1_out_boundary_wrapper_0__ap_done),
    .ap_idle(C_drain_IO_L1_out_boundary_wrapper_0__ap_idle),
    .ap_ready(C_drain_IO_L1_out_boundary_wrapper_0__ap_ready),
    .idx(64'd0),
    .idy(64'd17),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_0_17__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_0_17__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_0_17__write),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_17_0__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_17_0__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_17_0__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_17_0__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_17_0__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_boundary_wrapper
  C_drain_IO_L1_out_boundary_wrapper_1
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_boundary_wrapper_1__ap_start),
    .ap_done(C_drain_IO_L1_out_boundary_wrapper_1__ap_done),
    .ap_idle(C_drain_IO_L1_out_boundary_wrapper_1__ap_idle),
    .ap_ready(C_drain_IO_L1_out_boundary_wrapper_1__ap_ready),
    .idx(64'd1),
    .idy(64'd17),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_1_17__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_1_17__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_1_17__write),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_17_1__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_17_1__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_17_1__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_17_1__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_17_1__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_boundary_wrapper
  C_drain_IO_L1_out_boundary_wrapper_2
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_boundary_wrapper_2__ap_start),
    .ap_done(C_drain_IO_L1_out_boundary_wrapper_2__ap_done),
    .ap_idle(C_drain_IO_L1_out_boundary_wrapper_2__ap_idle),
    .ap_ready(C_drain_IO_L1_out_boundary_wrapper_2__ap_ready),
    .idy(64'd17),
    .idx(64'd2),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_2_17__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_2_17__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_2_17__write),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_17_2__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_17_2__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_17_2__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_17_2__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_17_2__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_boundary_wrapper
  C_drain_IO_L1_out_boundary_wrapper_3
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_boundary_wrapper_3__ap_start),
    .ap_done(C_drain_IO_L1_out_boundary_wrapper_3__ap_done),
    .ap_idle(C_drain_IO_L1_out_boundary_wrapper_3__ap_idle),
    .ap_ready(C_drain_IO_L1_out_boundary_wrapper_3__ap_ready),
    .idy(64'd17),
    .idx(64'd3),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_3_17__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_3_17__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_3_17__write),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_17_3__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_17_3__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_17_3__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_17_3__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_17_3__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_boundary_wrapper
  C_drain_IO_L1_out_boundary_wrapper_4
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_boundary_wrapper_4__ap_start),
    .ap_done(C_drain_IO_L1_out_boundary_wrapper_4__ap_done),
    .ap_idle(C_drain_IO_L1_out_boundary_wrapper_4__ap_idle),
    .ap_ready(C_drain_IO_L1_out_boundary_wrapper_4__ap_ready),
    .idy(64'd17),
    .idx(64'd4),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_4_17__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_4_17__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_4_17__write),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_17_4__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_17_4__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_17_4__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_17_4__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_17_4__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_boundary_wrapper
  C_drain_IO_L1_out_boundary_wrapper_5
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_boundary_wrapper_5__ap_start),
    .ap_done(C_drain_IO_L1_out_boundary_wrapper_5__ap_done),
    .ap_idle(C_drain_IO_L1_out_boundary_wrapper_5__ap_idle),
    .ap_ready(C_drain_IO_L1_out_boundary_wrapper_5__ap_ready),
    .idy(64'd17),
    .idx(64'd5),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_5_17__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_5_17__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_5_17__write),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_17_5__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_17_5__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_17_5__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_17_5__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_17_5__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_boundary_wrapper
  C_drain_IO_L1_out_boundary_wrapper_6
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_boundary_wrapper_6__ap_start),
    .ap_done(C_drain_IO_L1_out_boundary_wrapper_6__ap_done),
    .ap_idle(C_drain_IO_L1_out_boundary_wrapper_6__ap_idle),
    .ap_ready(C_drain_IO_L1_out_boundary_wrapper_6__ap_ready),
    .idy(64'd17),
    .idx(64'd6),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_6_17__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_6_17__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_6_17__write),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_17_6__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_17_6__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_17_6__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_17_6__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_17_6__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_boundary_wrapper
  C_drain_IO_L1_out_boundary_wrapper_7
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_boundary_wrapper_7__ap_start),
    .ap_done(C_drain_IO_L1_out_boundary_wrapper_7__ap_done),
    .ap_idle(C_drain_IO_L1_out_boundary_wrapper_7__ap_idle),
    .ap_ready(C_drain_IO_L1_out_boundary_wrapper_7__ap_ready),
    .idy(64'd17),
    .idx(64'd7),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_7_17__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_7_17__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_7_17__write),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_17_7__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_17_7__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_17_7__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_17_7__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_17_7__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_boundary_wrapper
  C_drain_IO_L1_out_boundary_wrapper_8
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_boundary_wrapper_8__ap_start),
    .ap_done(C_drain_IO_L1_out_boundary_wrapper_8__ap_done),
    .ap_idle(C_drain_IO_L1_out_boundary_wrapper_8__ap_idle),
    .ap_ready(C_drain_IO_L1_out_boundary_wrapper_8__ap_ready),
    .idy(64'd17),
    .idx(64'd8),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_8_17__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_8_17__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_8_17__write),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_17_8__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_17_8__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_17_8__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_17_8__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_17_8__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_boundary_wrapper
  C_drain_IO_L1_out_boundary_wrapper_9
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_boundary_wrapper_9__ap_start),
    .ap_done(C_drain_IO_L1_out_boundary_wrapper_9__ap_done),
    .ap_idle(C_drain_IO_L1_out_boundary_wrapper_9__ap_idle),
    .ap_ready(C_drain_IO_L1_out_boundary_wrapper_9__ap_ready),
    .idy(64'd17),
    .idx(64'd9),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_9_17__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_9_17__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_9_17__write),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_17_9__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_17_9__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_17_9__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_17_9__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_17_9__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_boundary_wrapper
  C_drain_IO_L1_out_boundary_wrapper_10
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_boundary_wrapper_10__ap_start),
    .ap_done(C_drain_IO_L1_out_boundary_wrapper_10__ap_done),
    .ap_idle(C_drain_IO_L1_out_boundary_wrapper_10__ap_idle),
    .ap_ready(C_drain_IO_L1_out_boundary_wrapper_10__ap_ready),
    .idx(64'd10),
    .idy(64'd17),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_10_17__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_10_17__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_10_17__write),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_17_10__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_17_10__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_17_10__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_17_10__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_17_10__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_boundary_wrapper
  C_drain_IO_L1_out_boundary_wrapper_11
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_boundary_wrapper_11__ap_start),
    .ap_done(C_drain_IO_L1_out_boundary_wrapper_11__ap_done),
    .ap_idle(C_drain_IO_L1_out_boundary_wrapper_11__ap_idle),
    .ap_ready(C_drain_IO_L1_out_boundary_wrapper_11__ap_ready),
    .idx(64'd11),
    .idy(64'd17),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_11_17__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_11_17__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_11_17__write),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_17_11__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_17_11__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_17_11__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_17_11__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_17_11__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_boundary_wrapper
  C_drain_IO_L1_out_boundary_wrapper_12
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_boundary_wrapper_12__ap_start),
    .ap_done(C_drain_IO_L1_out_boundary_wrapper_12__ap_done),
    .ap_idle(C_drain_IO_L1_out_boundary_wrapper_12__ap_idle),
    .ap_ready(C_drain_IO_L1_out_boundary_wrapper_12__ap_ready),
    .idx(64'd12),
    .idy(64'd17),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_12_17__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_12_17__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_12_17__write),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_17_12__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_17_12__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_17_12__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_17_12__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_17_12__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_boundary_wrapper
  C_drain_IO_L1_out_boundary_wrapper_13
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_boundary_wrapper_13__ap_start),
    .ap_done(C_drain_IO_L1_out_boundary_wrapper_13__ap_done),
    .ap_idle(C_drain_IO_L1_out_boundary_wrapper_13__ap_idle),
    .ap_ready(C_drain_IO_L1_out_boundary_wrapper_13__ap_ready),
    .idx(64'd13),
    .idy(64'd17),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_13_17__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_13_17__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_13_17__write),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_17_13__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_17_13__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_17_13__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_17_13__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_17_13__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_boundary_wrapper
  C_drain_IO_L1_out_boundary_wrapper_14
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_boundary_wrapper_14__ap_start),
    .ap_done(C_drain_IO_L1_out_boundary_wrapper_14__ap_done),
    .ap_idle(C_drain_IO_L1_out_boundary_wrapper_14__ap_idle),
    .ap_ready(C_drain_IO_L1_out_boundary_wrapper_14__ap_ready),
    .idx(64'd14),
    .idy(64'd17),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_14_17__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_14_17__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_14_17__write),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_17_14__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_17_14__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_17_14__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_17_14__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_17_14__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_boundary_wrapper
  C_drain_IO_L1_out_boundary_wrapper_15
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_boundary_wrapper_15__ap_start),
    .ap_done(C_drain_IO_L1_out_boundary_wrapper_15__ap_done),
    .ap_idle(C_drain_IO_L1_out_boundary_wrapper_15__ap_idle),
    .ap_ready(C_drain_IO_L1_out_boundary_wrapper_15__ap_ready),
    .idx(64'd15),
    .idy(64'd17),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_15_17__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_15_17__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_15_17__write),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_17_15__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_17_15__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_17_15__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_17_15__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_17_15__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_boundary_wrapper
  C_drain_IO_L1_out_boundary_wrapper_16
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_boundary_wrapper_16__ap_start),
    .ap_done(C_drain_IO_L1_out_boundary_wrapper_16__ap_done),
    .ap_idle(C_drain_IO_L1_out_boundary_wrapper_16__ap_idle),
    .ap_ready(C_drain_IO_L1_out_boundary_wrapper_16__ap_ready),
    .idx(64'd16),
    .idy(64'd17),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_16_17__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_16_17__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_16_17__write),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_17_16__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_17_16__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_17_16__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_17_16__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_17_16__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_0__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_0__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_0__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_0__ap_ready),
    .idx(64'd0),
    .idy(64'd0),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_0_0__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_0_0__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_0_0__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_0_1__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_0_1__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_1__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_1__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_0_1__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_0_0__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_0_0__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_0_0__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_0_0__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_0_0__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_1
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_1__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_1__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_1__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_1__ap_ready),
    .idx(64'd0),
    .idy(64'd1),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_0_1__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_0_1__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_0_1__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_0_2__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_0_2__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_2__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_2__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_0_2__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_1_0__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_1_0__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_1_0__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_1_0__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_1_0__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_2
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_2__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_2__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_2__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_2__ap_ready),
    .idx(64'd0),
    .idy(64'd2),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_0_2__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_0_2__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_0_2__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_0_3__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_0_3__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_3__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_3__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_0_3__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_2_0__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_2_0__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_2_0__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_2_0__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_2_0__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_3
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_3__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_3__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_3__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_3__ap_ready),
    .idx(64'd0),
    .idy(64'd3),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_0_3__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_0_3__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_0_3__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_0_4__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_0_4__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_4__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_4__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_0_4__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_3_0__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_3_0__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_3_0__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_3_0__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_3_0__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_4
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_4__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_4__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_4__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_4__ap_ready),
    .idx(64'd0),
    .idy(64'd4),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_0_4__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_0_4__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_0_4__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_0_5__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_0_5__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_5__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_5__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_0_5__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_4_0__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_4_0__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_4_0__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_4_0__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_4_0__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_5
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_5__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_5__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_5__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_5__ap_ready),
    .idx(64'd0),
    .idy(64'd5),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_0_5__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_0_5__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_0_5__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_0_6__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_0_6__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_6__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_6__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_0_6__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_5_0__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_5_0__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_5_0__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_5_0__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_5_0__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_6
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_6__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_6__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_6__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_6__ap_ready),
    .idx(64'd0),
    .idy(64'd6),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_0_6__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_0_6__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_0_6__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_0_7__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_0_7__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_7__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_7__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_0_7__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_6_0__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_6_0__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_6_0__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_6_0__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_6_0__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_7
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_7__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_7__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_7__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_7__ap_ready),
    .idx(64'd0),
    .idy(64'd7),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_0_7__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_0_7__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_0_7__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_0_8__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_0_8__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_8__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_8__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_0_8__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_7_0__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_7_0__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_7_0__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_7_0__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_7_0__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_8
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_8__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_8__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_8__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_8__ap_ready),
    .idx(64'd0),
    .idy(64'd8),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_0_8__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_0_8__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_0_8__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_0_9__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_0_9__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_9__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_9__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_0_9__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_8_0__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_8_0__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_8_0__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_8_0__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_8_0__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_9
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_9__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_9__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_9__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_9__ap_ready),
    .idx(64'd0),
    .idy(64'd9),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_0_10__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_0_10__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_10__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_10__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_0_10__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_0_9__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_0_9__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_0_9__write),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_9_0__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_9_0__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_9_0__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_9_0__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_9_0__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_10
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_10__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_10__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_10__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_10__ap_ready),
    .idx(64'd0),
    .idy(64'd10),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_0_10__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_0_10__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_0_10__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_0_11__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_0_11__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_11__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_11__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_0_11__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_10_0__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_10_0__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_10_0__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_10_0__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_10_0__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_11
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_11__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_11__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_11__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_11__ap_ready),
    .idx(64'd0),
    .idy(64'd11),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_0_11__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_0_11__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_0_11__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_0_12__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_0_12__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_12__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_12__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_0_12__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_11_0__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_11_0__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_11_0__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_11_0__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_11_0__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_12
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_12__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_12__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_12__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_12__ap_ready),
    .idx(64'd0),
    .idy(64'd12),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_0_12__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_0_12__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_0_12__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_0_13__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_0_13__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_13__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_13__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_0_13__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_12_0__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_12_0__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_12_0__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_12_0__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_12_0__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_13
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_13__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_13__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_13__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_13__ap_ready),
    .idx(64'd0),
    .idy(64'd13),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_0_13__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_0_13__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_0_13__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_0_14__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_0_14__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_14__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_14__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_0_14__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_13_0__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_13_0__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_13_0__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_13_0__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_13_0__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_14
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_14__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_14__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_14__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_14__ap_ready),
    .idx(64'd0),
    .idy(64'd14),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_0_14__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_0_14__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_0_14__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_0_15__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_0_15__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_15__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_15__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_0_15__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_14_0__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_14_0__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_14_0__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_14_0__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_14_0__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_15
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_15__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_15__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_15__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_15__ap_ready),
    .idx(64'd0),
    .idy(64'd15),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_0_15__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_0_15__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_0_15__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_0_16__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_0_16__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_16__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_16__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_0_16__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_15_0__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_15_0__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_15_0__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_15_0__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_15_0__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_16
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_16__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_16__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_16__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_16__ap_ready),
    .idx(64'd0),
    .idy(64'd16),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_0_16__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_0_16__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_0_16__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_0_17__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_0_17__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_17__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_17__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_0_17__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_16_0__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_16_0__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_16_0__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_16_0__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_16_0__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_17
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_17__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_17__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_17__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_17__ap_ready),
    .idy(64'd0),
    .idx(64'd1),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_1_0__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_1_0__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_1_0__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_1_1__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_1_1__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_1__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_1__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_1_1__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_0_1__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_0_1__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_0_1__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_0_1__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_0_1__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_18
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_18__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_18__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_18__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_18__ap_ready),
    .idx(64'd1),
    .idy(64'd1),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_1_1__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_1_1__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_1_1__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_1_2__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_1_2__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_2__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_2__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_1_2__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_1_1__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_1_1__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_1_1__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_1_1__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_1_1__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_19
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_19__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_19__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_19__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_19__ap_ready),
    .idx(64'd1),
    .idy(64'd2),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_1_2__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_1_2__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_1_2__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_1_3__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_1_3__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_3__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_3__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_1_3__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_2_1__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_2_1__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_2_1__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_2_1__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_2_1__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_20
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_20__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_20__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_20__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_20__ap_ready),
    .idx(64'd1),
    .idy(64'd3),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_1_3__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_1_3__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_1_3__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_1_4__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_1_4__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_4__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_4__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_1_4__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_3_1__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_3_1__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_3_1__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_3_1__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_3_1__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_21
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_21__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_21__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_21__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_21__ap_ready),
    .idx(64'd1),
    .idy(64'd4),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_1_4__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_1_4__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_1_4__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_1_5__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_1_5__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_5__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_5__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_1_5__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_4_1__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_4_1__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_4_1__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_4_1__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_4_1__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_22
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_22__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_22__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_22__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_22__ap_ready),
    .idx(64'd1),
    .idy(64'd5),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_1_5__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_1_5__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_1_5__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_1_6__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_1_6__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_6__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_6__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_1_6__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_5_1__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_5_1__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_5_1__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_5_1__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_5_1__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_23
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_23__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_23__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_23__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_23__ap_ready),
    .idx(64'd1),
    .idy(64'd6),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_1_6__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_1_6__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_1_6__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_1_7__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_1_7__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_7__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_7__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_1_7__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_6_1__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_6_1__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_6_1__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_6_1__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_6_1__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_24
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_24__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_24__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_24__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_24__ap_ready),
    .idx(64'd1),
    .idy(64'd7),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_1_7__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_1_7__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_1_7__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_1_8__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_1_8__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_8__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_8__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_1_8__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_7_1__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_7_1__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_7_1__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_7_1__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_7_1__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_25
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_25__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_25__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_25__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_25__ap_ready),
    .idx(64'd1),
    .idy(64'd8),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_1_8__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_1_8__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_1_8__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_1_9__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_1_9__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_9__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_9__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_1_9__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_8_1__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_8_1__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_8_1__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_8_1__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_8_1__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_26
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_26__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_26__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_26__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_26__ap_ready),
    .idx(64'd1),
    .idy(64'd9),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_1_10__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_1_10__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_10__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_10__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_1_10__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_1_9__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_1_9__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_1_9__write),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_9_1__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_9_1__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_9_1__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_9_1__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_9_1__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_27
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_27__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_27__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_27__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_27__ap_ready),
    .idx(64'd1),
    .idy(64'd10),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_1_10__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_1_10__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_1_10__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_1_11__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_1_11__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_11__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_11__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_1_11__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_10_1__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_10_1__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_10_1__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_10_1__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_10_1__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_28
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_28__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_28__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_28__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_28__ap_ready),
    .idx(64'd1),
    .idy(64'd11),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_1_11__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_1_11__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_1_11__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_1_12__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_1_12__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_12__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_12__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_1_12__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_11_1__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_11_1__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_11_1__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_11_1__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_11_1__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_29
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_29__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_29__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_29__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_29__ap_ready),
    .idx(64'd1),
    .idy(64'd12),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_1_12__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_1_12__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_1_12__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_1_13__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_1_13__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_13__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_13__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_1_13__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_12_1__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_12_1__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_12_1__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_12_1__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_12_1__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_30
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_30__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_30__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_30__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_30__ap_ready),
    .idx(64'd1),
    .idy(64'd13),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_1_13__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_1_13__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_1_13__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_1_14__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_1_14__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_14__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_14__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_1_14__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_13_1__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_13_1__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_13_1__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_13_1__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_13_1__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_31
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_31__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_31__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_31__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_31__ap_ready),
    .idx(64'd1),
    .idy(64'd14),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_1_14__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_1_14__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_1_14__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_1_15__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_1_15__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_15__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_15__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_1_15__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_14_1__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_14_1__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_14_1__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_14_1__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_14_1__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_32
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_32__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_32__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_32__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_32__ap_ready),
    .idx(64'd1),
    .idy(64'd15),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_1_15__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_1_15__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_1_15__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_1_16__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_1_16__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_16__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_16__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_1_16__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_15_1__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_15_1__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_15_1__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_15_1__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_15_1__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_33
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_33__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_33__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_33__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_33__ap_ready),
    .idx(64'd1),
    .idy(64'd16),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_1_16__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_1_16__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_1_16__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_1_17__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_1_17__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_17__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_17__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_1_17__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_16_1__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_16_1__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_16_1__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_16_1__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_16_1__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_34
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_34__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_34__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_34__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_34__ap_ready),
    .idy(64'd0),
    .idx(64'd2),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_2_0__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_2_0__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_2_0__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_2_1__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_2_1__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_1__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_1__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_2_1__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_0_2__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_0_2__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_0_2__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_0_2__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_0_2__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_35
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_35__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_35__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_35__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_35__ap_ready),
    .idy(64'd1),
    .idx(64'd2),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_2_1__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_2_1__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_2_1__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_2_2__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_2_2__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_2__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_2__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_2_2__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_1_2__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_1_2__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_1_2__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_1_2__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_1_2__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_36
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_36__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_36__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_36__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_36__ap_ready),
    .idx(64'd2),
    .idy(64'd2),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_2_2__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_2_2__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_2_2__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_2_3__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_2_3__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_3__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_3__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_2_3__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_2_2__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_2_2__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_2_2__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_2_2__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_2_2__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_37
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_37__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_37__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_37__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_37__ap_ready),
    .idx(64'd2),
    .idy(64'd3),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_2_3__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_2_3__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_2_3__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_2_4__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_2_4__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_4__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_4__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_2_4__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_3_2__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_3_2__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_3_2__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_3_2__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_3_2__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_38
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_38__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_38__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_38__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_38__ap_ready),
    .idx(64'd2),
    .idy(64'd4),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_2_4__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_2_4__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_2_4__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_2_5__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_2_5__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_5__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_5__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_2_5__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_4_2__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_4_2__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_4_2__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_4_2__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_4_2__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_39
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_39__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_39__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_39__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_39__ap_ready),
    .idx(64'd2),
    .idy(64'd5),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_2_5__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_2_5__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_2_5__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_2_6__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_2_6__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_6__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_6__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_2_6__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_5_2__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_5_2__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_5_2__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_5_2__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_5_2__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_40
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_40__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_40__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_40__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_40__ap_ready),
    .idx(64'd2),
    .idy(64'd6),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_2_6__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_2_6__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_2_6__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_2_7__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_2_7__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_7__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_7__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_2_7__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_6_2__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_6_2__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_6_2__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_6_2__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_6_2__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_41
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_41__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_41__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_41__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_41__ap_ready),
    .idx(64'd2),
    .idy(64'd7),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_2_7__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_2_7__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_2_7__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_2_8__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_2_8__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_8__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_8__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_2_8__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_7_2__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_7_2__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_7_2__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_7_2__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_7_2__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_42
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_42__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_42__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_42__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_42__ap_ready),
    .idx(64'd2),
    .idy(64'd8),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_2_8__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_2_8__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_2_8__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_2_9__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_2_9__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_9__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_9__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_2_9__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_8_2__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_8_2__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_8_2__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_8_2__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_8_2__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_43
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_43__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_43__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_43__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_43__ap_ready),
    .idx(64'd2),
    .idy(64'd9),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_2_10__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_2_10__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_10__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_10__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_2_10__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_2_9__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_2_9__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_2_9__write),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_9_2__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_9_2__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_9_2__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_9_2__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_9_2__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_44
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_44__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_44__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_44__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_44__ap_ready),
    .idy(64'd10),
    .idx(64'd2),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_2_10__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_2_10__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_2_10__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_2_11__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_2_11__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_11__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_11__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_2_11__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_10_2__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_10_2__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_10_2__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_10_2__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_10_2__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_45
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_45__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_45__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_45__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_45__ap_ready),
    .idy(64'd11),
    .idx(64'd2),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_2_11__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_2_11__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_2_11__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_2_12__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_2_12__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_12__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_12__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_2_12__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_11_2__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_11_2__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_11_2__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_11_2__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_11_2__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_46
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_46__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_46__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_46__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_46__ap_ready),
    .idy(64'd12),
    .idx(64'd2),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_2_12__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_2_12__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_2_12__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_2_13__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_2_13__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_13__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_13__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_2_13__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_12_2__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_12_2__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_12_2__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_12_2__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_12_2__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_47
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_47__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_47__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_47__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_47__ap_ready),
    .idy(64'd13),
    .idx(64'd2),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_2_13__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_2_13__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_2_13__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_2_14__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_2_14__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_14__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_14__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_2_14__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_13_2__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_13_2__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_13_2__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_13_2__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_13_2__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_48
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_48__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_48__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_48__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_48__ap_ready),
    .idy(64'd14),
    .idx(64'd2),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_2_14__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_2_14__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_2_14__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_2_15__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_2_15__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_15__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_15__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_2_15__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_14_2__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_14_2__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_14_2__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_14_2__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_14_2__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_49
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_49__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_49__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_49__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_49__ap_ready),
    .idy(64'd15),
    .idx(64'd2),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_2_15__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_2_15__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_2_15__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_2_16__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_2_16__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_16__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_16__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_2_16__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_15_2__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_15_2__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_15_2__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_15_2__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_15_2__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_50
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_50__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_50__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_50__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_50__ap_ready),
    .idy(64'd16),
    .idx(64'd2),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_2_16__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_2_16__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_2_16__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_2_17__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_2_17__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_17__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_17__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_2_17__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_16_2__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_16_2__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_16_2__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_16_2__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_16_2__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_51
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_51__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_51__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_51__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_51__ap_ready),
    .idy(64'd0),
    .idx(64'd3),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_3_0__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_3_0__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_3_0__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_3_1__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_3_1__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_1__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_1__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_3_1__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_0_3__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_0_3__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_0_3__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_0_3__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_0_3__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_52
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_52__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_52__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_52__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_52__ap_ready),
    .idy(64'd1),
    .idx(64'd3),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_3_1__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_3_1__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_3_1__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_3_2__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_3_2__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_2__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_2__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_3_2__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_1_3__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_1_3__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_1_3__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_1_3__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_1_3__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_53
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_53__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_53__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_53__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_53__ap_ready),
    .idy(64'd2),
    .idx(64'd3),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_3_2__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_3_2__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_3_2__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_3_3__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_3_3__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_3__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_3__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_3_3__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_2_3__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_2_3__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_2_3__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_2_3__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_2_3__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_54
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_54__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_54__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_54__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_54__ap_ready),
    .idx(64'd3),
    .idy(64'd3),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_3_3__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_3_3__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_3_3__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_3_4__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_3_4__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_4__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_4__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_3_4__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_3_3__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_3_3__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_3_3__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_3_3__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_3_3__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_55
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_55__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_55__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_55__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_55__ap_ready),
    .idx(64'd3),
    .idy(64'd4),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_3_4__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_3_4__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_3_4__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_3_5__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_3_5__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_5__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_5__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_3_5__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_4_3__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_4_3__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_4_3__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_4_3__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_4_3__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_56
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_56__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_56__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_56__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_56__ap_ready),
    .idx(64'd3),
    .idy(64'd5),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_3_5__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_3_5__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_3_5__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_3_6__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_3_6__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_6__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_6__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_3_6__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_5_3__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_5_3__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_5_3__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_5_3__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_5_3__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_57
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_57__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_57__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_57__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_57__ap_ready),
    .idx(64'd3),
    .idy(64'd6),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_3_6__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_3_6__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_3_6__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_3_7__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_3_7__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_7__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_7__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_3_7__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_6_3__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_6_3__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_6_3__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_6_3__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_6_3__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_58
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_58__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_58__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_58__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_58__ap_ready),
    .idx(64'd3),
    .idy(64'd7),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_3_7__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_3_7__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_3_7__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_3_8__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_3_8__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_8__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_8__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_3_8__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_7_3__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_7_3__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_7_3__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_7_3__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_7_3__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_59
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_59__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_59__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_59__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_59__ap_ready),
    .idx(64'd3),
    .idy(64'd8),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_3_8__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_3_8__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_3_8__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_3_9__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_3_9__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_9__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_9__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_3_9__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_8_3__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_8_3__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_8_3__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_8_3__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_8_3__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_60
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_60__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_60__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_60__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_60__ap_ready),
    .idx(64'd3),
    .idy(64'd9),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_3_10__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_3_10__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_10__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_10__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_3_10__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_3_9__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_3_9__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_3_9__write),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_9_3__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_9_3__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_9_3__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_9_3__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_9_3__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_61
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_61__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_61__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_61__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_61__ap_ready),
    .idy(64'd10),
    .idx(64'd3),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_3_10__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_3_10__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_3_10__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_3_11__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_3_11__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_11__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_11__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_3_11__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_10_3__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_10_3__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_10_3__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_10_3__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_10_3__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_62
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_62__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_62__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_62__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_62__ap_ready),
    .idy(64'd11),
    .idx(64'd3),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_3_11__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_3_11__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_3_11__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_3_12__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_3_12__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_12__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_12__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_3_12__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_11_3__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_11_3__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_11_3__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_11_3__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_11_3__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_63
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_63__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_63__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_63__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_63__ap_ready),
    .idy(64'd12),
    .idx(64'd3),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_3_12__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_3_12__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_3_12__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_3_13__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_3_13__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_13__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_13__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_3_13__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_12_3__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_12_3__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_12_3__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_12_3__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_12_3__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_64
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_64__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_64__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_64__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_64__ap_ready),
    .idy(64'd13),
    .idx(64'd3),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_3_13__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_3_13__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_3_13__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_3_14__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_3_14__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_14__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_14__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_3_14__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_13_3__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_13_3__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_13_3__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_13_3__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_13_3__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_65
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_65__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_65__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_65__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_65__ap_ready),
    .idy(64'd14),
    .idx(64'd3),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_3_14__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_3_14__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_3_14__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_3_15__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_3_15__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_15__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_15__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_3_15__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_14_3__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_14_3__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_14_3__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_14_3__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_14_3__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_66
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_66__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_66__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_66__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_66__ap_ready),
    .idy(64'd15),
    .idx(64'd3),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_3_15__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_3_15__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_3_15__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_3_16__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_3_16__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_16__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_16__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_3_16__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_15_3__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_15_3__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_15_3__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_15_3__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_15_3__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_67
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_67__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_67__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_67__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_67__ap_ready),
    .idy(64'd16),
    .idx(64'd3),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_3_16__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_3_16__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_3_16__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_3_17__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_3_17__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_17__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_17__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_3_17__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_16_3__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_16_3__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_16_3__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_16_3__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_16_3__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_68
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_68__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_68__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_68__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_68__ap_ready),
    .idy(64'd0),
    .idx(64'd4),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_4_0__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_4_0__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_4_0__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_4_1__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_4_1__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_1__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_1__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_4_1__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_0_4__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_0_4__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_0_4__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_0_4__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_0_4__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_69
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_69__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_69__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_69__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_69__ap_ready),
    .idy(64'd1),
    .idx(64'd4),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_4_1__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_4_1__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_4_1__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_4_2__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_4_2__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_2__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_2__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_4_2__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_1_4__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_1_4__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_1_4__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_1_4__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_1_4__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_70
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_70__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_70__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_70__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_70__ap_ready),
    .idy(64'd2),
    .idx(64'd4),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_4_2__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_4_2__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_4_2__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_4_3__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_4_3__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_3__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_3__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_4_3__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_2_4__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_2_4__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_2_4__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_2_4__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_2_4__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_71
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_71__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_71__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_71__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_71__ap_ready),
    .idy(64'd3),
    .idx(64'd4),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_4_3__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_4_3__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_4_3__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_4_4__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_4_4__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_4__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_4__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_4_4__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_3_4__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_3_4__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_3_4__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_3_4__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_3_4__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_72
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_72__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_72__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_72__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_72__ap_ready),
    .idx(64'd4),
    .idy(64'd4),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_4_4__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_4_4__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_4_4__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_4_5__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_4_5__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_5__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_5__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_4_5__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_4_4__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_4_4__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_4_4__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_4_4__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_4_4__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_73
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_73__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_73__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_73__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_73__ap_ready),
    .idx(64'd4),
    .idy(64'd5),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_4_5__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_4_5__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_4_5__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_4_6__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_4_6__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_6__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_6__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_4_6__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_5_4__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_5_4__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_5_4__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_5_4__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_5_4__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_74
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_74__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_74__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_74__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_74__ap_ready),
    .idx(64'd4),
    .idy(64'd6),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_4_6__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_4_6__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_4_6__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_4_7__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_4_7__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_7__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_7__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_4_7__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_6_4__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_6_4__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_6_4__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_6_4__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_6_4__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_75
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_75__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_75__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_75__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_75__ap_ready),
    .idx(64'd4),
    .idy(64'd7),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_4_7__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_4_7__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_4_7__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_4_8__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_4_8__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_8__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_8__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_4_8__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_7_4__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_7_4__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_7_4__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_7_4__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_7_4__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_76
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_76__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_76__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_76__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_76__ap_ready),
    .idx(64'd4),
    .idy(64'd8),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_4_8__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_4_8__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_4_8__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_4_9__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_4_9__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_9__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_9__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_4_9__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_8_4__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_8_4__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_8_4__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_8_4__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_8_4__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_77
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_77__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_77__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_77__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_77__ap_ready),
    .idx(64'd4),
    .idy(64'd9),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_4_10__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_4_10__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_10__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_10__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_4_10__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_4_9__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_4_9__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_4_9__write),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_9_4__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_9_4__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_9_4__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_9_4__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_9_4__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_78
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_78__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_78__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_78__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_78__ap_ready),
    .idy(64'd10),
    .idx(64'd4),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_4_10__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_4_10__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_4_10__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_4_11__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_4_11__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_11__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_11__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_4_11__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_10_4__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_10_4__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_10_4__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_10_4__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_10_4__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_79
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_79__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_79__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_79__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_79__ap_ready),
    .idy(64'd11),
    .idx(64'd4),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_4_11__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_4_11__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_4_11__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_4_12__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_4_12__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_12__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_12__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_4_12__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_11_4__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_11_4__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_11_4__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_11_4__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_11_4__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_80
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_80__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_80__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_80__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_80__ap_ready),
    .idy(64'd12),
    .idx(64'd4),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_4_12__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_4_12__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_4_12__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_4_13__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_4_13__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_13__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_13__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_4_13__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_12_4__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_12_4__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_12_4__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_12_4__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_12_4__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_81
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_81__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_81__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_81__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_81__ap_ready),
    .idy(64'd13),
    .idx(64'd4),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_4_13__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_4_13__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_4_13__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_4_14__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_4_14__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_14__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_14__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_4_14__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_13_4__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_13_4__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_13_4__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_13_4__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_13_4__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_82
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_82__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_82__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_82__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_82__ap_ready),
    .idy(64'd14),
    .idx(64'd4),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_4_14__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_4_14__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_4_14__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_4_15__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_4_15__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_15__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_15__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_4_15__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_14_4__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_14_4__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_14_4__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_14_4__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_14_4__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_83
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_83__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_83__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_83__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_83__ap_ready),
    .idy(64'd15),
    .idx(64'd4),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_4_15__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_4_15__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_4_15__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_4_16__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_4_16__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_16__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_16__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_4_16__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_15_4__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_15_4__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_15_4__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_15_4__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_15_4__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_84
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_84__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_84__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_84__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_84__ap_ready),
    .idy(64'd16),
    .idx(64'd4),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_4_16__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_4_16__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_4_16__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_4_17__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_4_17__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_17__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_17__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_4_17__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_16_4__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_16_4__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_16_4__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_16_4__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_16_4__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_85
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_85__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_85__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_85__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_85__ap_ready),
    .idy(64'd0),
    .idx(64'd5),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_5_0__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_5_0__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_5_0__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_5_1__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_5_1__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_1__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_1__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_5_1__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_0_5__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_0_5__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_0_5__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_0_5__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_0_5__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_86
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_86__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_86__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_86__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_86__ap_ready),
    .idy(64'd1),
    .idx(64'd5),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_5_1__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_5_1__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_5_1__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_5_2__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_5_2__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_2__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_2__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_5_2__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_1_5__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_1_5__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_1_5__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_1_5__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_1_5__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_87
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_87__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_87__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_87__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_87__ap_ready),
    .idy(64'd2),
    .idx(64'd5),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_5_2__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_5_2__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_5_2__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_5_3__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_5_3__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_3__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_3__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_5_3__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_2_5__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_2_5__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_2_5__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_2_5__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_2_5__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_88
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_88__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_88__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_88__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_88__ap_ready),
    .idy(64'd3),
    .idx(64'd5),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_5_3__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_5_3__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_5_3__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_5_4__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_5_4__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_4__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_4__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_5_4__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_3_5__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_3_5__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_3_5__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_3_5__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_3_5__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_89
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_89__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_89__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_89__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_89__ap_ready),
    .idy(64'd4),
    .idx(64'd5),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_5_4__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_5_4__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_5_4__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_5_5__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_5_5__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_5__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_5__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_5_5__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_4_5__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_4_5__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_4_5__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_4_5__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_4_5__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_90
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_90__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_90__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_90__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_90__ap_ready),
    .idx(64'd5),
    .idy(64'd5),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_5_5__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_5_5__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_5_5__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_5_6__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_5_6__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_6__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_6__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_5_6__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_5_5__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_5_5__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_5_5__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_5_5__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_5_5__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_91
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_91__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_91__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_91__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_91__ap_ready),
    .idx(64'd5),
    .idy(64'd6),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_5_6__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_5_6__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_5_6__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_5_7__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_5_7__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_7__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_7__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_5_7__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_6_5__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_6_5__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_6_5__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_6_5__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_6_5__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_92
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_92__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_92__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_92__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_92__ap_ready),
    .idx(64'd5),
    .idy(64'd7),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_5_7__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_5_7__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_5_7__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_5_8__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_5_8__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_8__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_8__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_5_8__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_7_5__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_7_5__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_7_5__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_7_5__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_7_5__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_93
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_93__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_93__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_93__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_93__ap_ready),
    .idx(64'd5),
    .idy(64'd8),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_5_8__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_5_8__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_5_8__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_5_9__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_5_9__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_9__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_9__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_5_9__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_8_5__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_8_5__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_8_5__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_8_5__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_8_5__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_94
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_94__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_94__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_94__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_94__ap_ready),
    .idx(64'd5),
    .idy(64'd9),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_5_10__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_5_10__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_10__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_10__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_5_10__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_5_9__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_5_9__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_5_9__write),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_9_5__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_9_5__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_9_5__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_9_5__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_9_5__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_95
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_95__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_95__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_95__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_95__ap_ready),
    .idy(64'd10),
    .idx(64'd5),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_5_10__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_5_10__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_5_10__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_5_11__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_5_11__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_11__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_11__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_5_11__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_10_5__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_10_5__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_10_5__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_10_5__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_10_5__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_96
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_96__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_96__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_96__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_96__ap_ready),
    .idy(64'd11),
    .idx(64'd5),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_5_11__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_5_11__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_5_11__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_5_12__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_5_12__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_12__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_12__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_5_12__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_11_5__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_11_5__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_11_5__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_11_5__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_11_5__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_97
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_97__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_97__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_97__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_97__ap_ready),
    .idy(64'd12),
    .idx(64'd5),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_5_12__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_5_12__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_5_12__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_5_13__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_5_13__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_13__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_13__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_5_13__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_12_5__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_12_5__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_12_5__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_12_5__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_12_5__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_98
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_98__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_98__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_98__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_98__ap_ready),
    .idy(64'd13),
    .idx(64'd5),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_5_13__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_5_13__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_5_13__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_5_14__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_5_14__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_14__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_14__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_5_14__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_13_5__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_13_5__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_13_5__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_13_5__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_13_5__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_99
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_99__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_99__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_99__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_99__ap_ready),
    .idy(64'd14),
    .idx(64'd5),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_5_14__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_5_14__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_5_14__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_5_15__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_5_15__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_15__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_15__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_5_15__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_14_5__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_14_5__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_14_5__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_14_5__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_14_5__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_100
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_100__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_100__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_100__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_100__ap_ready),
    .idy(64'd15),
    .idx(64'd5),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_5_15__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_5_15__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_5_15__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_5_16__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_5_16__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_16__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_16__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_5_16__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_15_5__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_15_5__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_15_5__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_15_5__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_15_5__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_101
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_101__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_101__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_101__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_101__ap_ready),
    .idy(64'd16),
    .idx(64'd5),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_5_16__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_5_16__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_5_16__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_5_17__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_5_17__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_17__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_17__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_5_17__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_16_5__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_16_5__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_16_5__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_16_5__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_16_5__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_102
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_102__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_102__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_102__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_102__ap_ready),
    .idy(64'd0),
    .idx(64'd6),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_6_0__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_6_0__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_6_0__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_6_1__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_6_1__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_1__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_1__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_6_1__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_0_6__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_0_6__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_0_6__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_0_6__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_0_6__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_103
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_103__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_103__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_103__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_103__ap_ready),
    .idy(64'd1),
    .idx(64'd6),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_6_1__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_6_1__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_6_1__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_6_2__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_6_2__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_2__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_2__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_6_2__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_1_6__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_1_6__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_1_6__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_1_6__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_1_6__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_104
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_104__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_104__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_104__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_104__ap_ready),
    .idy(64'd2),
    .idx(64'd6),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_6_2__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_6_2__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_6_2__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_6_3__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_6_3__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_3__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_3__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_6_3__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_2_6__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_2_6__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_2_6__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_2_6__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_2_6__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_105
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_105__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_105__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_105__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_105__ap_ready),
    .idy(64'd3),
    .idx(64'd6),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_6_3__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_6_3__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_6_3__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_6_4__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_6_4__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_4__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_4__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_6_4__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_3_6__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_3_6__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_3_6__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_3_6__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_3_6__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_106
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_106__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_106__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_106__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_106__ap_ready),
    .idy(64'd4),
    .idx(64'd6),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_6_4__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_6_4__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_6_4__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_6_5__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_6_5__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_5__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_5__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_6_5__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_4_6__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_4_6__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_4_6__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_4_6__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_4_6__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_107
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_107__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_107__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_107__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_107__ap_ready),
    .idy(64'd5),
    .idx(64'd6),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_6_5__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_6_5__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_6_5__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_6_6__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_6_6__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_6__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_6__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_6_6__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_5_6__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_5_6__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_5_6__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_5_6__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_5_6__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_108
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_108__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_108__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_108__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_108__ap_ready),
    .idx(64'd6),
    .idy(64'd6),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_6_6__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_6_6__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_6_6__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_6_7__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_6_7__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_7__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_7__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_6_7__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_6_6__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_6_6__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_6_6__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_6_6__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_6_6__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_109
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_109__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_109__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_109__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_109__ap_ready),
    .idx(64'd6),
    .idy(64'd7),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_6_7__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_6_7__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_6_7__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_6_8__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_6_8__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_8__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_8__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_6_8__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_7_6__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_7_6__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_7_6__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_7_6__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_7_6__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_110
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_110__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_110__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_110__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_110__ap_ready),
    .idx(64'd6),
    .idy(64'd8),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_6_8__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_6_8__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_6_8__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_6_9__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_6_9__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_9__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_9__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_6_9__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_8_6__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_8_6__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_8_6__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_8_6__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_8_6__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_111
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_111__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_111__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_111__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_111__ap_ready),
    .idx(64'd6),
    .idy(64'd9),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_6_10__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_6_10__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_10__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_10__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_6_10__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_6_9__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_6_9__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_6_9__write),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_9_6__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_9_6__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_9_6__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_9_6__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_9_6__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_112
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_112__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_112__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_112__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_112__ap_ready),
    .idy(64'd10),
    .idx(64'd6),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_6_10__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_6_10__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_6_10__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_6_11__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_6_11__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_11__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_11__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_6_11__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_10_6__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_10_6__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_10_6__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_10_6__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_10_6__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_113
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_113__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_113__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_113__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_113__ap_ready),
    .idy(64'd11),
    .idx(64'd6),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_6_11__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_6_11__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_6_11__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_6_12__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_6_12__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_12__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_12__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_6_12__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_11_6__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_11_6__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_11_6__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_11_6__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_11_6__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_114
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_114__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_114__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_114__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_114__ap_ready),
    .idy(64'd12),
    .idx(64'd6),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_6_12__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_6_12__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_6_12__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_6_13__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_6_13__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_13__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_13__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_6_13__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_12_6__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_12_6__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_12_6__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_12_6__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_12_6__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_115
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_115__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_115__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_115__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_115__ap_ready),
    .idy(64'd13),
    .idx(64'd6),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_6_13__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_6_13__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_6_13__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_6_14__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_6_14__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_14__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_14__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_6_14__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_13_6__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_13_6__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_13_6__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_13_6__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_13_6__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_116
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_116__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_116__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_116__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_116__ap_ready),
    .idy(64'd14),
    .idx(64'd6),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_6_14__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_6_14__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_6_14__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_6_15__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_6_15__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_15__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_15__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_6_15__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_14_6__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_14_6__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_14_6__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_14_6__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_14_6__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_117
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_117__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_117__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_117__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_117__ap_ready),
    .idy(64'd15),
    .idx(64'd6),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_6_15__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_6_15__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_6_15__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_6_16__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_6_16__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_16__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_16__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_6_16__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_15_6__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_15_6__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_15_6__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_15_6__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_15_6__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_118
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_118__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_118__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_118__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_118__ap_ready),
    .idy(64'd16),
    .idx(64'd6),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_6_16__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_6_16__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_6_16__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_6_17__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_6_17__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_17__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_17__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_6_17__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_16_6__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_16_6__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_16_6__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_16_6__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_16_6__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_119
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_119__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_119__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_119__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_119__ap_ready),
    .idy(64'd0),
    .idx(64'd7),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_7_0__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_7_0__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_7_0__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_7_1__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_7_1__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_1__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_1__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_7_1__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_0_7__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_0_7__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_0_7__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_0_7__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_0_7__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_120
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_120__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_120__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_120__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_120__ap_ready),
    .idy(64'd1),
    .idx(64'd7),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_7_1__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_7_1__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_7_1__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_7_2__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_7_2__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_2__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_2__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_7_2__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_1_7__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_1_7__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_1_7__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_1_7__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_1_7__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_121
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_121__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_121__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_121__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_121__ap_ready),
    .idy(64'd2),
    .idx(64'd7),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_7_2__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_7_2__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_7_2__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_7_3__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_7_3__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_3__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_3__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_7_3__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_2_7__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_2_7__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_2_7__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_2_7__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_2_7__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_122
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_122__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_122__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_122__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_122__ap_ready),
    .idy(64'd3),
    .idx(64'd7),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_7_3__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_7_3__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_7_3__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_7_4__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_7_4__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_4__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_4__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_7_4__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_3_7__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_3_7__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_3_7__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_3_7__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_3_7__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_123
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_123__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_123__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_123__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_123__ap_ready),
    .idy(64'd4),
    .idx(64'd7),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_7_4__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_7_4__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_7_4__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_7_5__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_7_5__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_5__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_5__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_7_5__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_4_7__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_4_7__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_4_7__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_4_7__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_4_7__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_124
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_124__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_124__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_124__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_124__ap_ready),
    .idy(64'd5),
    .idx(64'd7),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_7_5__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_7_5__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_7_5__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_7_6__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_7_6__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_6__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_6__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_7_6__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_5_7__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_5_7__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_5_7__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_5_7__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_5_7__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_125
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_125__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_125__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_125__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_125__ap_ready),
    .idy(64'd6),
    .idx(64'd7),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_7_6__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_7_6__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_7_6__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_7_7__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_7_7__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_7__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_7__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_7_7__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_6_7__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_6_7__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_6_7__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_6_7__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_6_7__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_126
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_126__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_126__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_126__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_126__ap_ready),
    .idx(64'd7),
    .idy(64'd7),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_7_7__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_7_7__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_7_7__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_7_8__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_7_8__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_8__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_8__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_7_8__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_7_7__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_7_7__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_7_7__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_7_7__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_7_7__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_127
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_127__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_127__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_127__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_127__ap_ready),
    .idx(64'd7),
    .idy(64'd8),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_7_8__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_7_8__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_7_8__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_7_9__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_7_9__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_9__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_9__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_7_9__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_8_7__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_8_7__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_8_7__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_8_7__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_8_7__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_128
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_128__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_128__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_128__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_128__ap_ready),
    .idx(64'd7),
    .idy(64'd9),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_7_10__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_7_10__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_10__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_10__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_7_10__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_7_9__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_7_9__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_7_9__write),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_9_7__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_9_7__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_9_7__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_9_7__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_9_7__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_129
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_129__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_129__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_129__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_129__ap_ready),
    .idy(64'd10),
    .idx(64'd7),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_7_10__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_7_10__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_7_10__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_7_11__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_7_11__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_11__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_11__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_7_11__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_10_7__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_10_7__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_10_7__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_10_7__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_10_7__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_130
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_130__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_130__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_130__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_130__ap_ready),
    .idy(64'd11),
    .idx(64'd7),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_7_11__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_7_11__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_7_11__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_7_12__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_7_12__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_12__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_12__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_7_12__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_11_7__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_11_7__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_11_7__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_11_7__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_11_7__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_131
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_131__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_131__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_131__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_131__ap_ready),
    .idy(64'd12),
    .idx(64'd7),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_7_12__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_7_12__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_7_12__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_7_13__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_7_13__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_13__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_13__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_7_13__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_12_7__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_12_7__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_12_7__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_12_7__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_12_7__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_132
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_132__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_132__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_132__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_132__ap_ready),
    .idy(64'd13),
    .idx(64'd7),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_7_13__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_7_13__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_7_13__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_7_14__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_7_14__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_14__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_14__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_7_14__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_13_7__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_13_7__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_13_7__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_13_7__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_13_7__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_133
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_133__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_133__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_133__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_133__ap_ready),
    .idy(64'd14),
    .idx(64'd7),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_7_14__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_7_14__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_7_14__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_7_15__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_7_15__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_15__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_15__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_7_15__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_14_7__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_14_7__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_14_7__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_14_7__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_14_7__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_134
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_134__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_134__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_134__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_134__ap_ready),
    .idy(64'd15),
    .idx(64'd7),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_7_15__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_7_15__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_7_15__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_7_16__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_7_16__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_16__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_16__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_7_16__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_15_7__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_15_7__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_15_7__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_15_7__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_15_7__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_135
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_135__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_135__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_135__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_135__ap_ready),
    .idy(64'd16),
    .idx(64'd7),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_7_16__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_7_16__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_7_16__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_7_17__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_7_17__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_17__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_17__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_7_17__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_16_7__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_16_7__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_16_7__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_16_7__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_16_7__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_136
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_136__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_136__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_136__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_136__ap_ready),
    .idy(64'd0),
    .idx(64'd8),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_8_0__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_8_0__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_8_0__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_8_1__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_8_1__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_1__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_1__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_8_1__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_0_8__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_0_8__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_0_8__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_0_8__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_0_8__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_137
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_137__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_137__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_137__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_137__ap_ready),
    .idy(64'd1),
    .idx(64'd8),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_8_1__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_8_1__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_8_1__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_8_2__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_8_2__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_2__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_2__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_8_2__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_1_8__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_1_8__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_1_8__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_1_8__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_1_8__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_138
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_138__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_138__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_138__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_138__ap_ready),
    .idy(64'd2),
    .idx(64'd8),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_8_2__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_8_2__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_8_2__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_8_3__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_8_3__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_3__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_3__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_8_3__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_2_8__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_2_8__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_2_8__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_2_8__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_2_8__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_139
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_139__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_139__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_139__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_139__ap_ready),
    .idy(64'd3),
    .idx(64'd8),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_8_3__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_8_3__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_8_3__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_8_4__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_8_4__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_4__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_4__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_8_4__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_3_8__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_3_8__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_3_8__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_3_8__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_3_8__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_140
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_140__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_140__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_140__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_140__ap_ready),
    .idy(64'd4),
    .idx(64'd8),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_8_4__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_8_4__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_8_4__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_8_5__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_8_5__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_5__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_5__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_8_5__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_4_8__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_4_8__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_4_8__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_4_8__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_4_8__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_141
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_141__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_141__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_141__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_141__ap_ready),
    .idy(64'd5),
    .idx(64'd8),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_8_5__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_8_5__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_8_5__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_8_6__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_8_6__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_6__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_6__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_8_6__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_5_8__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_5_8__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_5_8__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_5_8__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_5_8__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_142
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_142__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_142__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_142__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_142__ap_ready),
    .idy(64'd6),
    .idx(64'd8),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_8_6__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_8_6__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_8_6__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_8_7__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_8_7__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_7__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_7__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_8_7__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_6_8__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_6_8__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_6_8__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_6_8__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_6_8__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_143
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_143__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_143__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_143__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_143__ap_ready),
    .idy(64'd7),
    .idx(64'd8),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_8_7__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_8_7__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_8_7__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_8_8__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_8_8__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_8__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_8__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_8_8__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_7_8__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_7_8__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_7_8__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_7_8__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_7_8__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_144
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_144__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_144__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_144__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_144__ap_ready),
    .idx(64'd8),
    .idy(64'd8),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_8_8__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_8_8__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_8_8__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_8_9__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_8_9__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_9__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_9__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_8_9__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_8_8__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_8_8__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_8_8__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_8_8__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_8_8__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_145
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_145__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_145__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_145__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_145__ap_ready),
    .idx(64'd8),
    .idy(64'd9),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_8_10__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_8_10__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_10__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_10__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_8_10__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_8_9__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_8_9__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_8_9__write),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_9_8__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_9_8__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_9_8__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_9_8__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_9_8__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_146
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_146__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_146__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_146__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_146__ap_ready),
    .idy(64'd10),
    .idx(64'd8),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_8_10__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_8_10__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_8_10__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_8_11__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_8_11__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_11__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_11__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_8_11__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_10_8__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_10_8__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_10_8__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_10_8__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_10_8__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_147
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_147__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_147__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_147__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_147__ap_ready),
    .idy(64'd11),
    .idx(64'd8),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_8_11__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_8_11__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_8_11__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_8_12__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_8_12__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_12__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_12__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_8_12__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_11_8__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_11_8__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_11_8__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_11_8__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_11_8__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_148
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_148__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_148__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_148__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_148__ap_ready),
    .idy(64'd12),
    .idx(64'd8),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_8_12__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_8_12__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_8_12__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_8_13__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_8_13__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_13__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_13__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_8_13__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_12_8__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_12_8__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_12_8__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_12_8__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_12_8__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_149
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_149__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_149__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_149__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_149__ap_ready),
    .idy(64'd13),
    .idx(64'd8),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_8_13__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_8_13__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_8_13__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_8_14__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_8_14__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_14__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_14__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_8_14__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_13_8__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_13_8__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_13_8__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_13_8__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_13_8__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_150
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_150__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_150__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_150__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_150__ap_ready),
    .idy(64'd14),
    .idx(64'd8),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_8_14__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_8_14__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_8_14__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_8_15__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_8_15__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_15__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_15__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_8_15__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_14_8__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_14_8__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_14_8__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_14_8__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_14_8__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_151
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_151__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_151__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_151__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_151__ap_ready),
    .idy(64'd15),
    .idx(64'd8),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_8_15__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_8_15__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_8_15__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_8_16__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_8_16__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_16__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_16__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_8_16__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_15_8__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_15_8__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_15_8__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_15_8__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_15_8__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_152
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_152__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_152__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_152__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_152__ap_ready),
    .idy(64'd16),
    .idx(64'd8),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_8_16__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_8_16__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_8_16__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_8_17__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_8_17__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_17__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_17__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_8_17__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_16_8__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_16_8__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_16_8__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_16_8__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_16_8__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_153
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_153__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_153__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_153__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_153__ap_ready),
    .idy(64'd0),
    .idx(64'd9),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_9_0__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_9_0__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_9_0__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_9_1__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_9_1__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_1__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_1__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_9_1__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_0_9__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_0_9__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_0_9__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_0_9__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_0_9__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_154
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_154__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_154__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_154__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_154__ap_ready),
    .idy(64'd1),
    .idx(64'd9),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_9_1__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_9_1__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_9_1__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_9_2__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_9_2__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_2__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_2__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_9_2__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_1_9__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_1_9__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_1_9__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_1_9__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_1_9__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_155
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_155__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_155__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_155__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_155__ap_ready),
    .idy(64'd2),
    .idx(64'd9),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_9_2__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_9_2__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_9_2__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_9_3__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_9_3__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_3__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_3__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_9_3__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_2_9__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_2_9__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_2_9__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_2_9__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_2_9__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_156
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_156__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_156__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_156__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_156__ap_ready),
    .idy(64'd3),
    .idx(64'd9),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_9_3__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_9_3__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_9_3__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_9_4__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_9_4__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_4__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_4__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_9_4__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_3_9__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_3_9__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_3_9__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_3_9__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_3_9__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_157
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_157__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_157__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_157__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_157__ap_ready),
    .idy(64'd4),
    .idx(64'd9),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_9_4__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_9_4__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_9_4__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_9_5__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_9_5__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_5__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_5__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_9_5__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_4_9__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_4_9__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_4_9__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_4_9__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_4_9__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_158
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_158__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_158__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_158__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_158__ap_ready),
    .idy(64'd5),
    .idx(64'd9),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_9_5__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_9_5__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_9_5__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_9_6__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_9_6__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_6__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_6__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_9_6__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_5_9__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_5_9__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_5_9__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_5_9__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_5_9__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_159
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_159__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_159__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_159__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_159__ap_ready),
    .idy(64'd6),
    .idx(64'd9),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_9_6__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_9_6__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_9_6__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_9_7__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_9_7__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_7__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_7__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_9_7__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_6_9__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_6_9__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_6_9__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_6_9__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_6_9__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_160
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_160__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_160__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_160__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_160__ap_ready),
    .idy(64'd7),
    .idx(64'd9),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_9_7__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_9_7__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_9_7__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_9_8__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_9_8__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_8__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_8__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_9_8__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_7_9__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_7_9__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_7_9__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_7_9__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_7_9__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_161
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_161__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_161__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_161__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_161__ap_ready),
    .idy(64'd8),
    .idx(64'd9),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_9_8__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_9_8__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_9_8__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_9_9__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_9_9__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_9__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_9__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_9_9__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_8_9__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_8_9__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_8_9__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_8_9__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_8_9__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_162
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_162__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_162__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_162__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_162__ap_ready),
    .idx(64'd9),
    .idy(64'd9),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_9_10__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_9_10__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_10__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_10__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_9_10__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_9_9__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_9_9__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_9_9__write),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_9_9__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_9_9__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_9_9__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_9_9__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_9_9__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_163
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_163__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_163__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_163__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_163__ap_ready),
    .idy(64'd10),
    .idx(64'd9),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_9_10__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_9_10__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_9_10__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_9_11__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_9_11__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_11__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_11__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_9_11__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_10_9__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_10_9__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_10_9__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_10_9__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_10_9__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_164
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_164__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_164__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_164__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_164__ap_ready),
    .idy(64'd11),
    .idx(64'd9),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_9_11__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_9_11__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_9_11__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_9_12__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_9_12__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_12__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_12__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_9_12__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_11_9__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_11_9__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_11_9__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_11_9__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_11_9__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_165
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_165__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_165__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_165__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_165__ap_ready),
    .idy(64'd12),
    .idx(64'd9),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_9_12__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_9_12__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_9_12__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_9_13__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_9_13__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_13__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_13__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_9_13__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_12_9__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_12_9__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_12_9__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_12_9__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_12_9__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_166
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_166__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_166__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_166__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_166__ap_ready),
    .idy(64'd13),
    .idx(64'd9),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_9_13__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_9_13__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_9_13__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_9_14__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_9_14__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_14__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_14__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_9_14__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_13_9__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_13_9__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_13_9__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_13_9__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_13_9__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_167
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_167__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_167__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_167__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_167__ap_ready),
    .idy(64'd14),
    .idx(64'd9),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_9_14__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_9_14__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_9_14__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_9_15__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_9_15__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_15__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_15__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_9_15__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_14_9__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_14_9__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_14_9__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_14_9__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_14_9__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_168
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_168__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_168__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_168__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_168__ap_ready),
    .idy(64'd15),
    .idx(64'd9),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_9_15__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_9_15__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_9_15__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_9_16__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_9_16__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_16__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_16__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_9_16__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_15_9__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_15_9__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_15_9__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_15_9__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_15_9__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_169
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_169__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_169__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_169__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_169__ap_ready),
    .idy(64'd16),
    .idx(64'd9),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_9_16__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_9_16__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_9_16__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_9_17__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_9_17__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_17__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_17__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_9_17__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_16_9__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_16_9__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_16_9__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_16_9__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_16_9__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_170
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_170__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_170__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_170__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_170__ap_ready),
    .idy(64'd0),
    .idx(64'd10),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_10_0__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_10_0__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_10_0__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_10_1__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_10_1__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_1__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_1__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_10_1__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_0_10__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_0_10__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_0_10__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_0_10__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_0_10__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_171
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_171__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_171__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_171__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_171__ap_ready),
    .idy(64'd1),
    .idx(64'd10),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_10_1__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_10_1__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_10_1__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_10_2__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_10_2__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_2__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_2__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_10_2__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_1_10__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_1_10__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_1_10__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_1_10__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_1_10__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_172
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_172__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_172__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_172__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_172__ap_ready),
    .idx(64'd10),
    .idy(64'd2),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_10_2__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_10_2__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_10_2__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_10_3__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_10_3__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_3__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_3__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_10_3__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_2_10__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_2_10__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_2_10__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_2_10__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_2_10__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_173
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_173__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_173__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_173__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_173__ap_ready),
    .idx(64'd10),
    .idy(64'd3),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_10_3__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_10_3__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_10_3__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_10_4__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_10_4__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_4__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_4__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_10_4__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_3_10__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_3_10__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_3_10__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_3_10__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_3_10__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_174
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_174__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_174__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_174__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_174__ap_ready),
    .idx(64'd10),
    .idy(64'd4),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_10_4__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_10_4__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_10_4__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_10_5__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_10_5__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_5__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_5__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_10_5__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_4_10__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_4_10__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_4_10__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_4_10__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_4_10__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_175
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_175__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_175__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_175__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_175__ap_ready),
    .idx(64'd10),
    .idy(64'd5),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_10_5__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_10_5__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_10_5__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_10_6__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_10_6__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_6__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_6__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_10_6__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_5_10__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_5_10__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_5_10__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_5_10__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_5_10__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_176
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_176__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_176__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_176__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_176__ap_ready),
    .idx(64'd10),
    .idy(64'd6),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_10_6__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_10_6__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_10_6__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_10_7__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_10_7__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_7__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_7__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_10_7__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_6_10__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_6_10__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_6_10__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_6_10__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_6_10__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_177
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_177__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_177__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_177__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_177__ap_ready),
    .idx(64'd10),
    .idy(64'd7),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_10_7__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_10_7__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_10_7__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_10_8__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_10_8__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_8__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_8__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_10_8__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_7_10__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_7_10__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_7_10__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_7_10__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_7_10__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_178
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_178__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_178__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_178__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_178__ap_ready),
    .idx(64'd10),
    .idy(64'd8),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_10_8__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_10_8__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_10_8__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_10_9__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_10_9__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_9__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_9__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_10_9__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_8_10__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_8_10__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_8_10__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_8_10__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_8_10__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_179
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_179__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_179__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_179__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_179__ap_ready),
    .idx(64'd10),
    .idy(64'd9),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_10_10__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_10_10__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_10__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_10__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_10_10__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_10_9__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_10_9__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_10_9__write),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_9_10__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_9_10__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_9_10__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_9_10__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_9_10__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_180
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_180__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_180__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_180__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_180__ap_ready),
    .idx(64'd10),
    .idy(64'd10),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_10_10__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_10_10__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_10_10__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_10_11__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_10_11__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_11__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_11__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_10_11__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_10_10__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_10_10__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_10_10__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_10_10__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_10_10__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_181
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_181__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_181__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_181__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_181__ap_ready),
    .idx(64'd10),
    .idy(64'd11),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_10_11__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_10_11__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_10_11__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_10_12__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_10_12__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_12__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_12__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_10_12__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_11_10__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_11_10__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_11_10__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_11_10__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_11_10__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_182
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_182__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_182__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_182__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_182__ap_ready),
    .idx(64'd10),
    .idy(64'd12),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_10_12__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_10_12__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_10_12__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_10_13__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_10_13__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_13__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_13__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_10_13__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_12_10__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_12_10__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_12_10__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_12_10__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_12_10__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_183
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_183__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_183__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_183__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_183__ap_ready),
    .idx(64'd10),
    .idy(64'd13),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_10_13__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_10_13__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_10_13__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_10_14__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_10_14__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_14__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_14__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_10_14__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_13_10__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_13_10__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_13_10__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_13_10__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_13_10__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_184
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_184__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_184__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_184__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_184__ap_ready),
    .idx(64'd10),
    .idy(64'd14),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_10_14__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_10_14__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_10_14__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_10_15__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_10_15__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_15__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_15__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_10_15__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_14_10__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_14_10__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_14_10__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_14_10__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_14_10__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_185
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_185__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_185__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_185__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_185__ap_ready),
    .idx(64'd10),
    .idy(64'd15),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_10_15__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_10_15__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_10_15__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_10_16__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_10_16__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_16__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_16__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_10_16__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_15_10__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_15_10__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_15_10__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_15_10__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_15_10__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_186
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_186__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_186__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_186__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_186__ap_ready),
    .idx(64'd10),
    .idy(64'd16),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_10_16__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_10_16__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_10_16__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_10_17__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_10_17__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_17__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_17__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_10_17__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_16_10__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_16_10__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_16_10__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_16_10__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_16_10__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_187
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_187__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_187__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_187__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_187__ap_ready),
    .idy(64'd0),
    .idx(64'd11),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_11_0__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_11_0__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_11_0__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_11_1__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_11_1__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_1__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_1__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_11_1__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_0_11__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_0_11__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_0_11__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_0_11__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_0_11__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_188
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_188__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_188__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_188__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_188__ap_ready),
    .idy(64'd1),
    .idx(64'd11),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_11_1__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_11_1__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_11_1__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_11_2__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_11_2__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_2__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_2__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_11_2__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_1_11__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_1_11__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_1_11__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_1_11__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_1_11__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_189
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_189__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_189__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_189__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_189__ap_ready),
    .idx(64'd11),
    .idy(64'd2),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_11_2__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_11_2__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_11_2__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_11_3__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_11_3__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_3__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_3__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_11_3__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_2_11__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_2_11__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_2_11__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_2_11__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_2_11__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_190
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_190__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_190__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_190__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_190__ap_ready),
    .idx(64'd11),
    .idy(64'd3),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_11_3__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_11_3__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_11_3__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_11_4__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_11_4__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_4__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_4__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_11_4__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_3_11__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_3_11__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_3_11__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_3_11__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_3_11__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_191
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_191__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_191__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_191__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_191__ap_ready),
    .idx(64'd11),
    .idy(64'd4),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_11_4__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_11_4__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_11_4__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_11_5__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_11_5__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_5__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_5__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_11_5__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_4_11__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_4_11__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_4_11__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_4_11__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_4_11__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_192
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_192__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_192__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_192__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_192__ap_ready),
    .idx(64'd11),
    .idy(64'd5),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_11_5__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_11_5__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_11_5__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_11_6__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_11_6__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_6__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_6__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_11_6__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_5_11__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_5_11__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_5_11__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_5_11__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_5_11__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_193
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_193__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_193__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_193__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_193__ap_ready),
    .idx(64'd11),
    .idy(64'd6),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_11_6__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_11_6__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_11_6__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_11_7__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_11_7__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_7__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_7__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_11_7__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_6_11__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_6_11__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_6_11__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_6_11__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_6_11__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_194
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_194__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_194__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_194__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_194__ap_ready),
    .idx(64'd11),
    .idy(64'd7),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_11_7__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_11_7__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_11_7__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_11_8__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_11_8__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_8__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_8__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_11_8__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_7_11__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_7_11__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_7_11__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_7_11__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_7_11__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_195
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_195__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_195__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_195__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_195__ap_ready),
    .idx(64'd11),
    .idy(64'd8),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_11_8__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_11_8__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_11_8__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_11_9__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_11_9__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_9__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_9__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_11_9__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_8_11__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_8_11__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_8_11__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_8_11__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_8_11__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_196
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_196__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_196__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_196__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_196__ap_ready),
    .idx(64'd11),
    .idy(64'd9),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_11_10__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_11_10__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_10__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_10__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_11_10__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_11_9__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_11_9__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_11_9__write),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_9_11__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_9_11__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_9_11__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_9_11__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_9_11__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_197
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_197__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_197__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_197__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_197__ap_ready),
    .idy(64'd10),
    .idx(64'd11),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_11_10__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_11_10__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_11_10__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_11_11__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_11_11__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_11__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_11__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_11_11__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_10_11__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_10_11__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_10_11__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_10_11__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_10_11__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_198
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_198__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_198__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_198__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_198__ap_ready),
    .idx(64'd11),
    .idy(64'd11),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_11_11__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_11_11__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_11_11__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_11_12__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_11_12__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_12__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_12__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_11_12__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_11_11__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_11_11__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_11_11__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_11_11__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_11_11__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_199
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_199__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_199__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_199__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_199__ap_ready),
    .idx(64'd11),
    .idy(64'd12),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_11_12__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_11_12__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_11_12__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_11_13__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_11_13__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_13__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_13__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_11_13__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_12_11__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_12_11__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_12_11__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_12_11__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_12_11__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_200
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_200__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_200__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_200__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_200__ap_ready),
    .idx(64'd11),
    .idy(64'd13),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_11_13__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_11_13__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_11_13__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_11_14__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_11_14__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_14__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_14__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_11_14__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_13_11__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_13_11__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_13_11__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_13_11__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_13_11__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_201
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_201__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_201__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_201__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_201__ap_ready),
    .idx(64'd11),
    .idy(64'd14),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_11_14__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_11_14__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_11_14__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_11_15__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_11_15__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_15__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_15__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_11_15__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_14_11__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_14_11__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_14_11__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_14_11__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_14_11__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_202
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_202__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_202__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_202__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_202__ap_ready),
    .idx(64'd11),
    .idy(64'd15),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_11_15__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_11_15__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_11_15__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_11_16__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_11_16__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_16__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_16__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_11_16__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_15_11__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_15_11__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_15_11__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_15_11__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_15_11__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_203
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_203__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_203__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_203__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_203__ap_ready),
    .idx(64'd11),
    .idy(64'd16),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_11_16__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_11_16__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_11_16__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_11_17__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_11_17__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_17__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_17__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_11_17__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_16_11__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_16_11__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_16_11__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_16_11__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_16_11__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_204
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_204__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_204__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_204__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_204__ap_ready),
    .idy(64'd0),
    .idx(64'd12),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_12_0__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_12_0__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_12_0__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_12_1__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_12_1__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_1__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_1__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_12_1__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_0_12__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_0_12__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_0_12__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_0_12__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_0_12__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_205
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_205__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_205__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_205__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_205__ap_ready),
    .idy(64'd1),
    .idx(64'd12),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_12_1__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_12_1__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_12_1__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_12_2__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_12_2__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_2__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_2__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_12_2__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_1_12__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_1_12__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_1_12__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_1_12__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_1_12__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_206
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_206__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_206__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_206__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_206__ap_ready),
    .idx(64'd12),
    .idy(64'd2),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_12_2__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_12_2__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_12_2__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_12_3__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_12_3__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_3__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_3__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_12_3__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_2_12__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_2_12__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_2_12__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_2_12__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_2_12__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_207
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_207__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_207__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_207__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_207__ap_ready),
    .idx(64'd12),
    .idy(64'd3),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_12_3__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_12_3__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_12_3__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_12_4__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_12_4__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_4__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_4__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_12_4__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_3_12__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_3_12__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_3_12__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_3_12__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_3_12__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_208
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_208__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_208__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_208__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_208__ap_ready),
    .idx(64'd12),
    .idy(64'd4),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_12_4__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_12_4__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_12_4__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_12_5__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_12_5__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_5__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_5__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_12_5__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_4_12__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_4_12__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_4_12__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_4_12__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_4_12__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_209
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_209__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_209__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_209__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_209__ap_ready),
    .idx(64'd12),
    .idy(64'd5),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_12_5__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_12_5__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_12_5__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_12_6__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_12_6__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_6__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_6__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_12_6__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_5_12__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_5_12__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_5_12__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_5_12__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_5_12__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_210
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_210__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_210__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_210__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_210__ap_ready),
    .idx(64'd12),
    .idy(64'd6),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_12_6__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_12_6__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_12_6__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_12_7__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_12_7__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_7__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_7__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_12_7__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_6_12__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_6_12__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_6_12__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_6_12__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_6_12__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_211
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_211__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_211__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_211__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_211__ap_ready),
    .idx(64'd12),
    .idy(64'd7),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_12_7__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_12_7__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_12_7__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_12_8__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_12_8__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_8__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_8__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_12_8__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_7_12__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_7_12__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_7_12__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_7_12__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_7_12__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_212
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_212__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_212__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_212__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_212__ap_ready),
    .idx(64'd12),
    .idy(64'd8),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_12_8__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_12_8__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_12_8__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_12_9__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_12_9__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_9__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_9__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_12_9__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_8_12__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_8_12__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_8_12__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_8_12__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_8_12__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_213
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_213__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_213__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_213__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_213__ap_ready),
    .idx(64'd12),
    .idy(64'd9),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_12_10__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_12_10__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_10__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_10__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_12_10__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_12_9__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_12_9__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_12_9__write),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_9_12__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_9_12__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_9_12__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_9_12__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_9_12__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_214
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_214__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_214__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_214__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_214__ap_ready),
    .idy(64'd10),
    .idx(64'd12),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_12_10__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_12_10__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_12_10__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_12_11__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_12_11__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_11__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_11__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_12_11__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_10_12__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_10_12__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_10_12__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_10_12__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_10_12__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_215
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_215__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_215__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_215__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_215__ap_ready),
    .idy(64'd11),
    .idx(64'd12),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_12_11__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_12_11__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_12_11__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_12_12__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_12_12__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_12__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_12__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_12_12__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_11_12__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_11_12__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_11_12__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_11_12__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_11_12__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_216
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_216__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_216__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_216__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_216__ap_ready),
    .idx(64'd12),
    .idy(64'd12),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_12_12__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_12_12__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_12_12__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_12_13__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_12_13__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_13__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_13__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_12_13__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_12_12__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_12_12__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_12_12__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_12_12__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_12_12__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_217
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_217__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_217__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_217__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_217__ap_ready),
    .idx(64'd12),
    .idy(64'd13),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_12_13__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_12_13__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_12_13__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_12_14__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_12_14__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_14__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_14__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_12_14__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_13_12__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_13_12__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_13_12__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_13_12__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_13_12__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_218
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_218__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_218__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_218__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_218__ap_ready),
    .idx(64'd12),
    .idy(64'd14),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_12_14__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_12_14__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_12_14__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_12_15__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_12_15__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_15__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_15__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_12_15__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_14_12__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_14_12__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_14_12__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_14_12__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_14_12__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_219
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_219__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_219__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_219__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_219__ap_ready),
    .idx(64'd12),
    .idy(64'd15),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_12_15__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_12_15__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_12_15__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_12_16__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_12_16__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_16__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_16__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_12_16__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_15_12__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_15_12__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_15_12__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_15_12__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_15_12__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_220
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_220__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_220__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_220__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_220__ap_ready),
    .idx(64'd12),
    .idy(64'd16),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_12_16__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_12_16__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_12_16__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_12_17__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_12_17__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_17__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_17__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_12_17__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_16_12__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_16_12__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_16_12__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_16_12__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_16_12__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_221
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_221__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_221__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_221__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_221__ap_ready),
    .idy(64'd0),
    .idx(64'd13),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_13_0__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_13_0__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_13_0__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_13_1__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_13_1__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_1__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_1__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_13_1__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_0_13__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_0_13__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_0_13__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_0_13__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_0_13__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_222
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_222__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_222__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_222__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_222__ap_ready),
    .idy(64'd1),
    .idx(64'd13),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_13_1__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_13_1__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_13_1__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_13_2__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_13_2__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_2__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_2__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_13_2__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_1_13__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_1_13__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_1_13__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_1_13__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_1_13__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_223
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_223__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_223__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_223__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_223__ap_ready),
    .idx(64'd13),
    .idy(64'd2),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_13_2__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_13_2__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_13_2__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_13_3__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_13_3__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_3__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_3__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_13_3__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_2_13__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_2_13__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_2_13__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_2_13__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_2_13__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_224
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_224__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_224__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_224__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_224__ap_ready),
    .idx(64'd13),
    .idy(64'd3),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_13_3__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_13_3__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_13_3__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_13_4__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_13_4__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_4__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_4__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_13_4__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_3_13__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_3_13__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_3_13__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_3_13__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_3_13__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_225
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_225__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_225__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_225__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_225__ap_ready),
    .idx(64'd13),
    .idy(64'd4),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_13_4__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_13_4__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_13_4__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_13_5__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_13_5__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_5__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_5__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_13_5__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_4_13__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_4_13__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_4_13__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_4_13__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_4_13__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_226
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_226__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_226__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_226__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_226__ap_ready),
    .idx(64'd13),
    .idy(64'd5),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_13_5__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_13_5__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_13_5__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_13_6__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_13_6__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_6__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_6__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_13_6__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_5_13__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_5_13__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_5_13__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_5_13__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_5_13__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_227
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_227__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_227__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_227__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_227__ap_ready),
    .idx(64'd13),
    .idy(64'd6),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_13_6__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_13_6__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_13_6__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_13_7__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_13_7__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_7__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_7__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_13_7__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_6_13__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_6_13__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_6_13__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_6_13__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_6_13__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_228
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_228__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_228__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_228__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_228__ap_ready),
    .idx(64'd13),
    .idy(64'd7),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_13_7__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_13_7__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_13_7__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_13_8__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_13_8__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_8__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_8__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_13_8__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_7_13__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_7_13__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_7_13__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_7_13__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_7_13__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_229
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_229__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_229__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_229__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_229__ap_ready),
    .idx(64'd13),
    .idy(64'd8),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_13_8__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_13_8__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_13_8__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_13_9__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_13_9__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_9__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_9__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_13_9__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_8_13__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_8_13__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_8_13__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_8_13__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_8_13__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_230
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_230__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_230__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_230__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_230__ap_ready),
    .idx(64'd13),
    .idy(64'd9),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_13_10__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_13_10__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_10__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_10__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_13_10__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_13_9__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_13_9__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_13_9__write),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_9_13__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_9_13__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_9_13__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_9_13__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_9_13__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_231
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_231__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_231__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_231__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_231__ap_ready),
    .idy(64'd10),
    .idx(64'd13),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_13_10__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_13_10__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_13_10__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_13_11__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_13_11__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_11__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_11__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_13_11__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_10_13__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_10_13__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_10_13__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_10_13__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_10_13__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_232
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_232__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_232__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_232__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_232__ap_ready),
    .idy(64'd11),
    .idx(64'd13),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_13_11__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_13_11__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_13_11__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_13_12__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_13_12__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_12__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_12__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_13_12__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_11_13__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_11_13__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_11_13__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_11_13__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_11_13__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_233
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_233__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_233__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_233__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_233__ap_ready),
    .idy(64'd12),
    .idx(64'd13),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_13_12__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_13_12__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_13_12__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_13_13__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_13_13__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_13__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_13__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_13_13__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_12_13__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_12_13__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_12_13__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_12_13__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_12_13__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_234
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_234__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_234__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_234__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_234__ap_ready),
    .idx(64'd13),
    .idy(64'd13),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_13_13__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_13_13__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_13_13__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_13_14__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_13_14__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_14__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_14__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_13_14__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_13_13__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_13_13__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_13_13__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_13_13__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_13_13__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_235
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_235__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_235__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_235__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_235__ap_ready),
    .idx(64'd13),
    .idy(64'd14),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_13_14__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_13_14__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_13_14__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_13_15__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_13_15__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_15__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_15__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_13_15__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_14_13__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_14_13__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_14_13__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_14_13__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_14_13__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_236
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_236__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_236__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_236__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_236__ap_ready),
    .idx(64'd13),
    .idy(64'd15),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_13_15__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_13_15__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_13_15__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_13_16__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_13_16__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_16__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_16__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_13_16__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_15_13__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_15_13__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_15_13__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_15_13__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_15_13__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_237
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_237__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_237__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_237__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_237__ap_ready),
    .idx(64'd13),
    .idy(64'd16),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_13_16__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_13_16__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_13_16__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_13_17__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_13_17__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_17__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_17__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_13_17__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_16_13__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_16_13__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_16_13__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_16_13__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_16_13__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_238
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_238__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_238__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_238__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_238__ap_ready),
    .idy(64'd0),
    .idx(64'd14),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_14_0__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_14_0__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_14_0__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_14_1__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_14_1__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_1__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_1__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_14_1__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_0_14__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_0_14__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_0_14__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_0_14__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_0_14__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_239
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_239__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_239__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_239__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_239__ap_ready),
    .idy(64'd1),
    .idx(64'd14),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_14_1__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_14_1__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_14_1__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_14_2__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_14_2__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_2__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_2__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_14_2__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_1_14__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_1_14__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_1_14__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_1_14__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_1_14__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_240
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_240__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_240__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_240__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_240__ap_ready),
    .idx(64'd14),
    .idy(64'd2),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_14_2__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_14_2__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_14_2__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_14_3__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_14_3__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_3__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_3__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_14_3__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_2_14__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_2_14__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_2_14__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_2_14__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_2_14__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_241
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_241__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_241__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_241__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_241__ap_ready),
    .idx(64'd14),
    .idy(64'd3),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_14_3__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_14_3__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_14_3__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_14_4__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_14_4__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_4__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_4__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_14_4__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_3_14__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_3_14__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_3_14__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_3_14__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_3_14__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_242
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_242__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_242__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_242__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_242__ap_ready),
    .idx(64'd14),
    .idy(64'd4),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_14_4__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_14_4__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_14_4__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_14_5__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_14_5__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_5__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_5__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_14_5__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_4_14__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_4_14__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_4_14__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_4_14__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_4_14__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_243
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_243__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_243__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_243__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_243__ap_ready),
    .idx(64'd14),
    .idy(64'd5),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_14_5__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_14_5__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_14_5__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_14_6__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_14_6__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_6__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_6__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_14_6__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_5_14__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_5_14__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_5_14__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_5_14__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_5_14__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_244
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_244__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_244__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_244__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_244__ap_ready),
    .idx(64'd14),
    .idy(64'd6),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_14_6__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_14_6__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_14_6__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_14_7__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_14_7__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_7__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_7__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_14_7__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_6_14__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_6_14__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_6_14__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_6_14__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_6_14__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_245
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_245__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_245__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_245__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_245__ap_ready),
    .idx(64'd14),
    .idy(64'd7),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_14_7__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_14_7__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_14_7__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_14_8__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_14_8__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_8__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_8__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_14_8__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_7_14__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_7_14__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_7_14__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_7_14__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_7_14__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_246
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_246__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_246__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_246__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_246__ap_ready),
    .idx(64'd14),
    .idy(64'd8),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_14_8__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_14_8__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_14_8__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_14_9__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_14_9__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_9__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_9__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_14_9__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_8_14__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_8_14__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_8_14__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_8_14__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_8_14__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_247
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_247__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_247__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_247__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_247__ap_ready),
    .idx(64'd14),
    .idy(64'd9),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_14_10__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_14_10__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_10__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_10__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_14_10__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_14_9__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_14_9__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_14_9__write),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_9_14__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_9_14__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_9_14__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_9_14__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_9_14__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_248
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_248__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_248__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_248__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_248__ap_ready),
    .idy(64'd10),
    .idx(64'd14),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_14_10__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_14_10__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_14_10__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_14_11__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_14_11__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_11__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_11__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_14_11__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_10_14__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_10_14__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_10_14__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_10_14__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_10_14__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_249
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_249__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_249__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_249__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_249__ap_ready),
    .idy(64'd11),
    .idx(64'd14),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_14_11__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_14_11__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_14_11__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_14_12__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_14_12__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_12__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_12__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_14_12__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_11_14__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_11_14__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_11_14__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_11_14__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_11_14__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_250
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_250__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_250__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_250__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_250__ap_ready),
    .idy(64'd12),
    .idx(64'd14),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_14_12__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_14_12__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_14_12__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_14_13__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_14_13__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_13__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_13__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_14_13__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_12_14__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_12_14__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_12_14__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_12_14__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_12_14__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_251
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_251__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_251__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_251__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_251__ap_ready),
    .idy(64'd13),
    .idx(64'd14),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_14_13__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_14_13__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_14_13__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_14_14__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_14_14__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_14__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_14__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_14_14__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_13_14__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_13_14__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_13_14__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_13_14__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_13_14__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_252
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_252__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_252__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_252__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_252__ap_ready),
    .idx(64'd14),
    .idy(64'd14),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_14_14__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_14_14__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_14_14__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_14_15__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_14_15__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_15__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_15__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_14_15__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_14_14__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_14_14__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_14_14__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_14_14__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_14_14__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_253
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_253__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_253__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_253__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_253__ap_ready),
    .idx(64'd14),
    .idy(64'd15),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_14_15__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_14_15__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_14_15__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_14_16__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_14_16__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_16__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_16__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_14_16__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_15_14__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_15_14__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_15_14__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_15_14__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_15_14__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_254
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_254__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_254__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_254__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_254__ap_ready),
    .idx(64'd14),
    .idy(64'd16),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_14_16__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_14_16__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_14_16__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_14_17__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_14_17__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_17__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_17__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_14_17__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_16_14__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_16_14__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_16_14__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_16_14__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_16_14__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_255
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_255__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_255__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_255__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_255__ap_ready),
    .idy(64'd0),
    .idx(64'd15),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_15_0__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_15_0__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_15_0__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_15_1__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_15_1__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_1__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_1__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_15_1__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_0_15__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_0_15__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_0_15__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_0_15__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_0_15__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_256
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_256__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_256__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_256__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_256__ap_ready),
    .idy(64'd1),
    .idx(64'd15),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_15_1__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_15_1__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_15_1__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_15_2__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_15_2__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_2__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_2__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_15_2__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_1_15__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_1_15__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_1_15__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_1_15__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_1_15__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_257
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_257__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_257__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_257__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_257__ap_ready),
    .idx(64'd15),
    .idy(64'd2),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_15_2__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_15_2__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_15_2__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_15_3__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_15_3__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_3__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_3__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_15_3__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_2_15__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_2_15__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_2_15__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_2_15__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_2_15__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_258
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_258__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_258__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_258__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_258__ap_ready),
    .idx(64'd15),
    .idy(64'd3),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_15_3__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_15_3__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_15_3__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_15_4__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_15_4__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_4__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_4__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_15_4__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_3_15__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_3_15__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_3_15__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_3_15__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_3_15__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_259
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_259__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_259__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_259__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_259__ap_ready),
    .idx(64'd15),
    .idy(64'd4),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_15_4__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_15_4__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_15_4__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_15_5__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_15_5__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_5__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_5__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_15_5__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_4_15__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_4_15__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_4_15__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_4_15__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_4_15__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_260
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_260__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_260__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_260__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_260__ap_ready),
    .idx(64'd15),
    .idy(64'd5),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_15_5__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_15_5__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_15_5__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_15_6__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_15_6__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_6__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_6__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_15_6__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_5_15__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_5_15__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_5_15__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_5_15__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_5_15__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_261
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_261__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_261__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_261__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_261__ap_ready),
    .idx(64'd15),
    .idy(64'd6),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_15_6__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_15_6__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_15_6__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_15_7__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_15_7__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_7__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_7__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_15_7__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_6_15__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_6_15__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_6_15__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_6_15__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_6_15__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_262
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_262__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_262__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_262__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_262__ap_ready),
    .idx(64'd15),
    .idy(64'd7),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_15_7__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_15_7__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_15_7__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_15_8__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_15_8__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_8__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_8__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_15_8__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_7_15__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_7_15__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_7_15__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_7_15__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_7_15__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_263
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_263__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_263__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_263__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_263__ap_ready),
    .idx(64'd15),
    .idy(64'd8),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_15_8__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_15_8__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_15_8__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_15_9__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_15_9__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_9__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_9__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_15_9__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_8_15__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_8_15__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_8_15__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_8_15__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_8_15__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_264
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_264__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_264__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_264__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_264__ap_ready),
    .idx(64'd15),
    .idy(64'd9),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_15_10__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_15_10__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_10__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_10__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_15_10__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_15_9__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_15_9__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_15_9__write),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_9_15__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_9_15__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_9_15__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_9_15__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_9_15__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_265
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_265__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_265__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_265__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_265__ap_ready),
    .idy(64'd10),
    .idx(64'd15),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_15_10__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_15_10__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_15_10__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_15_11__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_15_11__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_11__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_11__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_15_11__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_10_15__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_10_15__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_10_15__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_10_15__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_10_15__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_266
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_266__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_266__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_266__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_266__ap_ready),
    .idy(64'd11),
    .idx(64'd15),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_15_11__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_15_11__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_15_11__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_15_12__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_15_12__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_12__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_12__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_15_12__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_11_15__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_11_15__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_11_15__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_11_15__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_11_15__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_267
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_267__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_267__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_267__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_267__ap_ready),
    .idy(64'd12),
    .idx(64'd15),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_15_12__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_15_12__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_15_12__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_15_13__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_15_13__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_13__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_13__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_15_13__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_12_15__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_12_15__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_12_15__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_12_15__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_12_15__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_268
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_268__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_268__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_268__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_268__ap_ready),
    .idy(64'd13),
    .idx(64'd15),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_15_13__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_15_13__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_15_13__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_15_14__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_15_14__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_14__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_14__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_15_14__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_13_15__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_13_15__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_13_15__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_13_15__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_13_15__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_269
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_269__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_269__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_269__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_269__ap_ready),
    .idy(64'd14),
    .idx(64'd15),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_15_14__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_15_14__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_15_14__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_15_15__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_15_15__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_15__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_15__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_15_15__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_14_15__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_14_15__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_14_15__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_14_15__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_14_15__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_270
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_270__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_270__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_270__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_270__ap_ready),
    .idx(64'd15),
    .idy(64'd15),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_15_15__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_15_15__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_15_15__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_15_16__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_15_16__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_16__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_16__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_15_16__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_15_15__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_15_15__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_15_15__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_15_15__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_15_15__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_271
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_271__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_271__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_271__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_271__ap_ready),
    .idx(64'd15),
    .idy(64'd16),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_15_16__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_15_16__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_15_16__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_15_17__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_15_17__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_17__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_17__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_15_17__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_16_15__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_16_15__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_16_15__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_16_15__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_16_15__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_272
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_272__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_272__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_272__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_272__ap_ready),
    .idy(64'd0),
    .idx(64'd16),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_16_0__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_16_0__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_16_0__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_16_1__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_16_1__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_1__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_1__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_16_1__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_0_16__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_0_16__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_0_16__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_0_16__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_0_16__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_273
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_273__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_273__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_273__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_273__ap_ready),
    .idy(64'd1),
    .idx(64'd16),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_16_1__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_16_1__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_16_1__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_16_2__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_16_2__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_2__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_2__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_16_2__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_1_16__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_1_16__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_1_16__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_1_16__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_1_16__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_274
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_274__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_274__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_274__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_274__ap_ready),
    .idx(64'd16),
    .idy(64'd2),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_16_2__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_16_2__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_16_2__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_16_3__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_16_3__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_3__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_3__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_16_3__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_2_16__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_2_16__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_2_16__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_2_16__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_2_16__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_275
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_275__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_275__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_275__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_275__ap_ready),
    .idx(64'd16),
    .idy(64'd3),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_16_3__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_16_3__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_16_3__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_16_4__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_16_4__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_4__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_4__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_16_4__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_3_16__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_3_16__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_3_16__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_3_16__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_3_16__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_276
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_276__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_276__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_276__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_276__ap_ready),
    .idx(64'd16),
    .idy(64'd4),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_16_4__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_16_4__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_16_4__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_16_5__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_16_5__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_5__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_5__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_16_5__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_4_16__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_4_16__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_4_16__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_4_16__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_4_16__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_277
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_277__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_277__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_277__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_277__ap_ready),
    .idx(64'd16),
    .idy(64'd5),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_16_5__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_16_5__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_16_5__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_16_6__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_16_6__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_6__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_6__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_16_6__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_5_16__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_5_16__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_5_16__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_5_16__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_5_16__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_278
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_278__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_278__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_278__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_278__ap_ready),
    .idx(64'd16),
    .idy(64'd6),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_16_6__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_16_6__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_16_6__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_16_7__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_16_7__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_7__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_7__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_16_7__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_6_16__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_6_16__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_6_16__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_6_16__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_6_16__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_279
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_279__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_279__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_279__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_279__ap_ready),
    .idx(64'd16),
    .idy(64'd7),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_16_7__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_16_7__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_16_7__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_16_8__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_16_8__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_8__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_8__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_16_8__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_7_16__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_7_16__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_7_16__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_7_16__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_7_16__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_280
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_280__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_280__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_280__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_280__ap_ready),
    .idx(64'd16),
    .idy(64'd8),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_16_8__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_16_8__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_16_8__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_16_9__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_16_9__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_9__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_9__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_16_9__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_8_16__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_8_16__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_8_16__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_8_16__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_8_16__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_281
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_281__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_281__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_281__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_281__ap_ready),
    .idx(64'd16),
    .idy(64'd9),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_16_10__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_16_10__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_10__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_10__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_16_10__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_16_9__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_16_9__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_16_9__write),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_9_16__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_9_16__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_9_16__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_9_16__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_9_16__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_282
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_282__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_282__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_282__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_282__ap_ready),
    .idy(64'd10),
    .idx(64'd16),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_16_10__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_16_10__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_16_10__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_16_11__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_16_11__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_11__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_11__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_16_11__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_10_16__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_10_16__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_10_16__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_10_16__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_10_16__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_283
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_283__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_283__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_283__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_283__ap_ready),
    .idy(64'd11),
    .idx(64'd16),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_16_11__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_16_11__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_16_11__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_16_12__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_16_12__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_12__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_12__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_16_12__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_11_16__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_11_16__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_11_16__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_11_16__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_11_16__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_284
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_284__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_284__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_284__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_284__ap_ready),
    .idy(64'd12),
    .idx(64'd16),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_16_12__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_16_12__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_16_12__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_16_13__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_16_13__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_13__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_13__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_16_13__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_12_16__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_12_16__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_12_16__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_12_16__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_12_16__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_285
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_285__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_285__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_285__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_285__ap_ready),
    .idy(64'd13),
    .idx(64'd16),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_16_13__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_16_13__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_16_13__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_16_14__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_16_14__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_14__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_14__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_16_14__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_13_16__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_13_16__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_13_16__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_13_16__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_13_16__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_286
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_286__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_286__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_286__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_286__ap_ready),
    .idy(64'd14),
    .idx(64'd16),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_16_14__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_16_14__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_16_14__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_16_15__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_16_15__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_15__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_15__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_16_15__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_14_16__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_14_16__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_14_16__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_14_16__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_14_16__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_287
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_287__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_287__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_287__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_287__ap_ready),
    .idy(64'd15),
    .idx(64'd16),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_16_15__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_16_15__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_16_15__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_16_16__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_16_16__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_16__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_16__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_16_16__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_15_16__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_15_16__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_15_16__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_15_16__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_15_16__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L1_out_wrapper
  C_drain_IO_L1_out_wrapper_288
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L1_out_wrapper_288__ap_start),
    .ap_done(C_drain_IO_L1_out_wrapper_288__ap_done),
    .ap_idle(C_drain_IO_L1_out_wrapper_288__ap_idle),
    .ap_ready(C_drain_IO_L1_out_wrapper_288__ap_ready),
    .idx(64'd16),
    .idy(64'd16),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L1_out_16_16__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L1_out_16_16__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L1_out_16_16__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_16_17__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_16_17__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_17__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_17__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L1_out_16_17__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_PE_16_16__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_PE_16_16__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_PE_16_16__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_PE_16_16__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_PE_16_16__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L2_out
  C_drain_IO_L2_out_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L2_out_0__ap_start),
    .ap_done(C_drain_IO_L2_out_0__ap_done),
    .ap_idle(C_drain_IO_L2_out_0__ap_idle),
    .ap_ready(C_drain_IO_L2_out_0__ap_ready),
    .idx(64'd0),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_0_0__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_0_0__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_0__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_0_0__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_C_drain_IO_L1_out_0_0__read),
    .fifo_C_drain_local_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L2_out_0__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L2_out_0__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L2_out_0__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L2_out_1__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L2_out_1__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L2_out_1__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L2_out_1__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L2_out_1__read),
    .fifo_C_drain_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L2_out
  C_drain_IO_L2_out_1
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L2_out_1__ap_start),
    .ap_done(C_drain_IO_L2_out_1__ap_done),
    .ap_idle(C_drain_IO_L2_out_1__ap_idle),
    .ap_ready(C_drain_IO_L2_out_1__ap_ready),
    .idx(64'd1),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_1_0__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_1_0__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_0__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_1_0__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_C_drain_IO_L1_out_1_0__read),
    .fifo_C_drain_local_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L2_out_1__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L2_out_1__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L2_out_1__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L2_out_2__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L2_out_2__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L2_out_2__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L2_out_2__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L2_out_2__read),
    .fifo_C_drain_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L2_out
  C_drain_IO_L2_out_2
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L2_out_2__ap_start),
    .ap_done(C_drain_IO_L2_out_2__ap_done),
    .ap_idle(C_drain_IO_L2_out_2__ap_idle),
    .ap_ready(C_drain_IO_L2_out_2__ap_ready),
    .idx(64'd2),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_2_0__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_2_0__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_0__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_2_0__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_C_drain_IO_L1_out_2_0__read),
    .fifo_C_drain_local_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L2_out_2__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L2_out_2__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L2_out_2__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L2_out_3__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L2_out_3__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L2_out_3__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L2_out_3__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L2_out_3__read),
    .fifo_C_drain_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L2_out
  C_drain_IO_L2_out_3
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L2_out_3__ap_start),
    .ap_done(C_drain_IO_L2_out_3__ap_done),
    .ap_idle(C_drain_IO_L2_out_3__ap_idle),
    .ap_ready(C_drain_IO_L2_out_3__ap_ready),
    .idx(64'd3),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_3_0__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_3_0__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_0__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_3_0__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_C_drain_IO_L1_out_3_0__read),
    .fifo_C_drain_local_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L2_out_3__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L2_out_3__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L2_out_3__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L2_out_4__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L2_out_4__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L2_out_4__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L2_out_4__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L2_out_4__read),
    .fifo_C_drain_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L2_out
  C_drain_IO_L2_out_4
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L2_out_4__ap_start),
    .ap_done(C_drain_IO_L2_out_4__ap_done),
    .ap_idle(C_drain_IO_L2_out_4__ap_idle),
    .ap_ready(C_drain_IO_L2_out_4__ap_ready),
    .idx(64'd4),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_4_0__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_4_0__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_0__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_4_0__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_C_drain_IO_L1_out_4_0__read),
    .fifo_C_drain_local_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L2_out_4__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L2_out_4__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L2_out_4__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L2_out_5__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L2_out_5__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L2_out_5__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L2_out_5__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L2_out_5__read),
    .fifo_C_drain_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L2_out
  C_drain_IO_L2_out_5
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L2_out_5__ap_start),
    .ap_done(C_drain_IO_L2_out_5__ap_done),
    .ap_idle(C_drain_IO_L2_out_5__ap_idle),
    .ap_ready(C_drain_IO_L2_out_5__ap_ready),
    .idx(64'd5),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_5_0__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_5_0__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_0__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_5_0__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_C_drain_IO_L1_out_5_0__read),
    .fifo_C_drain_local_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L2_out_5__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L2_out_5__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L2_out_5__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L2_out_6__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L2_out_6__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L2_out_6__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L2_out_6__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L2_out_6__read),
    .fifo_C_drain_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L2_out
  C_drain_IO_L2_out_6
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L2_out_6__ap_start),
    .ap_done(C_drain_IO_L2_out_6__ap_done),
    .ap_idle(C_drain_IO_L2_out_6__ap_idle),
    .ap_ready(C_drain_IO_L2_out_6__ap_ready),
    .idx(64'd6),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_6_0__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_6_0__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_0__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_6_0__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_C_drain_IO_L1_out_6_0__read),
    .fifo_C_drain_local_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L2_out_6__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L2_out_6__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L2_out_6__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L2_out_7__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L2_out_7__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L2_out_7__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L2_out_7__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L2_out_7__read),
    .fifo_C_drain_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L2_out
  C_drain_IO_L2_out_7
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L2_out_7__ap_start),
    .ap_done(C_drain_IO_L2_out_7__ap_done),
    .ap_idle(C_drain_IO_L2_out_7__ap_idle),
    .ap_ready(C_drain_IO_L2_out_7__ap_ready),
    .idx(64'd7),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_7_0__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_7_0__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_0__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_7_0__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_C_drain_IO_L1_out_7_0__read),
    .fifo_C_drain_local_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L2_out_7__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L2_out_7__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L2_out_7__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L2_out_8__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L2_out_8__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L2_out_8__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L2_out_8__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L2_out_8__read),
    .fifo_C_drain_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L2_out
  C_drain_IO_L2_out_8
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L2_out_8__ap_start),
    .ap_done(C_drain_IO_L2_out_8__ap_done),
    .ap_idle(C_drain_IO_L2_out_8__ap_idle),
    .ap_ready(C_drain_IO_L2_out_8__ap_ready),
    .idx(64'd8),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_8_0__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_8_0__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_0__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_8_0__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_C_drain_IO_L1_out_8_0__read),
    .fifo_C_drain_local_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L2_out_8__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L2_out_8__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L2_out_8__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L2_out_9__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L2_out_9__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L2_out_9__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L2_out_9__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L2_out_9__read),
    .fifo_C_drain_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L2_out
  C_drain_IO_L2_out_9
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L2_out_9__ap_start),
    .ap_done(C_drain_IO_L2_out_9__ap_done),
    .ap_idle(C_drain_IO_L2_out_9__ap_idle),
    .ap_ready(C_drain_IO_L2_out_9__ap_ready),
    .idx(64'd9),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_9_0__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_9_0__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_0__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_9_0__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_C_drain_IO_L1_out_9_0__read),
    .fifo_C_drain_local_in_peek_read(),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L2_out_10__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L2_out_10__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L2_out_10__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L2_out_10__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L2_out_10__read),
    .fifo_C_drain_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L2_out_9__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L2_out_9__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L2_out_9__write)
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L2_out
  C_drain_IO_L2_out_10
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L2_out_10__ap_start),
    .ap_done(C_drain_IO_L2_out_10__ap_done),
    .ap_idle(C_drain_IO_L2_out_10__ap_idle),
    .ap_ready(C_drain_IO_L2_out_10__ap_ready),
    .idx(64'd10),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_10_0__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_10_0__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_0__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_10_0__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_C_drain_IO_L1_out_10_0__read),
    .fifo_C_drain_local_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L2_out_10__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L2_out_10__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L2_out_10__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L2_out_11__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L2_out_11__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L2_out_11__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L2_out_11__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L2_out_11__read),
    .fifo_C_drain_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L2_out
  C_drain_IO_L2_out_11
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L2_out_11__ap_start),
    .ap_done(C_drain_IO_L2_out_11__ap_done),
    .ap_idle(C_drain_IO_L2_out_11__ap_idle),
    .ap_ready(C_drain_IO_L2_out_11__ap_ready),
    .idx(64'd11),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_11_0__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_11_0__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_0__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_11_0__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_C_drain_IO_L1_out_11_0__read),
    .fifo_C_drain_local_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L2_out_11__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L2_out_11__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L2_out_11__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L2_out_12__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L2_out_12__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L2_out_12__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L2_out_12__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L2_out_12__read),
    .fifo_C_drain_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L2_out
  C_drain_IO_L2_out_12
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L2_out_12__ap_start),
    .ap_done(C_drain_IO_L2_out_12__ap_done),
    .ap_idle(C_drain_IO_L2_out_12__ap_idle),
    .ap_ready(C_drain_IO_L2_out_12__ap_ready),
    .idx(64'd12),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_12_0__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_12_0__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_0__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_12_0__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_C_drain_IO_L1_out_12_0__read),
    .fifo_C_drain_local_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L2_out_12__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L2_out_12__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L2_out_12__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L2_out_13__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L2_out_13__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L2_out_13__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L2_out_13__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L2_out_13__read),
    .fifo_C_drain_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L2_out
  C_drain_IO_L2_out_13
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L2_out_13__ap_start),
    .ap_done(C_drain_IO_L2_out_13__ap_done),
    .ap_idle(C_drain_IO_L2_out_13__ap_idle),
    .ap_ready(C_drain_IO_L2_out_13__ap_ready),
    .idx(64'd13),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_13_0__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_13_0__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_0__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_13_0__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_C_drain_IO_L1_out_13_0__read),
    .fifo_C_drain_local_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L2_out_13__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L2_out_13__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L2_out_13__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L2_out_14__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L2_out_14__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L2_out_14__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L2_out_14__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L2_out_14__read),
    .fifo_C_drain_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L2_out
  C_drain_IO_L2_out_14
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L2_out_14__ap_start),
    .ap_done(C_drain_IO_L2_out_14__ap_done),
    .ap_idle(C_drain_IO_L2_out_14__ap_idle),
    .ap_ready(C_drain_IO_L2_out_14__ap_ready),
    .idx(64'd14),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_14_0__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_14_0__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_0__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_14_0__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_C_drain_IO_L1_out_14_0__read),
    .fifo_C_drain_local_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L2_out_14__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L2_out_14__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L2_out_14__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L2_out_15__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L2_out_15__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L2_out_15__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L2_out_15__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L2_out_15__read),
    .fifo_C_drain_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L2_out
  C_drain_IO_L2_out_15
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L2_out_15__ap_start),
    .ap_done(C_drain_IO_L2_out_15__ap_done),
    .ap_idle(C_drain_IO_L2_out_15__ap_idle),
    .ap_ready(C_drain_IO_L2_out_15__ap_ready),
    .idx(64'd15),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_15_0__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_15_0__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_0__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_15_0__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_C_drain_IO_L1_out_15_0__read),
    .fifo_C_drain_local_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L2_out_15__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L2_out_15__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L2_out_15__write),
    .fifo_C_drain_in_s_dout(fifo_C_drain_C_drain_IO_L2_out_16__dout),
    .fifo_C_drain_in_peek_dout(fifo_C_drain_C_drain_IO_L2_out_16__dout),
    .fifo_C_drain_in_s_empty_n(fifo_C_drain_C_drain_IO_L2_out_16__empty_n),
    .fifo_C_drain_in_peek_empty_n(fifo_C_drain_C_drain_IO_L2_out_16__empty_n),
    .fifo_C_drain_in_s_read(fifo_C_drain_C_drain_IO_L2_out_16__read),
    .fifo_C_drain_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L2_out_boundary
  C_drain_IO_L2_out_boundary_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L2_out_boundary_0__ap_start),
    .ap_done(C_drain_IO_L2_out_boundary_0__ap_done),
    .ap_idle(C_drain_IO_L2_out_boundary_0__ap_idle),
    .ap_ready(C_drain_IO_L2_out_boundary_0__ap_ready),
    .idx(64'd16),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_C_drain_IO_L1_out_16_0__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_C_drain_IO_L1_out_16_0__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_0__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_C_drain_IO_L1_out_16_0__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_C_drain_IO_L1_out_16_0__read),
    .fifo_C_drain_local_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L2_out_16__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L2_out_16__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L2_out_16__write)
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L3_out
  C_drain_IO_L3_out_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L3_out_0__ap_start),
    .ap_done(C_drain_IO_L3_out_0__ap_done),
    .ap_idle(C_drain_IO_L3_out_0__ap_idle),
    .ap_ready(C_drain_IO_L3_out_0__ap_ready),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_C_drain_IO_L2_out_0__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_C_drain_IO_L2_out_0__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_C_drain_IO_L2_out_0__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_C_drain_IO_L2_out_0__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_C_drain_IO_L2_out_0__read),
    .fifo_C_drain_local_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_C_drain_IO_L3_out_serialize__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_C_drain_IO_L3_out_serialize__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_C_drain_IO_L3_out_serialize__write)
  );


  (* keep_hierarchy = "yes" *) C_drain_IO_L3_out_serialize
  C_drain_IO_L3_out_serialize_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(C_drain_IO_L3_out_serialize_0__ap_start),
    .ap_done(C_drain_IO_L3_out_serialize_0__ap_done),
    .ap_idle(C_drain_IO_L3_out_serialize_0__ap_idle),
    .ap_ready(C_drain_IO_L3_out_serialize_0__ap_ready),
    .m_axi_C_ARADDR(m_axi_C_ARADDR),
    .m_axi_C_ARBURST(m_axi_C_ARBURST),
    .m_axi_C_ARID(m_axi_C_ARID),
    .m_axi_C_ARLEN(m_axi_C_ARLEN),
    .m_axi_C_ARREADY(m_axi_C_ARREADY),
    .m_axi_C_ARSIZE(m_axi_C_ARSIZE),
    .m_axi_C_ARVALID(m_axi_C_ARVALID),
    .m_axi_C_AWADDR(m_axi_C_AWADDR),
    .m_axi_C_AWBURST(m_axi_C_AWBURST),
    .m_axi_C_AWID(m_axi_C_AWID),
    .m_axi_C_AWLEN(m_axi_C_AWLEN),
    .m_axi_C_AWREADY(m_axi_C_AWREADY),
    .m_axi_C_AWSIZE(m_axi_C_AWSIZE),
    .m_axi_C_AWVALID(m_axi_C_AWVALID),
    .m_axi_C_BID(m_axi_C_BID),
    .m_axi_C_BREADY(m_axi_C_BREADY),
    .m_axi_C_BRESP(m_axi_C_BRESP),
    .m_axi_C_BVALID(m_axi_C_BVALID),
    .m_axi_C_RDATA(m_axi_C_RDATA),
    .m_axi_C_RID(m_axi_C_RID),
    .m_axi_C_RLAST(m_axi_C_RLAST),
    .m_axi_C_RREADY(m_axi_C_RREADY),
    .m_axi_C_RRESP(m_axi_C_RRESP),
    .m_axi_C_RVALID(m_axi_C_RVALID),
    .m_axi_C_WDATA(m_axi_C_WDATA),
    .m_axi_C_WLAST(m_axi_C_WLAST),
    .m_axi_C_WREADY(m_axi_C_WREADY),
    .m_axi_C_WSTRB(m_axi_C_WSTRB),
    .m_axi_C_WVALID(m_axi_C_WVALID),
    .m_axi_C_ARLOCK(m_axi_C_ARLOCK),
    .m_axi_C_ARPROT(m_axi_C_ARPROT),
    .m_axi_C_ARQOS(m_axi_C_ARQOS),
    .m_axi_C_ARCACHE(m_axi_C_ARCACHE),
    .m_axi_C_AWCACHE(m_axi_C_AWCACHE),
    .m_axi_C_AWLOCK(m_axi_C_AWLOCK),
    .m_axi_C_AWPROT(m_axi_C_AWPROT),
    .m_axi_C_AWQOS(m_axi_C_AWQOS),
    .C_offset(C_drain_IO_L3_out_serialize_0___C__q0),
    .fifo_C_drain_local_in_s_dout(fifo_C_drain_C_drain_IO_L3_out_serialize__dout),
    .fifo_C_drain_local_in_peek_dout(fifo_C_drain_C_drain_IO_L3_out_serialize__dout),
    .fifo_C_drain_local_in_s_empty_n(fifo_C_drain_C_drain_IO_L3_out_serialize__empty_n),
    .fifo_C_drain_local_in_peek_empty_n(fifo_C_drain_C_drain_IO_L3_out_serialize__empty_n),
    .fifo_C_drain_local_in_s_read(fifo_C_drain_C_drain_IO_L3_out_serialize__read),
    .fifo_C_drain_local_in_peek_read()
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_0__ap_start),
    .ap_done(PE_wrapper_0__ap_done),
    .ap_idle(PE_wrapper_0__ap_idle),
    .ap_ready(PE_wrapper_0__ap_ready),
    .idx(64'd0),
    .idy(64'd0),
    .fifo_A_in_s_dout(fifo_A_PE_0_0__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_0_0__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_0_0__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_0_0__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_0_0__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_0_1__din),
    .fifo_A_out_full_n(fifo_A_PE_0_1__full_n),
    .fifo_A_out_write(fifo_A_PE_0_1__write),
    .fifo_B_in_s_dout(fifo_B_PE_0_0__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_0_0__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_0_0__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_0_0__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_0_0__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_1_0__din),
    .fifo_B_out_full_n(fifo_B_PE_1_0__full_n),
    .fifo_B_out_write(fifo_B_PE_1_0__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_0_0__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_0_0__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_0_0__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_1
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_1__ap_start),
    .ap_done(PE_wrapper_1__ap_done),
    .ap_idle(PE_wrapper_1__ap_idle),
    .ap_ready(PE_wrapper_1__ap_ready),
    .idx(64'd0),
    .idy(64'd1),
    .fifo_A_in_s_dout(fifo_A_PE_0_1__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_0_1__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_0_1__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_0_1__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_0_1__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_0_2__din),
    .fifo_A_out_full_n(fifo_A_PE_0_2__full_n),
    .fifo_A_out_write(fifo_A_PE_0_2__write),
    .fifo_B_in_s_dout(fifo_B_PE_0_1__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_0_1__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_0_1__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_0_1__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_0_1__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_1_1__din),
    .fifo_B_out_full_n(fifo_B_PE_1_1__full_n),
    .fifo_B_out_write(fifo_B_PE_1_1__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_0_1__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_0_1__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_0_1__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_2
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_2__ap_start),
    .ap_done(PE_wrapper_2__ap_done),
    .ap_idle(PE_wrapper_2__ap_idle),
    .ap_ready(PE_wrapper_2__ap_ready),
    .idx(64'd0),
    .idy(64'd2),
    .fifo_A_in_s_dout(fifo_A_PE_0_2__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_0_2__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_0_2__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_0_2__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_0_2__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_0_3__din),
    .fifo_A_out_full_n(fifo_A_PE_0_3__full_n),
    .fifo_A_out_write(fifo_A_PE_0_3__write),
    .fifo_B_in_s_dout(fifo_B_PE_0_2__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_0_2__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_0_2__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_0_2__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_0_2__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_1_2__din),
    .fifo_B_out_full_n(fifo_B_PE_1_2__full_n),
    .fifo_B_out_write(fifo_B_PE_1_2__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_0_2__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_0_2__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_0_2__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_3
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_3__ap_start),
    .ap_done(PE_wrapper_3__ap_done),
    .ap_idle(PE_wrapper_3__ap_idle),
    .ap_ready(PE_wrapper_3__ap_ready),
    .idx(64'd0),
    .idy(64'd3),
    .fifo_A_in_s_dout(fifo_A_PE_0_3__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_0_3__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_0_3__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_0_3__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_0_3__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_0_4__din),
    .fifo_A_out_full_n(fifo_A_PE_0_4__full_n),
    .fifo_A_out_write(fifo_A_PE_0_4__write),
    .fifo_B_in_s_dout(fifo_B_PE_0_3__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_0_3__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_0_3__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_0_3__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_0_3__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_1_3__din),
    .fifo_B_out_full_n(fifo_B_PE_1_3__full_n),
    .fifo_B_out_write(fifo_B_PE_1_3__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_0_3__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_0_3__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_0_3__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_4
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_4__ap_start),
    .ap_done(PE_wrapper_4__ap_done),
    .ap_idle(PE_wrapper_4__ap_idle),
    .ap_ready(PE_wrapper_4__ap_ready),
    .idx(64'd0),
    .idy(64'd4),
    .fifo_A_in_s_dout(fifo_A_PE_0_4__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_0_4__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_0_4__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_0_4__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_0_4__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_0_5__din),
    .fifo_A_out_full_n(fifo_A_PE_0_5__full_n),
    .fifo_A_out_write(fifo_A_PE_0_5__write),
    .fifo_B_in_s_dout(fifo_B_PE_0_4__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_0_4__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_0_4__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_0_4__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_0_4__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_1_4__din),
    .fifo_B_out_full_n(fifo_B_PE_1_4__full_n),
    .fifo_B_out_write(fifo_B_PE_1_4__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_0_4__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_0_4__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_0_4__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_5
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_5__ap_start),
    .ap_done(PE_wrapper_5__ap_done),
    .ap_idle(PE_wrapper_5__ap_idle),
    .ap_ready(PE_wrapper_5__ap_ready),
    .idx(64'd0),
    .idy(64'd5),
    .fifo_A_in_s_dout(fifo_A_PE_0_5__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_0_5__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_0_5__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_0_5__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_0_5__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_0_6__din),
    .fifo_A_out_full_n(fifo_A_PE_0_6__full_n),
    .fifo_A_out_write(fifo_A_PE_0_6__write),
    .fifo_B_in_s_dout(fifo_B_PE_0_5__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_0_5__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_0_5__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_0_5__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_0_5__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_1_5__din),
    .fifo_B_out_full_n(fifo_B_PE_1_5__full_n),
    .fifo_B_out_write(fifo_B_PE_1_5__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_0_5__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_0_5__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_0_5__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_6
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_6__ap_start),
    .ap_done(PE_wrapper_6__ap_done),
    .ap_idle(PE_wrapper_6__ap_idle),
    .ap_ready(PE_wrapper_6__ap_ready),
    .idx(64'd0),
    .idy(64'd6),
    .fifo_A_in_s_dout(fifo_A_PE_0_6__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_0_6__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_0_6__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_0_6__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_0_6__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_0_7__din),
    .fifo_A_out_full_n(fifo_A_PE_0_7__full_n),
    .fifo_A_out_write(fifo_A_PE_0_7__write),
    .fifo_B_in_s_dout(fifo_B_PE_0_6__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_0_6__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_0_6__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_0_6__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_0_6__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_1_6__din),
    .fifo_B_out_full_n(fifo_B_PE_1_6__full_n),
    .fifo_B_out_write(fifo_B_PE_1_6__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_0_6__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_0_6__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_0_6__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_7
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_7__ap_start),
    .ap_done(PE_wrapper_7__ap_done),
    .ap_idle(PE_wrapper_7__ap_idle),
    .ap_ready(PE_wrapper_7__ap_ready),
    .idx(64'd0),
    .idy(64'd7),
    .fifo_A_in_s_dout(fifo_A_PE_0_7__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_0_7__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_0_7__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_0_7__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_0_7__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_0_8__din),
    .fifo_A_out_full_n(fifo_A_PE_0_8__full_n),
    .fifo_A_out_write(fifo_A_PE_0_8__write),
    .fifo_B_in_s_dout(fifo_B_PE_0_7__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_0_7__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_0_7__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_0_7__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_0_7__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_1_7__din),
    .fifo_B_out_full_n(fifo_B_PE_1_7__full_n),
    .fifo_B_out_write(fifo_B_PE_1_7__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_0_7__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_0_7__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_0_7__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_8
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_8__ap_start),
    .ap_done(PE_wrapper_8__ap_done),
    .ap_idle(PE_wrapper_8__ap_idle),
    .ap_ready(PE_wrapper_8__ap_ready),
    .idx(64'd0),
    .idy(64'd8),
    .fifo_A_in_s_dout(fifo_A_PE_0_8__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_0_8__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_0_8__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_0_8__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_0_8__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_0_9__din),
    .fifo_A_out_full_n(fifo_A_PE_0_9__full_n),
    .fifo_A_out_write(fifo_A_PE_0_9__write),
    .fifo_B_in_s_dout(fifo_B_PE_0_8__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_0_8__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_0_8__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_0_8__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_0_8__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_1_8__din),
    .fifo_B_out_full_n(fifo_B_PE_1_8__full_n),
    .fifo_B_out_write(fifo_B_PE_1_8__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_0_8__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_0_8__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_0_8__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_9
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_9__ap_start),
    .ap_done(PE_wrapper_9__ap_done),
    .ap_idle(PE_wrapper_9__ap_idle),
    .ap_ready(PE_wrapper_9__ap_ready),
    .idx(64'd0),
    .idy(64'd9),
    .fifo_A_out_din(fifo_A_PE_0_10__din),
    .fifo_A_out_full_n(fifo_A_PE_0_10__full_n),
    .fifo_A_out_write(fifo_A_PE_0_10__write),
    .fifo_A_in_s_dout(fifo_A_PE_0_9__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_0_9__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_0_9__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_0_9__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_0_9__read),
    .fifo_A_in_peek_read(),
    .fifo_B_in_s_dout(fifo_B_PE_0_9__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_0_9__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_0_9__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_0_9__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_0_9__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_1_9__din),
    .fifo_B_out_full_n(fifo_B_PE_1_9__full_n),
    .fifo_B_out_write(fifo_B_PE_1_9__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_0_9__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_0_9__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_0_9__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_10
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_10__ap_start),
    .ap_done(PE_wrapper_10__ap_done),
    .ap_idle(PE_wrapper_10__ap_idle),
    .ap_ready(PE_wrapper_10__ap_ready),
    .idx(64'd0),
    .idy(64'd10),
    .fifo_A_in_s_dout(fifo_A_PE_0_10__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_0_10__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_0_10__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_0_10__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_0_10__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_0_11__din),
    .fifo_A_out_full_n(fifo_A_PE_0_11__full_n),
    .fifo_A_out_write(fifo_A_PE_0_11__write),
    .fifo_B_in_s_dout(fifo_B_PE_0_10__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_0_10__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_0_10__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_0_10__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_0_10__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_1_10__din),
    .fifo_B_out_full_n(fifo_B_PE_1_10__full_n),
    .fifo_B_out_write(fifo_B_PE_1_10__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_0_10__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_0_10__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_0_10__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_11
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_11__ap_start),
    .ap_done(PE_wrapper_11__ap_done),
    .ap_idle(PE_wrapper_11__ap_idle),
    .ap_ready(PE_wrapper_11__ap_ready),
    .idx(64'd0),
    .idy(64'd11),
    .fifo_A_in_s_dout(fifo_A_PE_0_11__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_0_11__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_0_11__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_0_11__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_0_11__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_0_12__din),
    .fifo_A_out_full_n(fifo_A_PE_0_12__full_n),
    .fifo_A_out_write(fifo_A_PE_0_12__write),
    .fifo_B_in_s_dout(fifo_B_PE_0_11__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_0_11__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_0_11__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_0_11__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_0_11__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_1_11__din),
    .fifo_B_out_full_n(fifo_B_PE_1_11__full_n),
    .fifo_B_out_write(fifo_B_PE_1_11__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_0_11__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_0_11__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_0_11__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_12
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_12__ap_start),
    .ap_done(PE_wrapper_12__ap_done),
    .ap_idle(PE_wrapper_12__ap_idle),
    .ap_ready(PE_wrapper_12__ap_ready),
    .idx(64'd0),
    .idy(64'd12),
    .fifo_A_in_s_dout(fifo_A_PE_0_12__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_0_12__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_0_12__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_0_12__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_0_12__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_0_13__din),
    .fifo_A_out_full_n(fifo_A_PE_0_13__full_n),
    .fifo_A_out_write(fifo_A_PE_0_13__write),
    .fifo_B_in_s_dout(fifo_B_PE_0_12__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_0_12__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_0_12__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_0_12__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_0_12__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_1_12__din),
    .fifo_B_out_full_n(fifo_B_PE_1_12__full_n),
    .fifo_B_out_write(fifo_B_PE_1_12__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_0_12__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_0_12__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_0_12__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_13
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_13__ap_start),
    .ap_done(PE_wrapper_13__ap_done),
    .ap_idle(PE_wrapper_13__ap_idle),
    .ap_ready(PE_wrapper_13__ap_ready),
    .idx(64'd0),
    .idy(64'd13),
    .fifo_A_in_s_dout(fifo_A_PE_0_13__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_0_13__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_0_13__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_0_13__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_0_13__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_0_14__din),
    .fifo_A_out_full_n(fifo_A_PE_0_14__full_n),
    .fifo_A_out_write(fifo_A_PE_0_14__write),
    .fifo_B_in_s_dout(fifo_B_PE_0_13__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_0_13__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_0_13__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_0_13__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_0_13__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_1_13__din),
    .fifo_B_out_full_n(fifo_B_PE_1_13__full_n),
    .fifo_B_out_write(fifo_B_PE_1_13__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_0_13__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_0_13__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_0_13__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_14
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_14__ap_start),
    .ap_done(PE_wrapper_14__ap_done),
    .ap_idle(PE_wrapper_14__ap_idle),
    .ap_ready(PE_wrapper_14__ap_ready),
    .idx(64'd0),
    .idy(64'd14),
    .fifo_A_in_s_dout(fifo_A_PE_0_14__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_0_14__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_0_14__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_0_14__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_0_14__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_0_15__din),
    .fifo_A_out_full_n(fifo_A_PE_0_15__full_n),
    .fifo_A_out_write(fifo_A_PE_0_15__write),
    .fifo_B_in_s_dout(fifo_B_PE_0_14__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_0_14__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_0_14__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_0_14__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_0_14__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_1_14__din),
    .fifo_B_out_full_n(fifo_B_PE_1_14__full_n),
    .fifo_B_out_write(fifo_B_PE_1_14__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_0_14__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_0_14__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_0_14__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_15
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_15__ap_start),
    .ap_done(PE_wrapper_15__ap_done),
    .ap_idle(PE_wrapper_15__ap_idle),
    .ap_ready(PE_wrapper_15__ap_ready),
    .idx(64'd0),
    .idy(64'd15),
    .fifo_A_in_s_dout(fifo_A_PE_0_15__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_0_15__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_0_15__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_0_15__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_0_15__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_0_16__din),
    .fifo_A_out_full_n(fifo_A_PE_0_16__full_n),
    .fifo_A_out_write(fifo_A_PE_0_16__write),
    .fifo_B_in_s_dout(fifo_B_PE_0_15__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_0_15__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_0_15__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_0_15__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_0_15__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_1_15__din),
    .fifo_B_out_full_n(fifo_B_PE_1_15__full_n),
    .fifo_B_out_write(fifo_B_PE_1_15__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_0_15__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_0_15__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_0_15__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_16
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_16__ap_start),
    .ap_done(PE_wrapper_16__ap_done),
    .ap_idle(PE_wrapper_16__ap_idle),
    .ap_ready(PE_wrapper_16__ap_ready),
    .idx(64'd0),
    .idy(64'd16),
    .fifo_A_in_s_dout(fifo_A_PE_0_16__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_0_16__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_0_16__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_0_16__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_0_16__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_0_17__din),
    .fifo_A_out_full_n(fifo_A_PE_0_17__full_n),
    .fifo_A_out_write(fifo_A_PE_0_17__write),
    .fifo_B_in_s_dout(fifo_B_PE_0_16__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_0_16__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_0_16__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_0_16__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_0_16__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_1_16__din),
    .fifo_B_out_full_n(fifo_B_PE_1_16__full_n),
    .fifo_B_out_write(fifo_B_PE_1_16__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_0_16__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_0_16__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_0_16__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_17
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_17__ap_start),
    .ap_done(PE_wrapper_17__ap_done),
    .ap_idle(PE_wrapper_17__ap_idle),
    .ap_ready(PE_wrapper_17__ap_ready),
    .idy(64'd0),
    .idx(64'd1),
    .fifo_A_in_s_dout(fifo_A_PE_1_0__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_1_0__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_1_0__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_1_0__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_1_0__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_1_1__din),
    .fifo_A_out_full_n(fifo_A_PE_1_1__full_n),
    .fifo_A_out_write(fifo_A_PE_1_1__write),
    .fifo_B_in_s_dout(fifo_B_PE_1_0__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_1_0__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_1_0__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_1_0__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_1_0__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_2_0__din),
    .fifo_B_out_full_n(fifo_B_PE_2_0__full_n),
    .fifo_B_out_write(fifo_B_PE_2_0__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_1_0__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_1_0__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_1_0__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_18
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_18__ap_start),
    .ap_done(PE_wrapper_18__ap_done),
    .ap_idle(PE_wrapper_18__ap_idle),
    .ap_ready(PE_wrapper_18__ap_ready),
    .idx(64'd1),
    .idy(64'd1),
    .fifo_A_in_s_dout(fifo_A_PE_1_1__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_1_1__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_1_1__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_1_1__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_1_1__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_1_2__din),
    .fifo_A_out_full_n(fifo_A_PE_1_2__full_n),
    .fifo_A_out_write(fifo_A_PE_1_2__write),
    .fifo_B_in_s_dout(fifo_B_PE_1_1__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_1_1__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_1_1__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_1_1__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_1_1__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_2_1__din),
    .fifo_B_out_full_n(fifo_B_PE_2_1__full_n),
    .fifo_B_out_write(fifo_B_PE_2_1__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_1_1__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_1_1__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_1_1__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_19
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_19__ap_start),
    .ap_done(PE_wrapper_19__ap_done),
    .ap_idle(PE_wrapper_19__ap_idle),
    .ap_ready(PE_wrapper_19__ap_ready),
    .idx(64'd1),
    .idy(64'd2),
    .fifo_A_in_s_dout(fifo_A_PE_1_2__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_1_2__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_1_2__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_1_2__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_1_2__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_1_3__din),
    .fifo_A_out_full_n(fifo_A_PE_1_3__full_n),
    .fifo_A_out_write(fifo_A_PE_1_3__write),
    .fifo_B_in_s_dout(fifo_B_PE_1_2__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_1_2__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_1_2__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_1_2__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_1_2__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_2_2__din),
    .fifo_B_out_full_n(fifo_B_PE_2_2__full_n),
    .fifo_B_out_write(fifo_B_PE_2_2__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_1_2__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_1_2__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_1_2__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_20
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_20__ap_start),
    .ap_done(PE_wrapper_20__ap_done),
    .ap_idle(PE_wrapper_20__ap_idle),
    .ap_ready(PE_wrapper_20__ap_ready),
    .idx(64'd1),
    .idy(64'd3),
    .fifo_A_in_s_dout(fifo_A_PE_1_3__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_1_3__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_1_3__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_1_3__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_1_3__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_1_4__din),
    .fifo_A_out_full_n(fifo_A_PE_1_4__full_n),
    .fifo_A_out_write(fifo_A_PE_1_4__write),
    .fifo_B_in_s_dout(fifo_B_PE_1_3__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_1_3__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_1_3__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_1_3__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_1_3__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_2_3__din),
    .fifo_B_out_full_n(fifo_B_PE_2_3__full_n),
    .fifo_B_out_write(fifo_B_PE_2_3__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_1_3__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_1_3__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_1_3__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_21
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_21__ap_start),
    .ap_done(PE_wrapper_21__ap_done),
    .ap_idle(PE_wrapper_21__ap_idle),
    .ap_ready(PE_wrapper_21__ap_ready),
    .idx(64'd1),
    .idy(64'd4),
    .fifo_A_in_s_dout(fifo_A_PE_1_4__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_1_4__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_1_4__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_1_4__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_1_4__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_1_5__din),
    .fifo_A_out_full_n(fifo_A_PE_1_5__full_n),
    .fifo_A_out_write(fifo_A_PE_1_5__write),
    .fifo_B_in_s_dout(fifo_B_PE_1_4__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_1_4__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_1_4__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_1_4__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_1_4__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_2_4__din),
    .fifo_B_out_full_n(fifo_B_PE_2_4__full_n),
    .fifo_B_out_write(fifo_B_PE_2_4__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_1_4__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_1_4__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_1_4__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_22
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_22__ap_start),
    .ap_done(PE_wrapper_22__ap_done),
    .ap_idle(PE_wrapper_22__ap_idle),
    .ap_ready(PE_wrapper_22__ap_ready),
    .idx(64'd1),
    .idy(64'd5),
    .fifo_A_in_s_dout(fifo_A_PE_1_5__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_1_5__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_1_5__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_1_5__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_1_5__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_1_6__din),
    .fifo_A_out_full_n(fifo_A_PE_1_6__full_n),
    .fifo_A_out_write(fifo_A_PE_1_6__write),
    .fifo_B_in_s_dout(fifo_B_PE_1_5__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_1_5__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_1_5__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_1_5__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_1_5__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_2_5__din),
    .fifo_B_out_full_n(fifo_B_PE_2_5__full_n),
    .fifo_B_out_write(fifo_B_PE_2_5__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_1_5__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_1_5__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_1_5__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_23
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_23__ap_start),
    .ap_done(PE_wrapper_23__ap_done),
    .ap_idle(PE_wrapper_23__ap_idle),
    .ap_ready(PE_wrapper_23__ap_ready),
    .idx(64'd1),
    .idy(64'd6),
    .fifo_A_in_s_dout(fifo_A_PE_1_6__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_1_6__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_1_6__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_1_6__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_1_6__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_1_7__din),
    .fifo_A_out_full_n(fifo_A_PE_1_7__full_n),
    .fifo_A_out_write(fifo_A_PE_1_7__write),
    .fifo_B_in_s_dout(fifo_B_PE_1_6__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_1_6__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_1_6__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_1_6__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_1_6__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_2_6__din),
    .fifo_B_out_full_n(fifo_B_PE_2_6__full_n),
    .fifo_B_out_write(fifo_B_PE_2_6__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_1_6__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_1_6__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_1_6__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_24
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_24__ap_start),
    .ap_done(PE_wrapper_24__ap_done),
    .ap_idle(PE_wrapper_24__ap_idle),
    .ap_ready(PE_wrapper_24__ap_ready),
    .idx(64'd1),
    .idy(64'd7),
    .fifo_A_in_s_dout(fifo_A_PE_1_7__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_1_7__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_1_7__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_1_7__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_1_7__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_1_8__din),
    .fifo_A_out_full_n(fifo_A_PE_1_8__full_n),
    .fifo_A_out_write(fifo_A_PE_1_8__write),
    .fifo_B_in_s_dout(fifo_B_PE_1_7__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_1_7__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_1_7__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_1_7__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_1_7__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_2_7__din),
    .fifo_B_out_full_n(fifo_B_PE_2_7__full_n),
    .fifo_B_out_write(fifo_B_PE_2_7__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_1_7__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_1_7__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_1_7__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_25
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_25__ap_start),
    .ap_done(PE_wrapper_25__ap_done),
    .ap_idle(PE_wrapper_25__ap_idle),
    .ap_ready(PE_wrapper_25__ap_ready),
    .idx(64'd1),
    .idy(64'd8),
    .fifo_A_in_s_dout(fifo_A_PE_1_8__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_1_8__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_1_8__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_1_8__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_1_8__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_1_9__din),
    .fifo_A_out_full_n(fifo_A_PE_1_9__full_n),
    .fifo_A_out_write(fifo_A_PE_1_9__write),
    .fifo_B_in_s_dout(fifo_B_PE_1_8__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_1_8__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_1_8__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_1_8__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_1_8__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_2_8__din),
    .fifo_B_out_full_n(fifo_B_PE_2_8__full_n),
    .fifo_B_out_write(fifo_B_PE_2_8__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_1_8__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_1_8__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_1_8__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_26
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_26__ap_start),
    .ap_done(PE_wrapper_26__ap_done),
    .ap_idle(PE_wrapper_26__ap_idle),
    .ap_ready(PE_wrapper_26__ap_ready),
    .idx(64'd1),
    .idy(64'd9),
    .fifo_A_out_din(fifo_A_PE_1_10__din),
    .fifo_A_out_full_n(fifo_A_PE_1_10__full_n),
    .fifo_A_out_write(fifo_A_PE_1_10__write),
    .fifo_A_in_s_dout(fifo_A_PE_1_9__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_1_9__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_1_9__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_1_9__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_1_9__read),
    .fifo_A_in_peek_read(),
    .fifo_B_in_s_dout(fifo_B_PE_1_9__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_1_9__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_1_9__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_1_9__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_1_9__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_2_9__din),
    .fifo_B_out_full_n(fifo_B_PE_2_9__full_n),
    .fifo_B_out_write(fifo_B_PE_2_9__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_1_9__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_1_9__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_1_9__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_27
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_27__ap_start),
    .ap_done(PE_wrapper_27__ap_done),
    .ap_idle(PE_wrapper_27__ap_idle),
    .ap_ready(PE_wrapper_27__ap_ready),
    .idx(64'd1),
    .idy(64'd10),
    .fifo_A_in_s_dout(fifo_A_PE_1_10__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_1_10__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_1_10__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_1_10__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_1_10__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_1_11__din),
    .fifo_A_out_full_n(fifo_A_PE_1_11__full_n),
    .fifo_A_out_write(fifo_A_PE_1_11__write),
    .fifo_B_in_s_dout(fifo_B_PE_1_10__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_1_10__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_1_10__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_1_10__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_1_10__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_2_10__din),
    .fifo_B_out_full_n(fifo_B_PE_2_10__full_n),
    .fifo_B_out_write(fifo_B_PE_2_10__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_1_10__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_1_10__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_1_10__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_28
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_28__ap_start),
    .ap_done(PE_wrapper_28__ap_done),
    .ap_idle(PE_wrapper_28__ap_idle),
    .ap_ready(PE_wrapper_28__ap_ready),
    .idx(64'd1),
    .idy(64'd11),
    .fifo_A_in_s_dout(fifo_A_PE_1_11__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_1_11__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_1_11__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_1_11__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_1_11__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_1_12__din),
    .fifo_A_out_full_n(fifo_A_PE_1_12__full_n),
    .fifo_A_out_write(fifo_A_PE_1_12__write),
    .fifo_B_in_s_dout(fifo_B_PE_1_11__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_1_11__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_1_11__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_1_11__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_1_11__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_2_11__din),
    .fifo_B_out_full_n(fifo_B_PE_2_11__full_n),
    .fifo_B_out_write(fifo_B_PE_2_11__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_1_11__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_1_11__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_1_11__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_29
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_29__ap_start),
    .ap_done(PE_wrapper_29__ap_done),
    .ap_idle(PE_wrapper_29__ap_idle),
    .ap_ready(PE_wrapper_29__ap_ready),
    .idx(64'd1),
    .idy(64'd12),
    .fifo_A_in_s_dout(fifo_A_PE_1_12__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_1_12__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_1_12__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_1_12__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_1_12__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_1_13__din),
    .fifo_A_out_full_n(fifo_A_PE_1_13__full_n),
    .fifo_A_out_write(fifo_A_PE_1_13__write),
    .fifo_B_in_s_dout(fifo_B_PE_1_12__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_1_12__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_1_12__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_1_12__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_1_12__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_2_12__din),
    .fifo_B_out_full_n(fifo_B_PE_2_12__full_n),
    .fifo_B_out_write(fifo_B_PE_2_12__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_1_12__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_1_12__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_1_12__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_30
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_30__ap_start),
    .ap_done(PE_wrapper_30__ap_done),
    .ap_idle(PE_wrapper_30__ap_idle),
    .ap_ready(PE_wrapper_30__ap_ready),
    .idx(64'd1),
    .idy(64'd13),
    .fifo_A_in_s_dout(fifo_A_PE_1_13__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_1_13__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_1_13__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_1_13__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_1_13__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_1_14__din),
    .fifo_A_out_full_n(fifo_A_PE_1_14__full_n),
    .fifo_A_out_write(fifo_A_PE_1_14__write),
    .fifo_B_in_s_dout(fifo_B_PE_1_13__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_1_13__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_1_13__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_1_13__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_1_13__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_2_13__din),
    .fifo_B_out_full_n(fifo_B_PE_2_13__full_n),
    .fifo_B_out_write(fifo_B_PE_2_13__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_1_13__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_1_13__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_1_13__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_31
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_31__ap_start),
    .ap_done(PE_wrapper_31__ap_done),
    .ap_idle(PE_wrapper_31__ap_idle),
    .ap_ready(PE_wrapper_31__ap_ready),
    .idx(64'd1),
    .idy(64'd14),
    .fifo_A_in_s_dout(fifo_A_PE_1_14__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_1_14__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_1_14__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_1_14__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_1_14__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_1_15__din),
    .fifo_A_out_full_n(fifo_A_PE_1_15__full_n),
    .fifo_A_out_write(fifo_A_PE_1_15__write),
    .fifo_B_in_s_dout(fifo_B_PE_1_14__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_1_14__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_1_14__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_1_14__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_1_14__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_2_14__din),
    .fifo_B_out_full_n(fifo_B_PE_2_14__full_n),
    .fifo_B_out_write(fifo_B_PE_2_14__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_1_14__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_1_14__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_1_14__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_32
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_32__ap_start),
    .ap_done(PE_wrapper_32__ap_done),
    .ap_idle(PE_wrapper_32__ap_idle),
    .ap_ready(PE_wrapper_32__ap_ready),
    .idx(64'd1),
    .idy(64'd15),
    .fifo_A_in_s_dout(fifo_A_PE_1_15__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_1_15__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_1_15__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_1_15__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_1_15__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_1_16__din),
    .fifo_A_out_full_n(fifo_A_PE_1_16__full_n),
    .fifo_A_out_write(fifo_A_PE_1_16__write),
    .fifo_B_in_s_dout(fifo_B_PE_1_15__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_1_15__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_1_15__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_1_15__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_1_15__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_2_15__din),
    .fifo_B_out_full_n(fifo_B_PE_2_15__full_n),
    .fifo_B_out_write(fifo_B_PE_2_15__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_1_15__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_1_15__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_1_15__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_33
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_33__ap_start),
    .ap_done(PE_wrapper_33__ap_done),
    .ap_idle(PE_wrapper_33__ap_idle),
    .ap_ready(PE_wrapper_33__ap_ready),
    .idx(64'd1),
    .idy(64'd16),
    .fifo_A_in_s_dout(fifo_A_PE_1_16__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_1_16__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_1_16__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_1_16__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_1_16__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_1_17__din),
    .fifo_A_out_full_n(fifo_A_PE_1_17__full_n),
    .fifo_A_out_write(fifo_A_PE_1_17__write),
    .fifo_B_in_s_dout(fifo_B_PE_1_16__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_1_16__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_1_16__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_1_16__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_1_16__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_2_16__din),
    .fifo_B_out_full_n(fifo_B_PE_2_16__full_n),
    .fifo_B_out_write(fifo_B_PE_2_16__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_1_16__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_1_16__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_1_16__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_34
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_34__ap_start),
    .ap_done(PE_wrapper_34__ap_done),
    .ap_idle(PE_wrapper_34__ap_idle),
    .ap_ready(PE_wrapper_34__ap_ready),
    .idy(64'd0),
    .idx(64'd2),
    .fifo_A_in_s_dout(fifo_A_PE_2_0__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_2_0__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_2_0__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_2_0__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_2_0__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_2_1__din),
    .fifo_A_out_full_n(fifo_A_PE_2_1__full_n),
    .fifo_A_out_write(fifo_A_PE_2_1__write),
    .fifo_B_in_s_dout(fifo_B_PE_2_0__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_2_0__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_2_0__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_2_0__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_2_0__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_3_0__din),
    .fifo_B_out_full_n(fifo_B_PE_3_0__full_n),
    .fifo_B_out_write(fifo_B_PE_3_0__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_2_0__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_2_0__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_2_0__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_35
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_35__ap_start),
    .ap_done(PE_wrapper_35__ap_done),
    .ap_idle(PE_wrapper_35__ap_idle),
    .ap_ready(PE_wrapper_35__ap_ready),
    .idy(64'd1),
    .idx(64'd2),
    .fifo_A_in_s_dout(fifo_A_PE_2_1__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_2_1__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_2_1__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_2_1__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_2_1__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_2_2__din),
    .fifo_A_out_full_n(fifo_A_PE_2_2__full_n),
    .fifo_A_out_write(fifo_A_PE_2_2__write),
    .fifo_B_in_s_dout(fifo_B_PE_2_1__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_2_1__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_2_1__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_2_1__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_2_1__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_3_1__din),
    .fifo_B_out_full_n(fifo_B_PE_3_1__full_n),
    .fifo_B_out_write(fifo_B_PE_3_1__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_2_1__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_2_1__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_2_1__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_36
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_36__ap_start),
    .ap_done(PE_wrapper_36__ap_done),
    .ap_idle(PE_wrapper_36__ap_idle),
    .ap_ready(PE_wrapper_36__ap_ready),
    .idx(64'd2),
    .idy(64'd2),
    .fifo_A_in_s_dout(fifo_A_PE_2_2__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_2_2__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_2_2__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_2_2__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_2_2__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_2_3__din),
    .fifo_A_out_full_n(fifo_A_PE_2_3__full_n),
    .fifo_A_out_write(fifo_A_PE_2_3__write),
    .fifo_B_in_s_dout(fifo_B_PE_2_2__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_2_2__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_2_2__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_2_2__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_2_2__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_3_2__din),
    .fifo_B_out_full_n(fifo_B_PE_3_2__full_n),
    .fifo_B_out_write(fifo_B_PE_3_2__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_2_2__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_2_2__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_2_2__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_37
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_37__ap_start),
    .ap_done(PE_wrapper_37__ap_done),
    .ap_idle(PE_wrapper_37__ap_idle),
    .ap_ready(PE_wrapper_37__ap_ready),
    .idx(64'd2),
    .idy(64'd3),
    .fifo_A_in_s_dout(fifo_A_PE_2_3__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_2_3__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_2_3__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_2_3__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_2_3__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_2_4__din),
    .fifo_A_out_full_n(fifo_A_PE_2_4__full_n),
    .fifo_A_out_write(fifo_A_PE_2_4__write),
    .fifo_B_in_s_dout(fifo_B_PE_2_3__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_2_3__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_2_3__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_2_3__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_2_3__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_3_3__din),
    .fifo_B_out_full_n(fifo_B_PE_3_3__full_n),
    .fifo_B_out_write(fifo_B_PE_3_3__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_2_3__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_2_3__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_2_3__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_38
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_38__ap_start),
    .ap_done(PE_wrapper_38__ap_done),
    .ap_idle(PE_wrapper_38__ap_idle),
    .ap_ready(PE_wrapper_38__ap_ready),
    .idx(64'd2),
    .idy(64'd4),
    .fifo_A_in_s_dout(fifo_A_PE_2_4__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_2_4__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_2_4__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_2_4__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_2_4__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_2_5__din),
    .fifo_A_out_full_n(fifo_A_PE_2_5__full_n),
    .fifo_A_out_write(fifo_A_PE_2_5__write),
    .fifo_B_in_s_dout(fifo_B_PE_2_4__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_2_4__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_2_4__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_2_4__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_2_4__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_3_4__din),
    .fifo_B_out_full_n(fifo_B_PE_3_4__full_n),
    .fifo_B_out_write(fifo_B_PE_3_4__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_2_4__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_2_4__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_2_4__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_39
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_39__ap_start),
    .ap_done(PE_wrapper_39__ap_done),
    .ap_idle(PE_wrapper_39__ap_idle),
    .ap_ready(PE_wrapper_39__ap_ready),
    .idx(64'd2),
    .idy(64'd5),
    .fifo_A_in_s_dout(fifo_A_PE_2_5__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_2_5__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_2_5__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_2_5__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_2_5__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_2_6__din),
    .fifo_A_out_full_n(fifo_A_PE_2_6__full_n),
    .fifo_A_out_write(fifo_A_PE_2_6__write),
    .fifo_B_in_s_dout(fifo_B_PE_2_5__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_2_5__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_2_5__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_2_5__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_2_5__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_3_5__din),
    .fifo_B_out_full_n(fifo_B_PE_3_5__full_n),
    .fifo_B_out_write(fifo_B_PE_3_5__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_2_5__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_2_5__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_2_5__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_40
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_40__ap_start),
    .ap_done(PE_wrapper_40__ap_done),
    .ap_idle(PE_wrapper_40__ap_idle),
    .ap_ready(PE_wrapper_40__ap_ready),
    .idx(64'd2),
    .idy(64'd6),
    .fifo_A_in_s_dout(fifo_A_PE_2_6__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_2_6__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_2_6__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_2_6__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_2_6__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_2_7__din),
    .fifo_A_out_full_n(fifo_A_PE_2_7__full_n),
    .fifo_A_out_write(fifo_A_PE_2_7__write),
    .fifo_B_in_s_dout(fifo_B_PE_2_6__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_2_6__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_2_6__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_2_6__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_2_6__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_3_6__din),
    .fifo_B_out_full_n(fifo_B_PE_3_6__full_n),
    .fifo_B_out_write(fifo_B_PE_3_6__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_2_6__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_2_6__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_2_6__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_41
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_41__ap_start),
    .ap_done(PE_wrapper_41__ap_done),
    .ap_idle(PE_wrapper_41__ap_idle),
    .ap_ready(PE_wrapper_41__ap_ready),
    .idx(64'd2),
    .idy(64'd7),
    .fifo_A_in_s_dout(fifo_A_PE_2_7__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_2_7__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_2_7__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_2_7__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_2_7__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_2_8__din),
    .fifo_A_out_full_n(fifo_A_PE_2_8__full_n),
    .fifo_A_out_write(fifo_A_PE_2_8__write),
    .fifo_B_in_s_dout(fifo_B_PE_2_7__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_2_7__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_2_7__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_2_7__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_2_7__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_3_7__din),
    .fifo_B_out_full_n(fifo_B_PE_3_7__full_n),
    .fifo_B_out_write(fifo_B_PE_3_7__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_2_7__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_2_7__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_2_7__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_42
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_42__ap_start),
    .ap_done(PE_wrapper_42__ap_done),
    .ap_idle(PE_wrapper_42__ap_idle),
    .ap_ready(PE_wrapper_42__ap_ready),
    .idx(64'd2),
    .idy(64'd8),
    .fifo_A_in_s_dout(fifo_A_PE_2_8__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_2_8__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_2_8__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_2_8__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_2_8__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_2_9__din),
    .fifo_A_out_full_n(fifo_A_PE_2_9__full_n),
    .fifo_A_out_write(fifo_A_PE_2_9__write),
    .fifo_B_in_s_dout(fifo_B_PE_2_8__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_2_8__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_2_8__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_2_8__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_2_8__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_3_8__din),
    .fifo_B_out_full_n(fifo_B_PE_3_8__full_n),
    .fifo_B_out_write(fifo_B_PE_3_8__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_2_8__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_2_8__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_2_8__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_43
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_43__ap_start),
    .ap_done(PE_wrapper_43__ap_done),
    .ap_idle(PE_wrapper_43__ap_idle),
    .ap_ready(PE_wrapper_43__ap_ready),
    .idx(64'd2),
    .idy(64'd9),
    .fifo_A_out_din(fifo_A_PE_2_10__din),
    .fifo_A_out_full_n(fifo_A_PE_2_10__full_n),
    .fifo_A_out_write(fifo_A_PE_2_10__write),
    .fifo_A_in_s_dout(fifo_A_PE_2_9__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_2_9__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_2_9__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_2_9__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_2_9__read),
    .fifo_A_in_peek_read(),
    .fifo_B_in_s_dout(fifo_B_PE_2_9__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_2_9__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_2_9__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_2_9__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_2_9__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_3_9__din),
    .fifo_B_out_full_n(fifo_B_PE_3_9__full_n),
    .fifo_B_out_write(fifo_B_PE_3_9__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_2_9__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_2_9__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_2_9__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_44
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_44__ap_start),
    .ap_done(PE_wrapper_44__ap_done),
    .ap_idle(PE_wrapper_44__ap_idle),
    .ap_ready(PE_wrapper_44__ap_ready),
    .idy(64'd10),
    .idx(64'd2),
    .fifo_A_in_s_dout(fifo_A_PE_2_10__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_2_10__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_2_10__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_2_10__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_2_10__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_2_11__din),
    .fifo_A_out_full_n(fifo_A_PE_2_11__full_n),
    .fifo_A_out_write(fifo_A_PE_2_11__write),
    .fifo_B_in_s_dout(fifo_B_PE_2_10__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_2_10__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_2_10__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_2_10__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_2_10__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_3_10__din),
    .fifo_B_out_full_n(fifo_B_PE_3_10__full_n),
    .fifo_B_out_write(fifo_B_PE_3_10__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_2_10__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_2_10__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_2_10__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_45
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_45__ap_start),
    .ap_done(PE_wrapper_45__ap_done),
    .ap_idle(PE_wrapper_45__ap_idle),
    .ap_ready(PE_wrapper_45__ap_ready),
    .idy(64'd11),
    .idx(64'd2),
    .fifo_A_in_s_dout(fifo_A_PE_2_11__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_2_11__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_2_11__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_2_11__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_2_11__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_2_12__din),
    .fifo_A_out_full_n(fifo_A_PE_2_12__full_n),
    .fifo_A_out_write(fifo_A_PE_2_12__write),
    .fifo_B_in_s_dout(fifo_B_PE_2_11__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_2_11__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_2_11__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_2_11__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_2_11__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_3_11__din),
    .fifo_B_out_full_n(fifo_B_PE_3_11__full_n),
    .fifo_B_out_write(fifo_B_PE_3_11__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_2_11__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_2_11__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_2_11__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_46
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_46__ap_start),
    .ap_done(PE_wrapper_46__ap_done),
    .ap_idle(PE_wrapper_46__ap_idle),
    .ap_ready(PE_wrapper_46__ap_ready),
    .idy(64'd12),
    .idx(64'd2),
    .fifo_A_in_s_dout(fifo_A_PE_2_12__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_2_12__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_2_12__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_2_12__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_2_12__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_2_13__din),
    .fifo_A_out_full_n(fifo_A_PE_2_13__full_n),
    .fifo_A_out_write(fifo_A_PE_2_13__write),
    .fifo_B_in_s_dout(fifo_B_PE_2_12__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_2_12__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_2_12__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_2_12__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_2_12__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_3_12__din),
    .fifo_B_out_full_n(fifo_B_PE_3_12__full_n),
    .fifo_B_out_write(fifo_B_PE_3_12__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_2_12__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_2_12__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_2_12__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_47
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_47__ap_start),
    .ap_done(PE_wrapper_47__ap_done),
    .ap_idle(PE_wrapper_47__ap_idle),
    .ap_ready(PE_wrapper_47__ap_ready),
    .idy(64'd13),
    .idx(64'd2),
    .fifo_A_in_s_dout(fifo_A_PE_2_13__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_2_13__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_2_13__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_2_13__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_2_13__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_2_14__din),
    .fifo_A_out_full_n(fifo_A_PE_2_14__full_n),
    .fifo_A_out_write(fifo_A_PE_2_14__write),
    .fifo_B_in_s_dout(fifo_B_PE_2_13__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_2_13__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_2_13__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_2_13__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_2_13__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_3_13__din),
    .fifo_B_out_full_n(fifo_B_PE_3_13__full_n),
    .fifo_B_out_write(fifo_B_PE_3_13__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_2_13__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_2_13__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_2_13__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_48
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_48__ap_start),
    .ap_done(PE_wrapper_48__ap_done),
    .ap_idle(PE_wrapper_48__ap_idle),
    .ap_ready(PE_wrapper_48__ap_ready),
    .idy(64'd14),
    .idx(64'd2),
    .fifo_A_in_s_dout(fifo_A_PE_2_14__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_2_14__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_2_14__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_2_14__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_2_14__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_2_15__din),
    .fifo_A_out_full_n(fifo_A_PE_2_15__full_n),
    .fifo_A_out_write(fifo_A_PE_2_15__write),
    .fifo_B_in_s_dout(fifo_B_PE_2_14__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_2_14__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_2_14__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_2_14__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_2_14__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_3_14__din),
    .fifo_B_out_full_n(fifo_B_PE_3_14__full_n),
    .fifo_B_out_write(fifo_B_PE_3_14__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_2_14__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_2_14__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_2_14__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_49
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_49__ap_start),
    .ap_done(PE_wrapper_49__ap_done),
    .ap_idle(PE_wrapper_49__ap_idle),
    .ap_ready(PE_wrapper_49__ap_ready),
    .idy(64'd15),
    .idx(64'd2),
    .fifo_A_in_s_dout(fifo_A_PE_2_15__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_2_15__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_2_15__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_2_15__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_2_15__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_2_16__din),
    .fifo_A_out_full_n(fifo_A_PE_2_16__full_n),
    .fifo_A_out_write(fifo_A_PE_2_16__write),
    .fifo_B_in_s_dout(fifo_B_PE_2_15__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_2_15__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_2_15__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_2_15__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_2_15__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_3_15__din),
    .fifo_B_out_full_n(fifo_B_PE_3_15__full_n),
    .fifo_B_out_write(fifo_B_PE_3_15__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_2_15__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_2_15__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_2_15__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_50
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_50__ap_start),
    .ap_done(PE_wrapper_50__ap_done),
    .ap_idle(PE_wrapper_50__ap_idle),
    .ap_ready(PE_wrapper_50__ap_ready),
    .idy(64'd16),
    .idx(64'd2),
    .fifo_A_in_s_dout(fifo_A_PE_2_16__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_2_16__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_2_16__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_2_16__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_2_16__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_2_17__din),
    .fifo_A_out_full_n(fifo_A_PE_2_17__full_n),
    .fifo_A_out_write(fifo_A_PE_2_17__write),
    .fifo_B_in_s_dout(fifo_B_PE_2_16__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_2_16__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_2_16__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_2_16__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_2_16__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_3_16__din),
    .fifo_B_out_full_n(fifo_B_PE_3_16__full_n),
    .fifo_B_out_write(fifo_B_PE_3_16__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_2_16__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_2_16__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_2_16__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_51
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_51__ap_start),
    .ap_done(PE_wrapper_51__ap_done),
    .ap_idle(PE_wrapper_51__ap_idle),
    .ap_ready(PE_wrapper_51__ap_ready),
    .idy(64'd0),
    .idx(64'd3),
    .fifo_A_in_s_dout(fifo_A_PE_3_0__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_3_0__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_3_0__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_3_0__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_3_0__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_3_1__din),
    .fifo_A_out_full_n(fifo_A_PE_3_1__full_n),
    .fifo_A_out_write(fifo_A_PE_3_1__write),
    .fifo_B_in_s_dout(fifo_B_PE_3_0__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_3_0__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_3_0__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_3_0__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_3_0__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_4_0__din),
    .fifo_B_out_full_n(fifo_B_PE_4_0__full_n),
    .fifo_B_out_write(fifo_B_PE_4_0__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_3_0__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_3_0__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_3_0__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_52
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_52__ap_start),
    .ap_done(PE_wrapper_52__ap_done),
    .ap_idle(PE_wrapper_52__ap_idle),
    .ap_ready(PE_wrapper_52__ap_ready),
    .idy(64'd1),
    .idx(64'd3),
    .fifo_A_in_s_dout(fifo_A_PE_3_1__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_3_1__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_3_1__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_3_1__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_3_1__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_3_2__din),
    .fifo_A_out_full_n(fifo_A_PE_3_2__full_n),
    .fifo_A_out_write(fifo_A_PE_3_2__write),
    .fifo_B_in_s_dout(fifo_B_PE_3_1__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_3_1__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_3_1__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_3_1__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_3_1__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_4_1__din),
    .fifo_B_out_full_n(fifo_B_PE_4_1__full_n),
    .fifo_B_out_write(fifo_B_PE_4_1__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_3_1__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_3_1__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_3_1__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_53
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_53__ap_start),
    .ap_done(PE_wrapper_53__ap_done),
    .ap_idle(PE_wrapper_53__ap_idle),
    .ap_ready(PE_wrapper_53__ap_ready),
    .idy(64'd2),
    .idx(64'd3),
    .fifo_A_in_s_dout(fifo_A_PE_3_2__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_3_2__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_3_2__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_3_2__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_3_2__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_3_3__din),
    .fifo_A_out_full_n(fifo_A_PE_3_3__full_n),
    .fifo_A_out_write(fifo_A_PE_3_3__write),
    .fifo_B_in_s_dout(fifo_B_PE_3_2__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_3_2__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_3_2__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_3_2__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_3_2__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_4_2__din),
    .fifo_B_out_full_n(fifo_B_PE_4_2__full_n),
    .fifo_B_out_write(fifo_B_PE_4_2__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_3_2__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_3_2__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_3_2__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_54
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_54__ap_start),
    .ap_done(PE_wrapper_54__ap_done),
    .ap_idle(PE_wrapper_54__ap_idle),
    .ap_ready(PE_wrapper_54__ap_ready),
    .idx(64'd3),
    .idy(64'd3),
    .fifo_A_in_s_dout(fifo_A_PE_3_3__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_3_3__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_3_3__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_3_3__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_3_3__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_3_4__din),
    .fifo_A_out_full_n(fifo_A_PE_3_4__full_n),
    .fifo_A_out_write(fifo_A_PE_3_4__write),
    .fifo_B_in_s_dout(fifo_B_PE_3_3__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_3_3__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_3_3__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_3_3__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_3_3__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_4_3__din),
    .fifo_B_out_full_n(fifo_B_PE_4_3__full_n),
    .fifo_B_out_write(fifo_B_PE_4_3__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_3_3__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_3_3__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_3_3__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_55
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_55__ap_start),
    .ap_done(PE_wrapper_55__ap_done),
    .ap_idle(PE_wrapper_55__ap_idle),
    .ap_ready(PE_wrapper_55__ap_ready),
    .idx(64'd3),
    .idy(64'd4),
    .fifo_A_in_s_dout(fifo_A_PE_3_4__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_3_4__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_3_4__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_3_4__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_3_4__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_3_5__din),
    .fifo_A_out_full_n(fifo_A_PE_3_5__full_n),
    .fifo_A_out_write(fifo_A_PE_3_5__write),
    .fifo_B_in_s_dout(fifo_B_PE_3_4__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_3_4__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_3_4__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_3_4__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_3_4__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_4_4__din),
    .fifo_B_out_full_n(fifo_B_PE_4_4__full_n),
    .fifo_B_out_write(fifo_B_PE_4_4__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_3_4__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_3_4__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_3_4__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_56
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_56__ap_start),
    .ap_done(PE_wrapper_56__ap_done),
    .ap_idle(PE_wrapper_56__ap_idle),
    .ap_ready(PE_wrapper_56__ap_ready),
    .idx(64'd3),
    .idy(64'd5),
    .fifo_A_in_s_dout(fifo_A_PE_3_5__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_3_5__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_3_5__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_3_5__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_3_5__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_3_6__din),
    .fifo_A_out_full_n(fifo_A_PE_3_6__full_n),
    .fifo_A_out_write(fifo_A_PE_3_6__write),
    .fifo_B_in_s_dout(fifo_B_PE_3_5__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_3_5__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_3_5__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_3_5__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_3_5__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_4_5__din),
    .fifo_B_out_full_n(fifo_B_PE_4_5__full_n),
    .fifo_B_out_write(fifo_B_PE_4_5__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_3_5__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_3_5__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_3_5__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_57
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_57__ap_start),
    .ap_done(PE_wrapper_57__ap_done),
    .ap_idle(PE_wrapper_57__ap_idle),
    .ap_ready(PE_wrapper_57__ap_ready),
    .idx(64'd3),
    .idy(64'd6),
    .fifo_A_in_s_dout(fifo_A_PE_3_6__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_3_6__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_3_6__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_3_6__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_3_6__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_3_7__din),
    .fifo_A_out_full_n(fifo_A_PE_3_7__full_n),
    .fifo_A_out_write(fifo_A_PE_3_7__write),
    .fifo_B_in_s_dout(fifo_B_PE_3_6__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_3_6__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_3_6__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_3_6__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_3_6__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_4_6__din),
    .fifo_B_out_full_n(fifo_B_PE_4_6__full_n),
    .fifo_B_out_write(fifo_B_PE_4_6__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_3_6__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_3_6__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_3_6__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_58
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_58__ap_start),
    .ap_done(PE_wrapper_58__ap_done),
    .ap_idle(PE_wrapper_58__ap_idle),
    .ap_ready(PE_wrapper_58__ap_ready),
    .idx(64'd3),
    .idy(64'd7),
    .fifo_A_in_s_dout(fifo_A_PE_3_7__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_3_7__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_3_7__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_3_7__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_3_7__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_3_8__din),
    .fifo_A_out_full_n(fifo_A_PE_3_8__full_n),
    .fifo_A_out_write(fifo_A_PE_3_8__write),
    .fifo_B_in_s_dout(fifo_B_PE_3_7__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_3_7__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_3_7__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_3_7__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_3_7__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_4_7__din),
    .fifo_B_out_full_n(fifo_B_PE_4_7__full_n),
    .fifo_B_out_write(fifo_B_PE_4_7__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_3_7__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_3_7__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_3_7__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_59
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_59__ap_start),
    .ap_done(PE_wrapper_59__ap_done),
    .ap_idle(PE_wrapper_59__ap_idle),
    .ap_ready(PE_wrapper_59__ap_ready),
    .idx(64'd3),
    .idy(64'd8),
    .fifo_A_in_s_dout(fifo_A_PE_3_8__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_3_8__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_3_8__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_3_8__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_3_8__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_3_9__din),
    .fifo_A_out_full_n(fifo_A_PE_3_9__full_n),
    .fifo_A_out_write(fifo_A_PE_3_9__write),
    .fifo_B_in_s_dout(fifo_B_PE_3_8__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_3_8__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_3_8__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_3_8__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_3_8__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_4_8__din),
    .fifo_B_out_full_n(fifo_B_PE_4_8__full_n),
    .fifo_B_out_write(fifo_B_PE_4_8__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_3_8__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_3_8__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_3_8__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_60
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_60__ap_start),
    .ap_done(PE_wrapper_60__ap_done),
    .ap_idle(PE_wrapper_60__ap_idle),
    .ap_ready(PE_wrapper_60__ap_ready),
    .idx(64'd3),
    .idy(64'd9),
    .fifo_A_out_din(fifo_A_PE_3_10__din),
    .fifo_A_out_full_n(fifo_A_PE_3_10__full_n),
    .fifo_A_out_write(fifo_A_PE_3_10__write),
    .fifo_A_in_s_dout(fifo_A_PE_3_9__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_3_9__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_3_9__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_3_9__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_3_9__read),
    .fifo_A_in_peek_read(),
    .fifo_B_in_s_dout(fifo_B_PE_3_9__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_3_9__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_3_9__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_3_9__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_3_9__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_4_9__din),
    .fifo_B_out_full_n(fifo_B_PE_4_9__full_n),
    .fifo_B_out_write(fifo_B_PE_4_9__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_3_9__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_3_9__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_3_9__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_61
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_61__ap_start),
    .ap_done(PE_wrapper_61__ap_done),
    .ap_idle(PE_wrapper_61__ap_idle),
    .ap_ready(PE_wrapper_61__ap_ready),
    .idy(64'd10),
    .idx(64'd3),
    .fifo_A_in_s_dout(fifo_A_PE_3_10__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_3_10__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_3_10__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_3_10__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_3_10__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_3_11__din),
    .fifo_A_out_full_n(fifo_A_PE_3_11__full_n),
    .fifo_A_out_write(fifo_A_PE_3_11__write),
    .fifo_B_in_s_dout(fifo_B_PE_3_10__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_3_10__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_3_10__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_3_10__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_3_10__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_4_10__din),
    .fifo_B_out_full_n(fifo_B_PE_4_10__full_n),
    .fifo_B_out_write(fifo_B_PE_4_10__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_3_10__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_3_10__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_3_10__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_62
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_62__ap_start),
    .ap_done(PE_wrapper_62__ap_done),
    .ap_idle(PE_wrapper_62__ap_idle),
    .ap_ready(PE_wrapper_62__ap_ready),
    .idy(64'd11),
    .idx(64'd3),
    .fifo_A_in_s_dout(fifo_A_PE_3_11__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_3_11__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_3_11__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_3_11__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_3_11__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_3_12__din),
    .fifo_A_out_full_n(fifo_A_PE_3_12__full_n),
    .fifo_A_out_write(fifo_A_PE_3_12__write),
    .fifo_B_in_s_dout(fifo_B_PE_3_11__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_3_11__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_3_11__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_3_11__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_3_11__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_4_11__din),
    .fifo_B_out_full_n(fifo_B_PE_4_11__full_n),
    .fifo_B_out_write(fifo_B_PE_4_11__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_3_11__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_3_11__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_3_11__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_63
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_63__ap_start),
    .ap_done(PE_wrapper_63__ap_done),
    .ap_idle(PE_wrapper_63__ap_idle),
    .ap_ready(PE_wrapper_63__ap_ready),
    .idy(64'd12),
    .idx(64'd3),
    .fifo_A_in_s_dout(fifo_A_PE_3_12__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_3_12__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_3_12__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_3_12__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_3_12__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_3_13__din),
    .fifo_A_out_full_n(fifo_A_PE_3_13__full_n),
    .fifo_A_out_write(fifo_A_PE_3_13__write),
    .fifo_B_in_s_dout(fifo_B_PE_3_12__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_3_12__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_3_12__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_3_12__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_3_12__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_4_12__din),
    .fifo_B_out_full_n(fifo_B_PE_4_12__full_n),
    .fifo_B_out_write(fifo_B_PE_4_12__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_3_12__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_3_12__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_3_12__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_64
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_64__ap_start),
    .ap_done(PE_wrapper_64__ap_done),
    .ap_idle(PE_wrapper_64__ap_idle),
    .ap_ready(PE_wrapper_64__ap_ready),
    .idy(64'd13),
    .idx(64'd3),
    .fifo_A_in_s_dout(fifo_A_PE_3_13__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_3_13__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_3_13__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_3_13__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_3_13__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_3_14__din),
    .fifo_A_out_full_n(fifo_A_PE_3_14__full_n),
    .fifo_A_out_write(fifo_A_PE_3_14__write),
    .fifo_B_in_s_dout(fifo_B_PE_3_13__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_3_13__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_3_13__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_3_13__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_3_13__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_4_13__din),
    .fifo_B_out_full_n(fifo_B_PE_4_13__full_n),
    .fifo_B_out_write(fifo_B_PE_4_13__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_3_13__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_3_13__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_3_13__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_65
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_65__ap_start),
    .ap_done(PE_wrapper_65__ap_done),
    .ap_idle(PE_wrapper_65__ap_idle),
    .ap_ready(PE_wrapper_65__ap_ready),
    .idy(64'd14),
    .idx(64'd3),
    .fifo_A_in_s_dout(fifo_A_PE_3_14__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_3_14__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_3_14__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_3_14__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_3_14__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_3_15__din),
    .fifo_A_out_full_n(fifo_A_PE_3_15__full_n),
    .fifo_A_out_write(fifo_A_PE_3_15__write),
    .fifo_B_in_s_dout(fifo_B_PE_3_14__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_3_14__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_3_14__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_3_14__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_3_14__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_4_14__din),
    .fifo_B_out_full_n(fifo_B_PE_4_14__full_n),
    .fifo_B_out_write(fifo_B_PE_4_14__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_3_14__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_3_14__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_3_14__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_66
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_66__ap_start),
    .ap_done(PE_wrapper_66__ap_done),
    .ap_idle(PE_wrapper_66__ap_idle),
    .ap_ready(PE_wrapper_66__ap_ready),
    .idy(64'd15),
    .idx(64'd3),
    .fifo_A_in_s_dout(fifo_A_PE_3_15__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_3_15__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_3_15__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_3_15__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_3_15__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_3_16__din),
    .fifo_A_out_full_n(fifo_A_PE_3_16__full_n),
    .fifo_A_out_write(fifo_A_PE_3_16__write),
    .fifo_B_in_s_dout(fifo_B_PE_3_15__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_3_15__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_3_15__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_3_15__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_3_15__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_4_15__din),
    .fifo_B_out_full_n(fifo_B_PE_4_15__full_n),
    .fifo_B_out_write(fifo_B_PE_4_15__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_3_15__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_3_15__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_3_15__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_67
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_67__ap_start),
    .ap_done(PE_wrapper_67__ap_done),
    .ap_idle(PE_wrapper_67__ap_idle),
    .ap_ready(PE_wrapper_67__ap_ready),
    .idy(64'd16),
    .idx(64'd3),
    .fifo_A_in_s_dout(fifo_A_PE_3_16__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_3_16__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_3_16__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_3_16__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_3_16__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_3_17__din),
    .fifo_A_out_full_n(fifo_A_PE_3_17__full_n),
    .fifo_A_out_write(fifo_A_PE_3_17__write),
    .fifo_B_in_s_dout(fifo_B_PE_3_16__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_3_16__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_3_16__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_3_16__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_3_16__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_4_16__din),
    .fifo_B_out_full_n(fifo_B_PE_4_16__full_n),
    .fifo_B_out_write(fifo_B_PE_4_16__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_3_16__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_3_16__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_3_16__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_68
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_68__ap_start),
    .ap_done(PE_wrapper_68__ap_done),
    .ap_idle(PE_wrapper_68__ap_idle),
    .ap_ready(PE_wrapper_68__ap_ready),
    .idy(64'd0),
    .idx(64'd4),
    .fifo_A_in_s_dout(fifo_A_PE_4_0__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_4_0__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_4_0__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_4_0__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_4_0__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_4_1__din),
    .fifo_A_out_full_n(fifo_A_PE_4_1__full_n),
    .fifo_A_out_write(fifo_A_PE_4_1__write),
    .fifo_B_in_s_dout(fifo_B_PE_4_0__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_4_0__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_4_0__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_4_0__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_4_0__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_5_0__din),
    .fifo_B_out_full_n(fifo_B_PE_5_0__full_n),
    .fifo_B_out_write(fifo_B_PE_5_0__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_4_0__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_4_0__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_4_0__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_69
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_69__ap_start),
    .ap_done(PE_wrapper_69__ap_done),
    .ap_idle(PE_wrapper_69__ap_idle),
    .ap_ready(PE_wrapper_69__ap_ready),
    .idy(64'd1),
    .idx(64'd4),
    .fifo_A_in_s_dout(fifo_A_PE_4_1__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_4_1__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_4_1__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_4_1__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_4_1__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_4_2__din),
    .fifo_A_out_full_n(fifo_A_PE_4_2__full_n),
    .fifo_A_out_write(fifo_A_PE_4_2__write),
    .fifo_B_in_s_dout(fifo_B_PE_4_1__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_4_1__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_4_1__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_4_1__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_4_1__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_5_1__din),
    .fifo_B_out_full_n(fifo_B_PE_5_1__full_n),
    .fifo_B_out_write(fifo_B_PE_5_1__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_4_1__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_4_1__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_4_1__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_70
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_70__ap_start),
    .ap_done(PE_wrapper_70__ap_done),
    .ap_idle(PE_wrapper_70__ap_idle),
    .ap_ready(PE_wrapper_70__ap_ready),
    .idy(64'd2),
    .idx(64'd4),
    .fifo_A_in_s_dout(fifo_A_PE_4_2__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_4_2__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_4_2__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_4_2__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_4_2__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_4_3__din),
    .fifo_A_out_full_n(fifo_A_PE_4_3__full_n),
    .fifo_A_out_write(fifo_A_PE_4_3__write),
    .fifo_B_in_s_dout(fifo_B_PE_4_2__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_4_2__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_4_2__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_4_2__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_4_2__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_5_2__din),
    .fifo_B_out_full_n(fifo_B_PE_5_2__full_n),
    .fifo_B_out_write(fifo_B_PE_5_2__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_4_2__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_4_2__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_4_2__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_71
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_71__ap_start),
    .ap_done(PE_wrapper_71__ap_done),
    .ap_idle(PE_wrapper_71__ap_idle),
    .ap_ready(PE_wrapper_71__ap_ready),
    .idy(64'd3),
    .idx(64'd4),
    .fifo_A_in_s_dout(fifo_A_PE_4_3__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_4_3__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_4_3__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_4_3__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_4_3__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_4_4__din),
    .fifo_A_out_full_n(fifo_A_PE_4_4__full_n),
    .fifo_A_out_write(fifo_A_PE_4_4__write),
    .fifo_B_in_s_dout(fifo_B_PE_4_3__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_4_3__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_4_3__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_4_3__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_4_3__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_5_3__din),
    .fifo_B_out_full_n(fifo_B_PE_5_3__full_n),
    .fifo_B_out_write(fifo_B_PE_5_3__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_4_3__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_4_3__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_4_3__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_72
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_72__ap_start),
    .ap_done(PE_wrapper_72__ap_done),
    .ap_idle(PE_wrapper_72__ap_idle),
    .ap_ready(PE_wrapper_72__ap_ready),
    .idx(64'd4),
    .idy(64'd4),
    .fifo_A_in_s_dout(fifo_A_PE_4_4__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_4_4__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_4_4__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_4_4__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_4_4__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_4_5__din),
    .fifo_A_out_full_n(fifo_A_PE_4_5__full_n),
    .fifo_A_out_write(fifo_A_PE_4_5__write),
    .fifo_B_in_s_dout(fifo_B_PE_4_4__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_4_4__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_4_4__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_4_4__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_4_4__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_5_4__din),
    .fifo_B_out_full_n(fifo_B_PE_5_4__full_n),
    .fifo_B_out_write(fifo_B_PE_5_4__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_4_4__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_4_4__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_4_4__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_73
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_73__ap_start),
    .ap_done(PE_wrapper_73__ap_done),
    .ap_idle(PE_wrapper_73__ap_idle),
    .ap_ready(PE_wrapper_73__ap_ready),
    .idx(64'd4),
    .idy(64'd5),
    .fifo_A_in_s_dout(fifo_A_PE_4_5__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_4_5__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_4_5__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_4_5__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_4_5__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_4_6__din),
    .fifo_A_out_full_n(fifo_A_PE_4_6__full_n),
    .fifo_A_out_write(fifo_A_PE_4_6__write),
    .fifo_B_in_s_dout(fifo_B_PE_4_5__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_4_5__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_4_5__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_4_5__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_4_5__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_5_5__din),
    .fifo_B_out_full_n(fifo_B_PE_5_5__full_n),
    .fifo_B_out_write(fifo_B_PE_5_5__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_4_5__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_4_5__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_4_5__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_74
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_74__ap_start),
    .ap_done(PE_wrapper_74__ap_done),
    .ap_idle(PE_wrapper_74__ap_idle),
    .ap_ready(PE_wrapper_74__ap_ready),
    .idx(64'd4),
    .idy(64'd6),
    .fifo_A_in_s_dout(fifo_A_PE_4_6__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_4_6__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_4_6__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_4_6__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_4_6__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_4_7__din),
    .fifo_A_out_full_n(fifo_A_PE_4_7__full_n),
    .fifo_A_out_write(fifo_A_PE_4_7__write),
    .fifo_B_in_s_dout(fifo_B_PE_4_6__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_4_6__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_4_6__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_4_6__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_4_6__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_5_6__din),
    .fifo_B_out_full_n(fifo_B_PE_5_6__full_n),
    .fifo_B_out_write(fifo_B_PE_5_6__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_4_6__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_4_6__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_4_6__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_75
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_75__ap_start),
    .ap_done(PE_wrapper_75__ap_done),
    .ap_idle(PE_wrapper_75__ap_idle),
    .ap_ready(PE_wrapper_75__ap_ready),
    .idx(64'd4),
    .idy(64'd7),
    .fifo_A_in_s_dout(fifo_A_PE_4_7__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_4_7__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_4_7__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_4_7__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_4_7__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_4_8__din),
    .fifo_A_out_full_n(fifo_A_PE_4_8__full_n),
    .fifo_A_out_write(fifo_A_PE_4_8__write),
    .fifo_B_in_s_dout(fifo_B_PE_4_7__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_4_7__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_4_7__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_4_7__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_4_7__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_5_7__din),
    .fifo_B_out_full_n(fifo_B_PE_5_7__full_n),
    .fifo_B_out_write(fifo_B_PE_5_7__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_4_7__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_4_7__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_4_7__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_76
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_76__ap_start),
    .ap_done(PE_wrapper_76__ap_done),
    .ap_idle(PE_wrapper_76__ap_idle),
    .ap_ready(PE_wrapper_76__ap_ready),
    .idx(64'd4),
    .idy(64'd8),
    .fifo_A_in_s_dout(fifo_A_PE_4_8__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_4_8__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_4_8__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_4_8__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_4_8__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_4_9__din),
    .fifo_A_out_full_n(fifo_A_PE_4_9__full_n),
    .fifo_A_out_write(fifo_A_PE_4_9__write),
    .fifo_B_in_s_dout(fifo_B_PE_4_8__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_4_8__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_4_8__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_4_8__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_4_8__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_5_8__din),
    .fifo_B_out_full_n(fifo_B_PE_5_8__full_n),
    .fifo_B_out_write(fifo_B_PE_5_8__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_4_8__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_4_8__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_4_8__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_77
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_77__ap_start),
    .ap_done(PE_wrapper_77__ap_done),
    .ap_idle(PE_wrapper_77__ap_idle),
    .ap_ready(PE_wrapper_77__ap_ready),
    .idx(64'd4),
    .idy(64'd9),
    .fifo_A_out_din(fifo_A_PE_4_10__din),
    .fifo_A_out_full_n(fifo_A_PE_4_10__full_n),
    .fifo_A_out_write(fifo_A_PE_4_10__write),
    .fifo_A_in_s_dout(fifo_A_PE_4_9__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_4_9__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_4_9__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_4_9__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_4_9__read),
    .fifo_A_in_peek_read(),
    .fifo_B_in_s_dout(fifo_B_PE_4_9__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_4_9__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_4_9__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_4_9__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_4_9__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_5_9__din),
    .fifo_B_out_full_n(fifo_B_PE_5_9__full_n),
    .fifo_B_out_write(fifo_B_PE_5_9__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_4_9__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_4_9__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_4_9__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_78
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_78__ap_start),
    .ap_done(PE_wrapper_78__ap_done),
    .ap_idle(PE_wrapper_78__ap_idle),
    .ap_ready(PE_wrapper_78__ap_ready),
    .idy(64'd10),
    .idx(64'd4),
    .fifo_A_in_s_dout(fifo_A_PE_4_10__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_4_10__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_4_10__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_4_10__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_4_10__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_4_11__din),
    .fifo_A_out_full_n(fifo_A_PE_4_11__full_n),
    .fifo_A_out_write(fifo_A_PE_4_11__write),
    .fifo_B_in_s_dout(fifo_B_PE_4_10__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_4_10__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_4_10__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_4_10__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_4_10__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_5_10__din),
    .fifo_B_out_full_n(fifo_B_PE_5_10__full_n),
    .fifo_B_out_write(fifo_B_PE_5_10__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_4_10__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_4_10__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_4_10__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_79
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_79__ap_start),
    .ap_done(PE_wrapper_79__ap_done),
    .ap_idle(PE_wrapper_79__ap_idle),
    .ap_ready(PE_wrapper_79__ap_ready),
    .idy(64'd11),
    .idx(64'd4),
    .fifo_A_in_s_dout(fifo_A_PE_4_11__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_4_11__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_4_11__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_4_11__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_4_11__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_4_12__din),
    .fifo_A_out_full_n(fifo_A_PE_4_12__full_n),
    .fifo_A_out_write(fifo_A_PE_4_12__write),
    .fifo_B_in_s_dout(fifo_B_PE_4_11__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_4_11__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_4_11__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_4_11__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_4_11__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_5_11__din),
    .fifo_B_out_full_n(fifo_B_PE_5_11__full_n),
    .fifo_B_out_write(fifo_B_PE_5_11__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_4_11__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_4_11__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_4_11__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_80
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_80__ap_start),
    .ap_done(PE_wrapper_80__ap_done),
    .ap_idle(PE_wrapper_80__ap_idle),
    .ap_ready(PE_wrapper_80__ap_ready),
    .idy(64'd12),
    .idx(64'd4),
    .fifo_A_in_s_dout(fifo_A_PE_4_12__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_4_12__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_4_12__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_4_12__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_4_12__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_4_13__din),
    .fifo_A_out_full_n(fifo_A_PE_4_13__full_n),
    .fifo_A_out_write(fifo_A_PE_4_13__write),
    .fifo_B_in_s_dout(fifo_B_PE_4_12__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_4_12__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_4_12__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_4_12__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_4_12__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_5_12__din),
    .fifo_B_out_full_n(fifo_B_PE_5_12__full_n),
    .fifo_B_out_write(fifo_B_PE_5_12__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_4_12__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_4_12__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_4_12__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_81
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_81__ap_start),
    .ap_done(PE_wrapper_81__ap_done),
    .ap_idle(PE_wrapper_81__ap_idle),
    .ap_ready(PE_wrapper_81__ap_ready),
    .idy(64'd13),
    .idx(64'd4),
    .fifo_A_in_s_dout(fifo_A_PE_4_13__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_4_13__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_4_13__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_4_13__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_4_13__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_4_14__din),
    .fifo_A_out_full_n(fifo_A_PE_4_14__full_n),
    .fifo_A_out_write(fifo_A_PE_4_14__write),
    .fifo_B_in_s_dout(fifo_B_PE_4_13__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_4_13__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_4_13__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_4_13__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_4_13__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_5_13__din),
    .fifo_B_out_full_n(fifo_B_PE_5_13__full_n),
    .fifo_B_out_write(fifo_B_PE_5_13__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_4_13__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_4_13__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_4_13__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_82
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_82__ap_start),
    .ap_done(PE_wrapper_82__ap_done),
    .ap_idle(PE_wrapper_82__ap_idle),
    .ap_ready(PE_wrapper_82__ap_ready),
    .idy(64'd14),
    .idx(64'd4),
    .fifo_A_in_s_dout(fifo_A_PE_4_14__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_4_14__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_4_14__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_4_14__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_4_14__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_4_15__din),
    .fifo_A_out_full_n(fifo_A_PE_4_15__full_n),
    .fifo_A_out_write(fifo_A_PE_4_15__write),
    .fifo_B_in_s_dout(fifo_B_PE_4_14__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_4_14__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_4_14__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_4_14__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_4_14__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_5_14__din),
    .fifo_B_out_full_n(fifo_B_PE_5_14__full_n),
    .fifo_B_out_write(fifo_B_PE_5_14__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_4_14__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_4_14__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_4_14__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_83
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_83__ap_start),
    .ap_done(PE_wrapper_83__ap_done),
    .ap_idle(PE_wrapper_83__ap_idle),
    .ap_ready(PE_wrapper_83__ap_ready),
    .idy(64'd15),
    .idx(64'd4),
    .fifo_A_in_s_dout(fifo_A_PE_4_15__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_4_15__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_4_15__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_4_15__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_4_15__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_4_16__din),
    .fifo_A_out_full_n(fifo_A_PE_4_16__full_n),
    .fifo_A_out_write(fifo_A_PE_4_16__write),
    .fifo_B_in_s_dout(fifo_B_PE_4_15__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_4_15__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_4_15__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_4_15__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_4_15__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_5_15__din),
    .fifo_B_out_full_n(fifo_B_PE_5_15__full_n),
    .fifo_B_out_write(fifo_B_PE_5_15__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_4_15__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_4_15__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_4_15__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_84
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_84__ap_start),
    .ap_done(PE_wrapper_84__ap_done),
    .ap_idle(PE_wrapper_84__ap_idle),
    .ap_ready(PE_wrapper_84__ap_ready),
    .idy(64'd16),
    .idx(64'd4),
    .fifo_A_in_s_dout(fifo_A_PE_4_16__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_4_16__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_4_16__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_4_16__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_4_16__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_4_17__din),
    .fifo_A_out_full_n(fifo_A_PE_4_17__full_n),
    .fifo_A_out_write(fifo_A_PE_4_17__write),
    .fifo_B_in_s_dout(fifo_B_PE_4_16__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_4_16__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_4_16__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_4_16__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_4_16__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_5_16__din),
    .fifo_B_out_full_n(fifo_B_PE_5_16__full_n),
    .fifo_B_out_write(fifo_B_PE_5_16__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_4_16__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_4_16__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_4_16__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_85
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_85__ap_start),
    .ap_done(PE_wrapper_85__ap_done),
    .ap_idle(PE_wrapper_85__ap_idle),
    .ap_ready(PE_wrapper_85__ap_ready),
    .idy(64'd0),
    .idx(64'd5),
    .fifo_A_in_s_dout(fifo_A_PE_5_0__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_5_0__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_5_0__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_5_0__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_5_0__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_5_1__din),
    .fifo_A_out_full_n(fifo_A_PE_5_1__full_n),
    .fifo_A_out_write(fifo_A_PE_5_1__write),
    .fifo_B_in_s_dout(fifo_B_PE_5_0__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_5_0__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_5_0__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_5_0__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_5_0__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_6_0__din),
    .fifo_B_out_full_n(fifo_B_PE_6_0__full_n),
    .fifo_B_out_write(fifo_B_PE_6_0__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_5_0__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_5_0__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_5_0__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_86
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_86__ap_start),
    .ap_done(PE_wrapper_86__ap_done),
    .ap_idle(PE_wrapper_86__ap_idle),
    .ap_ready(PE_wrapper_86__ap_ready),
    .idy(64'd1),
    .idx(64'd5),
    .fifo_A_in_s_dout(fifo_A_PE_5_1__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_5_1__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_5_1__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_5_1__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_5_1__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_5_2__din),
    .fifo_A_out_full_n(fifo_A_PE_5_2__full_n),
    .fifo_A_out_write(fifo_A_PE_5_2__write),
    .fifo_B_in_s_dout(fifo_B_PE_5_1__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_5_1__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_5_1__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_5_1__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_5_1__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_6_1__din),
    .fifo_B_out_full_n(fifo_B_PE_6_1__full_n),
    .fifo_B_out_write(fifo_B_PE_6_1__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_5_1__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_5_1__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_5_1__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_87
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_87__ap_start),
    .ap_done(PE_wrapper_87__ap_done),
    .ap_idle(PE_wrapper_87__ap_idle),
    .ap_ready(PE_wrapper_87__ap_ready),
    .idy(64'd2),
    .idx(64'd5),
    .fifo_A_in_s_dout(fifo_A_PE_5_2__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_5_2__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_5_2__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_5_2__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_5_2__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_5_3__din),
    .fifo_A_out_full_n(fifo_A_PE_5_3__full_n),
    .fifo_A_out_write(fifo_A_PE_5_3__write),
    .fifo_B_in_s_dout(fifo_B_PE_5_2__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_5_2__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_5_2__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_5_2__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_5_2__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_6_2__din),
    .fifo_B_out_full_n(fifo_B_PE_6_2__full_n),
    .fifo_B_out_write(fifo_B_PE_6_2__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_5_2__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_5_2__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_5_2__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_88
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_88__ap_start),
    .ap_done(PE_wrapper_88__ap_done),
    .ap_idle(PE_wrapper_88__ap_idle),
    .ap_ready(PE_wrapper_88__ap_ready),
    .idy(64'd3),
    .idx(64'd5),
    .fifo_A_in_s_dout(fifo_A_PE_5_3__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_5_3__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_5_3__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_5_3__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_5_3__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_5_4__din),
    .fifo_A_out_full_n(fifo_A_PE_5_4__full_n),
    .fifo_A_out_write(fifo_A_PE_5_4__write),
    .fifo_B_in_s_dout(fifo_B_PE_5_3__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_5_3__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_5_3__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_5_3__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_5_3__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_6_3__din),
    .fifo_B_out_full_n(fifo_B_PE_6_3__full_n),
    .fifo_B_out_write(fifo_B_PE_6_3__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_5_3__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_5_3__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_5_3__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_89
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_89__ap_start),
    .ap_done(PE_wrapper_89__ap_done),
    .ap_idle(PE_wrapper_89__ap_idle),
    .ap_ready(PE_wrapper_89__ap_ready),
    .idy(64'd4),
    .idx(64'd5),
    .fifo_A_in_s_dout(fifo_A_PE_5_4__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_5_4__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_5_4__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_5_4__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_5_4__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_5_5__din),
    .fifo_A_out_full_n(fifo_A_PE_5_5__full_n),
    .fifo_A_out_write(fifo_A_PE_5_5__write),
    .fifo_B_in_s_dout(fifo_B_PE_5_4__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_5_4__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_5_4__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_5_4__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_5_4__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_6_4__din),
    .fifo_B_out_full_n(fifo_B_PE_6_4__full_n),
    .fifo_B_out_write(fifo_B_PE_6_4__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_5_4__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_5_4__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_5_4__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_90
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_90__ap_start),
    .ap_done(PE_wrapper_90__ap_done),
    .ap_idle(PE_wrapper_90__ap_idle),
    .ap_ready(PE_wrapper_90__ap_ready),
    .idx(64'd5),
    .idy(64'd5),
    .fifo_A_in_s_dout(fifo_A_PE_5_5__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_5_5__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_5_5__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_5_5__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_5_5__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_5_6__din),
    .fifo_A_out_full_n(fifo_A_PE_5_6__full_n),
    .fifo_A_out_write(fifo_A_PE_5_6__write),
    .fifo_B_in_s_dout(fifo_B_PE_5_5__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_5_5__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_5_5__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_5_5__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_5_5__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_6_5__din),
    .fifo_B_out_full_n(fifo_B_PE_6_5__full_n),
    .fifo_B_out_write(fifo_B_PE_6_5__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_5_5__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_5_5__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_5_5__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_91
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_91__ap_start),
    .ap_done(PE_wrapper_91__ap_done),
    .ap_idle(PE_wrapper_91__ap_idle),
    .ap_ready(PE_wrapper_91__ap_ready),
    .idx(64'd5),
    .idy(64'd6),
    .fifo_A_in_s_dout(fifo_A_PE_5_6__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_5_6__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_5_6__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_5_6__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_5_6__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_5_7__din),
    .fifo_A_out_full_n(fifo_A_PE_5_7__full_n),
    .fifo_A_out_write(fifo_A_PE_5_7__write),
    .fifo_B_in_s_dout(fifo_B_PE_5_6__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_5_6__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_5_6__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_5_6__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_5_6__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_6_6__din),
    .fifo_B_out_full_n(fifo_B_PE_6_6__full_n),
    .fifo_B_out_write(fifo_B_PE_6_6__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_5_6__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_5_6__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_5_6__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_92
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_92__ap_start),
    .ap_done(PE_wrapper_92__ap_done),
    .ap_idle(PE_wrapper_92__ap_idle),
    .ap_ready(PE_wrapper_92__ap_ready),
    .idx(64'd5),
    .idy(64'd7),
    .fifo_A_in_s_dout(fifo_A_PE_5_7__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_5_7__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_5_7__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_5_7__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_5_7__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_5_8__din),
    .fifo_A_out_full_n(fifo_A_PE_5_8__full_n),
    .fifo_A_out_write(fifo_A_PE_5_8__write),
    .fifo_B_in_s_dout(fifo_B_PE_5_7__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_5_7__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_5_7__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_5_7__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_5_7__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_6_7__din),
    .fifo_B_out_full_n(fifo_B_PE_6_7__full_n),
    .fifo_B_out_write(fifo_B_PE_6_7__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_5_7__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_5_7__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_5_7__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_93
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_93__ap_start),
    .ap_done(PE_wrapper_93__ap_done),
    .ap_idle(PE_wrapper_93__ap_idle),
    .ap_ready(PE_wrapper_93__ap_ready),
    .idx(64'd5),
    .idy(64'd8),
    .fifo_A_in_s_dout(fifo_A_PE_5_8__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_5_8__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_5_8__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_5_8__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_5_8__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_5_9__din),
    .fifo_A_out_full_n(fifo_A_PE_5_9__full_n),
    .fifo_A_out_write(fifo_A_PE_5_9__write),
    .fifo_B_in_s_dout(fifo_B_PE_5_8__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_5_8__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_5_8__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_5_8__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_5_8__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_6_8__din),
    .fifo_B_out_full_n(fifo_B_PE_6_8__full_n),
    .fifo_B_out_write(fifo_B_PE_6_8__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_5_8__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_5_8__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_5_8__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_94
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_94__ap_start),
    .ap_done(PE_wrapper_94__ap_done),
    .ap_idle(PE_wrapper_94__ap_idle),
    .ap_ready(PE_wrapper_94__ap_ready),
    .idx(64'd5),
    .idy(64'd9),
    .fifo_A_out_din(fifo_A_PE_5_10__din),
    .fifo_A_out_full_n(fifo_A_PE_5_10__full_n),
    .fifo_A_out_write(fifo_A_PE_5_10__write),
    .fifo_A_in_s_dout(fifo_A_PE_5_9__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_5_9__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_5_9__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_5_9__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_5_9__read),
    .fifo_A_in_peek_read(),
    .fifo_B_in_s_dout(fifo_B_PE_5_9__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_5_9__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_5_9__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_5_9__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_5_9__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_6_9__din),
    .fifo_B_out_full_n(fifo_B_PE_6_9__full_n),
    .fifo_B_out_write(fifo_B_PE_6_9__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_5_9__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_5_9__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_5_9__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_95
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_95__ap_start),
    .ap_done(PE_wrapper_95__ap_done),
    .ap_idle(PE_wrapper_95__ap_idle),
    .ap_ready(PE_wrapper_95__ap_ready),
    .idy(64'd10),
    .idx(64'd5),
    .fifo_A_in_s_dout(fifo_A_PE_5_10__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_5_10__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_5_10__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_5_10__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_5_10__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_5_11__din),
    .fifo_A_out_full_n(fifo_A_PE_5_11__full_n),
    .fifo_A_out_write(fifo_A_PE_5_11__write),
    .fifo_B_in_s_dout(fifo_B_PE_5_10__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_5_10__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_5_10__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_5_10__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_5_10__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_6_10__din),
    .fifo_B_out_full_n(fifo_B_PE_6_10__full_n),
    .fifo_B_out_write(fifo_B_PE_6_10__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_5_10__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_5_10__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_5_10__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_96
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_96__ap_start),
    .ap_done(PE_wrapper_96__ap_done),
    .ap_idle(PE_wrapper_96__ap_idle),
    .ap_ready(PE_wrapper_96__ap_ready),
    .idy(64'd11),
    .idx(64'd5),
    .fifo_A_in_s_dout(fifo_A_PE_5_11__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_5_11__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_5_11__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_5_11__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_5_11__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_5_12__din),
    .fifo_A_out_full_n(fifo_A_PE_5_12__full_n),
    .fifo_A_out_write(fifo_A_PE_5_12__write),
    .fifo_B_in_s_dout(fifo_B_PE_5_11__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_5_11__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_5_11__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_5_11__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_5_11__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_6_11__din),
    .fifo_B_out_full_n(fifo_B_PE_6_11__full_n),
    .fifo_B_out_write(fifo_B_PE_6_11__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_5_11__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_5_11__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_5_11__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_97
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_97__ap_start),
    .ap_done(PE_wrapper_97__ap_done),
    .ap_idle(PE_wrapper_97__ap_idle),
    .ap_ready(PE_wrapper_97__ap_ready),
    .idy(64'd12),
    .idx(64'd5),
    .fifo_A_in_s_dout(fifo_A_PE_5_12__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_5_12__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_5_12__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_5_12__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_5_12__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_5_13__din),
    .fifo_A_out_full_n(fifo_A_PE_5_13__full_n),
    .fifo_A_out_write(fifo_A_PE_5_13__write),
    .fifo_B_in_s_dout(fifo_B_PE_5_12__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_5_12__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_5_12__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_5_12__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_5_12__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_6_12__din),
    .fifo_B_out_full_n(fifo_B_PE_6_12__full_n),
    .fifo_B_out_write(fifo_B_PE_6_12__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_5_12__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_5_12__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_5_12__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_98
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_98__ap_start),
    .ap_done(PE_wrapper_98__ap_done),
    .ap_idle(PE_wrapper_98__ap_idle),
    .ap_ready(PE_wrapper_98__ap_ready),
    .idy(64'd13),
    .idx(64'd5),
    .fifo_A_in_s_dout(fifo_A_PE_5_13__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_5_13__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_5_13__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_5_13__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_5_13__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_5_14__din),
    .fifo_A_out_full_n(fifo_A_PE_5_14__full_n),
    .fifo_A_out_write(fifo_A_PE_5_14__write),
    .fifo_B_in_s_dout(fifo_B_PE_5_13__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_5_13__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_5_13__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_5_13__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_5_13__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_6_13__din),
    .fifo_B_out_full_n(fifo_B_PE_6_13__full_n),
    .fifo_B_out_write(fifo_B_PE_6_13__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_5_13__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_5_13__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_5_13__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_99
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_99__ap_start),
    .ap_done(PE_wrapper_99__ap_done),
    .ap_idle(PE_wrapper_99__ap_idle),
    .ap_ready(PE_wrapper_99__ap_ready),
    .idy(64'd14),
    .idx(64'd5),
    .fifo_A_in_s_dout(fifo_A_PE_5_14__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_5_14__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_5_14__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_5_14__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_5_14__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_5_15__din),
    .fifo_A_out_full_n(fifo_A_PE_5_15__full_n),
    .fifo_A_out_write(fifo_A_PE_5_15__write),
    .fifo_B_in_s_dout(fifo_B_PE_5_14__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_5_14__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_5_14__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_5_14__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_5_14__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_6_14__din),
    .fifo_B_out_full_n(fifo_B_PE_6_14__full_n),
    .fifo_B_out_write(fifo_B_PE_6_14__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_5_14__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_5_14__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_5_14__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_100
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_100__ap_start),
    .ap_done(PE_wrapper_100__ap_done),
    .ap_idle(PE_wrapper_100__ap_idle),
    .ap_ready(PE_wrapper_100__ap_ready),
    .idy(64'd15),
    .idx(64'd5),
    .fifo_A_in_s_dout(fifo_A_PE_5_15__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_5_15__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_5_15__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_5_15__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_5_15__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_5_16__din),
    .fifo_A_out_full_n(fifo_A_PE_5_16__full_n),
    .fifo_A_out_write(fifo_A_PE_5_16__write),
    .fifo_B_in_s_dout(fifo_B_PE_5_15__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_5_15__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_5_15__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_5_15__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_5_15__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_6_15__din),
    .fifo_B_out_full_n(fifo_B_PE_6_15__full_n),
    .fifo_B_out_write(fifo_B_PE_6_15__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_5_15__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_5_15__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_5_15__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_101
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_101__ap_start),
    .ap_done(PE_wrapper_101__ap_done),
    .ap_idle(PE_wrapper_101__ap_idle),
    .ap_ready(PE_wrapper_101__ap_ready),
    .idy(64'd16),
    .idx(64'd5),
    .fifo_A_in_s_dout(fifo_A_PE_5_16__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_5_16__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_5_16__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_5_16__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_5_16__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_5_17__din),
    .fifo_A_out_full_n(fifo_A_PE_5_17__full_n),
    .fifo_A_out_write(fifo_A_PE_5_17__write),
    .fifo_B_in_s_dout(fifo_B_PE_5_16__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_5_16__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_5_16__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_5_16__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_5_16__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_6_16__din),
    .fifo_B_out_full_n(fifo_B_PE_6_16__full_n),
    .fifo_B_out_write(fifo_B_PE_6_16__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_5_16__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_5_16__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_5_16__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_102
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_102__ap_start),
    .ap_done(PE_wrapper_102__ap_done),
    .ap_idle(PE_wrapper_102__ap_idle),
    .ap_ready(PE_wrapper_102__ap_ready),
    .idy(64'd0),
    .idx(64'd6),
    .fifo_A_in_s_dout(fifo_A_PE_6_0__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_6_0__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_6_0__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_6_0__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_6_0__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_6_1__din),
    .fifo_A_out_full_n(fifo_A_PE_6_1__full_n),
    .fifo_A_out_write(fifo_A_PE_6_1__write),
    .fifo_B_in_s_dout(fifo_B_PE_6_0__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_6_0__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_6_0__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_6_0__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_6_0__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_7_0__din),
    .fifo_B_out_full_n(fifo_B_PE_7_0__full_n),
    .fifo_B_out_write(fifo_B_PE_7_0__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_6_0__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_6_0__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_6_0__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_103
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_103__ap_start),
    .ap_done(PE_wrapper_103__ap_done),
    .ap_idle(PE_wrapper_103__ap_idle),
    .ap_ready(PE_wrapper_103__ap_ready),
    .idy(64'd1),
    .idx(64'd6),
    .fifo_A_in_s_dout(fifo_A_PE_6_1__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_6_1__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_6_1__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_6_1__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_6_1__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_6_2__din),
    .fifo_A_out_full_n(fifo_A_PE_6_2__full_n),
    .fifo_A_out_write(fifo_A_PE_6_2__write),
    .fifo_B_in_s_dout(fifo_B_PE_6_1__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_6_1__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_6_1__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_6_1__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_6_1__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_7_1__din),
    .fifo_B_out_full_n(fifo_B_PE_7_1__full_n),
    .fifo_B_out_write(fifo_B_PE_7_1__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_6_1__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_6_1__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_6_1__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_104
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_104__ap_start),
    .ap_done(PE_wrapper_104__ap_done),
    .ap_idle(PE_wrapper_104__ap_idle),
    .ap_ready(PE_wrapper_104__ap_ready),
    .idy(64'd2),
    .idx(64'd6),
    .fifo_A_in_s_dout(fifo_A_PE_6_2__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_6_2__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_6_2__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_6_2__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_6_2__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_6_3__din),
    .fifo_A_out_full_n(fifo_A_PE_6_3__full_n),
    .fifo_A_out_write(fifo_A_PE_6_3__write),
    .fifo_B_in_s_dout(fifo_B_PE_6_2__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_6_2__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_6_2__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_6_2__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_6_2__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_7_2__din),
    .fifo_B_out_full_n(fifo_B_PE_7_2__full_n),
    .fifo_B_out_write(fifo_B_PE_7_2__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_6_2__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_6_2__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_6_2__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_105
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_105__ap_start),
    .ap_done(PE_wrapper_105__ap_done),
    .ap_idle(PE_wrapper_105__ap_idle),
    .ap_ready(PE_wrapper_105__ap_ready),
    .idy(64'd3),
    .idx(64'd6),
    .fifo_A_in_s_dout(fifo_A_PE_6_3__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_6_3__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_6_3__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_6_3__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_6_3__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_6_4__din),
    .fifo_A_out_full_n(fifo_A_PE_6_4__full_n),
    .fifo_A_out_write(fifo_A_PE_6_4__write),
    .fifo_B_in_s_dout(fifo_B_PE_6_3__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_6_3__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_6_3__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_6_3__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_6_3__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_7_3__din),
    .fifo_B_out_full_n(fifo_B_PE_7_3__full_n),
    .fifo_B_out_write(fifo_B_PE_7_3__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_6_3__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_6_3__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_6_3__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_106
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_106__ap_start),
    .ap_done(PE_wrapper_106__ap_done),
    .ap_idle(PE_wrapper_106__ap_idle),
    .ap_ready(PE_wrapper_106__ap_ready),
    .idy(64'd4),
    .idx(64'd6),
    .fifo_A_in_s_dout(fifo_A_PE_6_4__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_6_4__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_6_4__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_6_4__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_6_4__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_6_5__din),
    .fifo_A_out_full_n(fifo_A_PE_6_5__full_n),
    .fifo_A_out_write(fifo_A_PE_6_5__write),
    .fifo_B_in_s_dout(fifo_B_PE_6_4__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_6_4__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_6_4__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_6_4__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_6_4__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_7_4__din),
    .fifo_B_out_full_n(fifo_B_PE_7_4__full_n),
    .fifo_B_out_write(fifo_B_PE_7_4__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_6_4__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_6_4__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_6_4__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_107
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_107__ap_start),
    .ap_done(PE_wrapper_107__ap_done),
    .ap_idle(PE_wrapper_107__ap_idle),
    .ap_ready(PE_wrapper_107__ap_ready),
    .idy(64'd5),
    .idx(64'd6),
    .fifo_A_in_s_dout(fifo_A_PE_6_5__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_6_5__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_6_5__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_6_5__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_6_5__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_6_6__din),
    .fifo_A_out_full_n(fifo_A_PE_6_6__full_n),
    .fifo_A_out_write(fifo_A_PE_6_6__write),
    .fifo_B_in_s_dout(fifo_B_PE_6_5__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_6_5__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_6_5__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_6_5__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_6_5__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_7_5__din),
    .fifo_B_out_full_n(fifo_B_PE_7_5__full_n),
    .fifo_B_out_write(fifo_B_PE_7_5__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_6_5__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_6_5__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_6_5__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_108
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_108__ap_start),
    .ap_done(PE_wrapper_108__ap_done),
    .ap_idle(PE_wrapper_108__ap_idle),
    .ap_ready(PE_wrapper_108__ap_ready),
    .idx(64'd6),
    .idy(64'd6),
    .fifo_A_in_s_dout(fifo_A_PE_6_6__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_6_6__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_6_6__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_6_6__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_6_6__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_6_7__din),
    .fifo_A_out_full_n(fifo_A_PE_6_7__full_n),
    .fifo_A_out_write(fifo_A_PE_6_7__write),
    .fifo_B_in_s_dout(fifo_B_PE_6_6__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_6_6__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_6_6__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_6_6__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_6_6__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_7_6__din),
    .fifo_B_out_full_n(fifo_B_PE_7_6__full_n),
    .fifo_B_out_write(fifo_B_PE_7_6__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_6_6__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_6_6__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_6_6__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_109
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_109__ap_start),
    .ap_done(PE_wrapper_109__ap_done),
    .ap_idle(PE_wrapper_109__ap_idle),
    .ap_ready(PE_wrapper_109__ap_ready),
    .idx(64'd6),
    .idy(64'd7),
    .fifo_A_in_s_dout(fifo_A_PE_6_7__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_6_7__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_6_7__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_6_7__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_6_7__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_6_8__din),
    .fifo_A_out_full_n(fifo_A_PE_6_8__full_n),
    .fifo_A_out_write(fifo_A_PE_6_8__write),
    .fifo_B_in_s_dout(fifo_B_PE_6_7__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_6_7__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_6_7__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_6_7__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_6_7__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_7_7__din),
    .fifo_B_out_full_n(fifo_B_PE_7_7__full_n),
    .fifo_B_out_write(fifo_B_PE_7_7__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_6_7__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_6_7__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_6_7__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_110
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_110__ap_start),
    .ap_done(PE_wrapper_110__ap_done),
    .ap_idle(PE_wrapper_110__ap_idle),
    .ap_ready(PE_wrapper_110__ap_ready),
    .idx(64'd6),
    .idy(64'd8),
    .fifo_A_in_s_dout(fifo_A_PE_6_8__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_6_8__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_6_8__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_6_8__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_6_8__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_6_9__din),
    .fifo_A_out_full_n(fifo_A_PE_6_9__full_n),
    .fifo_A_out_write(fifo_A_PE_6_9__write),
    .fifo_B_in_s_dout(fifo_B_PE_6_8__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_6_8__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_6_8__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_6_8__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_6_8__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_7_8__din),
    .fifo_B_out_full_n(fifo_B_PE_7_8__full_n),
    .fifo_B_out_write(fifo_B_PE_7_8__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_6_8__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_6_8__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_6_8__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_111
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_111__ap_start),
    .ap_done(PE_wrapper_111__ap_done),
    .ap_idle(PE_wrapper_111__ap_idle),
    .ap_ready(PE_wrapper_111__ap_ready),
    .idx(64'd6),
    .idy(64'd9),
    .fifo_A_out_din(fifo_A_PE_6_10__din),
    .fifo_A_out_full_n(fifo_A_PE_6_10__full_n),
    .fifo_A_out_write(fifo_A_PE_6_10__write),
    .fifo_A_in_s_dout(fifo_A_PE_6_9__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_6_9__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_6_9__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_6_9__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_6_9__read),
    .fifo_A_in_peek_read(),
    .fifo_B_in_s_dout(fifo_B_PE_6_9__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_6_9__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_6_9__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_6_9__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_6_9__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_7_9__din),
    .fifo_B_out_full_n(fifo_B_PE_7_9__full_n),
    .fifo_B_out_write(fifo_B_PE_7_9__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_6_9__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_6_9__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_6_9__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_112
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_112__ap_start),
    .ap_done(PE_wrapper_112__ap_done),
    .ap_idle(PE_wrapper_112__ap_idle),
    .ap_ready(PE_wrapper_112__ap_ready),
    .idy(64'd10),
    .idx(64'd6),
    .fifo_A_in_s_dout(fifo_A_PE_6_10__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_6_10__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_6_10__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_6_10__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_6_10__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_6_11__din),
    .fifo_A_out_full_n(fifo_A_PE_6_11__full_n),
    .fifo_A_out_write(fifo_A_PE_6_11__write),
    .fifo_B_in_s_dout(fifo_B_PE_6_10__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_6_10__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_6_10__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_6_10__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_6_10__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_7_10__din),
    .fifo_B_out_full_n(fifo_B_PE_7_10__full_n),
    .fifo_B_out_write(fifo_B_PE_7_10__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_6_10__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_6_10__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_6_10__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_113
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_113__ap_start),
    .ap_done(PE_wrapper_113__ap_done),
    .ap_idle(PE_wrapper_113__ap_idle),
    .ap_ready(PE_wrapper_113__ap_ready),
    .idy(64'd11),
    .idx(64'd6),
    .fifo_A_in_s_dout(fifo_A_PE_6_11__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_6_11__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_6_11__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_6_11__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_6_11__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_6_12__din),
    .fifo_A_out_full_n(fifo_A_PE_6_12__full_n),
    .fifo_A_out_write(fifo_A_PE_6_12__write),
    .fifo_B_in_s_dout(fifo_B_PE_6_11__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_6_11__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_6_11__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_6_11__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_6_11__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_7_11__din),
    .fifo_B_out_full_n(fifo_B_PE_7_11__full_n),
    .fifo_B_out_write(fifo_B_PE_7_11__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_6_11__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_6_11__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_6_11__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_114
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_114__ap_start),
    .ap_done(PE_wrapper_114__ap_done),
    .ap_idle(PE_wrapper_114__ap_idle),
    .ap_ready(PE_wrapper_114__ap_ready),
    .idy(64'd12),
    .idx(64'd6),
    .fifo_A_in_s_dout(fifo_A_PE_6_12__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_6_12__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_6_12__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_6_12__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_6_12__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_6_13__din),
    .fifo_A_out_full_n(fifo_A_PE_6_13__full_n),
    .fifo_A_out_write(fifo_A_PE_6_13__write),
    .fifo_B_in_s_dout(fifo_B_PE_6_12__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_6_12__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_6_12__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_6_12__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_6_12__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_7_12__din),
    .fifo_B_out_full_n(fifo_B_PE_7_12__full_n),
    .fifo_B_out_write(fifo_B_PE_7_12__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_6_12__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_6_12__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_6_12__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_115
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_115__ap_start),
    .ap_done(PE_wrapper_115__ap_done),
    .ap_idle(PE_wrapper_115__ap_idle),
    .ap_ready(PE_wrapper_115__ap_ready),
    .idy(64'd13),
    .idx(64'd6),
    .fifo_A_in_s_dout(fifo_A_PE_6_13__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_6_13__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_6_13__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_6_13__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_6_13__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_6_14__din),
    .fifo_A_out_full_n(fifo_A_PE_6_14__full_n),
    .fifo_A_out_write(fifo_A_PE_6_14__write),
    .fifo_B_in_s_dout(fifo_B_PE_6_13__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_6_13__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_6_13__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_6_13__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_6_13__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_7_13__din),
    .fifo_B_out_full_n(fifo_B_PE_7_13__full_n),
    .fifo_B_out_write(fifo_B_PE_7_13__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_6_13__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_6_13__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_6_13__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_116
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_116__ap_start),
    .ap_done(PE_wrapper_116__ap_done),
    .ap_idle(PE_wrapper_116__ap_idle),
    .ap_ready(PE_wrapper_116__ap_ready),
    .idy(64'd14),
    .idx(64'd6),
    .fifo_A_in_s_dout(fifo_A_PE_6_14__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_6_14__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_6_14__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_6_14__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_6_14__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_6_15__din),
    .fifo_A_out_full_n(fifo_A_PE_6_15__full_n),
    .fifo_A_out_write(fifo_A_PE_6_15__write),
    .fifo_B_in_s_dout(fifo_B_PE_6_14__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_6_14__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_6_14__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_6_14__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_6_14__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_7_14__din),
    .fifo_B_out_full_n(fifo_B_PE_7_14__full_n),
    .fifo_B_out_write(fifo_B_PE_7_14__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_6_14__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_6_14__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_6_14__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_117
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_117__ap_start),
    .ap_done(PE_wrapper_117__ap_done),
    .ap_idle(PE_wrapper_117__ap_idle),
    .ap_ready(PE_wrapper_117__ap_ready),
    .idy(64'd15),
    .idx(64'd6),
    .fifo_A_in_s_dout(fifo_A_PE_6_15__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_6_15__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_6_15__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_6_15__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_6_15__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_6_16__din),
    .fifo_A_out_full_n(fifo_A_PE_6_16__full_n),
    .fifo_A_out_write(fifo_A_PE_6_16__write),
    .fifo_B_in_s_dout(fifo_B_PE_6_15__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_6_15__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_6_15__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_6_15__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_6_15__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_7_15__din),
    .fifo_B_out_full_n(fifo_B_PE_7_15__full_n),
    .fifo_B_out_write(fifo_B_PE_7_15__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_6_15__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_6_15__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_6_15__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_118
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_118__ap_start),
    .ap_done(PE_wrapper_118__ap_done),
    .ap_idle(PE_wrapper_118__ap_idle),
    .ap_ready(PE_wrapper_118__ap_ready),
    .idy(64'd16),
    .idx(64'd6),
    .fifo_A_in_s_dout(fifo_A_PE_6_16__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_6_16__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_6_16__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_6_16__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_6_16__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_6_17__din),
    .fifo_A_out_full_n(fifo_A_PE_6_17__full_n),
    .fifo_A_out_write(fifo_A_PE_6_17__write),
    .fifo_B_in_s_dout(fifo_B_PE_6_16__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_6_16__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_6_16__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_6_16__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_6_16__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_7_16__din),
    .fifo_B_out_full_n(fifo_B_PE_7_16__full_n),
    .fifo_B_out_write(fifo_B_PE_7_16__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_6_16__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_6_16__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_6_16__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_119
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_119__ap_start),
    .ap_done(PE_wrapper_119__ap_done),
    .ap_idle(PE_wrapper_119__ap_idle),
    .ap_ready(PE_wrapper_119__ap_ready),
    .idy(64'd0),
    .idx(64'd7),
    .fifo_A_in_s_dout(fifo_A_PE_7_0__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_7_0__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_7_0__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_7_0__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_7_0__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_7_1__din),
    .fifo_A_out_full_n(fifo_A_PE_7_1__full_n),
    .fifo_A_out_write(fifo_A_PE_7_1__write),
    .fifo_B_in_s_dout(fifo_B_PE_7_0__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_7_0__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_7_0__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_7_0__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_7_0__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_8_0__din),
    .fifo_B_out_full_n(fifo_B_PE_8_0__full_n),
    .fifo_B_out_write(fifo_B_PE_8_0__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_7_0__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_7_0__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_7_0__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_120
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_120__ap_start),
    .ap_done(PE_wrapper_120__ap_done),
    .ap_idle(PE_wrapper_120__ap_idle),
    .ap_ready(PE_wrapper_120__ap_ready),
    .idy(64'd1),
    .idx(64'd7),
    .fifo_A_in_s_dout(fifo_A_PE_7_1__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_7_1__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_7_1__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_7_1__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_7_1__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_7_2__din),
    .fifo_A_out_full_n(fifo_A_PE_7_2__full_n),
    .fifo_A_out_write(fifo_A_PE_7_2__write),
    .fifo_B_in_s_dout(fifo_B_PE_7_1__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_7_1__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_7_1__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_7_1__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_7_1__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_8_1__din),
    .fifo_B_out_full_n(fifo_B_PE_8_1__full_n),
    .fifo_B_out_write(fifo_B_PE_8_1__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_7_1__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_7_1__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_7_1__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_121
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_121__ap_start),
    .ap_done(PE_wrapper_121__ap_done),
    .ap_idle(PE_wrapper_121__ap_idle),
    .ap_ready(PE_wrapper_121__ap_ready),
    .idy(64'd2),
    .idx(64'd7),
    .fifo_A_in_s_dout(fifo_A_PE_7_2__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_7_2__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_7_2__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_7_2__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_7_2__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_7_3__din),
    .fifo_A_out_full_n(fifo_A_PE_7_3__full_n),
    .fifo_A_out_write(fifo_A_PE_7_3__write),
    .fifo_B_in_s_dout(fifo_B_PE_7_2__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_7_2__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_7_2__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_7_2__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_7_2__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_8_2__din),
    .fifo_B_out_full_n(fifo_B_PE_8_2__full_n),
    .fifo_B_out_write(fifo_B_PE_8_2__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_7_2__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_7_2__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_7_2__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_122
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_122__ap_start),
    .ap_done(PE_wrapper_122__ap_done),
    .ap_idle(PE_wrapper_122__ap_idle),
    .ap_ready(PE_wrapper_122__ap_ready),
    .idy(64'd3),
    .idx(64'd7),
    .fifo_A_in_s_dout(fifo_A_PE_7_3__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_7_3__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_7_3__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_7_3__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_7_3__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_7_4__din),
    .fifo_A_out_full_n(fifo_A_PE_7_4__full_n),
    .fifo_A_out_write(fifo_A_PE_7_4__write),
    .fifo_B_in_s_dout(fifo_B_PE_7_3__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_7_3__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_7_3__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_7_3__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_7_3__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_8_3__din),
    .fifo_B_out_full_n(fifo_B_PE_8_3__full_n),
    .fifo_B_out_write(fifo_B_PE_8_3__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_7_3__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_7_3__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_7_3__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_123
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_123__ap_start),
    .ap_done(PE_wrapper_123__ap_done),
    .ap_idle(PE_wrapper_123__ap_idle),
    .ap_ready(PE_wrapper_123__ap_ready),
    .idy(64'd4),
    .idx(64'd7),
    .fifo_A_in_s_dout(fifo_A_PE_7_4__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_7_4__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_7_4__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_7_4__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_7_4__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_7_5__din),
    .fifo_A_out_full_n(fifo_A_PE_7_5__full_n),
    .fifo_A_out_write(fifo_A_PE_7_5__write),
    .fifo_B_in_s_dout(fifo_B_PE_7_4__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_7_4__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_7_4__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_7_4__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_7_4__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_8_4__din),
    .fifo_B_out_full_n(fifo_B_PE_8_4__full_n),
    .fifo_B_out_write(fifo_B_PE_8_4__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_7_4__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_7_4__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_7_4__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_124
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_124__ap_start),
    .ap_done(PE_wrapper_124__ap_done),
    .ap_idle(PE_wrapper_124__ap_idle),
    .ap_ready(PE_wrapper_124__ap_ready),
    .idy(64'd5),
    .idx(64'd7),
    .fifo_A_in_s_dout(fifo_A_PE_7_5__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_7_5__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_7_5__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_7_5__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_7_5__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_7_6__din),
    .fifo_A_out_full_n(fifo_A_PE_7_6__full_n),
    .fifo_A_out_write(fifo_A_PE_7_6__write),
    .fifo_B_in_s_dout(fifo_B_PE_7_5__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_7_5__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_7_5__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_7_5__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_7_5__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_8_5__din),
    .fifo_B_out_full_n(fifo_B_PE_8_5__full_n),
    .fifo_B_out_write(fifo_B_PE_8_5__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_7_5__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_7_5__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_7_5__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_125
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_125__ap_start),
    .ap_done(PE_wrapper_125__ap_done),
    .ap_idle(PE_wrapper_125__ap_idle),
    .ap_ready(PE_wrapper_125__ap_ready),
    .idy(64'd6),
    .idx(64'd7),
    .fifo_A_in_s_dout(fifo_A_PE_7_6__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_7_6__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_7_6__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_7_6__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_7_6__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_7_7__din),
    .fifo_A_out_full_n(fifo_A_PE_7_7__full_n),
    .fifo_A_out_write(fifo_A_PE_7_7__write),
    .fifo_B_in_s_dout(fifo_B_PE_7_6__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_7_6__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_7_6__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_7_6__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_7_6__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_8_6__din),
    .fifo_B_out_full_n(fifo_B_PE_8_6__full_n),
    .fifo_B_out_write(fifo_B_PE_8_6__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_7_6__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_7_6__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_7_6__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_126
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_126__ap_start),
    .ap_done(PE_wrapper_126__ap_done),
    .ap_idle(PE_wrapper_126__ap_idle),
    .ap_ready(PE_wrapper_126__ap_ready),
    .idx(64'd7),
    .idy(64'd7),
    .fifo_A_in_s_dout(fifo_A_PE_7_7__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_7_7__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_7_7__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_7_7__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_7_7__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_7_8__din),
    .fifo_A_out_full_n(fifo_A_PE_7_8__full_n),
    .fifo_A_out_write(fifo_A_PE_7_8__write),
    .fifo_B_in_s_dout(fifo_B_PE_7_7__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_7_7__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_7_7__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_7_7__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_7_7__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_8_7__din),
    .fifo_B_out_full_n(fifo_B_PE_8_7__full_n),
    .fifo_B_out_write(fifo_B_PE_8_7__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_7_7__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_7_7__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_7_7__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_127
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_127__ap_start),
    .ap_done(PE_wrapper_127__ap_done),
    .ap_idle(PE_wrapper_127__ap_idle),
    .ap_ready(PE_wrapper_127__ap_ready),
    .idx(64'd7),
    .idy(64'd8),
    .fifo_A_in_s_dout(fifo_A_PE_7_8__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_7_8__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_7_8__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_7_8__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_7_8__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_7_9__din),
    .fifo_A_out_full_n(fifo_A_PE_7_9__full_n),
    .fifo_A_out_write(fifo_A_PE_7_9__write),
    .fifo_B_in_s_dout(fifo_B_PE_7_8__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_7_8__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_7_8__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_7_8__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_7_8__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_8_8__din),
    .fifo_B_out_full_n(fifo_B_PE_8_8__full_n),
    .fifo_B_out_write(fifo_B_PE_8_8__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_7_8__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_7_8__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_7_8__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_128
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_128__ap_start),
    .ap_done(PE_wrapper_128__ap_done),
    .ap_idle(PE_wrapper_128__ap_idle),
    .ap_ready(PE_wrapper_128__ap_ready),
    .idx(64'd7),
    .idy(64'd9),
    .fifo_A_out_din(fifo_A_PE_7_10__din),
    .fifo_A_out_full_n(fifo_A_PE_7_10__full_n),
    .fifo_A_out_write(fifo_A_PE_7_10__write),
    .fifo_A_in_s_dout(fifo_A_PE_7_9__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_7_9__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_7_9__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_7_9__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_7_9__read),
    .fifo_A_in_peek_read(),
    .fifo_B_in_s_dout(fifo_B_PE_7_9__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_7_9__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_7_9__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_7_9__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_7_9__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_8_9__din),
    .fifo_B_out_full_n(fifo_B_PE_8_9__full_n),
    .fifo_B_out_write(fifo_B_PE_8_9__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_7_9__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_7_9__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_7_9__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_129
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_129__ap_start),
    .ap_done(PE_wrapper_129__ap_done),
    .ap_idle(PE_wrapper_129__ap_idle),
    .ap_ready(PE_wrapper_129__ap_ready),
    .idy(64'd10),
    .idx(64'd7),
    .fifo_A_in_s_dout(fifo_A_PE_7_10__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_7_10__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_7_10__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_7_10__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_7_10__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_7_11__din),
    .fifo_A_out_full_n(fifo_A_PE_7_11__full_n),
    .fifo_A_out_write(fifo_A_PE_7_11__write),
    .fifo_B_in_s_dout(fifo_B_PE_7_10__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_7_10__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_7_10__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_7_10__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_7_10__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_8_10__din),
    .fifo_B_out_full_n(fifo_B_PE_8_10__full_n),
    .fifo_B_out_write(fifo_B_PE_8_10__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_7_10__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_7_10__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_7_10__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_130
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_130__ap_start),
    .ap_done(PE_wrapper_130__ap_done),
    .ap_idle(PE_wrapper_130__ap_idle),
    .ap_ready(PE_wrapper_130__ap_ready),
    .idy(64'd11),
    .idx(64'd7),
    .fifo_A_in_s_dout(fifo_A_PE_7_11__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_7_11__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_7_11__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_7_11__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_7_11__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_7_12__din),
    .fifo_A_out_full_n(fifo_A_PE_7_12__full_n),
    .fifo_A_out_write(fifo_A_PE_7_12__write),
    .fifo_B_in_s_dout(fifo_B_PE_7_11__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_7_11__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_7_11__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_7_11__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_7_11__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_8_11__din),
    .fifo_B_out_full_n(fifo_B_PE_8_11__full_n),
    .fifo_B_out_write(fifo_B_PE_8_11__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_7_11__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_7_11__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_7_11__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_131
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_131__ap_start),
    .ap_done(PE_wrapper_131__ap_done),
    .ap_idle(PE_wrapper_131__ap_idle),
    .ap_ready(PE_wrapper_131__ap_ready),
    .idy(64'd12),
    .idx(64'd7),
    .fifo_A_in_s_dout(fifo_A_PE_7_12__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_7_12__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_7_12__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_7_12__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_7_12__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_7_13__din),
    .fifo_A_out_full_n(fifo_A_PE_7_13__full_n),
    .fifo_A_out_write(fifo_A_PE_7_13__write),
    .fifo_B_in_s_dout(fifo_B_PE_7_12__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_7_12__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_7_12__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_7_12__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_7_12__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_8_12__din),
    .fifo_B_out_full_n(fifo_B_PE_8_12__full_n),
    .fifo_B_out_write(fifo_B_PE_8_12__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_7_12__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_7_12__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_7_12__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_132
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_132__ap_start),
    .ap_done(PE_wrapper_132__ap_done),
    .ap_idle(PE_wrapper_132__ap_idle),
    .ap_ready(PE_wrapper_132__ap_ready),
    .idy(64'd13),
    .idx(64'd7),
    .fifo_A_in_s_dout(fifo_A_PE_7_13__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_7_13__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_7_13__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_7_13__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_7_13__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_7_14__din),
    .fifo_A_out_full_n(fifo_A_PE_7_14__full_n),
    .fifo_A_out_write(fifo_A_PE_7_14__write),
    .fifo_B_in_s_dout(fifo_B_PE_7_13__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_7_13__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_7_13__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_7_13__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_7_13__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_8_13__din),
    .fifo_B_out_full_n(fifo_B_PE_8_13__full_n),
    .fifo_B_out_write(fifo_B_PE_8_13__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_7_13__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_7_13__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_7_13__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_133
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_133__ap_start),
    .ap_done(PE_wrapper_133__ap_done),
    .ap_idle(PE_wrapper_133__ap_idle),
    .ap_ready(PE_wrapper_133__ap_ready),
    .idy(64'd14),
    .idx(64'd7),
    .fifo_A_in_s_dout(fifo_A_PE_7_14__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_7_14__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_7_14__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_7_14__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_7_14__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_7_15__din),
    .fifo_A_out_full_n(fifo_A_PE_7_15__full_n),
    .fifo_A_out_write(fifo_A_PE_7_15__write),
    .fifo_B_in_s_dout(fifo_B_PE_7_14__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_7_14__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_7_14__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_7_14__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_7_14__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_8_14__din),
    .fifo_B_out_full_n(fifo_B_PE_8_14__full_n),
    .fifo_B_out_write(fifo_B_PE_8_14__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_7_14__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_7_14__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_7_14__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_134
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_134__ap_start),
    .ap_done(PE_wrapper_134__ap_done),
    .ap_idle(PE_wrapper_134__ap_idle),
    .ap_ready(PE_wrapper_134__ap_ready),
    .idy(64'd15),
    .idx(64'd7),
    .fifo_A_in_s_dout(fifo_A_PE_7_15__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_7_15__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_7_15__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_7_15__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_7_15__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_7_16__din),
    .fifo_A_out_full_n(fifo_A_PE_7_16__full_n),
    .fifo_A_out_write(fifo_A_PE_7_16__write),
    .fifo_B_in_s_dout(fifo_B_PE_7_15__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_7_15__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_7_15__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_7_15__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_7_15__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_8_15__din),
    .fifo_B_out_full_n(fifo_B_PE_8_15__full_n),
    .fifo_B_out_write(fifo_B_PE_8_15__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_7_15__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_7_15__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_7_15__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_135
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_135__ap_start),
    .ap_done(PE_wrapper_135__ap_done),
    .ap_idle(PE_wrapper_135__ap_idle),
    .ap_ready(PE_wrapper_135__ap_ready),
    .idy(64'd16),
    .idx(64'd7),
    .fifo_A_in_s_dout(fifo_A_PE_7_16__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_7_16__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_7_16__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_7_16__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_7_16__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_7_17__din),
    .fifo_A_out_full_n(fifo_A_PE_7_17__full_n),
    .fifo_A_out_write(fifo_A_PE_7_17__write),
    .fifo_B_in_s_dout(fifo_B_PE_7_16__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_7_16__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_7_16__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_7_16__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_7_16__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_8_16__din),
    .fifo_B_out_full_n(fifo_B_PE_8_16__full_n),
    .fifo_B_out_write(fifo_B_PE_8_16__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_7_16__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_7_16__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_7_16__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_136
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_136__ap_start),
    .ap_done(PE_wrapper_136__ap_done),
    .ap_idle(PE_wrapper_136__ap_idle),
    .ap_ready(PE_wrapper_136__ap_ready),
    .idy(64'd0),
    .idx(64'd8),
    .fifo_A_in_s_dout(fifo_A_PE_8_0__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_8_0__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_8_0__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_8_0__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_8_0__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_8_1__din),
    .fifo_A_out_full_n(fifo_A_PE_8_1__full_n),
    .fifo_A_out_write(fifo_A_PE_8_1__write),
    .fifo_B_in_s_dout(fifo_B_PE_8_0__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_8_0__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_8_0__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_8_0__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_8_0__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_9_0__din),
    .fifo_B_out_full_n(fifo_B_PE_9_0__full_n),
    .fifo_B_out_write(fifo_B_PE_9_0__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_8_0__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_8_0__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_8_0__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_137
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_137__ap_start),
    .ap_done(PE_wrapper_137__ap_done),
    .ap_idle(PE_wrapper_137__ap_idle),
    .ap_ready(PE_wrapper_137__ap_ready),
    .idy(64'd1),
    .idx(64'd8),
    .fifo_A_in_s_dout(fifo_A_PE_8_1__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_8_1__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_8_1__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_8_1__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_8_1__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_8_2__din),
    .fifo_A_out_full_n(fifo_A_PE_8_2__full_n),
    .fifo_A_out_write(fifo_A_PE_8_2__write),
    .fifo_B_in_s_dout(fifo_B_PE_8_1__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_8_1__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_8_1__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_8_1__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_8_1__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_9_1__din),
    .fifo_B_out_full_n(fifo_B_PE_9_1__full_n),
    .fifo_B_out_write(fifo_B_PE_9_1__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_8_1__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_8_1__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_8_1__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_138
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_138__ap_start),
    .ap_done(PE_wrapper_138__ap_done),
    .ap_idle(PE_wrapper_138__ap_idle),
    .ap_ready(PE_wrapper_138__ap_ready),
    .idy(64'd2),
    .idx(64'd8),
    .fifo_A_in_s_dout(fifo_A_PE_8_2__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_8_2__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_8_2__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_8_2__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_8_2__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_8_3__din),
    .fifo_A_out_full_n(fifo_A_PE_8_3__full_n),
    .fifo_A_out_write(fifo_A_PE_8_3__write),
    .fifo_B_in_s_dout(fifo_B_PE_8_2__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_8_2__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_8_2__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_8_2__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_8_2__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_9_2__din),
    .fifo_B_out_full_n(fifo_B_PE_9_2__full_n),
    .fifo_B_out_write(fifo_B_PE_9_2__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_8_2__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_8_2__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_8_2__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_139
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_139__ap_start),
    .ap_done(PE_wrapper_139__ap_done),
    .ap_idle(PE_wrapper_139__ap_idle),
    .ap_ready(PE_wrapper_139__ap_ready),
    .idy(64'd3),
    .idx(64'd8),
    .fifo_A_in_s_dout(fifo_A_PE_8_3__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_8_3__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_8_3__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_8_3__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_8_3__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_8_4__din),
    .fifo_A_out_full_n(fifo_A_PE_8_4__full_n),
    .fifo_A_out_write(fifo_A_PE_8_4__write),
    .fifo_B_in_s_dout(fifo_B_PE_8_3__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_8_3__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_8_3__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_8_3__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_8_3__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_9_3__din),
    .fifo_B_out_full_n(fifo_B_PE_9_3__full_n),
    .fifo_B_out_write(fifo_B_PE_9_3__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_8_3__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_8_3__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_8_3__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_140
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_140__ap_start),
    .ap_done(PE_wrapper_140__ap_done),
    .ap_idle(PE_wrapper_140__ap_idle),
    .ap_ready(PE_wrapper_140__ap_ready),
    .idy(64'd4),
    .idx(64'd8),
    .fifo_A_in_s_dout(fifo_A_PE_8_4__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_8_4__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_8_4__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_8_4__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_8_4__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_8_5__din),
    .fifo_A_out_full_n(fifo_A_PE_8_5__full_n),
    .fifo_A_out_write(fifo_A_PE_8_5__write),
    .fifo_B_in_s_dout(fifo_B_PE_8_4__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_8_4__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_8_4__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_8_4__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_8_4__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_9_4__din),
    .fifo_B_out_full_n(fifo_B_PE_9_4__full_n),
    .fifo_B_out_write(fifo_B_PE_9_4__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_8_4__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_8_4__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_8_4__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_141
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_141__ap_start),
    .ap_done(PE_wrapper_141__ap_done),
    .ap_idle(PE_wrapper_141__ap_idle),
    .ap_ready(PE_wrapper_141__ap_ready),
    .idy(64'd5),
    .idx(64'd8),
    .fifo_A_in_s_dout(fifo_A_PE_8_5__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_8_5__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_8_5__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_8_5__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_8_5__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_8_6__din),
    .fifo_A_out_full_n(fifo_A_PE_8_6__full_n),
    .fifo_A_out_write(fifo_A_PE_8_6__write),
    .fifo_B_in_s_dout(fifo_B_PE_8_5__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_8_5__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_8_5__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_8_5__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_8_5__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_9_5__din),
    .fifo_B_out_full_n(fifo_B_PE_9_5__full_n),
    .fifo_B_out_write(fifo_B_PE_9_5__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_8_5__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_8_5__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_8_5__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_142
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_142__ap_start),
    .ap_done(PE_wrapper_142__ap_done),
    .ap_idle(PE_wrapper_142__ap_idle),
    .ap_ready(PE_wrapper_142__ap_ready),
    .idy(64'd6),
    .idx(64'd8),
    .fifo_A_in_s_dout(fifo_A_PE_8_6__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_8_6__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_8_6__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_8_6__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_8_6__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_8_7__din),
    .fifo_A_out_full_n(fifo_A_PE_8_7__full_n),
    .fifo_A_out_write(fifo_A_PE_8_7__write),
    .fifo_B_in_s_dout(fifo_B_PE_8_6__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_8_6__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_8_6__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_8_6__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_8_6__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_9_6__din),
    .fifo_B_out_full_n(fifo_B_PE_9_6__full_n),
    .fifo_B_out_write(fifo_B_PE_9_6__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_8_6__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_8_6__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_8_6__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_143
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_143__ap_start),
    .ap_done(PE_wrapper_143__ap_done),
    .ap_idle(PE_wrapper_143__ap_idle),
    .ap_ready(PE_wrapper_143__ap_ready),
    .idy(64'd7),
    .idx(64'd8),
    .fifo_A_in_s_dout(fifo_A_PE_8_7__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_8_7__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_8_7__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_8_7__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_8_7__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_8_8__din),
    .fifo_A_out_full_n(fifo_A_PE_8_8__full_n),
    .fifo_A_out_write(fifo_A_PE_8_8__write),
    .fifo_B_in_s_dout(fifo_B_PE_8_7__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_8_7__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_8_7__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_8_7__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_8_7__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_9_7__din),
    .fifo_B_out_full_n(fifo_B_PE_9_7__full_n),
    .fifo_B_out_write(fifo_B_PE_9_7__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_8_7__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_8_7__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_8_7__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_144
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_144__ap_start),
    .ap_done(PE_wrapper_144__ap_done),
    .ap_idle(PE_wrapper_144__ap_idle),
    .ap_ready(PE_wrapper_144__ap_ready),
    .idx(64'd8),
    .idy(64'd8),
    .fifo_A_in_s_dout(fifo_A_PE_8_8__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_8_8__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_8_8__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_8_8__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_8_8__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_8_9__din),
    .fifo_A_out_full_n(fifo_A_PE_8_9__full_n),
    .fifo_A_out_write(fifo_A_PE_8_9__write),
    .fifo_B_in_s_dout(fifo_B_PE_8_8__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_8_8__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_8_8__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_8_8__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_8_8__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_9_8__din),
    .fifo_B_out_full_n(fifo_B_PE_9_8__full_n),
    .fifo_B_out_write(fifo_B_PE_9_8__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_8_8__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_8_8__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_8_8__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_145
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_145__ap_start),
    .ap_done(PE_wrapper_145__ap_done),
    .ap_idle(PE_wrapper_145__ap_idle),
    .ap_ready(PE_wrapper_145__ap_ready),
    .idx(64'd8),
    .idy(64'd9),
    .fifo_A_out_din(fifo_A_PE_8_10__din),
    .fifo_A_out_full_n(fifo_A_PE_8_10__full_n),
    .fifo_A_out_write(fifo_A_PE_8_10__write),
    .fifo_A_in_s_dout(fifo_A_PE_8_9__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_8_9__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_8_9__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_8_9__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_8_9__read),
    .fifo_A_in_peek_read(),
    .fifo_B_in_s_dout(fifo_B_PE_8_9__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_8_9__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_8_9__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_8_9__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_8_9__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_9_9__din),
    .fifo_B_out_full_n(fifo_B_PE_9_9__full_n),
    .fifo_B_out_write(fifo_B_PE_9_9__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_8_9__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_8_9__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_8_9__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_146
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_146__ap_start),
    .ap_done(PE_wrapper_146__ap_done),
    .ap_idle(PE_wrapper_146__ap_idle),
    .ap_ready(PE_wrapper_146__ap_ready),
    .idy(64'd10),
    .idx(64'd8),
    .fifo_A_in_s_dout(fifo_A_PE_8_10__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_8_10__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_8_10__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_8_10__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_8_10__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_8_11__din),
    .fifo_A_out_full_n(fifo_A_PE_8_11__full_n),
    .fifo_A_out_write(fifo_A_PE_8_11__write),
    .fifo_B_in_s_dout(fifo_B_PE_8_10__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_8_10__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_8_10__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_8_10__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_8_10__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_9_10__din),
    .fifo_B_out_full_n(fifo_B_PE_9_10__full_n),
    .fifo_B_out_write(fifo_B_PE_9_10__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_8_10__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_8_10__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_8_10__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_147
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_147__ap_start),
    .ap_done(PE_wrapper_147__ap_done),
    .ap_idle(PE_wrapper_147__ap_idle),
    .ap_ready(PE_wrapper_147__ap_ready),
    .idy(64'd11),
    .idx(64'd8),
    .fifo_A_in_s_dout(fifo_A_PE_8_11__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_8_11__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_8_11__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_8_11__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_8_11__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_8_12__din),
    .fifo_A_out_full_n(fifo_A_PE_8_12__full_n),
    .fifo_A_out_write(fifo_A_PE_8_12__write),
    .fifo_B_in_s_dout(fifo_B_PE_8_11__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_8_11__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_8_11__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_8_11__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_8_11__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_9_11__din),
    .fifo_B_out_full_n(fifo_B_PE_9_11__full_n),
    .fifo_B_out_write(fifo_B_PE_9_11__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_8_11__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_8_11__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_8_11__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_148
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_148__ap_start),
    .ap_done(PE_wrapper_148__ap_done),
    .ap_idle(PE_wrapper_148__ap_idle),
    .ap_ready(PE_wrapper_148__ap_ready),
    .idy(64'd12),
    .idx(64'd8),
    .fifo_A_in_s_dout(fifo_A_PE_8_12__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_8_12__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_8_12__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_8_12__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_8_12__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_8_13__din),
    .fifo_A_out_full_n(fifo_A_PE_8_13__full_n),
    .fifo_A_out_write(fifo_A_PE_8_13__write),
    .fifo_B_in_s_dout(fifo_B_PE_8_12__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_8_12__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_8_12__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_8_12__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_8_12__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_9_12__din),
    .fifo_B_out_full_n(fifo_B_PE_9_12__full_n),
    .fifo_B_out_write(fifo_B_PE_9_12__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_8_12__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_8_12__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_8_12__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_149
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_149__ap_start),
    .ap_done(PE_wrapper_149__ap_done),
    .ap_idle(PE_wrapper_149__ap_idle),
    .ap_ready(PE_wrapper_149__ap_ready),
    .idy(64'd13),
    .idx(64'd8),
    .fifo_A_in_s_dout(fifo_A_PE_8_13__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_8_13__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_8_13__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_8_13__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_8_13__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_8_14__din),
    .fifo_A_out_full_n(fifo_A_PE_8_14__full_n),
    .fifo_A_out_write(fifo_A_PE_8_14__write),
    .fifo_B_in_s_dout(fifo_B_PE_8_13__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_8_13__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_8_13__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_8_13__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_8_13__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_9_13__din),
    .fifo_B_out_full_n(fifo_B_PE_9_13__full_n),
    .fifo_B_out_write(fifo_B_PE_9_13__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_8_13__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_8_13__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_8_13__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_150
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_150__ap_start),
    .ap_done(PE_wrapper_150__ap_done),
    .ap_idle(PE_wrapper_150__ap_idle),
    .ap_ready(PE_wrapper_150__ap_ready),
    .idy(64'd14),
    .idx(64'd8),
    .fifo_A_in_s_dout(fifo_A_PE_8_14__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_8_14__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_8_14__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_8_14__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_8_14__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_8_15__din),
    .fifo_A_out_full_n(fifo_A_PE_8_15__full_n),
    .fifo_A_out_write(fifo_A_PE_8_15__write),
    .fifo_B_in_s_dout(fifo_B_PE_8_14__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_8_14__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_8_14__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_8_14__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_8_14__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_9_14__din),
    .fifo_B_out_full_n(fifo_B_PE_9_14__full_n),
    .fifo_B_out_write(fifo_B_PE_9_14__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_8_14__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_8_14__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_8_14__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_151
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_151__ap_start),
    .ap_done(PE_wrapper_151__ap_done),
    .ap_idle(PE_wrapper_151__ap_idle),
    .ap_ready(PE_wrapper_151__ap_ready),
    .idy(64'd15),
    .idx(64'd8),
    .fifo_A_in_s_dout(fifo_A_PE_8_15__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_8_15__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_8_15__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_8_15__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_8_15__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_8_16__din),
    .fifo_A_out_full_n(fifo_A_PE_8_16__full_n),
    .fifo_A_out_write(fifo_A_PE_8_16__write),
    .fifo_B_in_s_dout(fifo_B_PE_8_15__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_8_15__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_8_15__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_8_15__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_8_15__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_9_15__din),
    .fifo_B_out_full_n(fifo_B_PE_9_15__full_n),
    .fifo_B_out_write(fifo_B_PE_9_15__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_8_15__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_8_15__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_8_15__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_152
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_152__ap_start),
    .ap_done(PE_wrapper_152__ap_done),
    .ap_idle(PE_wrapper_152__ap_idle),
    .ap_ready(PE_wrapper_152__ap_ready),
    .idy(64'd16),
    .idx(64'd8),
    .fifo_A_in_s_dout(fifo_A_PE_8_16__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_8_16__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_8_16__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_8_16__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_8_16__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_8_17__din),
    .fifo_A_out_full_n(fifo_A_PE_8_17__full_n),
    .fifo_A_out_write(fifo_A_PE_8_17__write),
    .fifo_B_in_s_dout(fifo_B_PE_8_16__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_8_16__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_8_16__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_8_16__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_8_16__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_9_16__din),
    .fifo_B_out_full_n(fifo_B_PE_9_16__full_n),
    .fifo_B_out_write(fifo_B_PE_9_16__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_8_16__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_8_16__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_8_16__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_153
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_153__ap_start),
    .ap_done(PE_wrapper_153__ap_done),
    .ap_idle(PE_wrapper_153__ap_idle),
    .ap_ready(PE_wrapper_153__ap_ready),
    .idy(64'd0),
    .idx(64'd9),
    .fifo_A_in_s_dout(fifo_A_PE_9_0__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_9_0__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_9_0__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_9_0__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_9_0__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_9_1__din),
    .fifo_A_out_full_n(fifo_A_PE_9_1__full_n),
    .fifo_A_out_write(fifo_A_PE_9_1__write),
    .fifo_B_out_din(fifo_B_PE_10_0__din),
    .fifo_B_out_full_n(fifo_B_PE_10_0__full_n),
    .fifo_B_out_write(fifo_B_PE_10_0__write),
    .fifo_B_in_s_dout(fifo_B_PE_9_0__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_9_0__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_9_0__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_9_0__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_9_0__read),
    .fifo_B_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_PE_9_0__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_9_0__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_9_0__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_154
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_154__ap_start),
    .ap_done(PE_wrapper_154__ap_done),
    .ap_idle(PE_wrapper_154__ap_idle),
    .ap_ready(PE_wrapper_154__ap_ready),
    .idy(64'd1),
    .idx(64'd9),
    .fifo_A_in_s_dout(fifo_A_PE_9_1__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_9_1__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_9_1__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_9_1__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_9_1__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_9_2__din),
    .fifo_A_out_full_n(fifo_A_PE_9_2__full_n),
    .fifo_A_out_write(fifo_A_PE_9_2__write),
    .fifo_B_out_din(fifo_B_PE_10_1__din),
    .fifo_B_out_full_n(fifo_B_PE_10_1__full_n),
    .fifo_B_out_write(fifo_B_PE_10_1__write),
    .fifo_B_in_s_dout(fifo_B_PE_9_1__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_9_1__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_9_1__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_9_1__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_9_1__read),
    .fifo_B_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_PE_9_1__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_9_1__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_9_1__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_155
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_155__ap_start),
    .ap_done(PE_wrapper_155__ap_done),
    .ap_idle(PE_wrapper_155__ap_idle),
    .ap_ready(PE_wrapper_155__ap_ready),
    .idy(64'd2),
    .idx(64'd9),
    .fifo_A_in_s_dout(fifo_A_PE_9_2__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_9_2__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_9_2__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_9_2__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_9_2__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_9_3__din),
    .fifo_A_out_full_n(fifo_A_PE_9_3__full_n),
    .fifo_A_out_write(fifo_A_PE_9_3__write),
    .fifo_B_out_din(fifo_B_PE_10_2__din),
    .fifo_B_out_full_n(fifo_B_PE_10_2__full_n),
    .fifo_B_out_write(fifo_B_PE_10_2__write),
    .fifo_B_in_s_dout(fifo_B_PE_9_2__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_9_2__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_9_2__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_9_2__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_9_2__read),
    .fifo_B_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_PE_9_2__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_9_2__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_9_2__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_156
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_156__ap_start),
    .ap_done(PE_wrapper_156__ap_done),
    .ap_idle(PE_wrapper_156__ap_idle),
    .ap_ready(PE_wrapper_156__ap_ready),
    .idy(64'd3),
    .idx(64'd9),
    .fifo_A_in_s_dout(fifo_A_PE_9_3__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_9_3__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_9_3__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_9_3__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_9_3__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_9_4__din),
    .fifo_A_out_full_n(fifo_A_PE_9_4__full_n),
    .fifo_A_out_write(fifo_A_PE_9_4__write),
    .fifo_B_out_din(fifo_B_PE_10_3__din),
    .fifo_B_out_full_n(fifo_B_PE_10_3__full_n),
    .fifo_B_out_write(fifo_B_PE_10_3__write),
    .fifo_B_in_s_dout(fifo_B_PE_9_3__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_9_3__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_9_3__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_9_3__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_9_3__read),
    .fifo_B_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_PE_9_3__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_9_3__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_9_3__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_157
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_157__ap_start),
    .ap_done(PE_wrapper_157__ap_done),
    .ap_idle(PE_wrapper_157__ap_idle),
    .ap_ready(PE_wrapper_157__ap_ready),
    .idy(64'd4),
    .idx(64'd9),
    .fifo_A_in_s_dout(fifo_A_PE_9_4__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_9_4__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_9_4__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_9_4__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_9_4__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_9_5__din),
    .fifo_A_out_full_n(fifo_A_PE_9_5__full_n),
    .fifo_A_out_write(fifo_A_PE_9_5__write),
    .fifo_B_out_din(fifo_B_PE_10_4__din),
    .fifo_B_out_full_n(fifo_B_PE_10_4__full_n),
    .fifo_B_out_write(fifo_B_PE_10_4__write),
    .fifo_B_in_s_dout(fifo_B_PE_9_4__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_9_4__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_9_4__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_9_4__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_9_4__read),
    .fifo_B_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_PE_9_4__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_9_4__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_9_4__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_158
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_158__ap_start),
    .ap_done(PE_wrapper_158__ap_done),
    .ap_idle(PE_wrapper_158__ap_idle),
    .ap_ready(PE_wrapper_158__ap_ready),
    .idy(64'd5),
    .idx(64'd9),
    .fifo_A_in_s_dout(fifo_A_PE_9_5__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_9_5__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_9_5__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_9_5__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_9_5__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_9_6__din),
    .fifo_A_out_full_n(fifo_A_PE_9_6__full_n),
    .fifo_A_out_write(fifo_A_PE_9_6__write),
    .fifo_B_out_din(fifo_B_PE_10_5__din),
    .fifo_B_out_full_n(fifo_B_PE_10_5__full_n),
    .fifo_B_out_write(fifo_B_PE_10_5__write),
    .fifo_B_in_s_dout(fifo_B_PE_9_5__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_9_5__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_9_5__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_9_5__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_9_5__read),
    .fifo_B_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_PE_9_5__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_9_5__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_9_5__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_159
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_159__ap_start),
    .ap_done(PE_wrapper_159__ap_done),
    .ap_idle(PE_wrapper_159__ap_idle),
    .ap_ready(PE_wrapper_159__ap_ready),
    .idy(64'd6),
    .idx(64'd9),
    .fifo_A_in_s_dout(fifo_A_PE_9_6__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_9_6__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_9_6__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_9_6__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_9_6__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_9_7__din),
    .fifo_A_out_full_n(fifo_A_PE_9_7__full_n),
    .fifo_A_out_write(fifo_A_PE_9_7__write),
    .fifo_B_out_din(fifo_B_PE_10_6__din),
    .fifo_B_out_full_n(fifo_B_PE_10_6__full_n),
    .fifo_B_out_write(fifo_B_PE_10_6__write),
    .fifo_B_in_s_dout(fifo_B_PE_9_6__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_9_6__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_9_6__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_9_6__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_9_6__read),
    .fifo_B_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_PE_9_6__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_9_6__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_9_6__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_160
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_160__ap_start),
    .ap_done(PE_wrapper_160__ap_done),
    .ap_idle(PE_wrapper_160__ap_idle),
    .ap_ready(PE_wrapper_160__ap_ready),
    .idy(64'd7),
    .idx(64'd9),
    .fifo_A_in_s_dout(fifo_A_PE_9_7__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_9_7__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_9_7__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_9_7__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_9_7__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_9_8__din),
    .fifo_A_out_full_n(fifo_A_PE_9_8__full_n),
    .fifo_A_out_write(fifo_A_PE_9_8__write),
    .fifo_B_out_din(fifo_B_PE_10_7__din),
    .fifo_B_out_full_n(fifo_B_PE_10_7__full_n),
    .fifo_B_out_write(fifo_B_PE_10_7__write),
    .fifo_B_in_s_dout(fifo_B_PE_9_7__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_9_7__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_9_7__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_9_7__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_9_7__read),
    .fifo_B_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_PE_9_7__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_9_7__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_9_7__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_161
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_161__ap_start),
    .ap_done(PE_wrapper_161__ap_done),
    .ap_idle(PE_wrapper_161__ap_idle),
    .ap_ready(PE_wrapper_161__ap_ready),
    .idy(64'd8),
    .idx(64'd9),
    .fifo_A_in_s_dout(fifo_A_PE_9_8__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_9_8__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_9_8__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_9_8__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_9_8__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_9_9__din),
    .fifo_A_out_full_n(fifo_A_PE_9_9__full_n),
    .fifo_A_out_write(fifo_A_PE_9_9__write),
    .fifo_B_out_din(fifo_B_PE_10_8__din),
    .fifo_B_out_full_n(fifo_B_PE_10_8__full_n),
    .fifo_B_out_write(fifo_B_PE_10_8__write),
    .fifo_B_in_s_dout(fifo_B_PE_9_8__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_9_8__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_9_8__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_9_8__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_9_8__read),
    .fifo_B_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_PE_9_8__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_9_8__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_9_8__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_162
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_162__ap_start),
    .ap_done(PE_wrapper_162__ap_done),
    .ap_idle(PE_wrapper_162__ap_idle),
    .ap_ready(PE_wrapper_162__ap_ready),
    .idx(64'd9),
    .idy(64'd9),
    .fifo_A_out_din(fifo_A_PE_9_10__din),
    .fifo_A_out_full_n(fifo_A_PE_9_10__full_n),
    .fifo_A_out_write(fifo_A_PE_9_10__write),
    .fifo_A_in_s_dout(fifo_A_PE_9_9__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_9_9__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_9_9__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_9_9__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_9_9__read),
    .fifo_A_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_10_9__din),
    .fifo_B_out_full_n(fifo_B_PE_10_9__full_n),
    .fifo_B_out_write(fifo_B_PE_10_9__write),
    .fifo_B_in_s_dout(fifo_B_PE_9_9__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_9_9__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_9_9__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_9_9__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_9_9__read),
    .fifo_B_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_PE_9_9__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_9_9__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_9_9__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_163
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_163__ap_start),
    .ap_done(PE_wrapper_163__ap_done),
    .ap_idle(PE_wrapper_163__ap_idle),
    .ap_ready(PE_wrapper_163__ap_ready),
    .idy(64'd10),
    .idx(64'd9),
    .fifo_A_in_s_dout(fifo_A_PE_9_10__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_9_10__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_9_10__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_9_10__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_9_10__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_9_11__din),
    .fifo_A_out_full_n(fifo_A_PE_9_11__full_n),
    .fifo_A_out_write(fifo_A_PE_9_11__write),
    .fifo_B_out_din(fifo_B_PE_10_10__din),
    .fifo_B_out_full_n(fifo_B_PE_10_10__full_n),
    .fifo_B_out_write(fifo_B_PE_10_10__write),
    .fifo_B_in_s_dout(fifo_B_PE_9_10__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_9_10__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_9_10__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_9_10__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_9_10__read),
    .fifo_B_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_PE_9_10__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_9_10__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_9_10__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_164
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_164__ap_start),
    .ap_done(PE_wrapper_164__ap_done),
    .ap_idle(PE_wrapper_164__ap_idle),
    .ap_ready(PE_wrapper_164__ap_ready),
    .idy(64'd11),
    .idx(64'd9),
    .fifo_A_in_s_dout(fifo_A_PE_9_11__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_9_11__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_9_11__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_9_11__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_9_11__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_9_12__din),
    .fifo_A_out_full_n(fifo_A_PE_9_12__full_n),
    .fifo_A_out_write(fifo_A_PE_9_12__write),
    .fifo_B_out_din(fifo_B_PE_10_11__din),
    .fifo_B_out_full_n(fifo_B_PE_10_11__full_n),
    .fifo_B_out_write(fifo_B_PE_10_11__write),
    .fifo_B_in_s_dout(fifo_B_PE_9_11__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_9_11__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_9_11__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_9_11__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_9_11__read),
    .fifo_B_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_PE_9_11__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_9_11__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_9_11__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_165
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_165__ap_start),
    .ap_done(PE_wrapper_165__ap_done),
    .ap_idle(PE_wrapper_165__ap_idle),
    .ap_ready(PE_wrapper_165__ap_ready),
    .idy(64'd12),
    .idx(64'd9),
    .fifo_A_in_s_dout(fifo_A_PE_9_12__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_9_12__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_9_12__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_9_12__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_9_12__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_9_13__din),
    .fifo_A_out_full_n(fifo_A_PE_9_13__full_n),
    .fifo_A_out_write(fifo_A_PE_9_13__write),
    .fifo_B_out_din(fifo_B_PE_10_12__din),
    .fifo_B_out_full_n(fifo_B_PE_10_12__full_n),
    .fifo_B_out_write(fifo_B_PE_10_12__write),
    .fifo_B_in_s_dout(fifo_B_PE_9_12__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_9_12__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_9_12__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_9_12__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_9_12__read),
    .fifo_B_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_PE_9_12__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_9_12__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_9_12__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_166
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_166__ap_start),
    .ap_done(PE_wrapper_166__ap_done),
    .ap_idle(PE_wrapper_166__ap_idle),
    .ap_ready(PE_wrapper_166__ap_ready),
    .idy(64'd13),
    .idx(64'd9),
    .fifo_A_in_s_dout(fifo_A_PE_9_13__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_9_13__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_9_13__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_9_13__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_9_13__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_9_14__din),
    .fifo_A_out_full_n(fifo_A_PE_9_14__full_n),
    .fifo_A_out_write(fifo_A_PE_9_14__write),
    .fifo_B_out_din(fifo_B_PE_10_13__din),
    .fifo_B_out_full_n(fifo_B_PE_10_13__full_n),
    .fifo_B_out_write(fifo_B_PE_10_13__write),
    .fifo_B_in_s_dout(fifo_B_PE_9_13__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_9_13__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_9_13__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_9_13__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_9_13__read),
    .fifo_B_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_PE_9_13__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_9_13__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_9_13__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_167
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_167__ap_start),
    .ap_done(PE_wrapper_167__ap_done),
    .ap_idle(PE_wrapper_167__ap_idle),
    .ap_ready(PE_wrapper_167__ap_ready),
    .idy(64'd14),
    .idx(64'd9),
    .fifo_A_in_s_dout(fifo_A_PE_9_14__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_9_14__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_9_14__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_9_14__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_9_14__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_9_15__din),
    .fifo_A_out_full_n(fifo_A_PE_9_15__full_n),
    .fifo_A_out_write(fifo_A_PE_9_15__write),
    .fifo_B_out_din(fifo_B_PE_10_14__din),
    .fifo_B_out_full_n(fifo_B_PE_10_14__full_n),
    .fifo_B_out_write(fifo_B_PE_10_14__write),
    .fifo_B_in_s_dout(fifo_B_PE_9_14__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_9_14__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_9_14__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_9_14__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_9_14__read),
    .fifo_B_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_PE_9_14__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_9_14__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_9_14__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_168
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_168__ap_start),
    .ap_done(PE_wrapper_168__ap_done),
    .ap_idle(PE_wrapper_168__ap_idle),
    .ap_ready(PE_wrapper_168__ap_ready),
    .idy(64'd15),
    .idx(64'd9),
    .fifo_A_in_s_dout(fifo_A_PE_9_15__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_9_15__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_9_15__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_9_15__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_9_15__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_9_16__din),
    .fifo_A_out_full_n(fifo_A_PE_9_16__full_n),
    .fifo_A_out_write(fifo_A_PE_9_16__write),
    .fifo_B_out_din(fifo_B_PE_10_15__din),
    .fifo_B_out_full_n(fifo_B_PE_10_15__full_n),
    .fifo_B_out_write(fifo_B_PE_10_15__write),
    .fifo_B_in_s_dout(fifo_B_PE_9_15__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_9_15__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_9_15__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_9_15__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_9_15__read),
    .fifo_B_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_PE_9_15__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_9_15__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_9_15__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_169
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_169__ap_start),
    .ap_done(PE_wrapper_169__ap_done),
    .ap_idle(PE_wrapper_169__ap_idle),
    .ap_ready(PE_wrapper_169__ap_ready),
    .idy(64'd16),
    .idx(64'd9),
    .fifo_A_in_s_dout(fifo_A_PE_9_16__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_9_16__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_9_16__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_9_16__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_9_16__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_9_17__din),
    .fifo_A_out_full_n(fifo_A_PE_9_17__full_n),
    .fifo_A_out_write(fifo_A_PE_9_17__write),
    .fifo_B_out_din(fifo_B_PE_10_16__din),
    .fifo_B_out_full_n(fifo_B_PE_10_16__full_n),
    .fifo_B_out_write(fifo_B_PE_10_16__write),
    .fifo_B_in_s_dout(fifo_B_PE_9_16__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_9_16__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_9_16__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_9_16__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_9_16__read),
    .fifo_B_in_peek_read(),
    .fifo_C_drain_out_din(fifo_C_drain_PE_9_16__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_9_16__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_9_16__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_170
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_170__ap_start),
    .ap_done(PE_wrapper_170__ap_done),
    .ap_idle(PE_wrapper_170__ap_idle),
    .ap_ready(PE_wrapper_170__ap_ready),
    .idy(64'd0),
    .idx(64'd10),
    .fifo_A_in_s_dout(fifo_A_PE_10_0__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_10_0__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_10_0__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_10_0__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_10_0__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_10_1__din),
    .fifo_A_out_full_n(fifo_A_PE_10_1__full_n),
    .fifo_A_out_write(fifo_A_PE_10_1__write),
    .fifo_B_in_s_dout(fifo_B_PE_10_0__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_10_0__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_10_0__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_10_0__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_10_0__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_11_0__din),
    .fifo_B_out_full_n(fifo_B_PE_11_0__full_n),
    .fifo_B_out_write(fifo_B_PE_11_0__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_10_0__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_10_0__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_10_0__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_171
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_171__ap_start),
    .ap_done(PE_wrapper_171__ap_done),
    .ap_idle(PE_wrapper_171__ap_idle),
    .ap_ready(PE_wrapper_171__ap_ready),
    .idy(64'd1),
    .idx(64'd10),
    .fifo_A_in_s_dout(fifo_A_PE_10_1__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_10_1__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_10_1__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_10_1__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_10_1__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_10_2__din),
    .fifo_A_out_full_n(fifo_A_PE_10_2__full_n),
    .fifo_A_out_write(fifo_A_PE_10_2__write),
    .fifo_B_in_s_dout(fifo_B_PE_10_1__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_10_1__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_10_1__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_10_1__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_10_1__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_11_1__din),
    .fifo_B_out_full_n(fifo_B_PE_11_1__full_n),
    .fifo_B_out_write(fifo_B_PE_11_1__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_10_1__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_10_1__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_10_1__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_172
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_172__ap_start),
    .ap_done(PE_wrapper_172__ap_done),
    .ap_idle(PE_wrapper_172__ap_idle),
    .ap_ready(PE_wrapper_172__ap_ready),
    .idx(64'd10),
    .idy(64'd2),
    .fifo_A_in_s_dout(fifo_A_PE_10_2__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_10_2__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_10_2__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_10_2__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_10_2__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_10_3__din),
    .fifo_A_out_full_n(fifo_A_PE_10_3__full_n),
    .fifo_A_out_write(fifo_A_PE_10_3__write),
    .fifo_B_in_s_dout(fifo_B_PE_10_2__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_10_2__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_10_2__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_10_2__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_10_2__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_11_2__din),
    .fifo_B_out_full_n(fifo_B_PE_11_2__full_n),
    .fifo_B_out_write(fifo_B_PE_11_2__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_10_2__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_10_2__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_10_2__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_173
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_173__ap_start),
    .ap_done(PE_wrapper_173__ap_done),
    .ap_idle(PE_wrapper_173__ap_idle),
    .ap_ready(PE_wrapper_173__ap_ready),
    .idx(64'd10),
    .idy(64'd3),
    .fifo_A_in_s_dout(fifo_A_PE_10_3__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_10_3__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_10_3__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_10_3__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_10_3__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_10_4__din),
    .fifo_A_out_full_n(fifo_A_PE_10_4__full_n),
    .fifo_A_out_write(fifo_A_PE_10_4__write),
    .fifo_B_in_s_dout(fifo_B_PE_10_3__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_10_3__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_10_3__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_10_3__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_10_3__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_11_3__din),
    .fifo_B_out_full_n(fifo_B_PE_11_3__full_n),
    .fifo_B_out_write(fifo_B_PE_11_3__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_10_3__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_10_3__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_10_3__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_174
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_174__ap_start),
    .ap_done(PE_wrapper_174__ap_done),
    .ap_idle(PE_wrapper_174__ap_idle),
    .ap_ready(PE_wrapper_174__ap_ready),
    .idx(64'd10),
    .idy(64'd4),
    .fifo_A_in_s_dout(fifo_A_PE_10_4__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_10_4__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_10_4__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_10_4__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_10_4__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_10_5__din),
    .fifo_A_out_full_n(fifo_A_PE_10_5__full_n),
    .fifo_A_out_write(fifo_A_PE_10_5__write),
    .fifo_B_in_s_dout(fifo_B_PE_10_4__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_10_4__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_10_4__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_10_4__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_10_4__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_11_4__din),
    .fifo_B_out_full_n(fifo_B_PE_11_4__full_n),
    .fifo_B_out_write(fifo_B_PE_11_4__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_10_4__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_10_4__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_10_4__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_175
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_175__ap_start),
    .ap_done(PE_wrapper_175__ap_done),
    .ap_idle(PE_wrapper_175__ap_idle),
    .ap_ready(PE_wrapper_175__ap_ready),
    .idx(64'd10),
    .idy(64'd5),
    .fifo_A_in_s_dout(fifo_A_PE_10_5__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_10_5__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_10_5__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_10_5__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_10_5__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_10_6__din),
    .fifo_A_out_full_n(fifo_A_PE_10_6__full_n),
    .fifo_A_out_write(fifo_A_PE_10_6__write),
    .fifo_B_in_s_dout(fifo_B_PE_10_5__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_10_5__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_10_5__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_10_5__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_10_5__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_11_5__din),
    .fifo_B_out_full_n(fifo_B_PE_11_5__full_n),
    .fifo_B_out_write(fifo_B_PE_11_5__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_10_5__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_10_5__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_10_5__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_176
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_176__ap_start),
    .ap_done(PE_wrapper_176__ap_done),
    .ap_idle(PE_wrapper_176__ap_idle),
    .ap_ready(PE_wrapper_176__ap_ready),
    .idx(64'd10),
    .idy(64'd6),
    .fifo_A_in_s_dout(fifo_A_PE_10_6__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_10_6__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_10_6__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_10_6__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_10_6__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_10_7__din),
    .fifo_A_out_full_n(fifo_A_PE_10_7__full_n),
    .fifo_A_out_write(fifo_A_PE_10_7__write),
    .fifo_B_in_s_dout(fifo_B_PE_10_6__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_10_6__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_10_6__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_10_6__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_10_6__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_11_6__din),
    .fifo_B_out_full_n(fifo_B_PE_11_6__full_n),
    .fifo_B_out_write(fifo_B_PE_11_6__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_10_6__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_10_6__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_10_6__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_177
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_177__ap_start),
    .ap_done(PE_wrapper_177__ap_done),
    .ap_idle(PE_wrapper_177__ap_idle),
    .ap_ready(PE_wrapper_177__ap_ready),
    .idx(64'd10),
    .idy(64'd7),
    .fifo_A_in_s_dout(fifo_A_PE_10_7__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_10_7__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_10_7__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_10_7__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_10_7__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_10_8__din),
    .fifo_A_out_full_n(fifo_A_PE_10_8__full_n),
    .fifo_A_out_write(fifo_A_PE_10_8__write),
    .fifo_B_in_s_dout(fifo_B_PE_10_7__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_10_7__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_10_7__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_10_7__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_10_7__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_11_7__din),
    .fifo_B_out_full_n(fifo_B_PE_11_7__full_n),
    .fifo_B_out_write(fifo_B_PE_11_7__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_10_7__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_10_7__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_10_7__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_178
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_178__ap_start),
    .ap_done(PE_wrapper_178__ap_done),
    .ap_idle(PE_wrapper_178__ap_idle),
    .ap_ready(PE_wrapper_178__ap_ready),
    .idx(64'd10),
    .idy(64'd8),
    .fifo_A_in_s_dout(fifo_A_PE_10_8__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_10_8__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_10_8__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_10_8__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_10_8__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_10_9__din),
    .fifo_A_out_full_n(fifo_A_PE_10_9__full_n),
    .fifo_A_out_write(fifo_A_PE_10_9__write),
    .fifo_B_in_s_dout(fifo_B_PE_10_8__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_10_8__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_10_8__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_10_8__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_10_8__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_11_8__din),
    .fifo_B_out_full_n(fifo_B_PE_11_8__full_n),
    .fifo_B_out_write(fifo_B_PE_11_8__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_10_8__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_10_8__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_10_8__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_179
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_179__ap_start),
    .ap_done(PE_wrapper_179__ap_done),
    .ap_idle(PE_wrapper_179__ap_idle),
    .ap_ready(PE_wrapper_179__ap_ready),
    .idx(64'd10),
    .idy(64'd9),
    .fifo_A_out_din(fifo_A_PE_10_10__din),
    .fifo_A_out_full_n(fifo_A_PE_10_10__full_n),
    .fifo_A_out_write(fifo_A_PE_10_10__write),
    .fifo_A_in_s_dout(fifo_A_PE_10_9__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_10_9__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_10_9__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_10_9__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_10_9__read),
    .fifo_A_in_peek_read(),
    .fifo_B_in_s_dout(fifo_B_PE_10_9__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_10_9__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_10_9__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_10_9__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_10_9__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_11_9__din),
    .fifo_B_out_full_n(fifo_B_PE_11_9__full_n),
    .fifo_B_out_write(fifo_B_PE_11_9__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_10_9__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_10_9__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_10_9__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_180
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_180__ap_start),
    .ap_done(PE_wrapper_180__ap_done),
    .ap_idle(PE_wrapper_180__ap_idle),
    .ap_ready(PE_wrapper_180__ap_ready),
    .idx(64'd10),
    .idy(64'd10),
    .fifo_A_in_s_dout(fifo_A_PE_10_10__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_10_10__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_10_10__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_10_10__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_10_10__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_10_11__din),
    .fifo_A_out_full_n(fifo_A_PE_10_11__full_n),
    .fifo_A_out_write(fifo_A_PE_10_11__write),
    .fifo_B_in_s_dout(fifo_B_PE_10_10__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_10_10__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_10_10__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_10_10__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_10_10__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_11_10__din),
    .fifo_B_out_full_n(fifo_B_PE_11_10__full_n),
    .fifo_B_out_write(fifo_B_PE_11_10__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_10_10__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_10_10__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_10_10__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_181
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_181__ap_start),
    .ap_done(PE_wrapper_181__ap_done),
    .ap_idle(PE_wrapper_181__ap_idle),
    .ap_ready(PE_wrapper_181__ap_ready),
    .idx(64'd10),
    .idy(64'd11),
    .fifo_A_in_s_dout(fifo_A_PE_10_11__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_10_11__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_10_11__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_10_11__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_10_11__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_10_12__din),
    .fifo_A_out_full_n(fifo_A_PE_10_12__full_n),
    .fifo_A_out_write(fifo_A_PE_10_12__write),
    .fifo_B_in_s_dout(fifo_B_PE_10_11__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_10_11__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_10_11__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_10_11__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_10_11__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_11_11__din),
    .fifo_B_out_full_n(fifo_B_PE_11_11__full_n),
    .fifo_B_out_write(fifo_B_PE_11_11__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_10_11__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_10_11__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_10_11__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_182
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_182__ap_start),
    .ap_done(PE_wrapper_182__ap_done),
    .ap_idle(PE_wrapper_182__ap_idle),
    .ap_ready(PE_wrapper_182__ap_ready),
    .idx(64'd10),
    .idy(64'd12),
    .fifo_A_in_s_dout(fifo_A_PE_10_12__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_10_12__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_10_12__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_10_12__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_10_12__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_10_13__din),
    .fifo_A_out_full_n(fifo_A_PE_10_13__full_n),
    .fifo_A_out_write(fifo_A_PE_10_13__write),
    .fifo_B_in_s_dout(fifo_B_PE_10_12__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_10_12__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_10_12__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_10_12__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_10_12__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_11_12__din),
    .fifo_B_out_full_n(fifo_B_PE_11_12__full_n),
    .fifo_B_out_write(fifo_B_PE_11_12__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_10_12__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_10_12__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_10_12__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_183
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_183__ap_start),
    .ap_done(PE_wrapper_183__ap_done),
    .ap_idle(PE_wrapper_183__ap_idle),
    .ap_ready(PE_wrapper_183__ap_ready),
    .idx(64'd10),
    .idy(64'd13),
    .fifo_A_in_s_dout(fifo_A_PE_10_13__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_10_13__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_10_13__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_10_13__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_10_13__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_10_14__din),
    .fifo_A_out_full_n(fifo_A_PE_10_14__full_n),
    .fifo_A_out_write(fifo_A_PE_10_14__write),
    .fifo_B_in_s_dout(fifo_B_PE_10_13__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_10_13__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_10_13__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_10_13__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_10_13__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_11_13__din),
    .fifo_B_out_full_n(fifo_B_PE_11_13__full_n),
    .fifo_B_out_write(fifo_B_PE_11_13__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_10_13__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_10_13__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_10_13__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_184
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_184__ap_start),
    .ap_done(PE_wrapper_184__ap_done),
    .ap_idle(PE_wrapper_184__ap_idle),
    .ap_ready(PE_wrapper_184__ap_ready),
    .idx(64'd10),
    .idy(64'd14),
    .fifo_A_in_s_dout(fifo_A_PE_10_14__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_10_14__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_10_14__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_10_14__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_10_14__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_10_15__din),
    .fifo_A_out_full_n(fifo_A_PE_10_15__full_n),
    .fifo_A_out_write(fifo_A_PE_10_15__write),
    .fifo_B_in_s_dout(fifo_B_PE_10_14__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_10_14__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_10_14__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_10_14__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_10_14__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_11_14__din),
    .fifo_B_out_full_n(fifo_B_PE_11_14__full_n),
    .fifo_B_out_write(fifo_B_PE_11_14__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_10_14__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_10_14__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_10_14__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_185
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_185__ap_start),
    .ap_done(PE_wrapper_185__ap_done),
    .ap_idle(PE_wrapper_185__ap_idle),
    .ap_ready(PE_wrapper_185__ap_ready),
    .idx(64'd10),
    .idy(64'd15),
    .fifo_A_in_s_dout(fifo_A_PE_10_15__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_10_15__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_10_15__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_10_15__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_10_15__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_10_16__din),
    .fifo_A_out_full_n(fifo_A_PE_10_16__full_n),
    .fifo_A_out_write(fifo_A_PE_10_16__write),
    .fifo_B_in_s_dout(fifo_B_PE_10_15__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_10_15__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_10_15__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_10_15__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_10_15__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_11_15__din),
    .fifo_B_out_full_n(fifo_B_PE_11_15__full_n),
    .fifo_B_out_write(fifo_B_PE_11_15__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_10_15__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_10_15__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_10_15__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_186
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_186__ap_start),
    .ap_done(PE_wrapper_186__ap_done),
    .ap_idle(PE_wrapper_186__ap_idle),
    .ap_ready(PE_wrapper_186__ap_ready),
    .idx(64'd10),
    .idy(64'd16),
    .fifo_A_in_s_dout(fifo_A_PE_10_16__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_10_16__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_10_16__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_10_16__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_10_16__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_10_17__din),
    .fifo_A_out_full_n(fifo_A_PE_10_17__full_n),
    .fifo_A_out_write(fifo_A_PE_10_17__write),
    .fifo_B_in_s_dout(fifo_B_PE_10_16__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_10_16__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_10_16__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_10_16__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_10_16__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_11_16__din),
    .fifo_B_out_full_n(fifo_B_PE_11_16__full_n),
    .fifo_B_out_write(fifo_B_PE_11_16__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_10_16__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_10_16__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_10_16__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_187
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_187__ap_start),
    .ap_done(PE_wrapper_187__ap_done),
    .ap_idle(PE_wrapper_187__ap_idle),
    .ap_ready(PE_wrapper_187__ap_ready),
    .idy(64'd0),
    .idx(64'd11),
    .fifo_A_in_s_dout(fifo_A_PE_11_0__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_11_0__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_11_0__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_11_0__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_11_0__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_11_1__din),
    .fifo_A_out_full_n(fifo_A_PE_11_1__full_n),
    .fifo_A_out_write(fifo_A_PE_11_1__write),
    .fifo_B_in_s_dout(fifo_B_PE_11_0__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_11_0__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_11_0__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_11_0__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_11_0__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_12_0__din),
    .fifo_B_out_full_n(fifo_B_PE_12_0__full_n),
    .fifo_B_out_write(fifo_B_PE_12_0__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_11_0__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_11_0__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_11_0__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_188
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_188__ap_start),
    .ap_done(PE_wrapper_188__ap_done),
    .ap_idle(PE_wrapper_188__ap_idle),
    .ap_ready(PE_wrapper_188__ap_ready),
    .idy(64'd1),
    .idx(64'd11),
    .fifo_A_in_s_dout(fifo_A_PE_11_1__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_11_1__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_11_1__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_11_1__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_11_1__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_11_2__din),
    .fifo_A_out_full_n(fifo_A_PE_11_2__full_n),
    .fifo_A_out_write(fifo_A_PE_11_2__write),
    .fifo_B_in_s_dout(fifo_B_PE_11_1__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_11_1__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_11_1__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_11_1__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_11_1__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_12_1__din),
    .fifo_B_out_full_n(fifo_B_PE_12_1__full_n),
    .fifo_B_out_write(fifo_B_PE_12_1__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_11_1__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_11_1__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_11_1__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_189
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_189__ap_start),
    .ap_done(PE_wrapper_189__ap_done),
    .ap_idle(PE_wrapper_189__ap_idle),
    .ap_ready(PE_wrapper_189__ap_ready),
    .idx(64'd11),
    .idy(64'd2),
    .fifo_A_in_s_dout(fifo_A_PE_11_2__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_11_2__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_11_2__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_11_2__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_11_2__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_11_3__din),
    .fifo_A_out_full_n(fifo_A_PE_11_3__full_n),
    .fifo_A_out_write(fifo_A_PE_11_3__write),
    .fifo_B_in_s_dout(fifo_B_PE_11_2__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_11_2__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_11_2__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_11_2__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_11_2__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_12_2__din),
    .fifo_B_out_full_n(fifo_B_PE_12_2__full_n),
    .fifo_B_out_write(fifo_B_PE_12_2__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_11_2__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_11_2__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_11_2__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_190
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_190__ap_start),
    .ap_done(PE_wrapper_190__ap_done),
    .ap_idle(PE_wrapper_190__ap_idle),
    .ap_ready(PE_wrapper_190__ap_ready),
    .idx(64'd11),
    .idy(64'd3),
    .fifo_A_in_s_dout(fifo_A_PE_11_3__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_11_3__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_11_3__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_11_3__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_11_3__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_11_4__din),
    .fifo_A_out_full_n(fifo_A_PE_11_4__full_n),
    .fifo_A_out_write(fifo_A_PE_11_4__write),
    .fifo_B_in_s_dout(fifo_B_PE_11_3__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_11_3__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_11_3__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_11_3__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_11_3__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_12_3__din),
    .fifo_B_out_full_n(fifo_B_PE_12_3__full_n),
    .fifo_B_out_write(fifo_B_PE_12_3__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_11_3__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_11_3__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_11_3__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_191
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_191__ap_start),
    .ap_done(PE_wrapper_191__ap_done),
    .ap_idle(PE_wrapper_191__ap_idle),
    .ap_ready(PE_wrapper_191__ap_ready),
    .idx(64'd11),
    .idy(64'd4),
    .fifo_A_in_s_dout(fifo_A_PE_11_4__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_11_4__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_11_4__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_11_4__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_11_4__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_11_5__din),
    .fifo_A_out_full_n(fifo_A_PE_11_5__full_n),
    .fifo_A_out_write(fifo_A_PE_11_5__write),
    .fifo_B_in_s_dout(fifo_B_PE_11_4__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_11_4__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_11_4__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_11_4__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_11_4__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_12_4__din),
    .fifo_B_out_full_n(fifo_B_PE_12_4__full_n),
    .fifo_B_out_write(fifo_B_PE_12_4__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_11_4__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_11_4__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_11_4__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_192
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_192__ap_start),
    .ap_done(PE_wrapper_192__ap_done),
    .ap_idle(PE_wrapper_192__ap_idle),
    .ap_ready(PE_wrapper_192__ap_ready),
    .idx(64'd11),
    .idy(64'd5),
    .fifo_A_in_s_dout(fifo_A_PE_11_5__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_11_5__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_11_5__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_11_5__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_11_5__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_11_6__din),
    .fifo_A_out_full_n(fifo_A_PE_11_6__full_n),
    .fifo_A_out_write(fifo_A_PE_11_6__write),
    .fifo_B_in_s_dout(fifo_B_PE_11_5__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_11_5__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_11_5__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_11_5__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_11_5__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_12_5__din),
    .fifo_B_out_full_n(fifo_B_PE_12_5__full_n),
    .fifo_B_out_write(fifo_B_PE_12_5__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_11_5__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_11_5__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_11_5__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_193
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_193__ap_start),
    .ap_done(PE_wrapper_193__ap_done),
    .ap_idle(PE_wrapper_193__ap_idle),
    .ap_ready(PE_wrapper_193__ap_ready),
    .idx(64'd11),
    .idy(64'd6),
    .fifo_A_in_s_dout(fifo_A_PE_11_6__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_11_6__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_11_6__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_11_6__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_11_6__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_11_7__din),
    .fifo_A_out_full_n(fifo_A_PE_11_7__full_n),
    .fifo_A_out_write(fifo_A_PE_11_7__write),
    .fifo_B_in_s_dout(fifo_B_PE_11_6__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_11_6__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_11_6__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_11_6__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_11_6__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_12_6__din),
    .fifo_B_out_full_n(fifo_B_PE_12_6__full_n),
    .fifo_B_out_write(fifo_B_PE_12_6__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_11_6__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_11_6__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_11_6__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_194
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_194__ap_start),
    .ap_done(PE_wrapper_194__ap_done),
    .ap_idle(PE_wrapper_194__ap_idle),
    .ap_ready(PE_wrapper_194__ap_ready),
    .idx(64'd11),
    .idy(64'd7),
    .fifo_A_in_s_dout(fifo_A_PE_11_7__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_11_7__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_11_7__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_11_7__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_11_7__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_11_8__din),
    .fifo_A_out_full_n(fifo_A_PE_11_8__full_n),
    .fifo_A_out_write(fifo_A_PE_11_8__write),
    .fifo_B_in_s_dout(fifo_B_PE_11_7__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_11_7__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_11_7__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_11_7__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_11_7__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_12_7__din),
    .fifo_B_out_full_n(fifo_B_PE_12_7__full_n),
    .fifo_B_out_write(fifo_B_PE_12_7__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_11_7__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_11_7__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_11_7__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_195
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_195__ap_start),
    .ap_done(PE_wrapper_195__ap_done),
    .ap_idle(PE_wrapper_195__ap_idle),
    .ap_ready(PE_wrapper_195__ap_ready),
    .idx(64'd11),
    .idy(64'd8),
    .fifo_A_in_s_dout(fifo_A_PE_11_8__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_11_8__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_11_8__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_11_8__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_11_8__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_11_9__din),
    .fifo_A_out_full_n(fifo_A_PE_11_9__full_n),
    .fifo_A_out_write(fifo_A_PE_11_9__write),
    .fifo_B_in_s_dout(fifo_B_PE_11_8__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_11_8__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_11_8__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_11_8__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_11_8__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_12_8__din),
    .fifo_B_out_full_n(fifo_B_PE_12_8__full_n),
    .fifo_B_out_write(fifo_B_PE_12_8__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_11_8__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_11_8__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_11_8__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_196
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_196__ap_start),
    .ap_done(PE_wrapper_196__ap_done),
    .ap_idle(PE_wrapper_196__ap_idle),
    .ap_ready(PE_wrapper_196__ap_ready),
    .idx(64'd11),
    .idy(64'd9),
    .fifo_A_out_din(fifo_A_PE_11_10__din),
    .fifo_A_out_full_n(fifo_A_PE_11_10__full_n),
    .fifo_A_out_write(fifo_A_PE_11_10__write),
    .fifo_A_in_s_dout(fifo_A_PE_11_9__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_11_9__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_11_9__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_11_9__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_11_9__read),
    .fifo_A_in_peek_read(),
    .fifo_B_in_s_dout(fifo_B_PE_11_9__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_11_9__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_11_9__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_11_9__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_11_9__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_12_9__din),
    .fifo_B_out_full_n(fifo_B_PE_12_9__full_n),
    .fifo_B_out_write(fifo_B_PE_12_9__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_11_9__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_11_9__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_11_9__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_197
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_197__ap_start),
    .ap_done(PE_wrapper_197__ap_done),
    .ap_idle(PE_wrapper_197__ap_idle),
    .ap_ready(PE_wrapper_197__ap_ready),
    .idy(64'd10),
    .idx(64'd11),
    .fifo_A_in_s_dout(fifo_A_PE_11_10__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_11_10__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_11_10__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_11_10__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_11_10__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_11_11__din),
    .fifo_A_out_full_n(fifo_A_PE_11_11__full_n),
    .fifo_A_out_write(fifo_A_PE_11_11__write),
    .fifo_B_in_s_dout(fifo_B_PE_11_10__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_11_10__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_11_10__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_11_10__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_11_10__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_12_10__din),
    .fifo_B_out_full_n(fifo_B_PE_12_10__full_n),
    .fifo_B_out_write(fifo_B_PE_12_10__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_11_10__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_11_10__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_11_10__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_198
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_198__ap_start),
    .ap_done(PE_wrapper_198__ap_done),
    .ap_idle(PE_wrapper_198__ap_idle),
    .ap_ready(PE_wrapper_198__ap_ready),
    .idx(64'd11),
    .idy(64'd11),
    .fifo_A_in_s_dout(fifo_A_PE_11_11__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_11_11__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_11_11__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_11_11__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_11_11__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_11_12__din),
    .fifo_A_out_full_n(fifo_A_PE_11_12__full_n),
    .fifo_A_out_write(fifo_A_PE_11_12__write),
    .fifo_B_in_s_dout(fifo_B_PE_11_11__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_11_11__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_11_11__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_11_11__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_11_11__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_12_11__din),
    .fifo_B_out_full_n(fifo_B_PE_12_11__full_n),
    .fifo_B_out_write(fifo_B_PE_12_11__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_11_11__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_11_11__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_11_11__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_199
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_199__ap_start),
    .ap_done(PE_wrapper_199__ap_done),
    .ap_idle(PE_wrapper_199__ap_idle),
    .ap_ready(PE_wrapper_199__ap_ready),
    .idx(64'd11),
    .idy(64'd12),
    .fifo_A_in_s_dout(fifo_A_PE_11_12__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_11_12__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_11_12__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_11_12__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_11_12__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_11_13__din),
    .fifo_A_out_full_n(fifo_A_PE_11_13__full_n),
    .fifo_A_out_write(fifo_A_PE_11_13__write),
    .fifo_B_in_s_dout(fifo_B_PE_11_12__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_11_12__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_11_12__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_11_12__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_11_12__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_12_12__din),
    .fifo_B_out_full_n(fifo_B_PE_12_12__full_n),
    .fifo_B_out_write(fifo_B_PE_12_12__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_11_12__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_11_12__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_11_12__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_200
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_200__ap_start),
    .ap_done(PE_wrapper_200__ap_done),
    .ap_idle(PE_wrapper_200__ap_idle),
    .ap_ready(PE_wrapper_200__ap_ready),
    .idx(64'd11),
    .idy(64'd13),
    .fifo_A_in_s_dout(fifo_A_PE_11_13__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_11_13__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_11_13__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_11_13__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_11_13__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_11_14__din),
    .fifo_A_out_full_n(fifo_A_PE_11_14__full_n),
    .fifo_A_out_write(fifo_A_PE_11_14__write),
    .fifo_B_in_s_dout(fifo_B_PE_11_13__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_11_13__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_11_13__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_11_13__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_11_13__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_12_13__din),
    .fifo_B_out_full_n(fifo_B_PE_12_13__full_n),
    .fifo_B_out_write(fifo_B_PE_12_13__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_11_13__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_11_13__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_11_13__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_201
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_201__ap_start),
    .ap_done(PE_wrapper_201__ap_done),
    .ap_idle(PE_wrapper_201__ap_idle),
    .ap_ready(PE_wrapper_201__ap_ready),
    .idx(64'd11),
    .idy(64'd14),
    .fifo_A_in_s_dout(fifo_A_PE_11_14__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_11_14__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_11_14__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_11_14__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_11_14__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_11_15__din),
    .fifo_A_out_full_n(fifo_A_PE_11_15__full_n),
    .fifo_A_out_write(fifo_A_PE_11_15__write),
    .fifo_B_in_s_dout(fifo_B_PE_11_14__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_11_14__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_11_14__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_11_14__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_11_14__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_12_14__din),
    .fifo_B_out_full_n(fifo_B_PE_12_14__full_n),
    .fifo_B_out_write(fifo_B_PE_12_14__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_11_14__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_11_14__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_11_14__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_202
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_202__ap_start),
    .ap_done(PE_wrapper_202__ap_done),
    .ap_idle(PE_wrapper_202__ap_idle),
    .ap_ready(PE_wrapper_202__ap_ready),
    .idx(64'd11),
    .idy(64'd15),
    .fifo_A_in_s_dout(fifo_A_PE_11_15__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_11_15__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_11_15__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_11_15__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_11_15__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_11_16__din),
    .fifo_A_out_full_n(fifo_A_PE_11_16__full_n),
    .fifo_A_out_write(fifo_A_PE_11_16__write),
    .fifo_B_in_s_dout(fifo_B_PE_11_15__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_11_15__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_11_15__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_11_15__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_11_15__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_12_15__din),
    .fifo_B_out_full_n(fifo_B_PE_12_15__full_n),
    .fifo_B_out_write(fifo_B_PE_12_15__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_11_15__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_11_15__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_11_15__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_203
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_203__ap_start),
    .ap_done(PE_wrapper_203__ap_done),
    .ap_idle(PE_wrapper_203__ap_idle),
    .ap_ready(PE_wrapper_203__ap_ready),
    .idx(64'd11),
    .idy(64'd16),
    .fifo_A_in_s_dout(fifo_A_PE_11_16__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_11_16__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_11_16__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_11_16__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_11_16__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_11_17__din),
    .fifo_A_out_full_n(fifo_A_PE_11_17__full_n),
    .fifo_A_out_write(fifo_A_PE_11_17__write),
    .fifo_B_in_s_dout(fifo_B_PE_11_16__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_11_16__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_11_16__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_11_16__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_11_16__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_12_16__din),
    .fifo_B_out_full_n(fifo_B_PE_12_16__full_n),
    .fifo_B_out_write(fifo_B_PE_12_16__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_11_16__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_11_16__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_11_16__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_204
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_204__ap_start),
    .ap_done(PE_wrapper_204__ap_done),
    .ap_idle(PE_wrapper_204__ap_idle),
    .ap_ready(PE_wrapper_204__ap_ready),
    .idy(64'd0),
    .idx(64'd12),
    .fifo_A_in_s_dout(fifo_A_PE_12_0__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_12_0__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_12_0__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_12_0__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_12_0__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_12_1__din),
    .fifo_A_out_full_n(fifo_A_PE_12_1__full_n),
    .fifo_A_out_write(fifo_A_PE_12_1__write),
    .fifo_B_in_s_dout(fifo_B_PE_12_0__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_12_0__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_12_0__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_12_0__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_12_0__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_13_0__din),
    .fifo_B_out_full_n(fifo_B_PE_13_0__full_n),
    .fifo_B_out_write(fifo_B_PE_13_0__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_12_0__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_12_0__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_12_0__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_205
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_205__ap_start),
    .ap_done(PE_wrapper_205__ap_done),
    .ap_idle(PE_wrapper_205__ap_idle),
    .ap_ready(PE_wrapper_205__ap_ready),
    .idy(64'd1),
    .idx(64'd12),
    .fifo_A_in_s_dout(fifo_A_PE_12_1__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_12_1__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_12_1__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_12_1__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_12_1__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_12_2__din),
    .fifo_A_out_full_n(fifo_A_PE_12_2__full_n),
    .fifo_A_out_write(fifo_A_PE_12_2__write),
    .fifo_B_in_s_dout(fifo_B_PE_12_1__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_12_1__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_12_1__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_12_1__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_12_1__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_13_1__din),
    .fifo_B_out_full_n(fifo_B_PE_13_1__full_n),
    .fifo_B_out_write(fifo_B_PE_13_1__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_12_1__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_12_1__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_12_1__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_206
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_206__ap_start),
    .ap_done(PE_wrapper_206__ap_done),
    .ap_idle(PE_wrapper_206__ap_idle),
    .ap_ready(PE_wrapper_206__ap_ready),
    .idx(64'd12),
    .idy(64'd2),
    .fifo_A_in_s_dout(fifo_A_PE_12_2__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_12_2__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_12_2__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_12_2__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_12_2__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_12_3__din),
    .fifo_A_out_full_n(fifo_A_PE_12_3__full_n),
    .fifo_A_out_write(fifo_A_PE_12_3__write),
    .fifo_B_in_s_dout(fifo_B_PE_12_2__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_12_2__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_12_2__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_12_2__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_12_2__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_13_2__din),
    .fifo_B_out_full_n(fifo_B_PE_13_2__full_n),
    .fifo_B_out_write(fifo_B_PE_13_2__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_12_2__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_12_2__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_12_2__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_207
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_207__ap_start),
    .ap_done(PE_wrapper_207__ap_done),
    .ap_idle(PE_wrapper_207__ap_idle),
    .ap_ready(PE_wrapper_207__ap_ready),
    .idx(64'd12),
    .idy(64'd3),
    .fifo_A_in_s_dout(fifo_A_PE_12_3__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_12_3__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_12_3__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_12_3__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_12_3__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_12_4__din),
    .fifo_A_out_full_n(fifo_A_PE_12_4__full_n),
    .fifo_A_out_write(fifo_A_PE_12_4__write),
    .fifo_B_in_s_dout(fifo_B_PE_12_3__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_12_3__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_12_3__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_12_3__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_12_3__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_13_3__din),
    .fifo_B_out_full_n(fifo_B_PE_13_3__full_n),
    .fifo_B_out_write(fifo_B_PE_13_3__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_12_3__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_12_3__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_12_3__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_208
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_208__ap_start),
    .ap_done(PE_wrapper_208__ap_done),
    .ap_idle(PE_wrapper_208__ap_idle),
    .ap_ready(PE_wrapper_208__ap_ready),
    .idx(64'd12),
    .idy(64'd4),
    .fifo_A_in_s_dout(fifo_A_PE_12_4__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_12_4__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_12_4__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_12_4__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_12_4__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_12_5__din),
    .fifo_A_out_full_n(fifo_A_PE_12_5__full_n),
    .fifo_A_out_write(fifo_A_PE_12_5__write),
    .fifo_B_in_s_dout(fifo_B_PE_12_4__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_12_4__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_12_4__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_12_4__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_12_4__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_13_4__din),
    .fifo_B_out_full_n(fifo_B_PE_13_4__full_n),
    .fifo_B_out_write(fifo_B_PE_13_4__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_12_4__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_12_4__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_12_4__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_209
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_209__ap_start),
    .ap_done(PE_wrapper_209__ap_done),
    .ap_idle(PE_wrapper_209__ap_idle),
    .ap_ready(PE_wrapper_209__ap_ready),
    .idx(64'd12),
    .idy(64'd5),
    .fifo_A_in_s_dout(fifo_A_PE_12_5__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_12_5__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_12_5__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_12_5__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_12_5__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_12_6__din),
    .fifo_A_out_full_n(fifo_A_PE_12_6__full_n),
    .fifo_A_out_write(fifo_A_PE_12_6__write),
    .fifo_B_in_s_dout(fifo_B_PE_12_5__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_12_5__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_12_5__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_12_5__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_12_5__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_13_5__din),
    .fifo_B_out_full_n(fifo_B_PE_13_5__full_n),
    .fifo_B_out_write(fifo_B_PE_13_5__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_12_5__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_12_5__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_12_5__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_210
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_210__ap_start),
    .ap_done(PE_wrapper_210__ap_done),
    .ap_idle(PE_wrapper_210__ap_idle),
    .ap_ready(PE_wrapper_210__ap_ready),
    .idx(64'd12),
    .idy(64'd6),
    .fifo_A_in_s_dout(fifo_A_PE_12_6__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_12_6__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_12_6__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_12_6__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_12_6__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_12_7__din),
    .fifo_A_out_full_n(fifo_A_PE_12_7__full_n),
    .fifo_A_out_write(fifo_A_PE_12_7__write),
    .fifo_B_in_s_dout(fifo_B_PE_12_6__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_12_6__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_12_6__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_12_6__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_12_6__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_13_6__din),
    .fifo_B_out_full_n(fifo_B_PE_13_6__full_n),
    .fifo_B_out_write(fifo_B_PE_13_6__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_12_6__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_12_6__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_12_6__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_211
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_211__ap_start),
    .ap_done(PE_wrapper_211__ap_done),
    .ap_idle(PE_wrapper_211__ap_idle),
    .ap_ready(PE_wrapper_211__ap_ready),
    .idx(64'd12),
    .idy(64'd7),
    .fifo_A_in_s_dout(fifo_A_PE_12_7__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_12_7__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_12_7__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_12_7__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_12_7__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_12_8__din),
    .fifo_A_out_full_n(fifo_A_PE_12_8__full_n),
    .fifo_A_out_write(fifo_A_PE_12_8__write),
    .fifo_B_in_s_dout(fifo_B_PE_12_7__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_12_7__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_12_7__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_12_7__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_12_7__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_13_7__din),
    .fifo_B_out_full_n(fifo_B_PE_13_7__full_n),
    .fifo_B_out_write(fifo_B_PE_13_7__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_12_7__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_12_7__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_12_7__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_212
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_212__ap_start),
    .ap_done(PE_wrapper_212__ap_done),
    .ap_idle(PE_wrapper_212__ap_idle),
    .ap_ready(PE_wrapper_212__ap_ready),
    .idx(64'd12),
    .idy(64'd8),
    .fifo_A_in_s_dout(fifo_A_PE_12_8__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_12_8__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_12_8__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_12_8__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_12_8__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_12_9__din),
    .fifo_A_out_full_n(fifo_A_PE_12_9__full_n),
    .fifo_A_out_write(fifo_A_PE_12_9__write),
    .fifo_B_in_s_dout(fifo_B_PE_12_8__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_12_8__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_12_8__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_12_8__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_12_8__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_13_8__din),
    .fifo_B_out_full_n(fifo_B_PE_13_8__full_n),
    .fifo_B_out_write(fifo_B_PE_13_8__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_12_8__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_12_8__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_12_8__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_213
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_213__ap_start),
    .ap_done(PE_wrapper_213__ap_done),
    .ap_idle(PE_wrapper_213__ap_idle),
    .ap_ready(PE_wrapper_213__ap_ready),
    .idx(64'd12),
    .idy(64'd9),
    .fifo_A_out_din(fifo_A_PE_12_10__din),
    .fifo_A_out_full_n(fifo_A_PE_12_10__full_n),
    .fifo_A_out_write(fifo_A_PE_12_10__write),
    .fifo_A_in_s_dout(fifo_A_PE_12_9__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_12_9__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_12_9__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_12_9__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_12_9__read),
    .fifo_A_in_peek_read(),
    .fifo_B_in_s_dout(fifo_B_PE_12_9__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_12_9__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_12_9__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_12_9__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_12_9__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_13_9__din),
    .fifo_B_out_full_n(fifo_B_PE_13_9__full_n),
    .fifo_B_out_write(fifo_B_PE_13_9__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_12_9__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_12_9__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_12_9__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_214
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_214__ap_start),
    .ap_done(PE_wrapper_214__ap_done),
    .ap_idle(PE_wrapper_214__ap_idle),
    .ap_ready(PE_wrapper_214__ap_ready),
    .idy(64'd10),
    .idx(64'd12),
    .fifo_A_in_s_dout(fifo_A_PE_12_10__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_12_10__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_12_10__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_12_10__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_12_10__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_12_11__din),
    .fifo_A_out_full_n(fifo_A_PE_12_11__full_n),
    .fifo_A_out_write(fifo_A_PE_12_11__write),
    .fifo_B_in_s_dout(fifo_B_PE_12_10__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_12_10__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_12_10__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_12_10__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_12_10__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_13_10__din),
    .fifo_B_out_full_n(fifo_B_PE_13_10__full_n),
    .fifo_B_out_write(fifo_B_PE_13_10__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_12_10__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_12_10__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_12_10__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_215
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_215__ap_start),
    .ap_done(PE_wrapper_215__ap_done),
    .ap_idle(PE_wrapper_215__ap_idle),
    .ap_ready(PE_wrapper_215__ap_ready),
    .idy(64'd11),
    .idx(64'd12),
    .fifo_A_in_s_dout(fifo_A_PE_12_11__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_12_11__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_12_11__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_12_11__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_12_11__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_12_12__din),
    .fifo_A_out_full_n(fifo_A_PE_12_12__full_n),
    .fifo_A_out_write(fifo_A_PE_12_12__write),
    .fifo_B_in_s_dout(fifo_B_PE_12_11__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_12_11__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_12_11__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_12_11__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_12_11__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_13_11__din),
    .fifo_B_out_full_n(fifo_B_PE_13_11__full_n),
    .fifo_B_out_write(fifo_B_PE_13_11__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_12_11__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_12_11__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_12_11__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_216
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_216__ap_start),
    .ap_done(PE_wrapper_216__ap_done),
    .ap_idle(PE_wrapper_216__ap_idle),
    .ap_ready(PE_wrapper_216__ap_ready),
    .idx(64'd12),
    .idy(64'd12),
    .fifo_A_in_s_dout(fifo_A_PE_12_12__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_12_12__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_12_12__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_12_12__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_12_12__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_12_13__din),
    .fifo_A_out_full_n(fifo_A_PE_12_13__full_n),
    .fifo_A_out_write(fifo_A_PE_12_13__write),
    .fifo_B_in_s_dout(fifo_B_PE_12_12__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_12_12__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_12_12__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_12_12__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_12_12__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_13_12__din),
    .fifo_B_out_full_n(fifo_B_PE_13_12__full_n),
    .fifo_B_out_write(fifo_B_PE_13_12__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_12_12__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_12_12__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_12_12__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_217
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_217__ap_start),
    .ap_done(PE_wrapper_217__ap_done),
    .ap_idle(PE_wrapper_217__ap_idle),
    .ap_ready(PE_wrapper_217__ap_ready),
    .idx(64'd12),
    .idy(64'd13),
    .fifo_A_in_s_dout(fifo_A_PE_12_13__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_12_13__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_12_13__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_12_13__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_12_13__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_12_14__din),
    .fifo_A_out_full_n(fifo_A_PE_12_14__full_n),
    .fifo_A_out_write(fifo_A_PE_12_14__write),
    .fifo_B_in_s_dout(fifo_B_PE_12_13__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_12_13__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_12_13__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_12_13__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_12_13__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_13_13__din),
    .fifo_B_out_full_n(fifo_B_PE_13_13__full_n),
    .fifo_B_out_write(fifo_B_PE_13_13__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_12_13__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_12_13__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_12_13__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_218
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_218__ap_start),
    .ap_done(PE_wrapper_218__ap_done),
    .ap_idle(PE_wrapper_218__ap_idle),
    .ap_ready(PE_wrapper_218__ap_ready),
    .idx(64'd12),
    .idy(64'd14),
    .fifo_A_in_s_dout(fifo_A_PE_12_14__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_12_14__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_12_14__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_12_14__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_12_14__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_12_15__din),
    .fifo_A_out_full_n(fifo_A_PE_12_15__full_n),
    .fifo_A_out_write(fifo_A_PE_12_15__write),
    .fifo_B_in_s_dout(fifo_B_PE_12_14__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_12_14__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_12_14__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_12_14__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_12_14__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_13_14__din),
    .fifo_B_out_full_n(fifo_B_PE_13_14__full_n),
    .fifo_B_out_write(fifo_B_PE_13_14__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_12_14__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_12_14__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_12_14__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_219
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_219__ap_start),
    .ap_done(PE_wrapper_219__ap_done),
    .ap_idle(PE_wrapper_219__ap_idle),
    .ap_ready(PE_wrapper_219__ap_ready),
    .idx(64'd12),
    .idy(64'd15),
    .fifo_A_in_s_dout(fifo_A_PE_12_15__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_12_15__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_12_15__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_12_15__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_12_15__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_12_16__din),
    .fifo_A_out_full_n(fifo_A_PE_12_16__full_n),
    .fifo_A_out_write(fifo_A_PE_12_16__write),
    .fifo_B_in_s_dout(fifo_B_PE_12_15__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_12_15__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_12_15__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_12_15__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_12_15__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_13_15__din),
    .fifo_B_out_full_n(fifo_B_PE_13_15__full_n),
    .fifo_B_out_write(fifo_B_PE_13_15__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_12_15__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_12_15__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_12_15__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_220
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_220__ap_start),
    .ap_done(PE_wrapper_220__ap_done),
    .ap_idle(PE_wrapper_220__ap_idle),
    .ap_ready(PE_wrapper_220__ap_ready),
    .idx(64'd12),
    .idy(64'd16),
    .fifo_A_in_s_dout(fifo_A_PE_12_16__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_12_16__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_12_16__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_12_16__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_12_16__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_12_17__din),
    .fifo_A_out_full_n(fifo_A_PE_12_17__full_n),
    .fifo_A_out_write(fifo_A_PE_12_17__write),
    .fifo_B_in_s_dout(fifo_B_PE_12_16__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_12_16__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_12_16__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_12_16__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_12_16__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_13_16__din),
    .fifo_B_out_full_n(fifo_B_PE_13_16__full_n),
    .fifo_B_out_write(fifo_B_PE_13_16__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_12_16__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_12_16__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_12_16__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_221
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_221__ap_start),
    .ap_done(PE_wrapper_221__ap_done),
    .ap_idle(PE_wrapper_221__ap_idle),
    .ap_ready(PE_wrapper_221__ap_ready),
    .idy(64'd0),
    .idx(64'd13),
    .fifo_A_in_s_dout(fifo_A_PE_13_0__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_13_0__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_13_0__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_13_0__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_13_0__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_13_1__din),
    .fifo_A_out_full_n(fifo_A_PE_13_1__full_n),
    .fifo_A_out_write(fifo_A_PE_13_1__write),
    .fifo_B_in_s_dout(fifo_B_PE_13_0__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_13_0__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_13_0__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_13_0__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_13_0__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_14_0__din),
    .fifo_B_out_full_n(fifo_B_PE_14_0__full_n),
    .fifo_B_out_write(fifo_B_PE_14_0__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_13_0__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_13_0__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_13_0__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_222
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_222__ap_start),
    .ap_done(PE_wrapper_222__ap_done),
    .ap_idle(PE_wrapper_222__ap_idle),
    .ap_ready(PE_wrapper_222__ap_ready),
    .idy(64'd1),
    .idx(64'd13),
    .fifo_A_in_s_dout(fifo_A_PE_13_1__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_13_1__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_13_1__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_13_1__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_13_1__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_13_2__din),
    .fifo_A_out_full_n(fifo_A_PE_13_2__full_n),
    .fifo_A_out_write(fifo_A_PE_13_2__write),
    .fifo_B_in_s_dout(fifo_B_PE_13_1__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_13_1__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_13_1__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_13_1__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_13_1__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_14_1__din),
    .fifo_B_out_full_n(fifo_B_PE_14_1__full_n),
    .fifo_B_out_write(fifo_B_PE_14_1__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_13_1__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_13_1__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_13_1__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_223
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_223__ap_start),
    .ap_done(PE_wrapper_223__ap_done),
    .ap_idle(PE_wrapper_223__ap_idle),
    .ap_ready(PE_wrapper_223__ap_ready),
    .idx(64'd13),
    .idy(64'd2),
    .fifo_A_in_s_dout(fifo_A_PE_13_2__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_13_2__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_13_2__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_13_2__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_13_2__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_13_3__din),
    .fifo_A_out_full_n(fifo_A_PE_13_3__full_n),
    .fifo_A_out_write(fifo_A_PE_13_3__write),
    .fifo_B_in_s_dout(fifo_B_PE_13_2__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_13_2__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_13_2__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_13_2__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_13_2__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_14_2__din),
    .fifo_B_out_full_n(fifo_B_PE_14_2__full_n),
    .fifo_B_out_write(fifo_B_PE_14_2__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_13_2__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_13_2__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_13_2__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_224
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_224__ap_start),
    .ap_done(PE_wrapper_224__ap_done),
    .ap_idle(PE_wrapper_224__ap_idle),
    .ap_ready(PE_wrapper_224__ap_ready),
    .idx(64'd13),
    .idy(64'd3),
    .fifo_A_in_s_dout(fifo_A_PE_13_3__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_13_3__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_13_3__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_13_3__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_13_3__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_13_4__din),
    .fifo_A_out_full_n(fifo_A_PE_13_4__full_n),
    .fifo_A_out_write(fifo_A_PE_13_4__write),
    .fifo_B_in_s_dout(fifo_B_PE_13_3__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_13_3__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_13_3__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_13_3__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_13_3__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_14_3__din),
    .fifo_B_out_full_n(fifo_B_PE_14_3__full_n),
    .fifo_B_out_write(fifo_B_PE_14_3__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_13_3__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_13_3__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_13_3__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_225
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_225__ap_start),
    .ap_done(PE_wrapper_225__ap_done),
    .ap_idle(PE_wrapper_225__ap_idle),
    .ap_ready(PE_wrapper_225__ap_ready),
    .idx(64'd13),
    .idy(64'd4),
    .fifo_A_in_s_dout(fifo_A_PE_13_4__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_13_4__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_13_4__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_13_4__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_13_4__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_13_5__din),
    .fifo_A_out_full_n(fifo_A_PE_13_5__full_n),
    .fifo_A_out_write(fifo_A_PE_13_5__write),
    .fifo_B_in_s_dout(fifo_B_PE_13_4__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_13_4__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_13_4__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_13_4__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_13_4__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_14_4__din),
    .fifo_B_out_full_n(fifo_B_PE_14_4__full_n),
    .fifo_B_out_write(fifo_B_PE_14_4__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_13_4__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_13_4__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_13_4__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_226
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_226__ap_start),
    .ap_done(PE_wrapper_226__ap_done),
    .ap_idle(PE_wrapper_226__ap_idle),
    .ap_ready(PE_wrapper_226__ap_ready),
    .idx(64'd13),
    .idy(64'd5),
    .fifo_A_in_s_dout(fifo_A_PE_13_5__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_13_5__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_13_5__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_13_5__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_13_5__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_13_6__din),
    .fifo_A_out_full_n(fifo_A_PE_13_6__full_n),
    .fifo_A_out_write(fifo_A_PE_13_6__write),
    .fifo_B_in_s_dout(fifo_B_PE_13_5__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_13_5__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_13_5__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_13_5__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_13_5__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_14_5__din),
    .fifo_B_out_full_n(fifo_B_PE_14_5__full_n),
    .fifo_B_out_write(fifo_B_PE_14_5__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_13_5__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_13_5__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_13_5__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_227
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_227__ap_start),
    .ap_done(PE_wrapper_227__ap_done),
    .ap_idle(PE_wrapper_227__ap_idle),
    .ap_ready(PE_wrapper_227__ap_ready),
    .idx(64'd13),
    .idy(64'd6),
    .fifo_A_in_s_dout(fifo_A_PE_13_6__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_13_6__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_13_6__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_13_6__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_13_6__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_13_7__din),
    .fifo_A_out_full_n(fifo_A_PE_13_7__full_n),
    .fifo_A_out_write(fifo_A_PE_13_7__write),
    .fifo_B_in_s_dout(fifo_B_PE_13_6__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_13_6__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_13_6__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_13_6__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_13_6__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_14_6__din),
    .fifo_B_out_full_n(fifo_B_PE_14_6__full_n),
    .fifo_B_out_write(fifo_B_PE_14_6__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_13_6__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_13_6__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_13_6__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_228
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_228__ap_start),
    .ap_done(PE_wrapper_228__ap_done),
    .ap_idle(PE_wrapper_228__ap_idle),
    .ap_ready(PE_wrapper_228__ap_ready),
    .idx(64'd13),
    .idy(64'd7),
    .fifo_A_in_s_dout(fifo_A_PE_13_7__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_13_7__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_13_7__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_13_7__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_13_7__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_13_8__din),
    .fifo_A_out_full_n(fifo_A_PE_13_8__full_n),
    .fifo_A_out_write(fifo_A_PE_13_8__write),
    .fifo_B_in_s_dout(fifo_B_PE_13_7__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_13_7__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_13_7__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_13_7__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_13_7__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_14_7__din),
    .fifo_B_out_full_n(fifo_B_PE_14_7__full_n),
    .fifo_B_out_write(fifo_B_PE_14_7__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_13_7__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_13_7__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_13_7__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_229
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_229__ap_start),
    .ap_done(PE_wrapper_229__ap_done),
    .ap_idle(PE_wrapper_229__ap_idle),
    .ap_ready(PE_wrapper_229__ap_ready),
    .idx(64'd13),
    .idy(64'd8),
    .fifo_A_in_s_dout(fifo_A_PE_13_8__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_13_8__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_13_8__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_13_8__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_13_8__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_13_9__din),
    .fifo_A_out_full_n(fifo_A_PE_13_9__full_n),
    .fifo_A_out_write(fifo_A_PE_13_9__write),
    .fifo_B_in_s_dout(fifo_B_PE_13_8__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_13_8__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_13_8__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_13_8__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_13_8__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_14_8__din),
    .fifo_B_out_full_n(fifo_B_PE_14_8__full_n),
    .fifo_B_out_write(fifo_B_PE_14_8__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_13_8__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_13_8__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_13_8__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_230
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_230__ap_start),
    .ap_done(PE_wrapper_230__ap_done),
    .ap_idle(PE_wrapper_230__ap_idle),
    .ap_ready(PE_wrapper_230__ap_ready),
    .idx(64'd13),
    .idy(64'd9),
    .fifo_A_out_din(fifo_A_PE_13_10__din),
    .fifo_A_out_full_n(fifo_A_PE_13_10__full_n),
    .fifo_A_out_write(fifo_A_PE_13_10__write),
    .fifo_A_in_s_dout(fifo_A_PE_13_9__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_13_9__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_13_9__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_13_9__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_13_9__read),
    .fifo_A_in_peek_read(),
    .fifo_B_in_s_dout(fifo_B_PE_13_9__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_13_9__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_13_9__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_13_9__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_13_9__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_14_9__din),
    .fifo_B_out_full_n(fifo_B_PE_14_9__full_n),
    .fifo_B_out_write(fifo_B_PE_14_9__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_13_9__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_13_9__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_13_9__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_231
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_231__ap_start),
    .ap_done(PE_wrapper_231__ap_done),
    .ap_idle(PE_wrapper_231__ap_idle),
    .ap_ready(PE_wrapper_231__ap_ready),
    .idy(64'd10),
    .idx(64'd13),
    .fifo_A_in_s_dout(fifo_A_PE_13_10__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_13_10__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_13_10__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_13_10__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_13_10__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_13_11__din),
    .fifo_A_out_full_n(fifo_A_PE_13_11__full_n),
    .fifo_A_out_write(fifo_A_PE_13_11__write),
    .fifo_B_in_s_dout(fifo_B_PE_13_10__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_13_10__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_13_10__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_13_10__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_13_10__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_14_10__din),
    .fifo_B_out_full_n(fifo_B_PE_14_10__full_n),
    .fifo_B_out_write(fifo_B_PE_14_10__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_13_10__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_13_10__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_13_10__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_232
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_232__ap_start),
    .ap_done(PE_wrapper_232__ap_done),
    .ap_idle(PE_wrapper_232__ap_idle),
    .ap_ready(PE_wrapper_232__ap_ready),
    .idy(64'd11),
    .idx(64'd13),
    .fifo_A_in_s_dout(fifo_A_PE_13_11__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_13_11__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_13_11__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_13_11__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_13_11__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_13_12__din),
    .fifo_A_out_full_n(fifo_A_PE_13_12__full_n),
    .fifo_A_out_write(fifo_A_PE_13_12__write),
    .fifo_B_in_s_dout(fifo_B_PE_13_11__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_13_11__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_13_11__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_13_11__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_13_11__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_14_11__din),
    .fifo_B_out_full_n(fifo_B_PE_14_11__full_n),
    .fifo_B_out_write(fifo_B_PE_14_11__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_13_11__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_13_11__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_13_11__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_233
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_233__ap_start),
    .ap_done(PE_wrapper_233__ap_done),
    .ap_idle(PE_wrapper_233__ap_idle),
    .ap_ready(PE_wrapper_233__ap_ready),
    .idy(64'd12),
    .idx(64'd13),
    .fifo_A_in_s_dout(fifo_A_PE_13_12__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_13_12__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_13_12__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_13_12__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_13_12__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_13_13__din),
    .fifo_A_out_full_n(fifo_A_PE_13_13__full_n),
    .fifo_A_out_write(fifo_A_PE_13_13__write),
    .fifo_B_in_s_dout(fifo_B_PE_13_12__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_13_12__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_13_12__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_13_12__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_13_12__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_14_12__din),
    .fifo_B_out_full_n(fifo_B_PE_14_12__full_n),
    .fifo_B_out_write(fifo_B_PE_14_12__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_13_12__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_13_12__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_13_12__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_234
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_234__ap_start),
    .ap_done(PE_wrapper_234__ap_done),
    .ap_idle(PE_wrapper_234__ap_idle),
    .ap_ready(PE_wrapper_234__ap_ready),
    .idx(64'd13),
    .idy(64'd13),
    .fifo_A_in_s_dout(fifo_A_PE_13_13__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_13_13__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_13_13__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_13_13__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_13_13__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_13_14__din),
    .fifo_A_out_full_n(fifo_A_PE_13_14__full_n),
    .fifo_A_out_write(fifo_A_PE_13_14__write),
    .fifo_B_in_s_dout(fifo_B_PE_13_13__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_13_13__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_13_13__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_13_13__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_13_13__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_14_13__din),
    .fifo_B_out_full_n(fifo_B_PE_14_13__full_n),
    .fifo_B_out_write(fifo_B_PE_14_13__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_13_13__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_13_13__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_13_13__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_235
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_235__ap_start),
    .ap_done(PE_wrapper_235__ap_done),
    .ap_idle(PE_wrapper_235__ap_idle),
    .ap_ready(PE_wrapper_235__ap_ready),
    .idx(64'd13),
    .idy(64'd14),
    .fifo_A_in_s_dout(fifo_A_PE_13_14__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_13_14__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_13_14__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_13_14__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_13_14__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_13_15__din),
    .fifo_A_out_full_n(fifo_A_PE_13_15__full_n),
    .fifo_A_out_write(fifo_A_PE_13_15__write),
    .fifo_B_in_s_dout(fifo_B_PE_13_14__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_13_14__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_13_14__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_13_14__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_13_14__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_14_14__din),
    .fifo_B_out_full_n(fifo_B_PE_14_14__full_n),
    .fifo_B_out_write(fifo_B_PE_14_14__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_13_14__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_13_14__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_13_14__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_236
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_236__ap_start),
    .ap_done(PE_wrapper_236__ap_done),
    .ap_idle(PE_wrapper_236__ap_idle),
    .ap_ready(PE_wrapper_236__ap_ready),
    .idx(64'd13),
    .idy(64'd15),
    .fifo_A_in_s_dout(fifo_A_PE_13_15__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_13_15__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_13_15__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_13_15__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_13_15__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_13_16__din),
    .fifo_A_out_full_n(fifo_A_PE_13_16__full_n),
    .fifo_A_out_write(fifo_A_PE_13_16__write),
    .fifo_B_in_s_dout(fifo_B_PE_13_15__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_13_15__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_13_15__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_13_15__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_13_15__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_14_15__din),
    .fifo_B_out_full_n(fifo_B_PE_14_15__full_n),
    .fifo_B_out_write(fifo_B_PE_14_15__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_13_15__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_13_15__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_13_15__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_237
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_237__ap_start),
    .ap_done(PE_wrapper_237__ap_done),
    .ap_idle(PE_wrapper_237__ap_idle),
    .ap_ready(PE_wrapper_237__ap_ready),
    .idx(64'd13),
    .idy(64'd16),
    .fifo_A_in_s_dout(fifo_A_PE_13_16__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_13_16__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_13_16__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_13_16__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_13_16__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_13_17__din),
    .fifo_A_out_full_n(fifo_A_PE_13_17__full_n),
    .fifo_A_out_write(fifo_A_PE_13_17__write),
    .fifo_B_in_s_dout(fifo_B_PE_13_16__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_13_16__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_13_16__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_13_16__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_13_16__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_14_16__din),
    .fifo_B_out_full_n(fifo_B_PE_14_16__full_n),
    .fifo_B_out_write(fifo_B_PE_14_16__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_13_16__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_13_16__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_13_16__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_238
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_238__ap_start),
    .ap_done(PE_wrapper_238__ap_done),
    .ap_idle(PE_wrapper_238__ap_idle),
    .ap_ready(PE_wrapper_238__ap_ready),
    .idy(64'd0),
    .idx(64'd14),
    .fifo_A_in_s_dout(fifo_A_PE_14_0__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_14_0__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_14_0__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_14_0__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_14_0__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_14_1__din),
    .fifo_A_out_full_n(fifo_A_PE_14_1__full_n),
    .fifo_A_out_write(fifo_A_PE_14_1__write),
    .fifo_B_in_s_dout(fifo_B_PE_14_0__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_14_0__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_14_0__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_14_0__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_14_0__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_15_0__din),
    .fifo_B_out_full_n(fifo_B_PE_15_0__full_n),
    .fifo_B_out_write(fifo_B_PE_15_0__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_14_0__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_14_0__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_14_0__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_239
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_239__ap_start),
    .ap_done(PE_wrapper_239__ap_done),
    .ap_idle(PE_wrapper_239__ap_idle),
    .ap_ready(PE_wrapper_239__ap_ready),
    .idy(64'd1),
    .idx(64'd14),
    .fifo_A_in_s_dout(fifo_A_PE_14_1__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_14_1__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_14_1__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_14_1__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_14_1__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_14_2__din),
    .fifo_A_out_full_n(fifo_A_PE_14_2__full_n),
    .fifo_A_out_write(fifo_A_PE_14_2__write),
    .fifo_B_in_s_dout(fifo_B_PE_14_1__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_14_1__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_14_1__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_14_1__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_14_1__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_15_1__din),
    .fifo_B_out_full_n(fifo_B_PE_15_1__full_n),
    .fifo_B_out_write(fifo_B_PE_15_1__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_14_1__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_14_1__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_14_1__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_240
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_240__ap_start),
    .ap_done(PE_wrapper_240__ap_done),
    .ap_idle(PE_wrapper_240__ap_idle),
    .ap_ready(PE_wrapper_240__ap_ready),
    .idx(64'd14),
    .idy(64'd2),
    .fifo_A_in_s_dout(fifo_A_PE_14_2__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_14_2__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_14_2__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_14_2__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_14_2__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_14_3__din),
    .fifo_A_out_full_n(fifo_A_PE_14_3__full_n),
    .fifo_A_out_write(fifo_A_PE_14_3__write),
    .fifo_B_in_s_dout(fifo_B_PE_14_2__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_14_2__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_14_2__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_14_2__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_14_2__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_15_2__din),
    .fifo_B_out_full_n(fifo_B_PE_15_2__full_n),
    .fifo_B_out_write(fifo_B_PE_15_2__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_14_2__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_14_2__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_14_2__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_241
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_241__ap_start),
    .ap_done(PE_wrapper_241__ap_done),
    .ap_idle(PE_wrapper_241__ap_idle),
    .ap_ready(PE_wrapper_241__ap_ready),
    .idx(64'd14),
    .idy(64'd3),
    .fifo_A_in_s_dout(fifo_A_PE_14_3__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_14_3__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_14_3__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_14_3__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_14_3__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_14_4__din),
    .fifo_A_out_full_n(fifo_A_PE_14_4__full_n),
    .fifo_A_out_write(fifo_A_PE_14_4__write),
    .fifo_B_in_s_dout(fifo_B_PE_14_3__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_14_3__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_14_3__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_14_3__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_14_3__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_15_3__din),
    .fifo_B_out_full_n(fifo_B_PE_15_3__full_n),
    .fifo_B_out_write(fifo_B_PE_15_3__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_14_3__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_14_3__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_14_3__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_242
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_242__ap_start),
    .ap_done(PE_wrapper_242__ap_done),
    .ap_idle(PE_wrapper_242__ap_idle),
    .ap_ready(PE_wrapper_242__ap_ready),
    .idx(64'd14),
    .idy(64'd4),
    .fifo_A_in_s_dout(fifo_A_PE_14_4__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_14_4__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_14_4__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_14_4__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_14_4__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_14_5__din),
    .fifo_A_out_full_n(fifo_A_PE_14_5__full_n),
    .fifo_A_out_write(fifo_A_PE_14_5__write),
    .fifo_B_in_s_dout(fifo_B_PE_14_4__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_14_4__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_14_4__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_14_4__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_14_4__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_15_4__din),
    .fifo_B_out_full_n(fifo_B_PE_15_4__full_n),
    .fifo_B_out_write(fifo_B_PE_15_4__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_14_4__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_14_4__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_14_4__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_243
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_243__ap_start),
    .ap_done(PE_wrapper_243__ap_done),
    .ap_idle(PE_wrapper_243__ap_idle),
    .ap_ready(PE_wrapper_243__ap_ready),
    .idx(64'd14),
    .idy(64'd5),
    .fifo_A_in_s_dout(fifo_A_PE_14_5__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_14_5__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_14_5__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_14_5__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_14_5__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_14_6__din),
    .fifo_A_out_full_n(fifo_A_PE_14_6__full_n),
    .fifo_A_out_write(fifo_A_PE_14_6__write),
    .fifo_B_in_s_dout(fifo_B_PE_14_5__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_14_5__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_14_5__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_14_5__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_14_5__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_15_5__din),
    .fifo_B_out_full_n(fifo_B_PE_15_5__full_n),
    .fifo_B_out_write(fifo_B_PE_15_5__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_14_5__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_14_5__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_14_5__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_244
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_244__ap_start),
    .ap_done(PE_wrapper_244__ap_done),
    .ap_idle(PE_wrapper_244__ap_idle),
    .ap_ready(PE_wrapper_244__ap_ready),
    .idx(64'd14),
    .idy(64'd6),
    .fifo_A_in_s_dout(fifo_A_PE_14_6__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_14_6__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_14_6__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_14_6__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_14_6__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_14_7__din),
    .fifo_A_out_full_n(fifo_A_PE_14_7__full_n),
    .fifo_A_out_write(fifo_A_PE_14_7__write),
    .fifo_B_in_s_dout(fifo_B_PE_14_6__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_14_6__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_14_6__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_14_6__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_14_6__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_15_6__din),
    .fifo_B_out_full_n(fifo_B_PE_15_6__full_n),
    .fifo_B_out_write(fifo_B_PE_15_6__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_14_6__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_14_6__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_14_6__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_245
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_245__ap_start),
    .ap_done(PE_wrapper_245__ap_done),
    .ap_idle(PE_wrapper_245__ap_idle),
    .ap_ready(PE_wrapper_245__ap_ready),
    .idx(64'd14),
    .idy(64'd7),
    .fifo_A_in_s_dout(fifo_A_PE_14_7__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_14_7__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_14_7__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_14_7__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_14_7__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_14_8__din),
    .fifo_A_out_full_n(fifo_A_PE_14_8__full_n),
    .fifo_A_out_write(fifo_A_PE_14_8__write),
    .fifo_B_in_s_dout(fifo_B_PE_14_7__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_14_7__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_14_7__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_14_7__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_14_7__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_15_7__din),
    .fifo_B_out_full_n(fifo_B_PE_15_7__full_n),
    .fifo_B_out_write(fifo_B_PE_15_7__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_14_7__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_14_7__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_14_7__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_246
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_246__ap_start),
    .ap_done(PE_wrapper_246__ap_done),
    .ap_idle(PE_wrapper_246__ap_idle),
    .ap_ready(PE_wrapper_246__ap_ready),
    .idx(64'd14),
    .idy(64'd8),
    .fifo_A_in_s_dout(fifo_A_PE_14_8__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_14_8__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_14_8__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_14_8__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_14_8__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_14_9__din),
    .fifo_A_out_full_n(fifo_A_PE_14_9__full_n),
    .fifo_A_out_write(fifo_A_PE_14_9__write),
    .fifo_B_in_s_dout(fifo_B_PE_14_8__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_14_8__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_14_8__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_14_8__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_14_8__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_15_8__din),
    .fifo_B_out_full_n(fifo_B_PE_15_8__full_n),
    .fifo_B_out_write(fifo_B_PE_15_8__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_14_8__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_14_8__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_14_8__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_247
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_247__ap_start),
    .ap_done(PE_wrapper_247__ap_done),
    .ap_idle(PE_wrapper_247__ap_idle),
    .ap_ready(PE_wrapper_247__ap_ready),
    .idx(64'd14),
    .idy(64'd9),
    .fifo_A_out_din(fifo_A_PE_14_10__din),
    .fifo_A_out_full_n(fifo_A_PE_14_10__full_n),
    .fifo_A_out_write(fifo_A_PE_14_10__write),
    .fifo_A_in_s_dout(fifo_A_PE_14_9__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_14_9__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_14_9__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_14_9__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_14_9__read),
    .fifo_A_in_peek_read(),
    .fifo_B_in_s_dout(fifo_B_PE_14_9__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_14_9__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_14_9__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_14_9__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_14_9__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_15_9__din),
    .fifo_B_out_full_n(fifo_B_PE_15_9__full_n),
    .fifo_B_out_write(fifo_B_PE_15_9__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_14_9__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_14_9__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_14_9__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_248
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_248__ap_start),
    .ap_done(PE_wrapper_248__ap_done),
    .ap_idle(PE_wrapper_248__ap_idle),
    .ap_ready(PE_wrapper_248__ap_ready),
    .idy(64'd10),
    .idx(64'd14),
    .fifo_A_in_s_dout(fifo_A_PE_14_10__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_14_10__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_14_10__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_14_10__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_14_10__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_14_11__din),
    .fifo_A_out_full_n(fifo_A_PE_14_11__full_n),
    .fifo_A_out_write(fifo_A_PE_14_11__write),
    .fifo_B_in_s_dout(fifo_B_PE_14_10__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_14_10__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_14_10__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_14_10__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_14_10__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_15_10__din),
    .fifo_B_out_full_n(fifo_B_PE_15_10__full_n),
    .fifo_B_out_write(fifo_B_PE_15_10__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_14_10__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_14_10__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_14_10__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_249
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_249__ap_start),
    .ap_done(PE_wrapper_249__ap_done),
    .ap_idle(PE_wrapper_249__ap_idle),
    .ap_ready(PE_wrapper_249__ap_ready),
    .idy(64'd11),
    .idx(64'd14),
    .fifo_A_in_s_dout(fifo_A_PE_14_11__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_14_11__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_14_11__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_14_11__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_14_11__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_14_12__din),
    .fifo_A_out_full_n(fifo_A_PE_14_12__full_n),
    .fifo_A_out_write(fifo_A_PE_14_12__write),
    .fifo_B_in_s_dout(fifo_B_PE_14_11__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_14_11__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_14_11__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_14_11__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_14_11__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_15_11__din),
    .fifo_B_out_full_n(fifo_B_PE_15_11__full_n),
    .fifo_B_out_write(fifo_B_PE_15_11__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_14_11__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_14_11__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_14_11__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_250
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_250__ap_start),
    .ap_done(PE_wrapper_250__ap_done),
    .ap_idle(PE_wrapper_250__ap_idle),
    .ap_ready(PE_wrapper_250__ap_ready),
    .idy(64'd12),
    .idx(64'd14),
    .fifo_A_in_s_dout(fifo_A_PE_14_12__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_14_12__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_14_12__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_14_12__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_14_12__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_14_13__din),
    .fifo_A_out_full_n(fifo_A_PE_14_13__full_n),
    .fifo_A_out_write(fifo_A_PE_14_13__write),
    .fifo_B_in_s_dout(fifo_B_PE_14_12__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_14_12__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_14_12__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_14_12__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_14_12__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_15_12__din),
    .fifo_B_out_full_n(fifo_B_PE_15_12__full_n),
    .fifo_B_out_write(fifo_B_PE_15_12__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_14_12__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_14_12__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_14_12__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_251
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_251__ap_start),
    .ap_done(PE_wrapper_251__ap_done),
    .ap_idle(PE_wrapper_251__ap_idle),
    .ap_ready(PE_wrapper_251__ap_ready),
    .idy(64'd13),
    .idx(64'd14),
    .fifo_A_in_s_dout(fifo_A_PE_14_13__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_14_13__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_14_13__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_14_13__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_14_13__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_14_14__din),
    .fifo_A_out_full_n(fifo_A_PE_14_14__full_n),
    .fifo_A_out_write(fifo_A_PE_14_14__write),
    .fifo_B_in_s_dout(fifo_B_PE_14_13__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_14_13__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_14_13__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_14_13__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_14_13__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_15_13__din),
    .fifo_B_out_full_n(fifo_B_PE_15_13__full_n),
    .fifo_B_out_write(fifo_B_PE_15_13__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_14_13__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_14_13__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_14_13__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_252
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_252__ap_start),
    .ap_done(PE_wrapper_252__ap_done),
    .ap_idle(PE_wrapper_252__ap_idle),
    .ap_ready(PE_wrapper_252__ap_ready),
    .idx(64'd14),
    .idy(64'd14),
    .fifo_A_in_s_dout(fifo_A_PE_14_14__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_14_14__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_14_14__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_14_14__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_14_14__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_14_15__din),
    .fifo_A_out_full_n(fifo_A_PE_14_15__full_n),
    .fifo_A_out_write(fifo_A_PE_14_15__write),
    .fifo_B_in_s_dout(fifo_B_PE_14_14__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_14_14__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_14_14__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_14_14__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_14_14__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_15_14__din),
    .fifo_B_out_full_n(fifo_B_PE_15_14__full_n),
    .fifo_B_out_write(fifo_B_PE_15_14__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_14_14__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_14_14__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_14_14__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_253
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_253__ap_start),
    .ap_done(PE_wrapper_253__ap_done),
    .ap_idle(PE_wrapper_253__ap_idle),
    .ap_ready(PE_wrapper_253__ap_ready),
    .idx(64'd14),
    .idy(64'd15),
    .fifo_A_in_s_dout(fifo_A_PE_14_15__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_14_15__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_14_15__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_14_15__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_14_15__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_14_16__din),
    .fifo_A_out_full_n(fifo_A_PE_14_16__full_n),
    .fifo_A_out_write(fifo_A_PE_14_16__write),
    .fifo_B_in_s_dout(fifo_B_PE_14_15__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_14_15__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_14_15__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_14_15__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_14_15__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_15_15__din),
    .fifo_B_out_full_n(fifo_B_PE_15_15__full_n),
    .fifo_B_out_write(fifo_B_PE_15_15__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_14_15__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_14_15__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_14_15__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_254
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_254__ap_start),
    .ap_done(PE_wrapper_254__ap_done),
    .ap_idle(PE_wrapper_254__ap_idle),
    .ap_ready(PE_wrapper_254__ap_ready),
    .idx(64'd14),
    .idy(64'd16),
    .fifo_A_in_s_dout(fifo_A_PE_14_16__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_14_16__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_14_16__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_14_16__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_14_16__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_14_17__din),
    .fifo_A_out_full_n(fifo_A_PE_14_17__full_n),
    .fifo_A_out_write(fifo_A_PE_14_17__write),
    .fifo_B_in_s_dout(fifo_B_PE_14_16__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_14_16__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_14_16__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_14_16__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_14_16__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_15_16__din),
    .fifo_B_out_full_n(fifo_B_PE_15_16__full_n),
    .fifo_B_out_write(fifo_B_PE_15_16__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_14_16__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_14_16__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_14_16__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_255
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_255__ap_start),
    .ap_done(PE_wrapper_255__ap_done),
    .ap_idle(PE_wrapper_255__ap_idle),
    .ap_ready(PE_wrapper_255__ap_ready),
    .idy(64'd0),
    .idx(64'd15),
    .fifo_A_in_s_dout(fifo_A_PE_15_0__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_15_0__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_15_0__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_15_0__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_15_0__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_15_1__din),
    .fifo_A_out_full_n(fifo_A_PE_15_1__full_n),
    .fifo_A_out_write(fifo_A_PE_15_1__write),
    .fifo_B_in_s_dout(fifo_B_PE_15_0__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_15_0__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_15_0__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_15_0__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_15_0__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_16_0__din),
    .fifo_B_out_full_n(fifo_B_PE_16_0__full_n),
    .fifo_B_out_write(fifo_B_PE_16_0__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_15_0__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_15_0__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_15_0__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_256
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_256__ap_start),
    .ap_done(PE_wrapper_256__ap_done),
    .ap_idle(PE_wrapper_256__ap_idle),
    .ap_ready(PE_wrapper_256__ap_ready),
    .idy(64'd1),
    .idx(64'd15),
    .fifo_A_in_s_dout(fifo_A_PE_15_1__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_15_1__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_15_1__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_15_1__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_15_1__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_15_2__din),
    .fifo_A_out_full_n(fifo_A_PE_15_2__full_n),
    .fifo_A_out_write(fifo_A_PE_15_2__write),
    .fifo_B_in_s_dout(fifo_B_PE_15_1__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_15_1__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_15_1__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_15_1__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_15_1__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_16_1__din),
    .fifo_B_out_full_n(fifo_B_PE_16_1__full_n),
    .fifo_B_out_write(fifo_B_PE_16_1__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_15_1__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_15_1__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_15_1__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_257
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_257__ap_start),
    .ap_done(PE_wrapper_257__ap_done),
    .ap_idle(PE_wrapper_257__ap_idle),
    .ap_ready(PE_wrapper_257__ap_ready),
    .idx(64'd15),
    .idy(64'd2),
    .fifo_A_in_s_dout(fifo_A_PE_15_2__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_15_2__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_15_2__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_15_2__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_15_2__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_15_3__din),
    .fifo_A_out_full_n(fifo_A_PE_15_3__full_n),
    .fifo_A_out_write(fifo_A_PE_15_3__write),
    .fifo_B_in_s_dout(fifo_B_PE_15_2__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_15_2__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_15_2__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_15_2__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_15_2__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_16_2__din),
    .fifo_B_out_full_n(fifo_B_PE_16_2__full_n),
    .fifo_B_out_write(fifo_B_PE_16_2__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_15_2__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_15_2__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_15_2__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_258
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_258__ap_start),
    .ap_done(PE_wrapper_258__ap_done),
    .ap_idle(PE_wrapper_258__ap_idle),
    .ap_ready(PE_wrapper_258__ap_ready),
    .idx(64'd15),
    .idy(64'd3),
    .fifo_A_in_s_dout(fifo_A_PE_15_3__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_15_3__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_15_3__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_15_3__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_15_3__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_15_4__din),
    .fifo_A_out_full_n(fifo_A_PE_15_4__full_n),
    .fifo_A_out_write(fifo_A_PE_15_4__write),
    .fifo_B_in_s_dout(fifo_B_PE_15_3__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_15_3__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_15_3__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_15_3__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_15_3__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_16_3__din),
    .fifo_B_out_full_n(fifo_B_PE_16_3__full_n),
    .fifo_B_out_write(fifo_B_PE_16_3__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_15_3__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_15_3__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_15_3__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_259
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_259__ap_start),
    .ap_done(PE_wrapper_259__ap_done),
    .ap_idle(PE_wrapper_259__ap_idle),
    .ap_ready(PE_wrapper_259__ap_ready),
    .idx(64'd15),
    .idy(64'd4),
    .fifo_A_in_s_dout(fifo_A_PE_15_4__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_15_4__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_15_4__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_15_4__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_15_4__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_15_5__din),
    .fifo_A_out_full_n(fifo_A_PE_15_5__full_n),
    .fifo_A_out_write(fifo_A_PE_15_5__write),
    .fifo_B_in_s_dout(fifo_B_PE_15_4__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_15_4__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_15_4__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_15_4__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_15_4__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_16_4__din),
    .fifo_B_out_full_n(fifo_B_PE_16_4__full_n),
    .fifo_B_out_write(fifo_B_PE_16_4__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_15_4__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_15_4__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_15_4__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_260
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_260__ap_start),
    .ap_done(PE_wrapper_260__ap_done),
    .ap_idle(PE_wrapper_260__ap_idle),
    .ap_ready(PE_wrapper_260__ap_ready),
    .idx(64'd15),
    .idy(64'd5),
    .fifo_A_in_s_dout(fifo_A_PE_15_5__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_15_5__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_15_5__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_15_5__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_15_5__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_15_6__din),
    .fifo_A_out_full_n(fifo_A_PE_15_6__full_n),
    .fifo_A_out_write(fifo_A_PE_15_6__write),
    .fifo_B_in_s_dout(fifo_B_PE_15_5__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_15_5__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_15_5__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_15_5__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_15_5__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_16_5__din),
    .fifo_B_out_full_n(fifo_B_PE_16_5__full_n),
    .fifo_B_out_write(fifo_B_PE_16_5__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_15_5__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_15_5__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_15_5__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_261
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_261__ap_start),
    .ap_done(PE_wrapper_261__ap_done),
    .ap_idle(PE_wrapper_261__ap_idle),
    .ap_ready(PE_wrapper_261__ap_ready),
    .idx(64'd15),
    .idy(64'd6),
    .fifo_A_in_s_dout(fifo_A_PE_15_6__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_15_6__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_15_6__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_15_6__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_15_6__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_15_7__din),
    .fifo_A_out_full_n(fifo_A_PE_15_7__full_n),
    .fifo_A_out_write(fifo_A_PE_15_7__write),
    .fifo_B_in_s_dout(fifo_B_PE_15_6__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_15_6__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_15_6__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_15_6__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_15_6__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_16_6__din),
    .fifo_B_out_full_n(fifo_B_PE_16_6__full_n),
    .fifo_B_out_write(fifo_B_PE_16_6__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_15_6__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_15_6__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_15_6__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_262
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_262__ap_start),
    .ap_done(PE_wrapper_262__ap_done),
    .ap_idle(PE_wrapper_262__ap_idle),
    .ap_ready(PE_wrapper_262__ap_ready),
    .idx(64'd15),
    .idy(64'd7),
    .fifo_A_in_s_dout(fifo_A_PE_15_7__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_15_7__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_15_7__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_15_7__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_15_7__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_15_8__din),
    .fifo_A_out_full_n(fifo_A_PE_15_8__full_n),
    .fifo_A_out_write(fifo_A_PE_15_8__write),
    .fifo_B_in_s_dout(fifo_B_PE_15_7__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_15_7__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_15_7__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_15_7__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_15_7__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_16_7__din),
    .fifo_B_out_full_n(fifo_B_PE_16_7__full_n),
    .fifo_B_out_write(fifo_B_PE_16_7__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_15_7__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_15_7__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_15_7__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_263
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_263__ap_start),
    .ap_done(PE_wrapper_263__ap_done),
    .ap_idle(PE_wrapper_263__ap_idle),
    .ap_ready(PE_wrapper_263__ap_ready),
    .idx(64'd15),
    .idy(64'd8),
    .fifo_A_in_s_dout(fifo_A_PE_15_8__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_15_8__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_15_8__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_15_8__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_15_8__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_15_9__din),
    .fifo_A_out_full_n(fifo_A_PE_15_9__full_n),
    .fifo_A_out_write(fifo_A_PE_15_9__write),
    .fifo_B_in_s_dout(fifo_B_PE_15_8__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_15_8__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_15_8__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_15_8__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_15_8__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_16_8__din),
    .fifo_B_out_full_n(fifo_B_PE_16_8__full_n),
    .fifo_B_out_write(fifo_B_PE_16_8__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_15_8__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_15_8__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_15_8__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_264
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_264__ap_start),
    .ap_done(PE_wrapper_264__ap_done),
    .ap_idle(PE_wrapper_264__ap_idle),
    .ap_ready(PE_wrapper_264__ap_ready),
    .idx(64'd15),
    .idy(64'd9),
    .fifo_A_out_din(fifo_A_PE_15_10__din),
    .fifo_A_out_full_n(fifo_A_PE_15_10__full_n),
    .fifo_A_out_write(fifo_A_PE_15_10__write),
    .fifo_A_in_s_dout(fifo_A_PE_15_9__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_15_9__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_15_9__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_15_9__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_15_9__read),
    .fifo_A_in_peek_read(),
    .fifo_B_in_s_dout(fifo_B_PE_15_9__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_15_9__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_15_9__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_15_9__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_15_9__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_16_9__din),
    .fifo_B_out_full_n(fifo_B_PE_16_9__full_n),
    .fifo_B_out_write(fifo_B_PE_16_9__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_15_9__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_15_9__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_15_9__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_265
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_265__ap_start),
    .ap_done(PE_wrapper_265__ap_done),
    .ap_idle(PE_wrapper_265__ap_idle),
    .ap_ready(PE_wrapper_265__ap_ready),
    .idy(64'd10),
    .idx(64'd15),
    .fifo_A_in_s_dout(fifo_A_PE_15_10__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_15_10__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_15_10__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_15_10__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_15_10__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_15_11__din),
    .fifo_A_out_full_n(fifo_A_PE_15_11__full_n),
    .fifo_A_out_write(fifo_A_PE_15_11__write),
    .fifo_B_in_s_dout(fifo_B_PE_15_10__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_15_10__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_15_10__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_15_10__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_15_10__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_16_10__din),
    .fifo_B_out_full_n(fifo_B_PE_16_10__full_n),
    .fifo_B_out_write(fifo_B_PE_16_10__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_15_10__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_15_10__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_15_10__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_266
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_266__ap_start),
    .ap_done(PE_wrapper_266__ap_done),
    .ap_idle(PE_wrapper_266__ap_idle),
    .ap_ready(PE_wrapper_266__ap_ready),
    .idy(64'd11),
    .idx(64'd15),
    .fifo_A_in_s_dout(fifo_A_PE_15_11__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_15_11__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_15_11__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_15_11__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_15_11__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_15_12__din),
    .fifo_A_out_full_n(fifo_A_PE_15_12__full_n),
    .fifo_A_out_write(fifo_A_PE_15_12__write),
    .fifo_B_in_s_dout(fifo_B_PE_15_11__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_15_11__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_15_11__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_15_11__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_15_11__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_16_11__din),
    .fifo_B_out_full_n(fifo_B_PE_16_11__full_n),
    .fifo_B_out_write(fifo_B_PE_16_11__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_15_11__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_15_11__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_15_11__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_267
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_267__ap_start),
    .ap_done(PE_wrapper_267__ap_done),
    .ap_idle(PE_wrapper_267__ap_idle),
    .ap_ready(PE_wrapper_267__ap_ready),
    .idy(64'd12),
    .idx(64'd15),
    .fifo_A_in_s_dout(fifo_A_PE_15_12__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_15_12__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_15_12__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_15_12__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_15_12__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_15_13__din),
    .fifo_A_out_full_n(fifo_A_PE_15_13__full_n),
    .fifo_A_out_write(fifo_A_PE_15_13__write),
    .fifo_B_in_s_dout(fifo_B_PE_15_12__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_15_12__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_15_12__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_15_12__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_15_12__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_16_12__din),
    .fifo_B_out_full_n(fifo_B_PE_16_12__full_n),
    .fifo_B_out_write(fifo_B_PE_16_12__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_15_12__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_15_12__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_15_12__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_268
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_268__ap_start),
    .ap_done(PE_wrapper_268__ap_done),
    .ap_idle(PE_wrapper_268__ap_idle),
    .ap_ready(PE_wrapper_268__ap_ready),
    .idy(64'd13),
    .idx(64'd15),
    .fifo_A_in_s_dout(fifo_A_PE_15_13__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_15_13__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_15_13__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_15_13__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_15_13__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_15_14__din),
    .fifo_A_out_full_n(fifo_A_PE_15_14__full_n),
    .fifo_A_out_write(fifo_A_PE_15_14__write),
    .fifo_B_in_s_dout(fifo_B_PE_15_13__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_15_13__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_15_13__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_15_13__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_15_13__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_16_13__din),
    .fifo_B_out_full_n(fifo_B_PE_16_13__full_n),
    .fifo_B_out_write(fifo_B_PE_16_13__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_15_13__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_15_13__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_15_13__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_269
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_269__ap_start),
    .ap_done(PE_wrapper_269__ap_done),
    .ap_idle(PE_wrapper_269__ap_idle),
    .ap_ready(PE_wrapper_269__ap_ready),
    .idy(64'd14),
    .idx(64'd15),
    .fifo_A_in_s_dout(fifo_A_PE_15_14__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_15_14__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_15_14__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_15_14__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_15_14__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_15_15__din),
    .fifo_A_out_full_n(fifo_A_PE_15_15__full_n),
    .fifo_A_out_write(fifo_A_PE_15_15__write),
    .fifo_B_in_s_dout(fifo_B_PE_15_14__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_15_14__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_15_14__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_15_14__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_15_14__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_16_14__din),
    .fifo_B_out_full_n(fifo_B_PE_16_14__full_n),
    .fifo_B_out_write(fifo_B_PE_16_14__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_15_14__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_15_14__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_15_14__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_270
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_270__ap_start),
    .ap_done(PE_wrapper_270__ap_done),
    .ap_idle(PE_wrapper_270__ap_idle),
    .ap_ready(PE_wrapper_270__ap_ready),
    .idx(64'd15),
    .idy(64'd15),
    .fifo_A_in_s_dout(fifo_A_PE_15_15__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_15_15__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_15_15__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_15_15__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_15_15__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_15_16__din),
    .fifo_A_out_full_n(fifo_A_PE_15_16__full_n),
    .fifo_A_out_write(fifo_A_PE_15_16__write),
    .fifo_B_in_s_dout(fifo_B_PE_15_15__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_15_15__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_15_15__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_15_15__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_15_15__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_16_15__din),
    .fifo_B_out_full_n(fifo_B_PE_16_15__full_n),
    .fifo_B_out_write(fifo_B_PE_16_15__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_15_15__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_15_15__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_15_15__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_271
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_271__ap_start),
    .ap_done(PE_wrapper_271__ap_done),
    .ap_idle(PE_wrapper_271__ap_idle),
    .ap_ready(PE_wrapper_271__ap_ready),
    .idx(64'd15),
    .idy(64'd16),
    .fifo_A_in_s_dout(fifo_A_PE_15_16__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_15_16__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_15_16__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_15_16__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_15_16__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_15_17__din),
    .fifo_A_out_full_n(fifo_A_PE_15_17__full_n),
    .fifo_A_out_write(fifo_A_PE_15_17__write),
    .fifo_B_in_s_dout(fifo_B_PE_15_16__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_15_16__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_15_16__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_15_16__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_15_16__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_16_16__din),
    .fifo_B_out_full_n(fifo_B_PE_16_16__full_n),
    .fifo_B_out_write(fifo_B_PE_16_16__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_15_16__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_15_16__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_15_16__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_272
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_272__ap_start),
    .ap_done(PE_wrapper_272__ap_done),
    .ap_idle(PE_wrapper_272__ap_idle),
    .ap_ready(PE_wrapper_272__ap_ready),
    .idy(64'd0),
    .idx(64'd16),
    .fifo_A_in_s_dout(fifo_A_PE_16_0__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_16_0__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_16_0__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_16_0__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_16_0__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_16_1__din),
    .fifo_A_out_full_n(fifo_A_PE_16_1__full_n),
    .fifo_A_out_write(fifo_A_PE_16_1__write),
    .fifo_B_in_s_dout(fifo_B_PE_16_0__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_16_0__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_16_0__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_16_0__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_16_0__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_17_0__din),
    .fifo_B_out_full_n(fifo_B_PE_17_0__full_n),
    .fifo_B_out_write(fifo_B_PE_17_0__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_16_0__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_16_0__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_16_0__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_273
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_273__ap_start),
    .ap_done(PE_wrapper_273__ap_done),
    .ap_idle(PE_wrapper_273__ap_idle),
    .ap_ready(PE_wrapper_273__ap_ready),
    .idy(64'd1),
    .idx(64'd16),
    .fifo_A_in_s_dout(fifo_A_PE_16_1__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_16_1__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_16_1__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_16_1__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_16_1__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_16_2__din),
    .fifo_A_out_full_n(fifo_A_PE_16_2__full_n),
    .fifo_A_out_write(fifo_A_PE_16_2__write),
    .fifo_B_in_s_dout(fifo_B_PE_16_1__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_16_1__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_16_1__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_16_1__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_16_1__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_17_1__din),
    .fifo_B_out_full_n(fifo_B_PE_17_1__full_n),
    .fifo_B_out_write(fifo_B_PE_17_1__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_16_1__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_16_1__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_16_1__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_274
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_274__ap_start),
    .ap_done(PE_wrapper_274__ap_done),
    .ap_idle(PE_wrapper_274__ap_idle),
    .ap_ready(PE_wrapper_274__ap_ready),
    .idx(64'd16),
    .idy(64'd2),
    .fifo_A_in_s_dout(fifo_A_PE_16_2__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_16_2__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_16_2__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_16_2__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_16_2__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_16_3__din),
    .fifo_A_out_full_n(fifo_A_PE_16_3__full_n),
    .fifo_A_out_write(fifo_A_PE_16_3__write),
    .fifo_B_in_s_dout(fifo_B_PE_16_2__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_16_2__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_16_2__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_16_2__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_16_2__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_17_2__din),
    .fifo_B_out_full_n(fifo_B_PE_17_2__full_n),
    .fifo_B_out_write(fifo_B_PE_17_2__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_16_2__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_16_2__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_16_2__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_275
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_275__ap_start),
    .ap_done(PE_wrapper_275__ap_done),
    .ap_idle(PE_wrapper_275__ap_idle),
    .ap_ready(PE_wrapper_275__ap_ready),
    .idx(64'd16),
    .idy(64'd3),
    .fifo_A_in_s_dout(fifo_A_PE_16_3__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_16_3__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_16_3__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_16_3__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_16_3__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_16_4__din),
    .fifo_A_out_full_n(fifo_A_PE_16_4__full_n),
    .fifo_A_out_write(fifo_A_PE_16_4__write),
    .fifo_B_in_s_dout(fifo_B_PE_16_3__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_16_3__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_16_3__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_16_3__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_16_3__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_17_3__din),
    .fifo_B_out_full_n(fifo_B_PE_17_3__full_n),
    .fifo_B_out_write(fifo_B_PE_17_3__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_16_3__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_16_3__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_16_3__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_276
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_276__ap_start),
    .ap_done(PE_wrapper_276__ap_done),
    .ap_idle(PE_wrapper_276__ap_idle),
    .ap_ready(PE_wrapper_276__ap_ready),
    .idx(64'd16),
    .idy(64'd4),
    .fifo_A_in_s_dout(fifo_A_PE_16_4__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_16_4__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_16_4__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_16_4__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_16_4__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_16_5__din),
    .fifo_A_out_full_n(fifo_A_PE_16_5__full_n),
    .fifo_A_out_write(fifo_A_PE_16_5__write),
    .fifo_B_in_s_dout(fifo_B_PE_16_4__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_16_4__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_16_4__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_16_4__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_16_4__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_17_4__din),
    .fifo_B_out_full_n(fifo_B_PE_17_4__full_n),
    .fifo_B_out_write(fifo_B_PE_17_4__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_16_4__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_16_4__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_16_4__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_277
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_277__ap_start),
    .ap_done(PE_wrapper_277__ap_done),
    .ap_idle(PE_wrapper_277__ap_idle),
    .ap_ready(PE_wrapper_277__ap_ready),
    .idx(64'd16),
    .idy(64'd5),
    .fifo_A_in_s_dout(fifo_A_PE_16_5__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_16_5__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_16_5__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_16_5__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_16_5__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_16_6__din),
    .fifo_A_out_full_n(fifo_A_PE_16_6__full_n),
    .fifo_A_out_write(fifo_A_PE_16_6__write),
    .fifo_B_in_s_dout(fifo_B_PE_16_5__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_16_5__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_16_5__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_16_5__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_16_5__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_17_5__din),
    .fifo_B_out_full_n(fifo_B_PE_17_5__full_n),
    .fifo_B_out_write(fifo_B_PE_17_5__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_16_5__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_16_5__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_16_5__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_278
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_278__ap_start),
    .ap_done(PE_wrapper_278__ap_done),
    .ap_idle(PE_wrapper_278__ap_idle),
    .ap_ready(PE_wrapper_278__ap_ready),
    .idx(64'd16),
    .idy(64'd6),
    .fifo_A_in_s_dout(fifo_A_PE_16_6__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_16_6__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_16_6__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_16_6__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_16_6__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_16_7__din),
    .fifo_A_out_full_n(fifo_A_PE_16_7__full_n),
    .fifo_A_out_write(fifo_A_PE_16_7__write),
    .fifo_B_in_s_dout(fifo_B_PE_16_6__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_16_6__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_16_6__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_16_6__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_16_6__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_17_6__din),
    .fifo_B_out_full_n(fifo_B_PE_17_6__full_n),
    .fifo_B_out_write(fifo_B_PE_17_6__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_16_6__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_16_6__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_16_6__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_279
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_279__ap_start),
    .ap_done(PE_wrapper_279__ap_done),
    .ap_idle(PE_wrapper_279__ap_idle),
    .ap_ready(PE_wrapper_279__ap_ready),
    .idx(64'd16),
    .idy(64'd7),
    .fifo_A_in_s_dout(fifo_A_PE_16_7__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_16_7__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_16_7__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_16_7__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_16_7__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_16_8__din),
    .fifo_A_out_full_n(fifo_A_PE_16_8__full_n),
    .fifo_A_out_write(fifo_A_PE_16_8__write),
    .fifo_B_in_s_dout(fifo_B_PE_16_7__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_16_7__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_16_7__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_16_7__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_16_7__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_17_7__din),
    .fifo_B_out_full_n(fifo_B_PE_17_7__full_n),
    .fifo_B_out_write(fifo_B_PE_17_7__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_16_7__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_16_7__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_16_7__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_280
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_280__ap_start),
    .ap_done(PE_wrapper_280__ap_done),
    .ap_idle(PE_wrapper_280__ap_idle),
    .ap_ready(PE_wrapper_280__ap_ready),
    .idx(64'd16),
    .idy(64'd8),
    .fifo_A_in_s_dout(fifo_A_PE_16_8__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_16_8__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_16_8__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_16_8__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_16_8__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_16_9__din),
    .fifo_A_out_full_n(fifo_A_PE_16_9__full_n),
    .fifo_A_out_write(fifo_A_PE_16_9__write),
    .fifo_B_in_s_dout(fifo_B_PE_16_8__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_16_8__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_16_8__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_16_8__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_16_8__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_17_8__din),
    .fifo_B_out_full_n(fifo_B_PE_17_8__full_n),
    .fifo_B_out_write(fifo_B_PE_17_8__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_16_8__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_16_8__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_16_8__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_281
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_281__ap_start),
    .ap_done(PE_wrapper_281__ap_done),
    .ap_idle(PE_wrapper_281__ap_idle),
    .ap_ready(PE_wrapper_281__ap_ready),
    .idx(64'd16),
    .idy(64'd9),
    .fifo_A_out_din(fifo_A_PE_16_10__din),
    .fifo_A_out_full_n(fifo_A_PE_16_10__full_n),
    .fifo_A_out_write(fifo_A_PE_16_10__write),
    .fifo_A_in_s_dout(fifo_A_PE_16_9__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_16_9__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_16_9__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_16_9__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_16_9__read),
    .fifo_A_in_peek_read(),
    .fifo_B_in_s_dout(fifo_B_PE_16_9__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_16_9__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_16_9__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_16_9__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_16_9__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_17_9__din),
    .fifo_B_out_full_n(fifo_B_PE_17_9__full_n),
    .fifo_B_out_write(fifo_B_PE_17_9__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_16_9__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_16_9__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_16_9__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_282
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_282__ap_start),
    .ap_done(PE_wrapper_282__ap_done),
    .ap_idle(PE_wrapper_282__ap_idle),
    .ap_ready(PE_wrapper_282__ap_ready),
    .idy(64'd10),
    .idx(64'd16),
    .fifo_A_in_s_dout(fifo_A_PE_16_10__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_16_10__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_16_10__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_16_10__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_16_10__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_16_11__din),
    .fifo_A_out_full_n(fifo_A_PE_16_11__full_n),
    .fifo_A_out_write(fifo_A_PE_16_11__write),
    .fifo_B_in_s_dout(fifo_B_PE_16_10__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_16_10__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_16_10__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_16_10__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_16_10__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_17_10__din),
    .fifo_B_out_full_n(fifo_B_PE_17_10__full_n),
    .fifo_B_out_write(fifo_B_PE_17_10__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_16_10__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_16_10__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_16_10__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_283
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_283__ap_start),
    .ap_done(PE_wrapper_283__ap_done),
    .ap_idle(PE_wrapper_283__ap_idle),
    .ap_ready(PE_wrapper_283__ap_ready),
    .idy(64'd11),
    .idx(64'd16),
    .fifo_A_in_s_dout(fifo_A_PE_16_11__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_16_11__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_16_11__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_16_11__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_16_11__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_16_12__din),
    .fifo_A_out_full_n(fifo_A_PE_16_12__full_n),
    .fifo_A_out_write(fifo_A_PE_16_12__write),
    .fifo_B_in_s_dout(fifo_B_PE_16_11__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_16_11__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_16_11__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_16_11__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_16_11__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_17_11__din),
    .fifo_B_out_full_n(fifo_B_PE_17_11__full_n),
    .fifo_B_out_write(fifo_B_PE_17_11__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_16_11__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_16_11__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_16_11__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_284
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_284__ap_start),
    .ap_done(PE_wrapper_284__ap_done),
    .ap_idle(PE_wrapper_284__ap_idle),
    .ap_ready(PE_wrapper_284__ap_ready),
    .idy(64'd12),
    .idx(64'd16),
    .fifo_A_in_s_dout(fifo_A_PE_16_12__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_16_12__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_16_12__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_16_12__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_16_12__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_16_13__din),
    .fifo_A_out_full_n(fifo_A_PE_16_13__full_n),
    .fifo_A_out_write(fifo_A_PE_16_13__write),
    .fifo_B_in_s_dout(fifo_B_PE_16_12__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_16_12__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_16_12__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_16_12__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_16_12__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_17_12__din),
    .fifo_B_out_full_n(fifo_B_PE_17_12__full_n),
    .fifo_B_out_write(fifo_B_PE_17_12__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_16_12__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_16_12__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_16_12__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_285
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_285__ap_start),
    .ap_done(PE_wrapper_285__ap_done),
    .ap_idle(PE_wrapper_285__ap_idle),
    .ap_ready(PE_wrapper_285__ap_ready),
    .idy(64'd13),
    .idx(64'd16),
    .fifo_A_in_s_dout(fifo_A_PE_16_13__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_16_13__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_16_13__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_16_13__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_16_13__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_16_14__din),
    .fifo_A_out_full_n(fifo_A_PE_16_14__full_n),
    .fifo_A_out_write(fifo_A_PE_16_14__write),
    .fifo_B_in_s_dout(fifo_B_PE_16_13__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_16_13__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_16_13__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_16_13__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_16_13__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_17_13__din),
    .fifo_B_out_full_n(fifo_B_PE_17_13__full_n),
    .fifo_B_out_write(fifo_B_PE_17_13__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_16_13__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_16_13__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_16_13__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_286
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_286__ap_start),
    .ap_done(PE_wrapper_286__ap_done),
    .ap_idle(PE_wrapper_286__ap_idle),
    .ap_ready(PE_wrapper_286__ap_ready),
    .idy(64'd14),
    .idx(64'd16),
    .fifo_A_in_s_dout(fifo_A_PE_16_14__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_16_14__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_16_14__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_16_14__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_16_14__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_16_15__din),
    .fifo_A_out_full_n(fifo_A_PE_16_15__full_n),
    .fifo_A_out_write(fifo_A_PE_16_15__write),
    .fifo_B_in_s_dout(fifo_B_PE_16_14__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_16_14__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_16_14__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_16_14__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_16_14__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_17_14__din),
    .fifo_B_out_full_n(fifo_B_PE_17_14__full_n),
    .fifo_B_out_write(fifo_B_PE_17_14__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_16_14__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_16_14__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_16_14__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_287
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_287__ap_start),
    .ap_done(PE_wrapper_287__ap_done),
    .ap_idle(PE_wrapper_287__ap_idle),
    .ap_ready(PE_wrapper_287__ap_ready),
    .idy(64'd15),
    .idx(64'd16),
    .fifo_A_in_s_dout(fifo_A_PE_16_15__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_16_15__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_16_15__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_16_15__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_16_15__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_16_16__din),
    .fifo_A_out_full_n(fifo_A_PE_16_16__full_n),
    .fifo_A_out_write(fifo_A_PE_16_16__write),
    .fifo_B_in_s_dout(fifo_B_PE_16_15__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_16_15__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_16_15__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_16_15__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_16_15__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_17_15__din),
    .fifo_B_out_full_n(fifo_B_PE_17_15__full_n),
    .fifo_B_out_write(fifo_B_PE_17_15__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_16_15__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_16_15__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_16_15__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_288
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_288__ap_start),
    .ap_done(PE_wrapper_288__ap_done),
    .ap_idle(PE_wrapper_288__ap_idle),
    .ap_ready(PE_wrapper_288__ap_ready),
    .idx(64'd16),
    .idy(64'd16),
    .fifo_A_in_s_dout(fifo_A_PE_16_16__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_16_16__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_16_16__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_16_16__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_16_16__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_16_17__din),
    .fifo_A_out_full_n(fifo_A_PE_16_17__full_n),
    .fifo_A_out_write(fifo_A_PE_16_17__write),
    .fifo_B_in_s_dout(fifo_B_PE_16_16__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_16_16__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_16_16__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_16_16__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_16_16__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_17_16__din),
    .fifo_B_out_full_n(fifo_B_PE_17_16__full_n),
    .fifo_B_out_write(fifo_B_PE_17_16__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_16_16__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_16_16__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_16_16__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_289
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_289__ap_start),
    .ap_done(PE_wrapper_289__ap_done),
    .ap_idle(PE_wrapper_289__ap_idle),
    .ap_ready(PE_wrapper_289__ap_ready),
    .idy(64'd0),
    .idx(64'd17),
    .fifo_A_in_s_dout(fifo_A_PE_17_0__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_17_0__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_17_0__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_17_0__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_17_0__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_17_1__din),
    .fifo_A_out_full_n(fifo_A_PE_17_1__full_n),
    .fifo_A_out_write(fifo_A_PE_17_1__write),
    .fifo_B_in_s_dout(fifo_B_PE_17_0__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_17_0__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_17_0__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_17_0__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_17_0__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_18_0__din),
    .fifo_B_out_full_n(fifo_B_PE_18_0__full_n),
    .fifo_B_out_write(fifo_B_PE_18_0__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_17_0__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_17_0__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_17_0__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_290
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_290__ap_start),
    .ap_done(PE_wrapper_290__ap_done),
    .ap_idle(PE_wrapper_290__ap_idle),
    .ap_ready(PE_wrapper_290__ap_ready),
    .idy(64'd1),
    .idx(64'd17),
    .fifo_A_in_s_dout(fifo_A_PE_17_1__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_17_1__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_17_1__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_17_1__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_17_1__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_17_2__din),
    .fifo_A_out_full_n(fifo_A_PE_17_2__full_n),
    .fifo_A_out_write(fifo_A_PE_17_2__write),
    .fifo_B_in_s_dout(fifo_B_PE_17_1__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_17_1__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_17_1__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_17_1__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_17_1__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_18_1__din),
    .fifo_B_out_full_n(fifo_B_PE_18_1__full_n),
    .fifo_B_out_write(fifo_B_PE_18_1__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_17_1__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_17_1__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_17_1__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_291
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_291__ap_start),
    .ap_done(PE_wrapper_291__ap_done),
    .ap_idle(PE_wrapper_291__ap_idle),
    .ap_ready(PE_wrapper_291__ap_ready),
    .idx(64'd17),
    .idy(64'd2),
    .fifo_A_in_s_dout(fifo_A_PE_17_2__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_17_2__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_17_2__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_17_2__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_17_2__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_17_3__din),
    .fifo_A_out_full_n(fifo_A_PE_17_3__full_n),
    .fifo_A_out_write(fifo_A_PE_17_3__write),
    .fifo_B_in_s_dout(fifo_B_PE_17_2__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_17_2__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_17_2__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_17_2__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_17_2__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_18_2__din),
    .fifo_B_out_full_n(fifo_B_PE_18_2__full_n),
    .fifo_B_out_write(fifo_B_PE_18_2__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_17_2__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_17_2__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_17_2__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_292
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_292__ap_start),
    .ap_done(PE_wrapper_292__ap_done),
    .ap_idle(PE_wrapper_292__ap_idle),
    .ap_ready(PE_wrapper_292__ap_ready),
    .idx(64'd17),
    .idy(64'd3),
    .fifo_A_in_s_dout(fifo_A_PE_17_3__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_17_3__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_17_3__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_17_3__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_17_3__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_17_4__din),
    .fifo_A_out_full_n(fifo_A_PE_17_4__full_n),
    .fifo_A_out_write(fifo_A_PE_17_4__write),
    .fifo_B_in_s_dout(fifo_B_PE_17_3__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_17_3__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_17_3__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_17_3__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_17_3__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_18_3__din),
    .fifo_B_out_full_n(fifo_B_PE_18_3__full_n),
    .fifo_B_out_write(fifo_B_PE_18_3__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_17_3__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_17_3__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_17_3__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_293
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_293__ap_start),
    .ap_done(PE_wrapper_293__ap_done),
    .ap_idle(PE_wrapper_293__ap_idle),
    .ap_ready(PE_wrapper_293__ap_ready),
    .idx(64'd17),
    .idy(64'd4),
    .fifo_A_in_s_dout(fifo_A_PE_17_4__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_17_4__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_17_4__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_17_4__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_17_4__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_17_5__din),
    .fifo_A_out_full_n(fifo_A_PE_17_5__full_n),
    .fifo_A_out_write(fifo_A_PE_17_5__write),
    .fifo_B_in_s_dout(fifo_B_PE_17_4__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_17_4__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_17_4__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_17_4__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_17_4__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_18_4__din),
    .fifo_B_out_full_n(fifo_B_PE_18_4__full_n),
    .fifo_B_out_write(fifo_B_PE_18_4__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_17_4__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_17_4__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_17_4__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_294
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_294__ap_start),
    .ap_done(PE_wrapper_294__ap_done),
    .ap_idle(PE_wrapper_294__ap_idle),
    .ap_ready(PE_wrapper_294__ap_ready),
    .idx(64'd17),
    .idy(64'd5),
    .fifo_A_in_s_dout(fifo_A_PE_17_5__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_17_5__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_17_5__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_17_5__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_17_5__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_17_6__din),
    .fifo_A_out_full_n(fifo_A_PE_17_6__full_n),
    .fifo_A_out_write(fifo_A_PE_17_6__write),
    .fifo_B_in_s_dout(fifo_B_PE_17_5__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_17_5__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_17_5__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_17_5__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_17_5__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_18_5__din),
    .fifo_B_out_full_n(fifo_B_PE_18_5__full_n),
    .fifo_B_out_write(fifo_B_PE_18_5__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_17_5__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_17_5__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_17_5__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_295
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_295__ap_start),
    .ap_done(PE_wrapper_295__ap_done),
    .ap_idle(PE_wrapper_295__ap_idle),
    .ap_ready(PE_wrapper_295__ap_ready),
    .idx(64'd17),
    .idy(64'd6),
    .fifo_A_in_s_dout(fifo_A_PE_17_6__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_17_6__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_17_6__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_17_6__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_17_6__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_17_7__din),
    .fifo_A_out_full_n(fifo_A_PE_17_7__full_n),
    .fifo_A_out_write(fifo_A_PE_17_7__write),
    .fifo_B_in_s_dout(fifo_B_PE_17_6__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_17_6__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_17_6__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_17_6__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_17_6__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_18_6__din),
    .fifo_B_out_full_n(fifo_B_PE_18_6__full_n),
    .fifo_B_out_write(fifo_B_PE_18_6__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_17_6__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_17_6__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_17_6__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_296
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_296__ap_start),
    .ap_done(PE_wrapper_296__ap_done),
    .ap_idle(PE_wrapper_296__ap_idle),
    .ap_ready(PE_wrapper_296__ap_ready),
    .idx(64'd17),
    .idy(64'd7),
    .fifo_A_in_s_dout(fifo_A_PE_17_7__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_17_7__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_17_7__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_17_7__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_17_7__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_17_8__din),
    .fifo_A_out_full_n(fifo_A_PE_17_8__full_n),
    .fifo_A_out_write(fifo_A_PE_17_8__write),
    .fifo_B_in_s_dout(fifo_B_PE_17_7__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_17_7__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_17_7__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_17_7__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_17_7__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_18_7__din),
    .fifo_B_out_full_n(fifo_B_PE_18_7__full_n),
    .fifo_B_out_write(fifo_B_PE_18_7__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_17_7__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_17_7__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_17_7__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_297
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_297__ap_start),
    .ap_done(PE_wrapper_297__ap_done),
    .ap_idle(PE_wrapper_297__ap_idle),
    .ap_ready(PE_wrapper_297__ap_ready),
    .idx(64'd17),
    .idy(64'd8),
    .fifo_A_in_s_dout(fifo_A_PE_17_8__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_17_8__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_17_8__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_17_8__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_17_8__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_17_9__din),
    .fifo_A_out_full_n(fifo_A_PE_17_9__full_n),
    .fifo_A_out_write(fifo_A_PE_17_9__write),
    .fifo_B_in_s_dout(fifo_B_PE_17_8__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_17_8__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_17_8__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_17_8__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_17_8__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_18_8__din),
    .fifo_B_out_full_n(fifo_B_PE_18_8__full_n),
    .fifo_B_out_write(fifo_B_PE_18_8__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_17_8__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_17_8__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_17_8__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_298
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_298__ap_start),
    .ap_done(PE_wrapper_298__ap_done),
    .ap_idle(PE_wrapper_298__ap_idle),
    .ap_ready(PE_wrapper_298__ap_ready),
    .idx(64'd17),
    .idy(64'd9),
    .fifo_A_out_din(fifo_A_PE_17_10__din),
    .fifo_A_out_full_n(fifo_A_PE_17_10__full_n),
    .fifo_A_out_write(fifo_A_PE_17_10__write),
    .fifo_A_in_s_dout(fifo_A_PE_17_9__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_17_9__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_17_9__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_17_9__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_17_9__read),
    .fifo_A_in_peek_read(),
    .fifo_B_in_s_dout(fifo_B_PE_17_9__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_17_9__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_17_9__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_17_9__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_17_9__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_18_9__din),
    .fifo_B_out_full_n(fifo_B_PE_18_9__full_n),
    .fifo_B_out_write(fifo_B_PE_18_9__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_17_9__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_17_9__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_17_9__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_299
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_299__ap_start),
    .ap_done(PE_wrapper_299__ap_done),
    .ap_idle(PE_wrapper_299__ap_idle),
    .ap_ready(PE_wrapper_299__ap_ready),
    .idy(64'd10),
    .idx(64'd17),
    .fifo_A_in_s_dout(fifo_A_PE_17_10__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_17_10__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_17_10__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_17_10__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_17_10__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_17_11__din),
    .fifo_A_out_full_n(fifo_A_PE_17_11__full_n),
    .fifo_A_out_write(fifo_A_PE_17_11__write),
    .fifo_B_in_s_dout(fifo_B_PE_17_10__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_17_10__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_17_10__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_17_10__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_17_10__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_18_10__din),
    .fifo_B_out_full_n(fifo_B_PE_18_10__full_n),
    .fifo_B_out_write(fifo_B_PE_18_10__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_17_10__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_17_10__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_17_10__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_300
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_300__ap_start),
    .ap_done(PE_wrapper_300__ap_done),
    .ap_idle(PE_wrapper_300__ap_idle),
    .ap_ready(PE_wrapper_300__ap_ready),
    .idy(64'd11),
    .idx(64'd17),
    .fifo_A_in_s_dout(fifo_A_PE_17_11__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_17_11__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_17_11__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_17_11__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_17_11__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_17_12__din),
    .fifo_A_out_full_n(fifo_A_PE_17_12__full_n),
    .fifo_A_out_write(fifo_A_PE_17_12__write),
    .fifo_B_in_s_dout(fifo_B_PE_17_11__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_17_11__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_17_11__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_17_11__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_17_11__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_18_11__din),
    .fifo_B_out_full_n(fifo_B_PE_18_11__full_n),
    .fifo_B_out_write(fifo_B_PE_18_11__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_17_11__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_17_11__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_17_11__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_301
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_301__ap_start),
    .ap_done(PE_wrapper_301__ap_done),
    .ap_idle(PE_wrapper_301__ap_idle),
    .ap_ready(PE_wrapper_301__ap_ready),
    .idy(64'd12),
    .idx(64'd17),
    .fifo_A_in_s_dout(fifo_A_PE_17_12__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_17_12__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_17_12__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_17_12__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_17_12__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_17_13__din),
    .fifo_A_out_full_n(fifo_A_PE_17_13__full_n),
    .fifo_A_out_write(fifo_A_PE_17_13__write),
    .fifo_B_in_s_dout(fifo_B_PE_17_12__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_17_12__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_17_12__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_17_12__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_17_12__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_18_12__din),
    .fifo_B_out_full_n(fifo_B_PE_18_12__full_n),
    .fifo_B_out_write(fifo_B_PE_18_12__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_17_12__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_17_12__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_17_12__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_302
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_302__ap_start),
    .ap_done(PE_wrapper_302__ap_done),
    .ap_idle(PE_wrapper_302__ap_idle),
    .ap_ready(PE_wrapper_302__ap_ready),
    .idy(64'd13),
    .idx(64'd17),
    .fifo_A_in_s_dout(fifo_A_PE_17_13__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_17_13__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_17_13__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_17_13__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_17_13__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_17_14__din),
    .fifo_A_out_full_n(fifo_A_PE_17_14__full_n),
    .fifo_A_out_write(fifo_A_PE_17_14__write),
    .fifo_B_in_s_dout(fifo_B_PE_17_13__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_17_13__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_17_13__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_17_13__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_17_13__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_18_13__din),
    .fifo_B_out_full_n(fifo_B_PE_18_13__full_n),
    .fifo_B_out_write(fifo_B_PE_18_13__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_17_13__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_17_13__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_17_13__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_303
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_303__ap_start),
    .ap_done(PE_wrapper_303__ap_done),
    .ap_idle(PE_wrapper_303__ap_idle),
    .ap_ready(PE_wrapper_303__ap_ready),
    .idy(64'd14),
    .idx(64'd17),
    .fifo_A_in_s_dout(fifo_A_PE_17_14__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_17_14__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_17_14__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_17_14__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_17_14__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_17_15__din),
    .fifo_A_out_full_n(fifo_A_PE_17_15__full_n),
    .fifo_A_out_write(fifo_A_PE_17_15__write),
    .fifo_B_in_s_dout(fifo_B_PE_17_14__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_17_14__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_17_14__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_17_14__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_17_14__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_18_14__din),
    .fifo_B_out_full_n(fifo_B_PE_18_14__full_n),
    .fifo_B_out_write(fifo_B_PE_18_14__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_17_14__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_17_14__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_17_14__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_304
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_304__ap_start),
    .ap_done(PE_wrapper_304__ap_done),
    .ap_idle(PE_wrapper_304__ap_idle),
    .ap_ready(PE_wrapper_304__ap_ready),
    .idy(64'd15),
    .idx(64'd17),
    .fifo_A_in_s_dout(fifo_A_PE_17_15__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_17_15__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_17_15__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_17_15__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_17_15__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_17_16__din),
    .fifo_A_out_full_n(fifo_A_PE_17_16__full_n),
    .fifo_A_out_write(fifo_A_PE_17_16__write),
    .fifo_B_in_s_dout(fifo_B_PE_17_15__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_17_15__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_17_15__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_17_15__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_17_15__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_18_15__din),
    .fifo_B_out_full_n(fifo_B_PE_18_15__full_n),
    .fifo_B_out_write(fifo_B_PE_18_15__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_17_15__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_17_15__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_17_15__write)
  );


  (* keep_hierarchy = "yes" *) PE_wrapper
  PE_wrapper_305
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(PE_wrapper_305__ap_start),
    .ap_done(PE_wrapper_305__ap_done),
    .ap_idle(PE_wrapper_305__ap_idle),
    .ap_ready(PE_wrapper_305__ap_ready),
    .idy(64'd16),
    .idx(64'd17),
    .fifo_A_in_s_dout(fifo_A_PE_17_16__dout),
    .fifo_A_in_peek_dout(fifo_A_PE_17_16__dout),
    .fifo_A_in_s_empty_n(fifo_A_PE_17_16__empty_n),
    .fifo_A_in_peek_empty_n(fifo_A_PE_17_16__empty_n),
    .fifo_A_in_s_read(fifo_A_PE_17_16__read),
    .fifo_A_in_peek_read(),
    .fifo_A_out_din(fifo_A_PE_17_17__din),
    .fifo_A_out_full_n(fifo_A_PE_17_17__full_n),
    .fifo_A_out_write(fifo_A_PE_17_17__write),
    .fifo_B_in_s_dout(fifo_B_PE_17_16__dout),
    .fifo_B_in_peek_dout(fifo_B_PE_17_16__dout),
    .fifo_B_in_s_empty_n(fifo_B_PE_17_16__empty_n),
    .fifo_B_in_peek_empty_n(fifo_B_PE_17_16__empty_n),
    .fifo_B_in_s_read(fifo_B_PE_17_16__read),
    .fifo_B_in_peek_read(),
    .fifo_B_out_din(fifo_B_PE_18_16__din),
    .fifo_B_out_full_n(fifo_B_PE_18_16__full_n),
    .fifo_B_out_write(fifo_B_PE_18_16__write),
    .fifo_C_drain_out_din(fifo_C_drain_PE_17_16__din),
    .fifo_C_drain_out_full_n(fifo_C_drain_PE_17_16__full_n),
    .fifo_C_drain_out_write(fifo_C_drain_PE_17_16__write)
  );


  (* keep_hierarchy = "yes" *) kernel0_fsm
  __tapa_fsm_unit
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(ap_start),
    .ap_done(ap_done),
    .ap_idle(ap_idle),
    .ap_ready(ap_ready),
    .A(A),
    .B(B),
    .C(C),
    .A_IO_L2_in_0__ap_start(A_IO_L2_in_0__ap_start),
    .A_IO_L2_in_0__ap_ready(A_IO_L2_in_0__ap_ready),
    .A_IO_L2_in_0__ap_done(A_IO_L2_in_0__ap_done),
    .A_IO_L2_in_0__ap_idle(A_IO_L2_in_0__ap_idle),
    .A_IO_L2_in_1__ap_start(A_IO_L2_in_1__ap_start),
    .A_IO_L2_in_1__ap_ready(A_IO_L2_in_1__ap_ready),
    .A_IO_L2_in_1__ap_done(A_IO_L2_in_1__ap_done),
    .A_IO_L2_in_1__ap_idle(A_IO_L2_in_1__ap_idle),
    .A_IO_L2_in_2__ap_start(A_IO_L2_in_2__ap_start),
    .A_IO_L2_in_2__ap_ready(A_IO_L2_in_2__ap_ready),
    .A_IO_L2_in_2__ap_done(A_IO_L2_in_2__ap_done),
    .A_IO_L2_in_2__ap_idle(A_IO_L2_in_2__ap_idle),
    .A_IO_L2_in_3__ap_start(A_IO_L2_in_3__ap_start),
    .A_IO_L2_in_3__ap_ready(A_IO_L2_in_3__ap_ready),
    .A_IO_L2_in_3__ap_done(A_IO_L2_in_3__ap_done),
    .A_IO_L2_in_3__ap_idle(A_IO_L2_in_3__ap_idle),
    .A_IO_L2_in_4__ap_start(A_IO_L2_in_4__ap_start),
    .A_IO_L2_in_4__ap_ready(A_IO_L2_in_4__ap_ready),
    .A_IO_L2_in_4__ap_done(A_IO_L2_in_4__ap_done),
    .A_IO_L2_in_4__ap_idle(A_IO_L2_in_4__ap_idle),
    .A_IO_L2_in_5__ap_start(A_IO_L2_in_5__ap_start),
    .A_IO_L2_in_5__ap_ready(A_IO_L2_in_5__ap_ready),
    .A_IO_L2_in_5__ap_done(A_IO_L2_in_5__ap_done),
    .A_IO_L2_in_5__ap_idle(A_IO_L2_in_5__ap_idle),
    .A_IO_L2_in_6__ap_start(A_IO_L2_in_6__ap_start),
    .A_IO_L2_in_6__ap_ready(A_IO_L2_in_6__ap_ready),
    .A_IO_L2_in_6__ap_done(A_IO_L2_in_6__ap_done),
    .A_IO_L2_in_6__ap_idle(A_IO_L2_in_6__ap_idle),
    .A_IO_L2_in_7__ap_start(A_IO_L2_in_7__ap_start),
    .A_IO_L2_in_7__ap_ready(A_IO_L2_in_7__ap_ready),
    .A_IO_L2_in_7__ap_done(A_IO_L2_in_7__ap_done),
    .A_IO_L2_in_7__ap_idle(A_IO_L2_in_7__ap_idle),
    .A_IO_L2_in_8__ap_start(A_IO_L2_in_8__ap_start),
    .A_IO_L2_in_8__ap_ready(A_IO_L2_in_8__ap_ready),
    .A_IO_L2_in_8__ap_done(A_IO_L2_in_8__ap_done),
    .A_IO_L2_in_8__ap_idle(A_IO_L2_in_8__ap_idle),
    .A_IO_L2_in_9__ap_start(A_IO_L2_in_9__ap_start),
    .A_IO_L2_in_9__ap_ready(A_IO_L2_in_9__ap_ready),
    .A_IO_L2_in_9__ap_done(A_IO_L2_in_9__ap_done),
    .A_IO_L2_in_9__ap_idle(A_IO_L2_in_9__ap_idle),
    .A_IO_L2_in_10__ap_start(A_IO_L2_in_10__ap_start),
    .A_IO_L2_in_10__ap_ready(A_IO_L2_in_10__ap_ready),
    .A_IO_L2_in_10__ap_done(A_IO_L2_in_10__ap_done),
    .A_IO_L2_in_10__ap_idle(A_IO_L2_in_10__ap_idle),
    .A_IO_L2_in_11__ap_start(A_IO_L2_in_11__ap_start),
    .A_IO_L2_in_11__ap_ready(A_IO_L2_in_11__ap_ready),
    .A_IO_L2_in_11__ap_done(A_IO_L2_in_11__ap_done),
    .A_IO_L2_in_11__ap_idle(A_IO_L2_in_11__ap_idle),
    .A_IO_L2_in_12__ap_start(A_IO_L2_in_12__ap_start),
    .A_IO_L2_in_12__ap_ready(A_IO_L2_in_12__ap_ready),
    .A_IO_L2_in_12__ap_done(A_IO_L2_in_12__ap_done),
    .A_IO_L2_in_12__ap_idle(A_IO_L2_in_12__ap_idle),
    .A_IO_L2_in_13__ap_start(A_IO_L2_in_13__ap_start),
    .A_IO_L2_in_13__ap_ready(A_IO_L2_in_13__ap_ready),
    .A_IO_L2_in_13__ap_done(A_IO_L2_in_13__ap_done),
    .A_IO_L2_in_13__ap_idle(A_IO_L2_in_13__ap_idle),
    .A_IO_L2_in_14__ap_start(A_IO_L2_in_14__ap_start),
    .A_IO_L2_in_14__ap_ready(A_IO_L2_in_14__ap_ready),
    .A_IO_L2_in_14__ap_done(A_IO_L2_in_14__ap_done),
    .A_IO_L2_in_14__ap_idle(A_IO_L2_in_14__ap_idle),
    .A_IO_L2_in_15__ap_start(A_IO_L2_in_15__ap_start),
    .A_IO_L2_in_15__ap_ready(A_IO_L2_in_15__ap_ready),
    .A_IO_L2_in_15__ap_done(A_IO_L2_in_15__ap_done),
    .A_IO_L2_in_15__ap_idle(A_IO_L2_in_15__ap_idle),
    .A_IO_L2_in_16__ap_start(A_IO_L2_in_16__ap_start),
    .A_IO_L2_in_16__ap_ready(A_IO_L2_in_16__ap_ready),
    .A_IO_L2_in_16__ap_done(A_IO_L2_in_16__ap_done),
    .A_IO_L2_in_16__ap_idle(A_IO_L2_in_16__ap_idle),
    .A_IO_L2_in_boundary_0__ap_start(A_IO_L2_in_boundary_0__ap_start),
    .A_IO_L2_in_boundary_0__ap_ready(A_IO_L2_in_boundary_0__ap_ready),
    .A_IO_L2_in_boundary_0__ap_done(A_IO_L2_in_boundary_0__ap_done),
    .A_IO_L2_in_boundary_0__ap_idle(A_IO_L2_in_boundary_0__ap_idle),
    .A_IO_L3_in_0__ap_start(A_IO_L3_in_0__ap_start),
    .A_IO_L3_in_0__ap_ready(A_IO_L3_in_0__ap_ready),
    .A_IO_L3_in_0__ap_done(A_IO_L3_in_0__ap_done),
    .A_IO_L3_in_0__ap_idle(A_IO_L3_in_0__ap_idle),
    .A_IO_L3_in_serialize_0___A__q0(A_IO_L3_in_serialize_0___A__q0),
    .A_IO_L3_in_serialize_0__ap_start(A_IO_L3_in_serialize_0__ap_start),
    .A_IO_L3_in_serialize_0__ap_ready(A_IO_L3_in_serialize_0__ap_ready),
    .A_IO_L3_in_serialize_0__ap_done(A_IO_L3_in_serialize_0__ap_done),
    .A_IO_L3_in_serialize_0__ap_idle(A_IO_L3_in_serialize_0__ap_idle),
    .A_PE_dummy_in_0__ap_start(A_PE_dummy_in_0__ap_start),
    .A_PE_dummy_in_0__ap_ready(A_PE_dummy_in_0__ap_ready),
    .A_PE_dummy_in_0__ap_done(A_PE_dummy_in_0__ap_done),
    .A_PE_dummy_in_0__ap_idle(A_PE_dummy_in_0__ap_idle),
    .A_PE_dummy_in_1__ap_start(A_PE_dummy_in_1__ap_start),
    .A_PE_dummy_in_1__ap_ready(A_PE_dummy_in_1__ap_ready),
    .A_PE_dummy_in_1__ap_done(A_PE_dummy_in_1__ap_done),
    .A_PE_dummy_in_1__ap_idle(A_PE_dummy_in_1__ap_idle),
    .A_PE_dummy_in_2__ap_start(A_PE_dummy_in_2__ap_start),
    .A_PE_dummy_in_2__ap_ready(A_PE_dummy_in_2__ap_ready),
    .A_PE_dummy_in_2__ap_done(A_PE_dummy_in_2__ap_done),
    .A_PE_dummy_in_2__ap_idle(A_PE_dummy_in_2__ap_idle),
    .A_PE_dummy_in_3__ap_start(A_PE_dummy_in_3__ap_start),
    .A_PE_dummy_in_3__ap_ready(A_PE_dummy_in_3__ap_ready),
    .A_PE_dummy_in_3__ap_done(A_PE_dummy_in_3__ap_done),
    .A_PE_dummy_in_3__ap_idle(A_PE_dummy_in_3__ap_idle),
    .A_PE_dummy_in_4__ap_start(A_PE_dummy_in_4__ap_start),
    .A_PE_dummy_in_4__ap_ready(A_PE_dummy_in_4__ap_ready),
    .A_PE_dummy_in_4__ap_done(A_PE_dummy_in_4__ap_done),
    .A_PE_dummy_in_4__ap_idle(A_PE_dummy_in_4__ap_idle),
    .A_PE_dummy_in_5__ap_start(A_PE_dummy_in_5__ap_start),
    .A_PE_dummy_in_5__ap_ready(A_PE_dummy_in_5__ap_ready),
    .A_PE_dummy_in_5__ap_done(A_PE_dummy_in_5__ap_done),
    .A_PE_dummy_in_5__ap_idle(A_PE_dummy_in_5__ap_idle),
    .A_PE_dummy_in_6__ap_start(A_PE_dummy_in_6__ap_start),
    .A_PE_dummy_in_6__ap_ready(A_PE_dummy_in_6__ap_ready),
    .A_PE_dummy_in_6__ap_done(A_PE_dummy_in_6__ap_done),
    .A_PE_dummy_in_6__ap_idle(A_PE_dummy_in_6__ap_idle),
    .A_PE_dummy_in_7__ap_start(A_PE_dummy_in_7__ap_start),
    .A_PE_dummy_in_7__ap_ready(A_PE_dummy_in_7__ap_ready),
    .A_PE_dummy_in_7__ap_done(A_PE_dummy_in_7__ap_done),
    .A_PE_dummy_in_7__ap_idle(A_PE_dummy_in_7__ap_idle),
    .A_PE_dummy_in_8__ap_start(A_PE_dummy_in_8__ap_start),
    .A_PE_dummy_in_8__ap_ready(A_PE_dummy_in_8__ap_ready),
    .A_PE_dummy_in_8__ap_done(A_PE_dummy_in_8__ap_done),
    .A_PE_dummy_in_8__ap_idle(A_PE_dummy_in_8__ap_idle),
    .A_PE_dummy_in_9__ap_start(A_PE_dummy_in_9__ap_start),
    .A_PE_dummy_in_9__ap_ready(A_PE_dummy_in_9__ap_ready),
    .A_PE_dummy_in_9__ap_done(A_PE_dummy_in_9__ap_done),
    .A_PE_dummy_in_9__ap_idle(A_PE_dummy_in_9__ap_idle),
    .A_PE_dummy_in_10__ap_start(A_PE_dummy_in_10__ap_start),
    .A_PE_dummy_in_10__ap_ready(A_PE_dummy_in_10__ap_ready),
    .A_PE_dummy_in_10__ap_done(A_PE_dummy_in_10__ap_done),
    .A_PE_dummy_in_10__ap_idle(A_PE_dummy_in_10__ap_idle),
    .A_PE_dummy_in_11__ap_start(A_PE_dummy_in_11__ap_start),
    .A_PE_dummy_in_11__ap_ready(A_PE_dummy_in_11__ap_ready),
    .A_PE_dummy_in_11__ap_done(A_PE_dummy_in_11__ap_done),
    .A_PE_dummy_in_11__ap_idle(A_PE_dummy_in_11__ap_idle),
    .A_PE_dummy_in_12__ap_start(A_PE_dummy_in_12__ap_start),
    .A_PE_dummy_in_12__ap_ready(A_PE_dummy_in_12__ap_ready),
    .A_PE_dummy_in_12__ap_done(A_PE_dummy_in_12__ap_done),
    .A_PE_dummy_in_12__ap_idle(A_PE_dummy_in_12__ap_idle),
    .A_PE_dummy_in_13__ap_start(A_PE_dummy_in_13__ap_start),
    .A_PE_dummy_in_13__ap_ready(A_PE_dummy_in_13__ap_ready),
    .A_PE_dummy_in_13__ap_done(A_PE_dummy_in_13__ap_done),
    .A_PE_dummy_in_13__ap_idle(A_PE_dummy_in_13__ap_idle),
    .A_PE_dummy_in_14__ap_start(A_PE_dummy_in_14__ap_start),
    .A_PE_dummy_in_14__ap_ready(A_PE_dummy_in_14__ap_ready),
    .A_PE_dummy_in_14__ap_done(A_PE_dummy_in_14__ap_done),
    .A_PE_dummy_in_14__ap_idle(A_PE_dummy_in_14__ap_idle),
    .A_PE_dummy_in_15__ap_start(A_PE_dummy_in_15__ap_start),
    .A_PE_dummy_in_15__ap_ready(A_PE_dummy_in_15__ap_ready),
    .A_PE_dummy_in_15__ap_done(A_PE_dummy_in_15__ap_done),
    .A_PE_dummy_in_15__ap_idle(A_PE_dummy_in_15__ap_idle),
    .A_PE_dummy_in_16__ap_start(A_PE_dummy_in_16__ap_start),
    .A_PE_dummy_in_16__ap_ready(A_PE_dummy_in_16__ap_ready),
    .A_PE_dummy_in_16__ap_done(A_PE_dummy_in_16__ap_done),
    .A_PE_dummy_in_16__ap_idle(A_PE_dummy_in_16__ap_idle),
    .A_PE_dummy_in_17__ap_start(A_PE_dummy_in_17__ap_start),
    .A_PE_dummy_in_17__ap_ready(A_PE_dummy_in_17__ap_ready),
    .A_PE_dummy_in_17__ap_done(A_PE_dummy_in_17__ap_done),
    .A_PE_dummy_in_17__ap_idle(A_PE_dummy_in_17__ap_idle),
    .B_IO_L2_in_0__ap_start(B_IO_L2_in_0__ap_start),
    .B_IO_L2_in_0__ap_ready(B_IO_L2_in_0__ap_ready),
    .B_IO_L2_in_0__ap_done(B_IO_L2_in_0__ap_done),
    .B_IO_L2_in_0__ap_idle(B_IO_L2_in_0__ap_idle),
    .B_IO_L2_in_1__ap_start(B_IO_L2_in_1__ap_start),
    .B_IO_L2_in_1__ap_ready(B_IO_L2_in_1__ap_ready),
    .B_IO_L2_in_1__ap_done(B_IO_L2_in_1__ap_done),
    .B_IO_L2_in_1__ap_idle(B_IO_L2_in_1__ap_idle),
    .B_IO_L2_in_2__ap_start(B_IO_L2_in_2__ap_start),
    .B_IO_L2_in_2__ap_ready(B_IO_L2_in_2__ap_ready),
    .B_IO_L2_in_2__ap_done(B_IO_L2_in_2__ap_done),
    .B_IO_L2_in_2__ap_idle(B_IO_L2_in_2__ap_idle),
    .B_IO_L2_in_3__ap_start(B_IO_L2_in_3__ap_start),
    .B_IO_L2_in_3__ap_ready(B_IO_L2_in_3__ap_ready),
    .B_IO_L2_in_3__ap_done(B_IO_L2_in_3__ap_done),
    .B_IO_L2_in_3__ap_idle(B_IO_L2_in_3__ap_idle),
    .B_IO_L2_in_4__ap_start(B_IO_L2_in_4__ap_start),
    .B_IO_L2_in_4__ap_ready(B_IO_L2_in_4__ap_ready),
    .B_IO_L2_in_4__ap_done(B_IO_L2_in_4__ap_done),
    .B_IO_L2_in_4__ap_idle(B_IO_L2_in_4__ap_idle),
    .B_IO_L2_in_5__ap_start(B_IO_L2_in_5__ap_start),
    .B_IO_L2_in_5__ap_ready(B_IO_L2_in_5__ap_ready),
    .B_IO_L2_in_5__ap_done(B_IO_L2_in_5__ap_done),
    .B_IO_L2_in_5__ap_idle(B_IO_L2_in_5__ap_idle),
    .B_IO_L2_in_6__ap_start(B_IO_L2_in_6__ap_start),
    .B_IO_L2_in_6__ap_ready(B_IO_L2_in_6__ap_ready),
    .B_IO_L2_in_6__ap_done(B_IO_L2_in_6__ap_done),
    .B_IO_L2_in_6__ap_idle(B_IO_L2_in_6__ap_idle),
    .B_IO_L2_in_7__ap_start(B_IO_L2_in_7__ap_start),
    .B_IO_L2_in_7__ap_ready(B_IO_L2_in_7__ap_ready),
    .B_IO_L2_in_7__ap_done(B_IO_L2_in_7__ap_done),
    .B_IO_L2_in_7__ap_idle(B_IO_L2_in_7__ap_idle),
    .B_IO_L2_in_8__ap_start(B_IO_L2_in_8__ap_start),
    .B_IO_L2_in_8__ap_ready(B_IO_L2_in_8__ap_ready),
    .B_IO_L2_in_8__ap_done(B_IO_L2_in_8__ap_done),
    .B_IO_L2_in_8__ap_idle(B_IO_L2_in_8__ap_idle),
    .B_IO_L2_in_9__ap_start(B_IO_L2_in_9__ap_start),
    .B_IO_L2_in_9__ap_ready(B_IO_L2_in_9__ap_ready),
    .B_IO_L2_in_9__ap_done(B_IO_L2_in_9__ap_done),
    .B_IO_L2_in_9__ap_idle(B_IO_L2_in_9__ap_idle),
    .B_IO_L2_in_10__ap_start(B_IO_L2_in_10__ap_start),
    .B_IO_L2_in_10__ap_ready(B_IO_L2_in_10__ap_ready),
    .B_IO_L2_in_10__ap_done(B_IO_L2_in_10__ap_done),
    .B_IO_L2_in_10__ap_idle(B_IO_L2_in_10__ap_idle),
    .B_IO_L2_in_11__ap_start(B_IO_L2_in_11__ap_start),
    .B_IO_L2_in_11__ap_ready(B_IO_L2_in_11__ap_ready),
    .B_IO_L2_in_11__ap_done(B_IO_L2_in_11__ap_done),
    .B_IO_L2_in_11__ap_idle(B_IO_L2_in_11__ap_idle),
    .B_IO_L2_in_12__ap_start(B_IO_L2_in_12__ap_start),
    .B_IO_L2_in_12__ap_ready(B_IO_L2_in_12__ap_ready),
    .B_IO_L2_in_12__ap_done(B_IO_L2_in_12__ap_done),
    .B_IO_L2_in_12__ap_idle(B_IO_L2_in_12__ap_idle),
    .B_IO_L2_in_13__ap_start(B_IO_L2_in_13__ap_start),
    .B_IO_L2_in_13__ap_ready(B_IO_L2_in_13__ap_ready),
    .B_IO_L2_in_13__ap_done(B_IO_L2_in_13__ap_done),
    .B_IO_L2_in_13__ap_idle(B_IO_L2_in_13__ap_idle),
    .B_IO_L2_in_14__ap_start(B_IO_L2_in_14__ap_start),
    .B_IO_L2_in_14__ap_ready(B_IO_L2_in_14__ap_ready),
    .B_IO_L2_in_14__ap_done(B_IO_L2_in_14__ap_done),
    .B_IO_L2_in_14__ap_idle(B_IO_L2_in_14__ap_idle),
    .B_IO_L2_in_15__ap_start(B_IO_L2_in_15__ap_start),
    .B_IO_L2_in_15__ap_ready(B_IO_L2_in_15__ap_ready),
    .B_IO_L2_in_15__ap_done(B_IO_L2_in_15__ap_done),
    .B_IO_L2_in_15__ap_idle(B_IO_L2_in_15__ap_idle),
    .B_IO_L2_in_boundary_0__ap_start(B_IO_L2_in_boundary_0__ap_start),
    .B_IO_L2_in_boundary_0__ap_ready(B_IO_L2_in_boundary_0__ap_ready),
    .B_IO_L2_in_boundary_0__ap_done(B_IO_L2_in_boundary_0__ap_done),
    .B_IO_L2_in_boundary_0__ap_idle(B_IO_L2_in_boundary_0__ap_idle),
    .B_IO_L3_in_0__ap_start(B_IO_L3_in_0__ap_start),
    .B_IO_L3_in_0__ap_ready(B_IO_L3_in_0__ap_ready),
    .B_IO_L3_in_0__ap_done(B_IO_L3_in_0__ap_done),
    .B_IO_L3_in_0__ap_idle(B_IO_L3_in_0__ap_idle),
    .B_IO_L3_in_serialize_0___B__q0(B_IO_L3_in_serialize_0___B__q0),
    .B_IO_L3_in_serialize_0__ap_start(B_IO_L3_in_serialize_0__ap_start),
    .B_IO_L3_in_serialize_0__ap_ready(B_IO_L3_in_serialize_0__ap_ready),
    .B_IO_L3_in_serialize_0__ap_done(B_IO_L3_in_serialize_0__ap_done),
    .B_IO_L3_in_serialize_0__ap_idle(B_IO_L3_in_serialize_0__ap_idle),
    .B_PE_dummy_in_0__ap_start(B_PE_dummy_in_0__ap_start),
    .B_PE_dummy_in_0__ap_ready(B_PE_dummy_in_0__ap_ready),
    .B_PE_dummy_in_0__ap_done(B_PE_dummy_in_0__ap_done),
    .B_PE_dummy_in_0__ap_idle(B_PE_dummy_in_0__ap_idle),
    .B_PE_dummy_in_1__ap_start(B_PE_dummy_in_1__ap_start),
    .B_PE_dummy_in_1__ap_ready(B_PE_dummy_in_1__ap_ready),
    .B_PE_dummy_in_1__ap_done(B_PE_dummy_in_1__ap_done),
    .B_PE_dummy_in_1__ap_idle(B_PE_dummy_in_1__ap_idle),
    .B_PE_dummy_in_2__ap_start(B_PE_dummy_in_2__ap_start),
    .B_PE_dummy_in_2__ap_ready(B_PE_dummy_in_2__ap_ready),
    .B_PE_dummy_in_2__ap_done(B_PE_dummy_in_2__ap_done),
    .B_PE_dummy_in_2__ap_idle(B_PE_dummy_in_2__ap_idle),
    .B_PE_dummy_in_3__ap_start(B_PE_dummy_in_3__ap_start),
    .B_PE_dummy_in_3__ap_ready(B_PE_dummy_in_3__ap_ready),
    .B_PE_dummy_in_3__ap_done(B_PE_dummy_in_3__ap_done),
    .B_PE_dummy_in_3__ap_idle(B_PE_dummy_in_3__ap_idle),
    .B_PE_dummy_in_4__ap_start(B_PE_dummy_in_4__ap_start),
    .B_PE_dummy_in_4__ap_ready(B_PE_dummy_in_4__ap_ready),
    .B_PE_dummy_in_4__ap_done(B_PE_dummy_in_4__ap_done),
    .B_PE_dummy_in_4__ap_idle(B_PE_dummy_in_4__ap_idle),
    .B_PE_dummy_in_5__ap_start(B_PE_dummy_in_5__ap_start),
    .B_PE_dummy_in_5__ap_ready(B_PE_dummy_in_5__ap_ready),
    .B_PE_dummy_in_5__ap_done(B_PE_dummy_in_5__ap_done),
    .B_PE_dummy_in_5__ap_idle(B_PE_dummy_in_5__ap_idle),
    .B_PE_dummy_in_6__ap_start(B_PE_dummy_in_6__ap_start),
    .B_PE_dummy_in_6__ap_ready(B_PE_dummy_in_6__ap_ready),
    .B_PE_dummy_in_6__ap_done(B_PE_dummy_in_6__ap_done),
    .B_PE_dummy_in_6__ap_idle(B_PE_dummy_in_6__ap_idle),
    .B_PE_dummy_in_7__ap_start(B_PE_dummy_in_7__ap_start),
    .B_PE_dummy_in_7__ap_ready(B_PE_dummy_in_7__ap_ready),
    .B_PE_dummy_in_7__ap_done(B_PE_dummy_in_7__ap_done),
    .B_PE_dummy_in_7__ap_idle(B_PE_dummy_in_7__ap_idle),
    .B_PE_dummy_in_8__ap_start(B_PE_dummy_in_8__ap_start),
    .B_PE_dummy_in_8__ap_ready(B_PE_dummy_in_8__ap_ready),
    .B_PE_dummy_in_8__ap_done(B_PE_dummy_in_8__ap_done),
    .B_PE_dummy_in_8__ap_idle(B_PE_dummy_in_8__ap_idle),
    .B_PE_dummy_in_9__ap_start(B_PE_dummy_in_9__ap_start),
    .B_PE_dummy_in_9__ap_ready(B_PE_dummy_in_9__ap_ready),
    .B_PE_dummy_in_9__ap_done(B_PE_dummy_in_9__ap_done),
    .B_PE_dummy_in_9__ap_idle(B_PE_dummy_in_9__ap_idle),
    .B_PE_dummy_in_10__ap_start(B_PE_dummy_in_10__ap_start),
    .B_PE_dummy_in_10__ap_ready(B_PE_dummy_in_10__ap_ready),
    .B_PE_dummy_in_10__ap_done(B_PE_dummy_in_10__ap_done),
    .B_PE_dummy_in_10__ap_idle(B_PE_dummy_in_10__ap_idle),
    .B_PE_dummy_in_11__ap_start(B_PE_dummy_in_11__ap_start),
    .B_PE_dummy_in_11__ap_ready(B_PE_dummy_in_11__ap_ready),
    .B_PE_dummy_in_11__ap_done(B_PE_dummy_in_11__ap_done),
    .B_PE_dummy_in_11__ap_idle(B_PE_dummy_in_11__ap_idle),
    .B_PE_dummy_in_12__ap_start(B_PE_dummy_in_12__ap_start),
    .B_PE_dummy_in_12__ap_ready(B_PE_dummy_in_12__ap_ready),
    .B_PE_dummy_in_12__ap_done(B_PE_dummy_in_12__ap_done),
    .B_PE_dummy_in_12__ap_idle(B_PE_dummy_in_12__ap_idle),
    .B_PE_dummy_in_13__ap_start(B_PE_dummy_in_13__ap_start),
    .B_PE_dummy_in_13__ap_ready(B_PE_dummy_in_13__ap_ready),
    .B_PE_dummy_in_13__ap_done(B_PE_dummy_in_13__ap_done),
    .B_PE_dummy_in_13__ap_idle(B_PE_dummy_in_13__ap_idle),
    .B_PE_dummy_in_14__ap_start(B_PE_dummy_in_14__ap_start),
    .B_PE_dummy_in_14__ap_ready(B_PE_dummy_in_14__ap_ready),
    .B_PE_dummy_in_14__ap_done(B_PE_dummy_in_14__ap_done),
    .B_PE_dummy_in_14__ap_idle(B_PE_dummy_in_14__ap_idle),
    .B_PE_dummy_in_15__ap_start(B_PE_dummy_in_15__ap_start),
    .B_PE_dummy_in_15__ap_ready(B_PE_dummy_in_15__ap_ready),
    .B_PE_dummy_in_15__ap_done(B_PE_dummy_in_15__ap_done),
    .B_PE_dummy_in_15__ap_idle(B_PE_dummy_in_15__ap_idle),
    .B_PE_dummy_in_16__ap_start(B_PE_dummy_in_16__ap_start),
    .B_PE_dummy_in_16__ap_ready(B_PE_dummy_in_16__ap_ready),
    .B_PE_dummy_in_16__ap_done(B_PE_dummy_in_16__ap_done),
    .B_PE_dummy_in_16__ap_idle(B_PE_dummy_in_16__ap_idle),
    .C_drain_IO_L1_out_boundary_wrapper_0__ap_start(C_drain_IO_L1_out_boundary_wrapper_0__ap_start),
    .C_drain_IO_L1_out_boundary_wrapper_0__ap_ready(C_drain_IO_L1_out_boundary_wrapper_0__ap_ready),
    .C_drain_IO_L1_out_boundary_wrapper_0__ap_done(C_drain_IO_L1_out_boundary_wrapper_0__ap_done),
    .C_drain_IO_L1_out_boundary_wrapper_0__ap_idle(C_drain_IO_L1_out_boundary_wrapper_0__ap_idle),
    .C_drain_IO_L1_out_boundary_wrapper_1__ap_start(C_drain_IO_L1_out_boundary_wrapper_1__ap_start),
    .C_drain_IO_L1_out_boundary_wrapper_1__ap_ready(C_drain_IO_L1_out_boundary_wrapper_1__ap_ready),
    .C_drain_IO_L1_out_boundary_wrapper_1__ap_done(C_drain_IO_L1_out_boundary_wrapper_1__ap_done),
    .C_drain_IO_L1_out_boundary_wrapper_1__ap_idle(C_drain_IO_L1_out_boundary_wrapper_1__ap_idle),
    .C_drain_IO_L1_out_boundary_wrapper_2__ap_start(C_drain_IO_L1_out_boundary_wrapper_2__ap_start),
    .C_drain_IO_L1_out_boundary_wrapper_2__ap_ready(C_drain_IO_L1_out_boundary_wrapper_2__ap_ready),
    .C_drain_IO_L1_out_boundary_wrapper_2__ap_done(C_drain_IO_L1_out_boundary_wrapper_2__ap_done),
    .C_drain_IO_L1_out_boundary_wrapper_2__ap_idle(C_drain_IO_L1_out_boundary_wrapper_2__ap_idle),
    .C_drain_IO_L1_out_boundary_wrapper_3__ap_start(C_drain_IO_L1_out_boundary_wrapper_3__ap_start),
    .C_drain_IO_L1_out_boundary_wrapper_3__ap_ready(C_drain_IO_L1_out_boundary_wrapper_3__ap_ready),
    .C_drain_IO_L1_out_boundary_wrapper_3__ap_done(C_drain_IO_L1_out_boundary_wrapper_3__ap_done),
    .C_drain_IO_L1_out_boundary_wrapper_3__ap_idle(C_drain_IO_L1_out_boundary_wrapper_3__ap_idle),
    .C_drain_IO_L1_out_boundary_wrapper_4__ap_start(C_drain_IO_L1_out_boundary_wrapper_4__ap_start),
    .C_drain_IO_L1_out_boundary_wrapper_4__ap_ready(C_drain_IO_L1_out_boundary_wrapper_4__ap_ready),
    .C_drain_IO_L1_out_boundary_wrapper_4__ap_done(C_drain_IO_L1_out_boundary_wrapper_4__ap_done),
    .C_drain_IO_L1_out_boundary_wrapper_4__ap_idle(C_drain_IO_L1_out_boundary_wrapper_4__ap_idle),
    .C_drain_IO_L1_out_boundary_wrapper_5__ap_start(C_drain_IO_L1_out_boundary_wrapper_5__ap_start),
    .C_drain_IO_L1_out_boundary_wrapper_5__ap_ready(C_drain_IO_L1_out_boundary_wrapper_5__ap_ready),
    .C_drain_IO_L1_out_boundary_wrapper_5__ap_done(C_drain_IO_L1_out_boundary_wrapper_5__ap_done),
    .C_drain_IO_L1_out_boundary_wrapper_5__ap_idle(C_drain_IO_L1_out_boundary_wrapper_5__ap_idle),
    .C_drain_IO_L1_out_boundary_wrapper_6__ap_start(C_drain_IO_L1_out_boundary_wrapper_6__ap_start),
    .C_drain_IO_L1_out_boundary_wrapper_6__ap_ready(C_drain_IO_L1_out_boundary_wrapper_6__ap_ready),
    .C_drain_IO_L1_out_boundary_wrapper_6__ap_done(C_drain_IO_L1_out_boundary_wrapper_6__ap_done),
    .C_drain_IO_L1_out_boundary_wrapper_6__ap_idle(C_drain_IO_L1_out_boundary_wrapper_6__ap_idle),
    .C_drain_IO_L1_out_boundary_wrapper_7__ap_start(C_drain_IO_L1_out_boundary_wrapper_7__ap_start),
    .C_drain_IO_L1_out_boundary_wrapper_7__ap_ready(C_drain_IO_L1_out_boundary_wrapper_7__ap_ready),
    .C_drain_IO_L1_out_boundary_wrapper_7__ap_done(C_drain_IO_L1_out_boundary_wrapper_7__ap_done),
    .C_drain_IO_L1_out_boundary_wrapper_7__ap_idle(C_drain_IO_L1_out_boundary_wrapper_7__ap_idle),
    .C_drain_IO_L1_out_boundary_wrapper_8__ap_start(C_drain_IO_L1_out_boundary_wrapper_8__ap_start),
    .C_drain_IO_L1_out_boundary_wrapper_8__ap_ready(C_drain_IO_L1_out_boundary_wrapper_8__ap_ready),
    .C_drain_IO_L1_out_boundary_wrapper_8__ap_done(C_drain_IO_L1_out_boundary_wrapper_8__ap_done),
    .C_drain_IO_L1_out_boundary_wrapper_8__ap_idle(C_drain_IO_L1_out_boundary_wrapper_8__ap_idle),
    .C_drain_IO_L1_out_boundary_wrapper_9__ap_start(C_drain_IO_L1_out_boundary_wrapper_9__ap_start),
    .C_drain_IO_L1_out_boundary_wrapper_9__ap_ready(C_drain_IO_L1_out_boundary_wrapper_9__ap_ready),
    .C_drain_IO_L1_out_boundary_wrapper_9__ap_done(C_drain_IO_L1_out_boundary_wrapper_9__ap_done),
    .C_drain_IO_L1_out_boundary_wrapper_9__ap_idle(C_drain_IO_L1_out_boundary_wrapper_9__ap_idle),
    .C_drain_IO_L1_out_boundary_wrapper_10__ap_start(C_drain_IO_L1_out_boundary_wrapper_10__ap_start),
    .C_drain_IO_L1_out_boundary_wrapper_10__ap_ready(C_drain_IO_L1_out_boundary_wrapper_10__ap_ready),
    .C_drain_IO_L1_out_boundary_wrapper_10__ap_done(C_drain_IO_L1_out_boundary_wrapper_10__ap_done),
    .C_drain_IO_L1_out_boundary_wrapper_10__ap_idle(C_drain_IO_L1_out_boundary_wrapper_10__ap_idle),
    .C_drain_IO_L1_out_boundary_wrapper_11__ap_start(C_drain_IO_L1_out_boundary_wrapper_11__ap_start),
    .C_drain_IO_L1_out_boundary_wrapper_11__ap_ready(C_drain_IO_L1_out_boundary_wrapper_11__ap_ready),
    .C_drain_IO_L1_out_boundary_wrapper_11__ap_done(C_drain_IO_L1_out_boundary_wrapper_11__ap_done),
    .C_drain_IO_L1_out_boundary_wrapper_11__ap_idle(C_drain_IO_L1_out_boundary_wrapper_11__ap_idle),
    .C_drain_IO_L1_out_boundary_wrapper_12__ap_start(C_drain_IO_L1_out_boundary_wrapper_12__ap_start),
    .C_drain_IO_L1_out_boundary_wrapper_12__ap_ready(C_drain_IO_L1_out_boundary_wrapper_12__ap_ready),
    .C_drain_IO_L1_out_boundary_wrapper_12__ap_done(C_drain_IO_L1_out_boundary_wrapper_12__ap_done),
    .C_drain_IO_L1_out_boundary_wrapper_12__ap_idle(C_drain_IO_L1_out_boundary_wrapper_12__ap_idle),
    .C_drain_IO_L1_out_boundary_wrapper_13__ap_start(C_drain_IO_L1_out_boundary_wrapper_13__ap_start),
    .C_drain_IO_L1_out_boundary_wrapper_13__ap_ready(C_drain_IO_L1_out_boundary_wrapper_13__ap_ready),
    .C_drain_IO_L1_out_boundary_wrapper_13__ap_done(C_drain_IO_L1_out_boundary_wrapper_13__ap_done),
    .C_drain_IO_L1_out_boundary_wrapper_13__ap_idle(C_drain_IO_L1_out_boundary_wrapper_13__ap_idle),
    .C_drain_IO_L1_out_boundary_wrapper_14__ap_start(C_drain_IO_L1_out_boundary_wrapper_14__ap_start),
    .C_drain_IO_L1_out_boundary_wrapper_14__ap_ready(C_drain_IO_L1_out_boundary_wrapper_14__ap_ready),
    .C_drain_IO_L1_out_boundary_wrapper_14__ap_done(C_drain_IO_L1_out_boundary_wrapper_14__ap_done),
    .C_drain_IO_L1_out_boundary_wrapper_14__ap_idle(C_drain_IO_L1_out_boundary_wrapper_14__ap_idle),
    .C_drain_IO_L1_out_boundary_wrapper_15__ap_start(C_drain_IO_L1_out_boundary_wrapper_15__ap_start),
    .C_drain_IO_L1_out_boundary_wrapper_15__ap_ready(C_drain_IO_L1_out_boundary_wrapper_15__ap_ready),
    .C_drain_IO_L1_out_boundary_wrapper_15__ap_done(C_drain_IO_L1_out_boundary_wrapper_15__ap_done),
    .C_drain_IO_L1_out_boundary_wrapper_15__ap_idle(C_drain_IO_L1_out_boundary_wrapper_15__ap_idle),
    .C_drain_IO_L1_out_boundary_wrapper_16__ap_start(C_drain_IO_L1_out_boundary_wrapper_16__ap_start),
    .C_drain_IO_L1_out_boundary_wrapper_16__ap_ready(C_drain_IO_L1_out_boundary_wrapper_16__ap_ready),
    .C_drain_IO_L1_out_boundary_wrapper_16__ap_done(C_drain_IO_L1_out_boundary_wrapper_16__ap_done),
    .C_drain_IO_L1_out_boundary_wrapper_16__ap_idle(C_drain_IO_L1_out_boundary_wrapper_16__ap_idle),
    .C_drain_IO_L1_out_wrapper_0__ap_start(C_drain_IO_L1_out_wrapper_0__ap_start),
    .C_drain_IO_L1_out_wrapper_0__ap_ready(C_drain_IO_L1_out_wrapper_0__ap_ready),
    .C_drain_IO_L1_out_wrapper_0__ap_done(C_drain_IO_L1_out_wrapper_0__ap_done),
    .C_drain_IO_L1_out_wrapper_0__ap_idle(C_drain_IO_L1_out_wrapper_0__ap_idle),
    .C_drain_IO_L1_out_wrapper_1__ap_start(C_drain_IO_L1_out_wrapper_1__ap_start),
    .C_drain_IO_L1_out_wrapper_1__ap_ready(C_drain_IO_L1_out_wrapper_1__ap_ready),
    .C_drain_IO_L1_out_wrapper_1__ap_done(C_drain_IO_L1_out_wrapper_1__ap_done),
    .C_drain_IO_L1_out_wrapper_1__ap_idle(C_drain_IO_L1_out_wrapper_1__ap_idle),
    .C_drain_IO_L1_out_wrapper_2__ap_start(C_drain_IO_L1_out_wrapper_2__ap_start),
    .C_drain_IO_L1_out_wrapper_2__ap_ready(C_drain_IO_L1_out_wrapper_2__ap_ready),
    .C_drain_IO_L1_out_wrapper_2__ap_done(C_drain_IO_L1_out_wrapper_2__ap_done),
    .C_drain_IO_L1_out_wrapper_2__ap_idle(C_drain_IO_L1_out_wrapper_2__ap_idle),
    .C_drain_IO_L1_out_wrapper_3__ap_start(C_drain_IO_L1_out_wrapper_3__ap_start),
    .C_drain_IO_L1_out_wrapper_3__ap_ready(C_drain_IO_L1_out_wrapper_3__ap_ready),
    .C_drain_IO_L1_out_wrapper_3__ap_done(C_drain_IO_L1_out_wrapper_3__ap_done),
    .C_drain_IO_L1_out_wrapper_3__ap_idle(C_drain_IO_L1_out_wrapper_3__ap_idle),
    .C_drain_IO_L1_out_wrapper_4__ap_start(C_drain_IO_L1_out_wrapper_4__ap_start),
    .C_drain_IO_L1_out_wrapper_4__ap_ready(C_drain_IO_L1_out_wrapper_4__ap_ready),
    .C_drain_IO_L1_out_wrapper_4__ap_done(C_drain_IO_L1_out_wrapper_4__ap_done),
    .C_drain_IO_L1_out_wrapper_4__ap_idle(C_drain_IO_L1_out_wrapper_4__ap_idle),
    .C_drain_IO_L1_out_wrapper_5__ap_start(C_drain_IO_L1_out_wrapper_5__ap_start),
    .C_drain_IO_L1_out_wrapper_5__ap_ready(C_drain_IO_L1_out_wrapper_5__ap_ready),
    .C_drain_IO_L1_out_wrapper_5__ap_done(C_drain_IO_L1_out_wrapper_5__ap_done),
    .C_drain_IO_L1_out_wrapper_5__ap_idle(C_drain_IO_L1_out_wrapper_5__ap_idle),
    .C_drain_IO_L1_out_wrapper_6__ap_start(C_drain_IO_L1_out_wrapper_6__ap_start),
    .C_drain_IO_L1_out_wrapper_6__ap_ready(C_drain_IO_L1_out_wrapper_6__ap_ready),
    .C_drain_IO_L1_out_wrapper_6__ap_done(C_drain_IO_L1_out_wrapper_6__ap_done),
    .C_drain_IO_L1_out_wrapper_6__ap_idle(C_drain_IO_L1_out_wrapper_6__ap_idle),
    .C_drain_IO_L1_out_wrapper_7__ap_start(C_drain_IO_L1_out_wrapper_7__ap_start),
    .C_drain_IO_L1_out_wrapper_7__ap_ready(C_drain_IO_L1_out_wrapper_7__ap_ready),
    .C_drain_IO_L1_out_wrapper_7__ap_done(C_drain_IO_L1_out_wrapper_7__ap_done),
    .C_drain_IO_L1_out_wrapper_7__ap_idle(C_drain_IO_L1_out_wrapper_7__ap_idle),
    .C_drain_IO_L1_out_wrapper_8__ap_start(C_drain_IO_L1_out_wrapper_8__ap_start),
    .C_drain_IO_L1_out_wrapper_8__ap_ready(C_drain_IO_L1_out_wrapper_8__ap_ready),
    .C_drain_IO_L1_out_wrapper_8__ap_done(C_drain_IO_L1_out_wrapper_8__ap_done),
    .C_drain_IO_L1_out_wrapper_8__ap_idle(C_drain_IO_L1_out_wrapper_8__ap_idle),
    .C_drain_IO_L1_out_wrapper_9__ap_start(C_drain_IO_L1_out_wrapper_9__ap_start),
    .C_drain_IO_L1_out_wrapper_9__ap_ready(C_drain_IO_L1_out_wrapper_9__ap_ready),
    .C_drain_IO_L1_out_wrapper_9__ap_done(C_drain_IO_L1_out_wrapper_9__ap_done),
    .C_drain_IO_L1_out_wrapper_9__ap_idle(C_drain_IO_L1_out_wrapper_9__ap_idle),
    .C_drain_IO_L1_out_wrapper_10__ap_start(C_drain_IO_L1_out_wrapper_10__ap_start),
    .C_drain_IO_L1_out_wrapper_10__ap_ready(C_drain_IO_L1_out_wrapper_10__ap_ready),
    .C_drain_IO_L1_out_wrapper_10__ap_done(C_drain_IO_L1_out_wrapper_10__ap_done),
    .C_drain_IO_L1_out_wrapper_10__ap_idle(C_drain_IO_L1_out_wrapper_10__ap_idle),
    .C_drain_IO_L1_out_wrapper_11__ap_start(C_drain_IO_L1_out_wrapper_11__ap_start),
    .C_drain_IO_L1_out_wrapper_11__ap_ready(C_drain_IO_L1_out_wrapper_11__ap_ready),
    .C_drain_IO_L1_out_wrapper_11__ap_done(C_drain_IO_L1_out_wrapper_11__ap_done),
    .C_drain_IO_L1_out_wrapper_11__ap_idle(C_drain_IO_L1_out_wrapper_11__ap_idle),
    .C_drain_IO_L1_out_wrapper_12__ap_start(C_drain_IO_L1_out_wrapper_12__ap_start),
    .C_drain_IO_L1_out_wrapper_12__ap_ready(C_drain_IO_L1_out_wrapper_12__ap_ready),
    .C_drain_IO_L1_out_wrapper_12__ap_done(C_drain_IO_L1_out_wrapper_12__ap_done),
    .C_drain_IO_L1_out_wrapper_12__ap_idle(C_drain_IO_L1_out_wrapper_12__ap_idle),
    .C_drain_IO_L1_out_wrapper_13__ap_start(C_drain_IO_L1_out_wrapper_13__ap_start),
    .C_drain_IO_L1_out_wrapper_13__ap_ready(C_drain_IO_L1_out_wrapper_13__ap_ready),
    .C_drain_IO_L1_out_wrapper_13__ap_done(C_drain_IO_L1_out_wrapper_13__ap_done),
    .C_drain_IO_L1_out_wrapper_13__ap_idle(C_drain_IO_L1_out_wrapper_13__ap_idle),
    .C_drain_IO_L1_out_wrapper_14__ap_start(C_drain_IO_L1_out_wrapper_14__ap_start),
    .C_drain_IO_L1_out_wrapper_14__ap_ready(C_drain_IO_L1_out_wrapper_14__ap_ready),
    .C_drain_IO_L1_out_wrapper_14__ap_done(C_drain_IO_L1_out_wrapper_14__ap_done),
    .C_drain_IO_L1_out_wrapper_14__ap_idle(C_drain_IO_L1_out_wrapper_14__ap_idle),
    .C_drain_IO_L1_out_wrapper_15__ap_start(C_drain_IO_L1_out_wrapper_15__ap_start),
    .C_drain_IO_L1_out_wrapper_15__ap_ready(C_drain_IO_L1_out_wrapper_15__ap_ready),
    .C_drain_IO_L1_out_wrapper_15__ap_done(C_drain_IO_L1_out_wrapper_15__ap_done),
    .C_drain_IO_L1_out_wrapper_15__ap_idle(C_drain_IO_L1_out_wrapper_15__ap_idle),
    .C_drain_IO_L1_out_wrapper_16__ap_start(C_drain_IO_L1_out_wrapper_16__ap_start),
    .C_drain_IO_L1_out_wrapper_16__ap_ready(C_drain_IO_L1_out_wrapper_16__ap_ready),
    .C_drain_IO_L1_out_wrapper_16__ap_done(C_drain_IO_L1_out_wrapper_16__ap_done),
    .C_drain_IO_L1_out_wrapper_16__ap_idle(C_drain_IO_L1_out_wrapper_16__ap_idle),
    .C_drain_IO_L1_out_wrapper_17__ap_start(C_drain_IO_L1_out_wrapper_17__ap_start),
    .C_drain_IO_L1_out_wrapper_17__ap_ready(C_drain_IO_L1_out_wrapper_17__ap_ready),
    .C_drain_IO_L1_out_wrapper_17__ap_done(C_drain_IO_L1_out_wrapper_17__ap_done),
    .C_drain_IO_L1_out_wrapper_17__ap_idle(C_drain_IO_L1_out_wrapper_17__ap_idle),
    .C_drain_IO_L1_out_wrapper_18__ap_start(C_drain_IO_L1_out_wrapper_18__ap_start),
    .C_drain_IO_L1_out_wrapper_18__ap_ready(C_drain_IO_L1_out_wrapper_18__ap_ready),
    .C_drain_IO_L1_out_wrapper_18__ap_done(C_drain_IO_L1_out_wrapper_18__ap_done),
    .C_drain_IO_L1_out_wrapper_18__ap_idle(C_drain_IO_L1_out_wrapper_18__ap_idle),
    .C_drain_IO_L1_out_wrapper_19__ap_start(C_drain_IO_L1_out_wrapper_19__ap_start),
    .C_drain_IO_L1_out_wrapper_19__ap_ready(C_drain_IO_L1_out_wrapper_19__ap_ready),
    .C_drain_IO_L1_out_wrapper_19__ap_done(C_drain_IO_L1_out_wrapper_19__ap_done),
    .C_drain_IO_L1_out_wrapper_19__ap_idle(C_drain_IO_L1_out_wrapper_19__ap_idle),
    .C_drain_IO_L1_out_wrapper_20__ap_start(C_drain_IO_L1_out_wrapper_20__ap_start),
    .C_drain_IO_L1_out_wrapper_20__ap_ready(C_drain_IO_L1_out_wrapper_20__ap_ready),
    .C_drain_IO_L1_out_wrapper_20__ap_done(C_drain_IO_L1_out_wrapper_20__ap_done),
    .C_drain_IO_L1_out_wrapper_20__ap_idle(C_drain_IO_L1_out_wrapper_20__ap_idle),
    .C_drain_IO_L1_out_wrapper_21__ap_start(C_drain_IO_L1_out_wrapper_21__ap_start),
    .C_drain_IO_L1_out_wrapper_21__ap_ready(C_drain_IO_L1_out_wrapper_21__ap_ready),
    .C_drain_IO_L1_out_wrapper_21__ap_done(C_drain_IO_L1_out_wrapper_21__ap_done),
    .C_drain_IO_L1_out_wrapper_21__ap_idle(C_drain_IO_L1_out_wrapper_21__ap_idle),
    .C_drain_IO_L1_out_wrapper_22__ap_start(C_drain_IO_L1_out_wrapper_22__ap_start),
    .C_drain_IO_L1_out_wrapper_22__ap_ready(C_drain_IO_L1_out_wrapper_22__ap_ready),
    .C_drain_IO_L1_out_wrapper_22__ap_done(C_drain_IO_L1_out_wrapper_22__ap_done),
    .C_drain_IO_L1_out_wrapper_22__ap_idle(C_drain_IO_L1_out_wrapper_22__ap_idle),
    .C_drain_IO_L1_out_wrapper_23__ap_start(C_drain_IO_L1_out_wrapper_23__ap_start),
    .C_drain_IO_L1_out_wrapper_23__ap_ready(C_drain_IO_L1_out_wrapper_23__ap_ready),
    .C_drain_IO_L1_out_wrapper_23__ap_done(C_drain_IO_L1_out_wrapper_23__ap_done),
    .C_drain_IO_L1_out_wrapper_23__ap_idle(C_drain_IO_L1_out_wrapper_23__ap_idle),
    .C_drain_IO_L1_out_wrapper_24__ap_start(C_drain_IO_L1_out_wrapper_24__ap_start),
    .C_drain_IO_L1_out_wrapper_24__ap_ready(C_drain_IO_L1_out_wrapper_24__ap_ready),
    .C_drain_IO_L1_out_wrapper_24__ap_done(C_drain_IO_L1_out_wrapper_24__ap_done),
    .C_drain_IO_L1_out_wrapper_24__ap_idle(C_drain_IO_L1_out_wrapper_24__ap_idle),
    .C_drain_IO_L1_out_wrapper_25__ap_start(C_drain_IO_L1_out_wrapper_25__ap_start),
    .C_drain_IO_L1_out_wrapper_25__ap_ready(C_drain_IO_L1_out_wrapper_25__ap_ready),
    .C_drain_IO_L1_out_wrapper_25__ap_done(C_drain_IO_L1_out_wrapper_25__ap_done),
    .C_drain_IO_L1_out_wrapper_25__ap_idle(C_drain_IO_L1_out_wrapper_25__ap_idle),
    .C_drain_IO_L1_out_wrapper_26__ap_start(C_drain_IO_L1_out_wrapper_26__ap_start),
    .C_drain_IO_L1_out_wrapper_26__ap_ready(C_drain_IO_L1_out_wrapper_26__ap_ready),
    .C_drain_IO_L1_out_wrapper_26__ap_done(C_drain_IO_L1_out_wrapper_26__ap_done),
    .C_drain_IO_L1_out_wrapper_26__ap_idle(C_drain_IO_L1_out_wrapper_26__ap_idle),
    .C_drain_IO_L1_out_wrapper_27__ap_start(C_drain_IO_L1_out_wrapper_27__ap_start),
    .C_drain_IO_L1_out_wrapper_27__ap_ready(C_drain_IO_L1_out_wrapper_27__ap_ready),
    .C_drain_IO_L1_out_wrapper_27__ap_done(C_drain_IO_L1_out_wrapper_27__ap_done),
    .C_drain_IO_L1_out_wrapper_27__ap_idle(C_drain_IO_L1_out_wrapper_27__ap_idle),
    .C_drain_IO_L1_out_wrapper_28__ap_start(C_drain_IO_L1_out_wrapper_28__ap_start),
    .C_drain_IO_L1_out_wrapper_28__ap_ready(C_drain_IO_L1_out_wrapper_28__ap_ready),
    .C_drain_IO_L1_out_wrapper_28__ap_done(C_drain_IO_L1_out_wrapper_28__ap_done),
    .C_drain_IO_L1_out_wrapper_28__ap_idle(C_drain_IO_L1_out_wrapper_28__ap_idle),
    .C_drain_IO_L1_out_wrapper_29__ap_start(C_drain_IO_L1_out_wrapper_29__ap_start),
    .C_drain_IO_L1_out_wrapper_29__ap_ready(C_drain_IO_L1_out_wrapper_29__ap_ready),
    .C_drain_IO_L1_out_wrapper_29__ap_done(C_drain_IO_L1_out_wrapper_29__ap_done),
    .C_drain_IO_L1_out_wrapper_29__ap_idle(C_drain_IO_L1_out_wrapper_29__ap_idle),
    .C_drain_IO_L1_out_wrapper_30__ap_start(C_drain_IO_L1_out_wrapper_30__ap_start),
    .C_drain_IO_L1_out_wrapper_30__ap_ready(C_drain_IO_L1_out_wrapper_30__ap_ready),
    .C_drain_IO_L1_out_wrapper_30__ap_done(C_drain_IO_L1_out_wrapper_30__ap_done),
    .C_drain_IO_L1_out_wrapper_30__ap_idle(C_drain_IO_L1_out_wrapper_30__ap_idle),
    .C_drain_IO_L1_out_wrapper_31__ap_start(C_drain_IO_L1_out_wrapper_31__ap_start),
    .C_drain_IO_L1_out_wrapper_31__ap_ready(C_drain_IO_L1_out_wrapper_31__ap_ready),
    .C_drain_IO_L1_out_wrapper_31__ap_done(C_drain_IO_L1_out_wrapper_31__ap_done),
    .C_drain_IO_L1_out_wrapper_31__ap_idle(C_drain_IO_L1_out_wrapper_31__ap_idle),
    .C_drain_IO_L1_out_wrapper_32__ap_start(C_drain_IO_L1_out_wrapper_32__ap_start),
    .C_drain_IO_L1_out_wrapper_32__ap_ready(C_drain_IO_L1_out_wrapper_32__ap_ready),
    .C_drain_IO_L1_out_wrapper_32__ap_done(C_drain_IO_L1_out_wrapper_32__ap_done),
    .C_drain_IO_L1_out_wrapper_32__ap_idle(C_drain_IO_L1_out_wrapper_32__ap_idle),
    .C_drain_IO_L1_out_wrapper_33__ap_start(C_drain_IO_L1_out_wrapper_33__ap_start),
    .C_drain_IO_L1_out_wrapper_33__ap_ready(C_drain_IO_L1_out_wrapper_33__ap_ready),
    .C_drain_IO_L1_out_wrapper_33__ap_done(C_drain_IO_L1_out_wrapper_33__ap_done),
    .C_drain_IO_L1_out_wrapper_33__ap_idle(C_drain_IO_L1_out_wrapper_33__ap_idle),
    .C_drain_IO_L1_out_wrapper_34__ap_start(C_drain_IO_L1_out_wrapper_34__ap_start),
    .C_drain_IO_L1_out_wrapper_34__ap_ready(C_drain_IO_L1_out_wrapper_34__ap_ready),
    .C_drain_IO_L1_out_wrapper_34__ap_done(C_drain_IO_L1_out_wrapper_34__ap_done),
    .C_drain_IO_L1_out_wrapper_34__ap_idle(C_drain_IO_L1_out_wrapper_34__ap_idle),
    .C_drain_IO_L1_out_wrapper_35__ap_start(C_drain_IO_L1_out_wrapper_35__ap_start),
    .C_drain_IO_L1_out_wrapper_35__ap_ready(C_drain_IO_L1_out_wrapper_35__ap_ready),
    .C_drain_IO_L1_out_wrapper_35__ap_done(C_drain_IO_L1_out_wrapper_35__ap_done),
    .C_drain_IO_L1_out_wrapper_35__ap_idle(C_drain_IO_L1_out_wrapper_35__ap_idle),
    .C_drain_IO_L1_out_wrapper_36__ap_start(C_drain_IO_L1_out_wrapper_36__ap_start),
    .C_drain_IO_L1_out_wrapper_36__ap_ready(C_drain_IO_L1_out_wrapper_36__ap_ready),
    .C_drain_IO_L1_out_wrapper_36__ap_done(C_drain_IO_L1_out_wrapper_36__ap_done),
    .C_drain_IO_L1_out_wrapper_36__ap_idle(C_drain_IO_L1_out_wrapper_36__ap_idle),
    .C_drain_IO_L1_out_wrapper_37__ap_start(C_drain_IO_L1_out_wrapper_37__ap_start),
    .C_drain_IO_L1_out_wrapper_37__ap_ready(C_drain_IO_L1_out_wrapper_37__ap_ready),
    .C_drain_IO_L1_out_wrapper_37__ap_done(C_drain_IO_L1_out_wrapper_37__ap_done),
    .C_drain_IO_L1_out_wrapper_37__ap_idle(C_drain_IO_L1_out_wrapper_37__ap_idle),
    .C_drain_IO_L1_out_wrapper_38__ap_start(C_drain_IO_L1_out_wrapper_38__ap_start),
    .C_drain_IO_L1_out_wrapper_38__ap_ready(C_drain_IO_L1_out_wrapper_38__ap_ready),
    .C_drain_IO_L1_out_wrapper_38__ap_done(C_drain_IO_L1_out_wrapper_38__ap_done),
    .C_drain_IO_L1_out_wrapper_38__ap_idle(C_drain_IO_L1_out_wrapper_38__ap_idle),
    .C_drain_IO_L1_out_wrapper_39__ap_start(C_drain_IO_L1_out_wrapper_39__ap_start),
    .C_drain_IO_L1_out_wrapper_39__ap_ready(C_drain_IO_L1_out_wrapper_39__ap_ready),
    .C_drain_IO_L1_out_wrapper_39__ap_done(C_drain_IO_L1_out_wrapper_39__ap_done),
    .C_drain_IO_L1_out_wrapper_39__ap_idle(C_drain_IO_L1_out_wrapper_39__ap_idle),
    .C_drain_IO_L1_out_wrapper_40__ap_start(C_drain_IO_L1_out_wrapper_40__ap_start),
    .C_drain_IO_L1_out_wrapper_40__ap_ready(C_drain_IO_L1_out_wrapper_40__ap_ready),
    .C_drain_IO_L1_out_wrapper_40__ap_done(C_drain_IO_L1_out_wrapper_40__ap_done),
    .C_drain_IO_L1_out_wrapper_40__ap_idle(C_drain_IO_L1_out_wrapper_40__ap_idle),
    .C_drain_IO_L1_out_wrapper_41__ap_start(C_drain_IO_L1_out_wrapper_41__ap_start),
    .C_drain_IO_L1_out_wrapper_41__ap_ready(C_drain_IO_L1_out_wrapper_41__ap_ready),
    .C_drain_IO_L1_out_wrapper_41__ap_done(C_drain_IO_L1_out_wrapper_41__ap_done),
    .C_drain_IO_L1_out_wrapper_41__ap_idle(C_drain_IO_L1_out_wrapper_41__ap_idle),
    .C_drain_IO_L1_out_wrapper_42__ap_start(C_drain_IO_L1_out_wrapper_42__ap_start),
    .C_drain_IO_L1_out_wrapper_42__ap_ready(C_drain_IO_L1_out_wrapper_42__ap_ready),
    .C_drain_IO_L1_out_wrapper_42__ap_done(C_drain_IO_L1_out_wrapper_42__ap_done),
    .C_drain_IO_L1_out_wrapper_42__ap_idle(C_drain_IO_L1_out_wrapper_42__ap_idle),
    .C_drain_IO_L1_out_wrapper_43__ap_start(C_drain_IO_L1_out_wrapper_43__ap_start),
    .C_drain_IO_L1_out_wrapper_43__ap_ready(C_drain_IO_L1_out_wrapper_43__ap_ready),
    .C_drain_IO_L1_out_wrapper_43__ap_done(C_drain_IO_L1_out_wrapper_43__ap_done),
    .C_drain_IO_L1_out_wrapper_43__ap_idle(C_drain_IO_L1_out_wrapper_43__ap_idle),
    .C_drain_IO_L1_out_wrapper_44__ap_start(C_drain_IO_L1_out_wrapper_44__ap_start),
    .C_drain_IO_L1_out_wrapper_44__ap_ready(C_drain_IO_L1_out_wrapper_44__ap_ready),
    .C_drain_IO_L1_out_wrapper_44__ap_done(C_drain_IO_L1_out_wrapper_44__ap_done),
    .C_drain_IO_L1_out_wrapper_44__ap_idle(C_drain_IO_L1_out_wrapper_44__ap_idle),
    .C_drain_IO_L1_out_wrapper_45__ap_start(C_drain_IO_L1_out_wrapper_45__ap_start),
    .C_drain_IO_L1_out_wrapper_45__ap_ready(C_drain_IO_L1_out_wrapper_45__ap_ready),
    .C_drain_IO_L1_out_wrapper_45__ap_done(C_drain_IO_L1_out_wrapper_45__ap_done),
    .C_drain_IO_L1_out_wrapper_45__ap_idle(C_drain_IO_L1_out_wrapper_45__ap_idle),
    .C_drain_IO_L1_out_wrapper_46__ap_start(C_drain_IO_L1_out_wrapper_46__ap_start),
    .C_drain_IO_L1_out_wrapper_46__ap_ready(C_drain_IO_L1_out_wrapper_46__ap_ready),
    .C_drain_IO_L1_out_wrapper_46__ap_done(C_drain_IO_L1_out_wrapper_46__ap_done),
    .C_drain_IO_L1_out_wrapper_46__ap_idle(C_drain_IO_L1_out_wrapper_46__ap_idle),
    .C_drain_IO_L1_out_wrapper_47__ap_start(C_drain_IO_L1_out_wrapper_47__ap_start),
    .C_drain_IO_L1_out_wrapper_47__ap_ready(C_drain_IO_L1_out_wrapper_47__ap_ready),
    .C_drain_IO_L1_out_wrapper_47__ap_done(C_drain_IO_L1_out_wrapper_47__ap_done),
    .C_drain_IO_L1_out_wrapper_47__ap_idle(C_drain_IO_L1_out_wrapper_47__ap_idle),
    .C_drain_IO_L1_out_wrapper_48__ap_start(C_drain_IO_L1_out_wrapper_48__ap_start),
    .C_drain_IO_L1_out_wrapper_48__ap_ready(C_drain_IO_L1_out_wrapper_48__ap_ready),
    .C_drain_IO_L1_out_wrapper_48__ap_done(C_drain_IO_L1_out_wrapper_48__ap_done),
    .C_drain_IO_L1_out_wrapper_48__ap_idle(C_drain_IO_L1_out_wrapper_48__ap_idle),
    .C_drain_IO_L1_out_wrapper_49__ap_start(C_drain_IO_L1_out_wrapper_49__ap_start),
    .C_drain_IO_L1_out_wrapper_49__ap_ready(C_drain_IO_L1_out_wrapper_49__ap_ready),
    .C_drain_IO_L1_out_wrapper_49__ap_done(C_drain_IO_L1_out_wrapper_49__ap_done),
    .C_drain_IO_L1_out_wrapper_49__ap_idle(C_drain_IO_L1_out_wrapper_49__ap_idle),
    .C_drain_IO_L1_out_wrapper_50__ap_start(C_drain_IO_L1_out_wrapper_50__ap_start),
    .C_drain_IO_L1_out_wrapper_50__ap_ready(C_drain_IO_L1_out_wrapper_50__ap_ready),
    .C_drain_IO_L1_out_wrapper_50__ap_done(C_drain_IO_L1_out_wrapper_50__ap_done),
    .C_drain_IO_L1_out_wrapper_50__ap_idle(C_drain_IO_L1_out_wrapper_50__ap_idle),
    .C_drain_IO_L1_out_wrapper_51__ap_start(C_drain_IO_L1_out_wrapper_51__ap_start),
    .C_drain_IO_L1_out_wrapper_51__ap_ready(C_drain_IO_L1_out_wrapper_51__ap_ready),
    .C_drain_IO_L1_out_wrapper_51__ap_done(C_drain_IO_L1_out_wrapper_51__ap_done),
    .C_drain_IO_L1_out_wrapper_51__ap_idle(C_drain_IO_L1_out_wrapper_51__ap_idle),
    .C_drain_IO_L1_out_wrapper_52__ap_start(C_drain_IO_L1_out_wrapper_52__ap_start),
    .C_drain_IO_L1_out_wrapper_52__ap_ready(C_drain_IO_L1_out_wrapper_52__ap_ready),
    .C_drain_IO_L1_out_wrapper_52__ap_done(C_drain_IO_L1_out_wrapper_52__ap_done),
    .C_drain_IO_L1_out_wrapper_52__ap_idle(C_drain_IO_L1_out_wrapper_52__ap_idle),
    .C_drain_IO_L1_out_wrapper_53__ap_start(C_drain_IO_L1_out_wrapper_53__ap_start),
    .C_drain_IO_L1_out_wrapper_53__ap_ready(C_drain_IO_L1_out_wrapper_53__ap_ready),
    .C_drain_IO_L1_out_wrapper_53__ap_done(C_drain_IO_L1_out_wrapper_53__ap_done),
    .C_drain_IO_L1_out_wrapper_53__ap_idle(C_drain_IO_L1_out_wrapper_53__ap_idle),
    .C_drain_IO_L1_out_wrapper_54__ap_start(C_drain_IO_L1_out_wrapper_54__ap_start),
    .C_drain_IO_L1_out_wrapper_54__ap_ready(C_drain_IO_L1_out_wrapper_54__ap_ready),
    .C_drain_IO_L1_out_wrapper_54__ap_done(C_drain_IO_L1_out_wrapper_54__ap_done),
    .C_drain_IO_L1_out_wrapper_54__ap_idle(C_drain_IO_L1_out_wrapper_54__ap_idle),
    .C_drain_IO_L1_out_wrapper_55__ap_start(C_drain_IO_L1_out_wrapper_55__ap_start),
    .C_drain_IO_L1_out_wrapper_55__ap_ready(C_drain_IO_L1_out_wrapper_55__ap_ready),
    .C_drain_IO_L1_out_wrapper_55__ap_done(C_drain_IO_L1_out_wrapper_55__ap_done),
    .C_drain_IO_L1_out_wrapper_55__ap_idle(C_drain_IO_L1_out_wrapper_55__ap_idle),
    .C_drain_IO_L1_out_wrapper_56__ap_start(C_drain_IO_L1_out_wrapper_56__ap_start),
    .C_drain_IO_L1_out_wrapper_56__ap_ready(C_drain_IO_L1_out_wrapper_56__ap_ready),
    .C_drain_IO_L1_out_wrapper_56__ap_done(C_drain_IO_L1_out_wrapper_56__ap_done),
    .C_drain_IO_L1_out_wrapper_56__ap_idle(C_drain_IO_L1_out_wrapper_56__ap_idle),
    .C_drain_IO_L1_out_wrapper_57__ap_start(C_drain_IO_L1_out_wrapper_57__ap_start),
    .C_drain_IO_L1_out_wrapper_57__ap_ready(C_drain_IO_L1_out_wrapper_57__ap_ready),
    .C_drain_IO_L1_out_wrapper_57__ap_done(C_drain_IO_L1_out_wrapper_57__ap_done),
    .C_drain_IO_L1_out_wrapper_57__ap_idle(C_drain_IO_L1_out_wrapper_57__ap_idle),
    .C_drain_IO_L1_out_wrapper_58__ap_start(C_drain_IO_L1_out_wrapper_58__ap_start),
    .C_drain_IO_L1_out_wrapper_58__ap_ready(C_drain_IO_L1_out_wrapper_58__ap_ready),
    .C_drain_IO_L1_out_wrapper_58__ap_done(C_drain_IO_L1_out_wrapper_58__ap_done),
    .C_drain_IO_L1_out_wrapper_58__ap_idle(C_drain_IO_L1_out_wrapper_58__ap_idle),
    .C_drain_IO_L1_out_wrapper_59__ap_start(C_drain_IO_L1_out_wrapper_59__ap_start),
    .C_drain_IO_L1_out_wrapper_59__ap_ready(C_drain_IO_L1_out_wrapper_59__ap_ready),
    .C_drain_IO_L1_out_wrapper_59__ap_done(C_drain_IO_L1_out_wrapper_59__ap_done),
    .C_drain_IO_L1_out_wrapper_59__ap_idle(C_drain_IO_L1_out_wrapper_59__ap_idle),
    .C_drain_IO_L1_out_wrapper_60__ap_start(C_drain_IO_L1_out_wrapper_60__ap_start),
    .C_drain_IO_L1_out_wrapper_60__ap_ready(C_drain_IO_L1_out_wrapper_60__ap_ready),
    .C_drain_IO_L1_out_wrapper_60__ap_done(C_drain_IO_L1_out_wrapper_60__ap_done),
    .C_drain_IO_L1_out_wrapper_60__ap_idle(C_drain_IO_L1_out_wrapper_60__ap_idle),
    .C_drain_IO_L1_out_wrapper_61__ap_start(C_drain_IO_L1_out_wrapper_61__ap_start),
    .C_drain_IO_L1_out_wrapper_61__ap_ready(C_drain_IO_L1_out_wrapper_61__ap_ready),
    .C_drain_IO_L1_out_wrapper_61__ap_done(C_drain_IO_L1_out_wrapper_61__ap_done),
    .C_drain_IO_L1_out_wrapper_61__ap_idle(C_drain_IO_L1_out_wrapper_61__ap_idle),
    .C_drain_IO_L1_out_wrapper_62__ap_start(C_drain_IO_L1_out_wrapper_62__ap_start),
    .C_drain_IO_L1_out_wrapper_62__ap_ready(C_drain_IO_L1_out_wrapper_62__ap_ready),
    .C_drain_IO_L1_out_wrapper_62__ap_done(C_drain_IO_L1_out_wrapper_62__ap_done),
    .C_drain_IO_L1_out_wrapper_62__ap_idle(C_drain_IO_L1_out_wrapper_62__ap_idle),
    .C_drain_IO_L1_out_wrapper_63__ap_start(C_drain_IO_L1_out_wrapper_63__ap_start),
    .C_drain_IO_L1_out_wrapper_63__ap_ready(C_drain_IO_L1_out_wrapper_63__ap_ready),
    .C_drain_IO_L1_out_wrapper_63__ap_done(C_drain_IO_L1_out_wrapper_63__ap_done),
    .C_drain_IO_L1_out_wrapper_63__ap_idle(C_drain_IO_L1_out_wrapper_63__ap_idle),
    .C_drain_IO_L1_out_wrapper_64__ap_start(C_drain_IO_L1_out_wrapper_64__ap_start),
    .C_drain_IO_L1_out_wrapper_64__ap_ready(C_drain_IO_L1_out_wrapper_64__ap_ready),
    .C_drain_IO_L1_out_wrapper_64__ap_done(C_drain_IO_L1_out_wrapper_64__ap_done),
    .C_drain_IO_L1_out_wrapper_64__ap_idle(C_drain_IO_L1_out_wrapper_64__ap_idle),
    .C_drain_IO_L1_out_wrapper_65__ap_start(C_drain_IO_L1_out_wrapper_65__ap_start),
    .C_drain_IO_L1_out_wrapper_65__ap_ready(C_drain_IO_L1_out_wrapper_65__ap_ready),
    .C_drain_IO_L1_out_wrapper_65__ap_done(C_drain_IO_L1_out_wrapper_65__ap_done),
    .C_drain_IO_L1_out_wrapper_65__ap_idle(C_drain_IO_L1_out_wrapper_65__ap_idle),
    .C_drain_IO_L1_out_wrapper_66__ap_start(C_drain_IO_L1_out_wrapper_66__ap_start),
    .C_drain_IO_L1_out_wrapper_66__ap_ready(C_drain_IO_L1_out_wrapper_66__ap_ready),
    .C_drain_IO_L1_out_wrapper_66__ap_done(C_drain_IO_L1_out_wrapper_66__ap_done),
    .C_drain_IO_L1_out_wrapper_66__ap_idle(C_drain_IO_L1_out_wrapper_66__ap_idle),
    .C_drain_IO_L1_out_wrapper_67__ap_start(C_drain_IO_L1_out_wrapper_67__ap_start),
    .C_drain_IO_L1_out_wrapper_67__ap_ready(C_drain_IO_L1_out_wrapper_67__ap_ready),
    .C_drain_IO_L1_out_wrapper_67__ap_done(C_drain_IO_L1_out_wrapper_67__ap_done),
    .C_drain_IO_L1_out_wrapper_67__ap_idle(C_drain_IO_L1_out_wrapper_67__ap_idle),
    .C_drain_IO_L1_out_wrapper_68__ap_start(C_drain_IO_L1_out_wrapper_68__ap_start),
    .C_drain_IO_L1_out_wrapper_68__ap_ready(C_drain_IO_L1_out_wrapper_68__ap_ready),
    .C_drain_IO_L1_out_wrapper_68__ap_done(C_drain_IO_L1_out_wrapper_68__ap_done),
    .C_drain_IO_L1_out_wrapper_68__ap_idle(C_drain_IO_L1_out_wrapper_68__ap_idle),
    .C_drain_IO_L1_out_wrapper_69__ap_start(C_drain_IO_L1_out_wrapper_69__ap_start),
    .C_drain_IO_L1_out_wrapper_69__ap_ready(C_drain_IO_L1_out_wrapper_69__ap_ready),
    .C_drain_IO_L1_out_wrapper_69__ap_done(C_drain_IO_L1_out_wrapper_69__ap_done),
    .C_drain_IO_L1_out_wrapper_69__ap_idle(C_drain_IO_L1_out_wrapper_69__ap_idle),
    .C_drain_IO_L1_out_wrapper_70__ap_start(C_drain_IO_L1_out_wrapper_70__ap_start),
    .C_drain_IO_L1_out_wrapper_70__ap_ready(C_drain_IO_L1_out_wrapper_70__ap_ready),
    .C_drain_IO_L1_out_wrapper_70__ap_done(C_drain_IO_L1_out_wrapper_70__ap_done),
    .C_drain_IO_L1_out_wrapper_70__ap_idle(C_drain_IO_L1_out_wrapper_70__ap_idle),
    .C_drain_IO_L1_out_wrapper_71__ap_start(C_drain_IO_L1_out_wrapper_71__ap_start),
    .C_drain_IO_L1_out_wrapper_71__ap_ready(C_drain_IO_L1_out_wrapper_71__ap_ready),
    .C_drain_IO_L1_out_wrapper_71__ap_done(C_drain_IO_L1_out_wrapper_71__ap_done),
    .C_drain_IO_L1_out_wrapper_71__ap_idle(C_drain_IO_L1_out_wrapper_71__ap_idle),
    .C_drain_IO_L1_out_wrapper_72__ap_start(C_drain_IO_L1_out_wrapper_72__ap_start),
    .C_drain_IO_L1_out_wrapper_72__ap_ready(C_drain_IO_L1_out_wrapper_72__ap_ready),
    .C_drain_IO_L1_out_wrapper_72__ap_done(C_drain_IO_L1_out_wrapper_72__ap_done),
    .C_drain_IO_L1_out_wrapper_72__ap_idle(C_drain_IO_L1_out_wrapper_72__ap_idle),
    .C_drain_IO_L1_out_wrapper_73__ap_start(C_drain_IO_L1_out_wrapper_73__ap_start),
    .C_drain_IO_L1_out_wrapper_73__ap_ready(C_drain_IO_L1_out_wrapper_73__ap_ready),
    .C_drain_IO_L1_out_wrapper_73__ap_done(C_drain_IO_L1_out_wrapper_73__ap_done),
    .C_drain_IO_L1_out_wrapper_73__ap_idle(C_drain_IO_L1_out_wrapper_73__ap_idle),
    .C_drain_IO_L1_out_wrapper_74__ap_start(C_drain_IO_L1_out_wrapper_74__ap_start),
    .C_drain_IO_L1_out_wrapper_74__ap_ready(C_drain_IO_L1_out_wrapper_74__ap_ready),
    .C_drain_IO_L1_out_wrapper_74__ap_done(C_drain_IO_L1_out_wrapper_74__ap_done),
    .C_drain_IO_L1_out_wrapper_74__ap_idle(C_drain_IO_L1_out_wrapper_74__ap_idle),
    .C_drain_IO_L1_out_wrapper_75__ap_start(C_drain_IO_L1_out_wrapper_75__ap_start),
    .C_drain_IO_L1_out_wrapper_75__ap_ready(C_drain_IO_L1_out_wrapper_75__ap_ready),
    .C_drain_IO_L1_out_wrapper_75__ap_done(C_drain_IO_L1_out_wrapper_75__ap_done),
    .C_drain_IO_L1_out_wrapper_75__ap_idle(C_drain_IO_L1_out_wrapper_75__ap_idle),
    .C_drain_IO_L1_out_wrapper_76__ap_start(C_drain_IO_L1_out_wrapper_76__ap_start),
    .C_drain_IO_L1_out_wrapper_76__ap_ready(C_drain_IO_L1_out_wrapper_76__ap_ready),
    .C_drain_IO_L1_out_wrapper_76__ap_done(C_drain_IO_L1_out_wrapper_76__ap_done),
    .C_drain_IO_L1_out_wrapper_76__ap_idle(C_drain_IO_L1_out_wrapper_76__ap_idle),
    .C_drain_IO_L1_out_wrapper_77__ap_start(C_drain_IO_L1_out_wrapper_77__ap_start),
    .C_drain_IO_L1_out_wrapper_77__ap_ready(C_drain_IO_L1_out_wrapper_77__ap_ready),
    .C_drain_IO_L1_out_wrapper_77__ap_done(C_drain_IO_L1_out_wrapper_77__ap_done),
    .C_drain_IO_L1_out_wrapper_77__ap_idle(C_drain_IO_L1_out_wrapper_77__ap_idle),
    .C_drain_IO_L1_out_wrapper_78__ap_start(C_drain_IO_L1_out_wrapper_78__ap_start),
    .C_drain_IO_L1_out_wrapper_78__ap_ready(C_drain_IO_L1_out_wrapper_78__ap_ready),
    .C_drain_IO_L1_out_wrapper_78__ap_done(C_drain_IO_L1_out_wrapper_78__ap_done),
    .C_drain_IO_L1_out_wrapper_78__ap_idle(C_drain_IO_L1_out_wrapper_78__ap_idle),
    .C_drain_IO_L1_out_wrapper_79__ap_start(C_drain_IO_L1_out_wrapper_79__ap_start),
    .C_drain_IO_L1_out_wrapper_79__ap_ready(C_drain_IO_L1_out_wrapper_79__ap_ready),
    .C_drain_IO_L1_out_wrapper_79__ap_done(C_drain_IO_L1_out_wrapper_79__ap_done),
    .C_drain_IO_L1_out_wrapper_79__ap_idle(C_drain_IO_L1_out_wrapper_79__ap_idle),
    .C_drain_IO_L1_out_wrapper_80__ap_start(C_drain_IO_L1_out_wrapper_80__ap_start),
    .C_drain_IO_L1_out_wrapper_80__ap_ready(C_drain_IO_L1_out_wrapper_80__ap_ready),
    .C_drain_IO_L1_out_wrapper_80__ap_done(C_drain_IO_L1_out_wrapper_80__ap_done),
    .C_drain_IO_L1_out_wrapper_80__ap_idle(C_drain_IO_L1_out_wrapper_80__ap_idle),
    .C_drain_IO_L1_out_wrapper_81__ap_start(C_drain_IO_L1_out_wrapper_81__ap_start),
    .C_drain_IO_L1_out_wrapper_81__ap_ready(C_drain_IO_L1_out_wrapper_81__ap_ready),
    .C_drain_IO_L1_out_wrapper_81__ap_done(C_drain_IO_L1_out_wrapper_81__ap_done),
    .C_drain_IO_L1_out_wrapper_81__ap_idle(C_drain_IO_L1_out_wrapper_81__ap_idle),
    .C_drain_IO_L1_out_wrapper_82__ap_start(C_drain_IO_L1_out_wrapper_82__ap_start),
    .C_drain_IO_L1_out_wrapper_82__ap_ready(C_drain_IO_L1_out_wrapper_82__ap_ready),
    .C_drain_IO_L1_out_wrapper_82__ap_done(C_drain_IO_L1_out_wrapper_82__ap_done),
    .C_drain_IO_L1_out_wrapper_82__ap_idle(C_drain_IO_L1_out_wrapper_82__ap_idle),
    .C_drain_IO_L1_out_wrapper_83__ap_start(C_drain_IO_L1_out_wrapper_83__ap_start),
    .C_drain_IO_L1_out_wrapper_83__ap_ready(C_drain_IO_L1_out_wrapper_83__ap_ready),
    .C_drain_IO_L1_out_wrapper_83__ap_done(C_drain_IO_L1_out_wrapper_83__ap_done),
    .C_drain_IO_L1_out_wrapper_83__ap_idle(C_drain_IO_L1_out_wrapper_83__ap_idle),
    .C_drain_IO_L1_out_wrapper_84__ap_start(C_drain_IO_L1_out_wrapper_84__ap_start),
    .C_drain_IO_L1_out_wrapper_84__ap_ready(C_drain_IO_L1_out_wrapper_84__ap_ready),
    .C_drain_IO_L1_out_wrapper_84__ap_done(C_drain_IO_L1_out_wrapper_84__ap_done),
    .C_drain_IO_L1_out_wrapper_84__ap_idle(C_drain_IO_L1_out_wrapper_84__ap_idle),
    .C_drain_IO_L1_out_wrapper_85__ap_start(C_drain_IO_L1_out_wrapper_85__ap_start),
    .C_drain_IO_L1_out_wrapper_85__ap_ready(C_drain_IO_L1_out_wrapper_85__ap_ready),
    .C_drain_IO_L1_out_wrapper_85__ap_done(C_drain_IO_L1_out_wrapper_85__ap_done),
    .C_drain_IO_L1_out_wrapper_85__ap_idle(C_drain_IO_L1_out_wrapper_85__ap_idle),
    .C_drain_IO_L1_out_wrapper_86__ap_start(C_drain_IO_L1_out_wrapper_86__ap_start),
    .C_drain_IO_L1_out_wrapper_86__ap_ready(C_drain_IO_L1_out_wrapper_86__ap_ready),
    .C_drain_IO_L1_out_wrapper_86__ap_done(C_drain_IO_L1_out_wrapper_86__ap_done),
    .C_drain_IO_L1_out_wrapper_86__ap_idle(C_drain_IO_L1_out_wrapper_86__ap_idle),
    .C_drain_IO_L1_out_wrapper_87__ap_start(C_drain_IO_L1_out_wrapper_87__ap_start),
    .C_drain_IO_L1_out_wrapper_87__ap_ready(C_drain_IO_L1_out_wrapper_87__ap_ready),
    .C_drain_IO_L1_out_wrapper_87__ap_done(C_drain_IO_L1_out_wrapper_87__ap_done),
    .C_drain_IO_L1_out_wrapper_87__ap_idle(C_drain_IO_L1_out_wrapper_87__ap_idle),
    .C_drain_IO_L1_out_wrapper_88__ap_start(C_drain_IO_L1_out_wrapper_88__ap_start),
    .C_drain_IO_L1_out_wrapper_88__ap_ready(C_drain_IO_L1_out_wrapper_88__ap_ready),
    .C_drain_IO_L1_out_wrapper_88__ap_done(C_drain_IO_L1_out_wrapper_88__ap_done),
    .C_drain_IO_L1_out_wrapper_88__ap_idle(C_drain_IO_L1_out_wrapper_88__ap_idle),
    .C_drain_IO_L1_out_wrapper_89__ap_start(C_drain_IO_L1_out_wrapper_89__ap_start),
    .C_drain_IO_L1_out_wrapper_89__ap_ready(C_drain_IO_L1_out_wrapper_89__ap_ready),
    .C_drain_IO_L1_out_wrapper_89__ap_done(C_drain_IO_L1_out_wrapper_89__ap_done),
    .C_drain_IO_L1_out_wrapper_89__ap_idle(C_drain_IO_L1_out_wrapper_89__ap_idle),
    .C_drain_IO_L1_out_wrapper_90__ap_start(C_drain_IO_L1_out_wrapper_90__ap_start),
    .C_drain_IO_L1_out_wrapper_90__ap_ready(C_drain_IO_L1_out_wrapper_90__ap_ready),
    .C_drain_IO_L1_out_wrapper_90__ap_done(C_drain_IO_L1_out_wrapper_90__ap_done),
    .C_drain_IO_L1_out_wrapper_90__ap_idle(C_drain_IO_L1_out_wrapper_90__ap_idle),
    .C_drain_IO_L1_out_wrapper_91__ap_start(C_drain_IO_L1_out_wrapper_91__ap_start),
    .C_drain_IO_L1_out_wrapper_91__ap_ready(C_drain_IO_L1_out_wrapper_91__ap_ready),
    .C_drain_IO_L1_out_wrapper_91__ap_done(C_drain_IO_L1_out_wrapper_91__ap_done),
    .C_drain_IO_L1_out_wrapper_91__ap_idle(C_drain_IO_L1_out_wrapper_91__ap_idle),
    .C_drain_IO_L1_out_wrapper_92__ap_start(C_drain_IO_L1_out_wrapper_92__ap_start),
    .C_drain_IO_L1_out_wrapper_92__ap_ready(C_drain_IO_L1_out_wrapper_92__ap_ready),
    .C_drain_IO_L1_out_wrapper_92__ap_done(C_drain_IO_L1_out_wrapper_92__ap_done),
    .C_drain_IO_L1_out_wrapper_92__ap_idle(C_drain_IO_L1_out_wrapper_92__ap_idle),
    .C_drain_IO_L1_out_wrapper_93__ap_start(C_drain_IO_L1_out_wrapper_93__ap_start),
    .C_drain_IO_L1_out_wrapper_93__ap_ready(C_drain_IO_L1_out_wrapper_93__ap_ready),
    .C_drain_IO_L1_out_wrapper_93__ap_done(C_drain_IO_L1_out_wrapper_93__ap_done),
    .C_drain_IO_L1_out_wrapper_93__ap_idle(C_drain_IO_L1_out_wrapper_93__ap_idle),
    .C_drain_IO_L1_out_wrapper_94__ap_start(C_drain_IO_L1_out_wrapper_94__ap_start),
    .C_drain_IO_L1_out_wrapper_94__ap_ready(C_drain_IO_L1_out_wrapper_94__ap_ready),
    .C_drain_IO_L1_out_wrapper_94__ap_done(C_drain_IO_L1_out_wrapper_94__ap_done),
    .C_drain_IO_L1_out_wrapper_94__ap_idle(C_drain_IO_L1_out_wrapper_94__ap_idle),
    .C_drain_IO_L1_out_wrapper_95__ap_start(C_drain_IO_L1_out_wrapper_95__ap_start),
    .C_drain_IO_L1_out_wrapper_95__ap_ready(C_drain_IO_L1_out_wrapper_95__ap_ready),
    .C_drain_IO_L1_out_wrapper_95__ap_done(C_drain_IO_L1_out_wrapper_95__ap_done),
    .C_drain_IO_L1_out_wrapper_95__ap_idle(C_drain_IO_L1_out_wrapper_95__ap_idle),
    .C_drain_IO_L1_out_wrapper_96__ap_start(C_drain_IO_L1_out_wrapper_96__ap_start),
    .C_drain_IO_L1_out_wrapper_96__ap_ready(C_drain_IO_L1_out_wrapper_96__ap_ready),
    .C_drain_IO_L1_out_wrapper_96__ap_done(C_drain_IO_L1_out_wrapper_96__ap_done),
    .C_drain_IO_L1_out_wrapper_96__ap_idle(C_drain_IO_L1_out_wrapper_96__ap_idle),
    .C_drain_IO_L1_out_wrapper_97__ap_start(C_drain_IO_L1_out_wrapper_97__ap_start),
    .C_drain_IO_L1_out_wrapper_97__ap_ready(C_drain_IO_L1_out_wrapper_97__ap_ready),
    .C_drain_IO_L1_out_wrapper_97__ap_done(C_drain_IO_L1_out_wrapper_97__ap_done),
    .C_drain_IO_L1_out_wrapper_97__ap_idle(C_drain_IO_L1_out_wrapper_97__ap_idle),
    .C_drain_IO_L1_out_wrapper_98__ap_start(C_drain_IO_L1_out_wrapper_98__ap_start),
    .C_drain_IO_L1_out_wrapper_98__ap_ready(C_drain_IO_L1_out_wrapper_98__ap_ready),
    .C_drain_IO_L1_out_wrapper_98__ap_done(C_drain_IO_L1_out_wrapper_98__ap_done),
    .C_drain_IO_L1_out_wrapper_98__ap_idle(C_drain_IO_L1_out_wrapper_98__ap_idle),
    .C_drain_IO_L1_out_wrapper_99__ap_start(C_drain_IO_L1_out_wrapper_99__ap_start),
    .C_drain_IO_L1_out_wrapper_99__ap_ready(C_drain_IO_L1_out_wrapper_99__ap_ready),
    .C_drain_IO_L1_out_wrapper_99__ap_done(C_drain_IO_L1_out_wrapper_99__ap_done),
    .C_drain_IO_L1_out_wrapper_99__ap_idle(C_drain_IO_L1_out_wrapper_99__ap_idle),
    .C_drain_IO_L1_out_wrapper_100__ap_start(C_drain_IO_L1_out_wrapper_100__ap_start),
    .C_drain_IO_L1_out_wrapper_100__ap_ready(C_drain_IO_L1_out_wrapper_100__ap_ready),
    .C_drain_IO_L1_out_wrapper_100__ap_done(C_drain_IO_L1_out_wrapper_100__ap_done),
    .C_drain_IO_L1_out_wrapper_100__ap_idle(C_drain_IO_L1_out_wrapper_100__ap_idle),
    .C_drain_IO_L1_out_wrapper_101__ap_start(C_drain_IO_L1_out_wrapper_101__ap_start),
    .C_drain_IO_L1_out_wrapper_101__ap_ready(C_drain_IO_L1_out_wrapper_101__ap_ready),
    .C_drain_IO_L1_out_wrapper_101__ap_done(C_drain_IO_L1_out_wrapper_101__ap_done),
    .C_drain_IO_L1_out_wrapper_101__ap_idle(C_drain_IO_L1_out_wrapper_101__ap_idle),
    .C_drain_IO_L1_out_wrapper_102__ap_start(C_drain_IO_L1_out_wrapper_102__ap_start),
    .C_drain_IO_L1_out_wrapper_102__ap_ready(C_drain_IO_L1_out_wrapper_102__ap_ready),
    .C_drain_IO_L1_out_wrapper_102__ap_done(C_drain_IO_L1_out_wrapper_102__ap_done),
    .C_drain_IO_L1_out_wrapper_102__ap_idle(C_drain_IO_L1_out_wrapper_102__ap_idle),
    .C_drain_IO_L1_out_wrapper_103__ap_start(C_drain_IO_L1_out_wrapper_103__ap_start),
    .C_drain_IO_L1_out_wrapper_103__ap_ready(C_drain_IO_L1_out_wrapper_103__ap_ready),
    .C_drain_IO_L1_out_wrapper_103__ap_done(C_drain_IO_L1_out_wrapper_103__ap_done),
    .C_drain_IO_L1_out_wrapper_103__ap_idle(C_drain_IO_L1_out_wrapper_103__ap_idle),
    .C_drain_IO_L1_out_wrapper_104__ap_start(C_drain_IO_L1_out_wrapper_104__ap_start),
    .C_drain_IO_L1_out_wrapper_104__ap_ready(C_drain_IO_L1_out_wrapper_104__ap_ready),
    .C_drain_IO_L1_out_wrapper_104__ap_done(C_drain_IO_L1_out_wrapper_104__ap_done),
    .C_drain_IO_L1_out_wrapper_104__ap_idle(C_drain_IO_L1_out_wrapper_104__ap_idle),
    .C_drain_IO_L1_out_wrapper_105__ap_start(C_drain_IO_L1_out_wrapper_105__ap_start),
    .C_drain_IO_L1_out_wrapper_105__ap_ready(C_drain_IO_L1_out_wrapper_105__ap_ready),
    .C_drain_IO_L1_out_wrapper_105__ap_done(C_drain_IO_L1_out_wrapper_105__ap_done),
    .C_drain_IO_L1_out_wrapper_105__ap_idle(C_drain_IO_L1_out_wrapper_105__ap_idle),
    .C_drain_IO_L1_out_wrapper_106__ap_start(C_drain_IO_L1_out_wrapper_106__ap_start),
    .C_drain_IO_L1_out_wrapper_106__ap_ready(C_drain_IO_L1_out_wrapper_106__ap_ready),
    .C_drain_IO_L1_out_wrapper_106__ap_done(C_drain_IO_L1_out_wrapper_106__ap_done),
    .C_drain_IO_L1_out_wrapper_106__ap_idle(C_drain_IO_L1_out_wrapper_106__ap_idle),
    .C_drain_IO_L1_out_wrapper_107__ap_start(C_drain_IO_L1_out_wrapper_107__ap_start),
    .C_drain_IO_L1_out_wrapper_107__ap_ready(C_drain_IO_L1_out_wrapper_107__ap_ready),
    .C_drain_IO_L1_out_wrapper_107__ap_done(C_drain_IO_L1_out_wrapper_107__ap_done),
    .C_drain_IO_L1_out_wrapper_107__ap_idle(C_drain_IO_L1_out_wrapper_107__ap_idle),
    .C_drain_IO_L1_out_wrapper_108__ap_start(C_drain_IO_L1_out_wrapper_108__ap_start),
    .C_drain_IO_L1_out_wrapper_108__ap_ready(C_drain_IO_L1_out_wrapper_108__ap_ready),
    .C_drain_IO_L1_out_wrapper_108__ap_done(C_drain_IO_L1_out_wrapper_108__ap_done),
    .C_drain_IO_L1_out_wrapper_108__ap_idle(C_drain_IO_L1_out_wrapper_108__ap_idle),
    .C_drain_IO_L1_out_wrapper_109__ap_start(C_drain_IO_L1_out_wrapper_109__ap_start),
    .C_drain_IO_L1_out_wrapper_109__ap_ready(C_drain_IO_L1_out_wrapper_109__ap_ready),
    .C_drain_IO_L1_out_wrapper_109__ap_done(C_drain_IO_L1_out_wrapper_109__ap_done),
    .C_drain_IO_L1_out_wrapper_109__ap_idle(C_drain_IO_L1_out_wrapper_109__ap_idle),
    .C_drain_IO_L1_out_wrapper_110__ap_start(C_drain_IO_L1_out_wrapper_110__ap_start),
    .C_drain_IO_L1_out_wrapper_110__ap_ready(C_drain_IO_L1_out_wrapper_110__ap_ready),
    .C_drain_IO_L1_out_wrapper_110__ap_done(C_drain_IO_L1_out_wrapper_110__ap_done),
    .C_drain_IO_L1_out_wrapper_110__ap_idle(C_drain_IO_L1_out_wrapper_110__ap_idle),
    .C_drain_IO_L1_out_wrapper_111__ap_start(C_drain_IO_L1_out_wrapper_111__ap_start),
    .C_drain_IO_L1_out_wrapper_111__ap_ready(C_drain_IO_L1_out_wrapper_111__ap_ready),
    .C_drain_IO_L1_out_wrapper_111__ap_done(C_drain_IO_L1_out_wrapper_111__ap_done),
    .C_drain_IO_L1_out_wrapper_111__ap_idle(C_drain_IO_L1_out_wrapper_111__ap_idle),
    .C_drain_IO_L1_out_wrapper_112__ap_start(C_drain_IO_L1_out_wrapper_112__ap_start),
    .C_drain_IO_L1_out_wrapper_112__ap_ready(C_drain_IO_L1_out_wrapper_112__ap_ready),
    .C_drain_IO_L1_out_wrapper_112__ap_done(C_drain_IO_L1_out_wrapper_112__ap_done),
    .C_drain_IO_L1_out_wrapper_112__ap_idle(C_drain_IO_L1_out_wrapper_112__ap_idle),
    .C_drain_IO_L1_out_wrapper_113__ap_start(C_drain_IO_L1_out_wrapper_113__ap_start),
    .C_drain_IO_L1_out_wrapper_113__ap_ready(C_drain_IO_L1_out_wrapper_113__ap_ready),
    .C_drain_IO_L1_out_wrapper_113__ap_done(C_drain_IO_L1_out_wrapper_113__ap_done),
    .C_drain_IO_L1_out_wrapper_113__ap_idle(C_drain_IO_L1_out_wrapper_113__ap_idle),
    .C_drain_IO_L1_out_wrapper_114__ap_start(C_drain_IO_L1_out_wrapper_114__ap_start),
    .C_drain_IO_L1_out_wrapper_114__ap_ready(C_drain_IO_L1_out_wrapper_114__ap_ready),
    .C_drain_IO_L1_out_wrapper_114__ap_done(C_drain_IO_L1_out_wrapper_114__ap_done),
    .C_drain_IO_L1_out_wrapper_114__ap_idle(C_drain_IO_L1_out_wrapper_114__ap_idle),
    .C_drain_IO_L1_out_wrapper_115__ap_start(C_drain_IO_L1_out_wrapper_115__ap_start),
    .C_drain_IO_L1_out_wrapper_115__ap_ready(C_drain_IO_L1_out_wrapper_115__ap_ready),
    .C_drain_IO_L1_out_wrapper_115__ap_done(C_drain_IO_L1_out_wrapper_115__ap_done),
    .C_drain_IO_L1_out_wrapper_115__ap_idle(C_drain_IO_L1_out_wrapper_115__ap_idle),
    .C_drain_IO_L1_out_wrapper_116__ap_start(C_drain_IO_L1_out_wrapper_116__ap_start),
    .C_drain_IO_L1_out_wrapper_116__ap_ready(C_drain_IO_L1_out_wrapper_116__ap_ready),
    .C_drain_IO_L1_out_wrapper_116__ap_done(C_drain_IO_L1_out_wrapper_116__ap_done),
    .C_drain_IO_L1_out_wrapper_116__ap_idle(C_drain_IO_L1_out_wrapper_116__ap_idle),
    .C_drain_IO_L1_out_wrapper_117__ap_start(C_drain_IO_L1_out_wrapper_117__ap_start),
    .C_drain_IO_L1_out_wrapper_117__ap_ready(C_drain_IO_L1_out_wrapper_117__ap_ready),
    .C_drain_IO_L1_out_wrapper_117__ap_done(C_drain_IO_L1_out_wrapper_117__ap_done),
    .C_drain_IO_L1_out_wrapper_117__ap_idle(C_drain_IO_L1_out_wrapper_117__ap_idle),
    .C_drain_IO_L1_out_wrapper_118__ap_start(C_drain_IO_L1_out_wrapper_118__ap_start),
    .C_drain_IO_L1_out_wrapper_118__ap_ready(C_drain_IO_L1_out_wrapper_118__ap_ready),
    .C_drain_IO_L1_out_wrapper_118__ap_done(C_drain_IO_L1_out_wrapper_118__ap_done),
    .C_drain_IO_L1_out_wrapper_118__ap_idle(C_drain_IO_L1_out_wrapper_118__ap_idle),
    .C_drain_IO_L1_out_wrapper_119__ap_start(C_drain_IO_L1_out_wrapper_119__ap_start),
    .C_drain_IO_L1_out_wrapper_119__ap_ready(C_drain_IO_L1_out_wrapper_119__ap_ready),
    .C_drain_IO_L1_out_wrapper_119__ap_done(C_drain_IO_L1_out_wrapper_119__ap_done),
    .C_drain_IO_L1_out_wrapper_119__ap_idle(C_drain_IO_L1_out_wrapper_119__ap_idle),
    .C_drain_IO_L1_out_wrapper_120__ap_start(C_drain_IO_L1_out_wrapper_120__ap_start),
    .C_drain_IO_L1_out_wrapper_120__ap_ready(C_drain_IO_L1_out_wrapper_120__ap_ready),
    .C_drain_IO_L1_out_wrapper_120__ap_done(C_drain_IO_L1_out_wrapper_120__ap_done),
    .C_drain_IO_L1_out_wrapper_120__ap_idle(C_drain_IO_L1_out_wrapper_120__ap_idle),
    .C_drain_IO_L1_out_wrapper_121__ap_start(C_drain_IO_L1_out_wrapper_121__ap_start),
    .C_drain_IO_L1_out_wrapper_121__ap_ready(C_drain_IO_L1_out_wrapper_121__ap_ready),
    .C_drain_IO_L1_out_wrapper_121__ap_done(C_drain_IO_L1_out_wrapper_121__ap_done),
    .C_drain_IO_L1_out_wrapper_121__ap_idle(C_drain_IO_L1_out_wrapper_121__ap_idle),
    .C_drain_IO_L1_out_wrapper_122__ap_start(C_drain_IO_L1_out_wrapper_122__ap_start),
    .C_drain_IO_L1_out_wrapper_122__ap_ready(C_drain_IO_L1_out_wrapper_122__ap_ready),
    .C_drain_IO_L1_out_wrapper_122__ap_done(C_drain_IO_L1_out_wrapper_122__ap_done),
    .C_drain_IO_L1_out_wrapper_122__ap_idle(C_drain_IO_L1_out_wrapper_122__ap_idle),
    .C_drain_IO_L1_out_wrapper_123__ap_start(C_drain_IO_L1_out_wrapper_123__ap_start),
    .C_drain_IO_L1_out_wrapper_123__ap_ready(C_drain_IO_L1_out_wrapper_123__ap_ready),
    .C_drain_IO_L1_out_wrapper_123__ap_done(C_drain_IO_L1_out_wrapper_123__ap_done),
    .C_drain_IO_L1_out_wrapper_123__ap_idle(C_drain_IO_L1_out_wrapper_123__ap_idle),
    .C_drain_IO_L1_out_wrapper_124__ap_start(C_drain_IO_L1_out_wrapper_124__ap_start),
    .C_drain_IO_L1_out_wrapper_124__ap_ready(C_drain_IO_L1_out_wrapper_124__ap_ready),
    .C_drain_IO_L1_out_wrapper_124__ap_done(C_drain_IO_L1_out_wrapper_124__ap_done),
    .C_drain_IO_L1_out_wrapper_124__ap_idle(C_drain_IO_L1_out_wrapper_124__ap_idle),
    .C_drain_IO_L1_out_wrapper_125__ap_start(C_drain_IO_L1_out_wrapper_125__ap_start),
    .C_drain_IO_L1_out_wrapper_125__ap_ready(C_drain_IO_L1_out_wrapper_125__ap_ready),
    .C_drain_IO_L1_out_wrapper_125__ap_done(C_drain_IO_L1_out_wrapper_125__ap_done),
    .C_drain_IO_L1_out_wrapper_125__ap_idle(C_drain_IO_L1_out_wrapper_125__ap_idle),
    .C_drain_IO_L1_out_wrapper_126__ap_start(C_drain_IO_L1_out_wrapper_126__ap_start),
    .C_drain_IO_L1_out_wrapper_126__ap_ready(C_drain_IO_L1_out_wrapper_126__ap_ready),
    .C_drain_IO_L1_out_wrapper_126__ap_done(C_drain_IO_L1_out_wrapper_126__ap_done),
    .C_drain_IO_L1_out_wrapper_126__ap_idle(C_drain_IO_L1_out_wrapper_126__ap_idle),
    .C_drain_IO_L1_out_wrapper_127__ap_start(C_drain_IO_L1_out_wrapper_127__ap_start),
    .C_drain_IO_L1_out_wrapper_127__ap_ready(C_drain_IO_L1_out_wrapper_127__ap_ready),
    .C_drain_IO_L1_out_wrapper_127__ap_done(C_drain_IO_L1_out_wrapper_127__ap_done),
    .C_drain_IO_L1_out_wrapper_127__ap_idle(C_drain_IO_L1_out_wrapper_127__ap_idle),
    .C_drain_IO_L1_out_wrapper_128__ap_start(C_drain_IO_L1_out_wrapper_128__ap_start),
    .C_drain_IO_L1_out_wrapper_128__ap_ready(C_drain_IO_L1_out_wrapper_128__ap_ready),
    .C_drain_IO_L1_out_wrapper_128__ap_done(C_drain_IO_L1_out_wrapper_128__ap_done),
    .C_drain_IO_L1_out_wrapper_128__ap_idle(C_drain_IO_L1_out_wrapper_128__ap_idle),
    .C_drain_IO_L1_out_wrapper_129__ap_start(C_drain_IO_L1_out_wrapper_129__ap_start),
    .C_drain_IO_L1_out_wrapper_129__ap_ready(C_drain_IO_L1_out_wrapper_129__ap_ready),
    .C_drain_IO_L1_out_wrapper_129__ap_done(C_drain_IO_L1_out_wrapper_129__ap_done),
    .C_drain_IO_L1_out_wrapper_129__ap_idle(C_drain_IO_L1_out_wrapper_129__ap_idle),
    .C_drain_IO_L1_out_wrapper_130__ap_start(C_drain_IO_L1_out_wrapper_130__ap_start),
    .C_drain_IO_L1_out_wrapper_130__ap_ready(C_drain_IO_L1_out_wrapper_130__ap_ready),
    .C_drain_IO_L1_out_wrapper_130__ap_done(C_drain_IO_L1_out_wrapper_130__ap_done),
    .C_drain_IO_L1_out_wrapper_130__ap_idle(C_drain_IO_L1_out_wrapper_130__ap_idle),
    .C_drain_IO_L1_out_wrapper_131__ap_start(C_drain_IO_L1_out_wrapper_131__ap_start),
    .C_drain_IO_L1_out_wrapper_131__ap_ready(C_drain_IO_L1_out_wrapper_131__ap_ready),
    .C_drain_IO_L1_out_wrapper_131__ap_done(C_drain_IO_L1_out_wrapper_131__ap_done),
    .C_drain_IO_L1_out_wrapper_131__ap_idle(C_drain_IO_L1_out_wrapper_131__ap_idle),
    .C_drain_IO_L1_out_wrapper_132__ap_start(C_drain_IO_L1_out_wrapper_132__ap_start),
    .C_drain_IO_L1_out_wrapper_132__ap_ready(C_drain_IO_L1_out_wrapper_132__ap_ready),
    .C_drain_IO_L1_out_wrapper_132__ap_done(C_drain_IO_L1_out_wrapper_132__ap_done),
    .C_drain_IO_L1_out_wrapper_132__ap_idle(C_drain_IO_L1_out_wrapper_132__ap_idle),
    .C_drain_IO_L1_out_wrapper_133__ap_start(C_drain_IO_L1_out_wrapper_133__ap_start),
    .C_drain_IO_L1_out_wrapper_133__ap_ready(C_drain_IO_L1_out_wrapper_133__ap_ready),
    .C_drain_IO_L1_out_wrapper_133__ap_done(C_drain_IO_L1_out_wrapper_133__ap_done),
    .C_drain_IO_L1_out_wrapper_133__ap_idle(C_drain_IO_L1_out_wrapper_133__ap_idle),
    .C_drain_IO_L1_out_wrapper_134__ap_start(C_drain_IO_L1_out_wrapper_134__ap_start),
    .C_drain_IO_L1_out_wrapper_134__ap_ready(C_drain_IO_L1_out_wrapper_134__ap_ready),
    .C_drain_IO_L1_out_wrapper_134__ap_done(C_drain_IO_L1_out_wrapper_134__ap_done),
    .C_drain_IO_L1_out_wrapper_134__ap_idle(C_drain_IO_L1_out_wrapper_134__ap_idle),
    .C_drain_IO_L1_out_wrapper_135__ap_start(C_drain_IO_L1_out_wrapper_135__ap_start),
    .C_drain_IO_L1_out_wrapper_135__ap_ready(C_drain_IO_L1_out_wrapper_135__ap_ready),
    .C_drain_IO_L1_out_wrapper_135__ap_done(C_drain_IO_L1_out_wrapper_135__ap_done),
    .C_drain_IO_L1_out_wrapper_135__ap_idle(C_drain_IO_L1_out_wrapper_135__ap_idle),
    .C_drain_IO_L1_out_wrapper_136__ap_start(C_drain_IO_L1_out_wrapper_136__ap_start),
    .C_drain_IO_L1_out_wrapper_136__ap_ready(C_drain_IO_L1_out_wrapper_136__ap_ready),
    .C_drain_IO_L1_out_wrapper_136__ap_done(C_drain_IO_L1_out_wrapper_136__ap_done),
    .C_drain_IO_L1_out_wrapper_136__ap_idle(C_drain_IO_L1_out_wrapper_136__ap_idle),
    .C_drain_IO_L1_out_wrapper_137__ap_start(C_drain_IO_L1_out_wrapper_137__ap_start),
    .C_drain_IO_L1_out_wrapper_137__ap_ready(C_drain_IO_L1_out_wrapper_137__ap_ready),
    .C_drain_IO_L1_out_wrapper_137__ap_done(C_drain_IO_L1_out_wrapper_137__ap_done),
    .C_drain_IO_L1_out_wrapper_137__ap_idle(C_drain_IO_L1_out_wrapper_137__ap_idle),
    .C_drain_IO_L1_out_wrapper_138__ap_start(C_drain_IO_L1_out_wrapper_138__ap_start),
    .C_drain_IO_L1_out_wrapper_138__ap_ready(C_drain_IO_L1_out_wrapper_138__ap_ready),
    .C_drain_IO_L1_out_wrapper_138__ap_done(C_drain_IO_L1_out_wrapper_138__ap_done),
    .C_drain_IO_L1_out_wrapper_138__ap_idle(C_drain_IO_L1_out_wrapper_138__ap_idle),
    .C_drain_IO_L1_out_wrapper_139__ap_start(C_drain_IO_L1_out_wrapper_139__ap_start),
    .C_drain_IO_L1_out_wrapper_139__ap_ready(C_drain_IO_L1_out_wrapper_139__ap_ready),
    .C_drain_IO_L1_out_wrapper_139__ap_done(C_drain_IO_L1_out_wrapper_139__ap_done),
    .C_drain_IO_L1_out_wrapper_139__ap_idle(C_drain_IO_L1_out_wrapper_139__ap_idle),
    .C_drain_IO_L1_out_wrapper_140__ap_start(C_drain_IO_L1_out_wrapper_140__ap_start),
    .C_drain_IO_L1_out_wrapper_140__ap_ready(C_drain_IO_L1_out_wrapper_140__ap_ready),
    .C_drain_IO_L1_out_wrapper_140__ap_done(C_drain_IO_L1_out_wrapper_140__ap_done),
    .C_drain_IO_L1_out_wrapper_140__ap_idle(C_drain_IO_L1_out_wrapper_140__ap_idle),
    .C_drain_IO_L1_out_wrapper_141__ap_start(C_drain_IO_L1_out_wrapper_141__ap_start),
    .C_drain_IO_L1_out_wrapper_141__ap_ready(C_drain_IO_L1_out_wrapper_141__ap_ready),
    .C_drain_IO_L1_out_wrapper_141__ap_done(C_drain_IO_L1_out_wrapper_141__ap_done),
    .C_drain_IO_L1_out_wrapper_141__ap_idle(C_drain_IO_L1_out_wrapper_141__ap_idle),
    .C_drain_IO_L1_out_wrapper_142__ap_start(C_drain_IO_L1_out_wrapper_142__ap_start),
    .C_drain_IO_L1_out_wrapper_142__ap_ready(C_drain_IO_L1_out_wrapper_142__ap_ready),
    .C_drain_IO_L1_out_wrapper_142__ap_done(C_drain_IO_L1_out_wrapper_142__ap_done),
    .C_drain_IO_L1_out_wrapper_142__ap_idle(C_drain_IO_L1_out_wrapper_142__ap_idle),
    .C_drain_IO_L1_out_wrapper_143__ap_start(C_drain_IO_L1_out_wrapper_143__ap_start),
    .C_drain_IO_L1_out_wrapper_143__ap_ready(C_drain_IO_L1_out_wrapper_143__ap_ready),
    .C_drain_IO_L1_out_wrapper_143__ap_done(C_drain_IO_L1_out_wrapper_143__ap_done),
    .C_drain_IO_L1_out_wrapper_143__ap_idle(C_drain_IO_L1_out_wrapper_143__ap_idle),
    .C_drain_IO_L1_out_wrapper_144__ap_start(C_drain_IO_L1_out_wrapper_144__ap_start),
    .C_drain_IO_L1_out_wrapper_144__ap_ready(C_drain_IO_L1_out_wrapper_144__ap_ready),
    .C_drain_IO_L1_out_wrapper_144__ap_done(C_drain_IO_L1_out_wrapper_144__ap_done),
    .C_drain_IO_L1_out_wrapper_144__ap_idle(C_drain_IO_L1_out_wrapper_144__ap_idle),
    .C_drain_IO_L1_out_wrapper_145__ap_start(C_drain_IO_L1_out_wrapper_145__ap_start),
    .C_drain_IO_L1_out_wrapper_145__ap_ready(C_drain_IO_L1_out_wrapper_145__ap_ready),
    .C_drain_IO_L1_out_wrapper_145__ap_done(C_drain_IO_L1_out_wrapper_145__ap_done),
    .C_drain_IO_L1_out_wrapper_145__ap_idle(C_drain_IO_L1_out_wrapper_145__ap_idle),
    .C_drain_IO_L1_out_wrapper_146__ap_start(C_drain_IO_L1_out_wrapper_146__ap_start),
    .C_drain_IO_L1_out_wrapper_146__ap_ready(C_drain_IO_L1_out_wrapper_146__ap_ready),
    .C_drain_IO_L1_out_wrapper_146__ap_done(C_drain_IO_L1_out_wrapper_146__ap_done),
    .C_drain_IO_L1_out_wrapper_146__ap_idle(C_drain_IO_L1_out_wrapper_146__ap_idle),
    .C_drain_IO_L1_out_wrapper_147__ap_start(C_drain_IO_L1_out_wrapper_147__ap_start),
    .C_drain_IO_L1_out_wrapper_147__ap_ready(C_drain_IO_L1_out_wrapper_147__ap_ready),
    .C_drain_IO_L1_out_wrapper_147__ap_done(C_drain_IO_L1_out_wrapper_147__ap_done),
    .C_drain_IO_L1_out_wrapper_147__ap_idle(C_drain_IO_L1_out_wrapper_147__ap_idle),
    .C_drain_IO_L1_out_wrapper_148__ap_start(C_drain_IO_L1_out_wrapper_148__ap_start),
    .C_drain_IO_L1_out_wrapper_148__ap_ready(C_drain_IO_L1_out_wrapper_148__ap_ready),
    .C_drain_IO_L1_out_wrapper_148__ap_done(C_drain_IO_L1_out_wrapper_148__ap_done),
    .C_drain_IO_L1_out_wrapper_148__ap_idle(C_drain_IO_L1_out_wrapper_148__ap_idle),
    .C_drain_IO_L1_out_wrapper_149__ap_start(C_drain_IO_L1_out_wrapper_149__ap_start),
    .C_drain_IO_L1_out_wrapper_149__ap_ready(C_drain_IO_L1_out_wrapper_149__ap_ready),
    .C_drain_IO_L1_out_wrapper_149__ap_done(C_drain_IO_L1_out_wrapper_149__ap_done),
    .C_drain_IO_L1_out_wrapper_149__ap_idle(C_drain_IO_L1_out_wrapper_149__ap_idle),
    .C_drain_IO_L1_out_wrapper_150__ap_start(C_drain_IO_L1_out_wrapper_150__ap_start),
    .C_drain_IO_L1_out_wrapper_150__ap_ready(C_drain_IO_L1_out_wrapper_150__ap_ready),
    .C_drain_IO_L1_out_wrapper_150__ap_done(C_drain_IO_L1_out_wrapper_150__ap_done),
    .C_drain_IO_L1_out_wrapper_150__ap_idle(C_drain_IO_L1_out_wrapper_150__ap_idle),
    .C_drain_IO_L1_out_wrapper_151__ap_start(C_drain_IO_L1_out_wrapper_151__ap_start),
    .C_drain_IO_L1_out_wrapper_151__ap_ready(C_drain_IO_L1_out_wrapper_151__ap_ready),
    .C_drain_IO_L1_out_wrapper_151__ap_done(C_drain_IO_L1_out_wrapper_151__ap_done),
    .C_drain_IO_L1_out_wrapper_151__ap_idle(C_drain_IO_L1_out_wrapper_151__ap_idle),
    .C_drain_IO_L1_out_wrapper_152__ap_start(C_drain_IO_L1_out_wrapper_152__ap_start),
    .C_drain_IO_L1_out_wrapper_152__ap_ready(C_drain_IO_L1_out_wrapper_152__ap_ready),
    .C_drain_IO_L1_out_wrapper_152__ap_done(C_drain_IO_L1_out_wrapper_152__ap_done),
    .C_drain_IO_L1_out_wrapper_152__ap_idle(C_drain_IO_L1_out_wrapper_152__ap_idle),
    .C_drain_IO_L1_out_wrapper_153__ap_start(C_drain_IO_L1_out_wrapper_153__ap_start),
    .C_drain_IO_L1_out_wrapper_153__ap_ready(C_drain_IO_L1_out_wrapper_153__ap_ready),
    .C_drain_IO_L1_out_wrapper_153__ap_done(C_drain_IO_L1_out_wrapper_153__ap_done),
    .C_drain_IO_L1_out_wrapper_153__ap_idle(C_drain_IO_L1_out_wrapper_153__ap_idle),
    .C_drain_IO_L1_out_wrapper_154__ap_start(C_drain_IO_L1_out_wrapper_154__ap_start),
    .C_drain_IO_L1_out_wrapper_154__ap_ready(C_drain_IO_L1_out_wrapper_154__ap_ready),
    .C_drain_IO_L1_out_wrapper_154__ap_done(C_drain_IO_L1_out_wrapper_154__ap_done),
    .C_drain_IO_L1_out_wrapper_154__ap_idle(C_drain_IO_L1_out_wrapper_154__ap_idle),
    .C_drain_IO_L1_out_wrapper_155__ap_start(C_drain_IO_L1_out_wrapper_155__ap_start),
    .C_drain_IO_L1_out_wrapper_155__ap_ready(C_drain_IO_L1_out_wrapper_155__ap_ready),
    .C_drain_IO_L1_out_wrapper_155__ap_done(C_drain_IO_L1_out_wrapper_155__ap_done),
    .C_drain_IO_L1_out_wrapper_155__ap_idle(C_drain_IO_L1_out_wrapper_155__ap_idle),
    .C_drain_IO_L1_out_wrapper_156__ap_start(C_drain_IO_L1_out_wrapper_156__ap_start),
    .C_drain_IO_L1_out_wrapper_156__ap_ready(C_drain_IO_L1_out_wrapper_156__ap_ready),
    .C_drain_IO_L1_out_wrapper_156__ap_done(C_drain_IO_L1_out_wrapper_156__ap_done),
    .C_drain_IO_L1_out_wrapper_156__ap_idle(C_drain_IO_L1_out_wrapper_156__ap_idle),
    .C_drain_IO_L1_out_wrapper_157__ap_start(C_drain_IO_L1_out_wrapper_157__ap_start),
    .C_drain_IO_L1_out_wrapper_157__ap_ready(C_drain_IO_L1_out_wrapper_157__ap_ready),
    .C_drain_IO_L1_out_wrapper_157__ap_done(C_drain_IO_L1_out_wrapper_157__ap_done),
    .C_drain_IO_L1_out_wrapper_157__ap_idle(C_drain_IO_L1_out_wrapper_157__ap_idle),
    .C_drain_IO_L1_out_wrapper_158__ap_start(C_drain_IO_L1_out_wrapper_158__ap_start),
    .C_drain_IO_L1_out_wrapper_158__ap_ready(C_drain_IO_L1_out_wrapper_158__ap_ready),
    .C_drain_IO_L1_out_wrapper_158__ap_done(C_drain_IO_L1_out_wrapper_158__ap_done),
    .C_drain_IO_L1_out_wrapper_158__ap_idle(C_drain_IO_L1_out_wrapper_158__ap_idle),
    .C_drain_IO_L1_out_wrapper_159__ap_start(C_drain_IO_L1_out_wrapper_159__ap_start),
    .C_drain_IO_L1_out_wrapper_159__ap_ready(C_drain_IO_L1_out_wrapper_159__ap_ready),
    .C_drain_IO_L1_out_wrapper_159__ap_done(C_drain_IO_L1_out_wrapper_159__ap_done),
    .C_drain_IO_L1_out_wrapper_159__ap_idle(C_drain_IO_L1_out_wrapper_159__ap_idle),
    .C_drain_IO_L1_out_wrapper_160__ap_start(C_drain_IO_L1_out_wrapper_160__ap_start),
    .C_drain_IO_L1_out_wrapper_160__ap_ready(C_drain_IO_L1_out_wrapper_160__ap_ready),
    .C_drain_IO_L1_out_wrapper_160__ap_done(C_drain_IO_L1_out_wrapper_160__ap_done),
    .C_drain_IO_L1_out_wrapper_160__ap_idle(C_drain_IO_L1_out_wrapper_160__ap_idle),
    .C_drain_IO_L1_out_wrapper_161__ap_start(C_drain_IO_L1_out_wrapper_161__ap_start),
    .C_drain_IO_L1_out_wrapper_161__ap_ready(C_drain_IO_L1_out_wrapper_161__ap_ready),
    .C_drain_IO_L1_out_wrapper_161__ap_done(C_drain_IO_L1_out_wrapper_161__ap_done),
    .C_drain_IO_L1_out_wrapper_161__ap_idle(C_drain_IO_L1_out_wrapper_161__ap_idle),
    .C_drain_IO_L1_out_wrapper_162__ap_start(C_drain_IO_L1_out_wrapper_162__ap_start),
    .C_drain_IO_L1_out_wrapper_162__ap_ready(C_drain_IO_L1_out_wrapper_162__ap_ready),
    .C_drain_IO_L1_out_wrapper_162__ap_done(C_drain_IO_L1_out_wrapper_162__ap_done),
    .C_drain_IO_L1_out_wrapper_162__ap_idle(C_drain_IO_L1_out_wrapper_162__ap_idle),
    .C_drain_IO_L1_out_wrapper_163__ap_start(C_drain_IO_L1_out_wrapper_163__ap_start),
    .C_drain_IO_L1_out_wrapper_163__ap_ready(C_drain_IO_L1_out_wrapper_163__ap_ready),
    .C_drain_IO_L1_out_wrapper_163__ap_done(C_drain_IO_L1_out_wrapper_163__ap_done),
    .C_drain_IO_L1_out_wrapper_163__ap_idle(C_drain_IO_L1_out_wrapper_163__ap_idle),
    .C_drain_IO_L1_out_wrapper_164__ap_start(C_drain_IO_L1_out_wrapper_164__ap_start),
    .C_drain_IO_L1_out_wrapper_164__ap_ready(C_drain_IO_L1_out_wrapper_164__ap_ready),
    .C_drain_IO_L1_out_wrapper_164__ap_done(C_drain_IO_L1_out_wrapper_164__ap_done),
    .C_drain_IO_L1_out_wrapper_164__ap_idle(C_drain_IO_L1_out_wrapper_164__ap_idle),
    .C_drain_IO_L1_out_wrapper_165__ap_start(C_drain_IO_L1_out_wrapper_165__ap_start),
    .C_drain_IO_L1_out_wrapper_165__ap_ready(C_drain_IO_L1_out_wrapper_165__ap_ready),
    .C_drain_IO_L1_out_wrapper_165__ap_done(C_drain_IO_L1_out_wrapper_165__ap_done),
    .C_drain_IO_L1_out_wrapper_165__ap_idle(C_drain_IO_L1_out_wrapper_165__ap_idle),
    .C_drain_IO_L1_out_wrapper_166__ap_start(C_drain_IO_L1_out_wrapper_166__ap_start),
    .C_drain_IO_L1_out_wrapper_166__ap_ready(C_drain_IO_L1_out_wrapper_166__ap_ready),
    .C_drain_IO_L1_out_wrapper_166__ap_done(C_drain_IO_L1_out_wrapper_166__ap_done),
    .C_drain_IO_L1_out_wrapper_166__ap_idle(C_drain_IO_L1_out_wrapper_166__ap_idle),
    .C_drain_IO_L1_out_wrapper_167__ap_start(C_drain_IO_L1_out_wrapper_167__ap_start),
    .C_drain_IO_L1_out_wrapper_167__ap_ready(C_drain_IO_L1_out_wrapper_167__ap_ready),
    .C_drain_IO_L1_out_wrapper_167__ap_done(C_drain_IO_L1_out_wrapper_167__ap_done),
    .C_drain_IO_L1_out_wrapper_167__ap_idle(C_drain_IO_L1_out_wrapper_167__ap_idle),
    .C_drain_IO_L1_out_wrapper_168__ap_start(C_drain_IO_L1_out_wrapper_168__ap_start),
    .C_drain_IO_L1_out_wrapper_168__ap_ready(C_drain_IO_L1_out_wrapper_168__ap_ready),
    .C_drain_IO_L1_out_wrapper_168__ap_done(C_drain_IO_L1_out_wrapper_168__ap_done),
    .C_drain_IO_L1_out_wrapper_168__ap_idle(C_drain_IO_L1_out_wrapper_168__ap_idle),
    .C_drain_IO_L1_out_wrapper_169__ap_start(C_drain_IO_L1_out_wrapper_169__ap_start),
    .C_drain_IO_L1_out_wrapper_169__ap_ready(C_drain_IO_L1_out_wrapper_169__ap_ready),
    .C_drain_IO_L1_out_wrapper_169__ap_done(C_drain_IO_L1_out_wrapper_169__ap_done),
    .C_drain_IO_L1_out_wrapper_169__ap_idle(C_drain_IO_L1_out_wrapper_169__ap_idle),
    .C_drain_IO_L1_out_wrapper_170__ap_start(C_drain_IO_L1_out_wrapper_170__ap_start),
    .C_drain_IO_L1_out_wrapper_170__ap_ready(C_drain_IO_L1_out_wrapper_170__ap_ready),
    .C_drain_IO_L1_out_wrapper_170__ap_done(C_drain_IO_L1_out_wrapper_170__ap_done),
    .C_drain_IO_L1_out_wrapper_170__ap_idle(C_drain_IO_L1_out_wrapper_170__ap_idle),
    .C_drain_IO_L1_out_wrapper_171__ap_start(C_drain_IO_L1_out_wrapper_171__ap_start),
    .C_drain_IO_L1_out_wrapper_171__ap_ready(C_drain_IO_L1_out_wrapper_171__ap_ready),
    .C_drain_IO_L1_out_wrapper_171__ap_done(C_drain_IO_L1_out_wrapper_171__ap_done),
    .C_drain_IO_L1_out_wrapper_171__ap_idle(C_drain_IO_L1_out_wrapper_171__ap_idle),
    .C_drain_IO_L1_out_wrapper_172__ap_start(C_drain_IO_L1_out_wrapper_172__ap_start),
    .C_drain_IO_L1_out_wrapper_172__ap_ready(C_drain_IO_L1_out_wrapper_172__ap_ready),
    .C_drain_IO_L1_out_wrapper_172__ap_done(C_drain_IO_L1_out_wrapper_172__ap_done),
    .C_drain_IO_L1_out_wrapper_172__ap_idle(C_drain_IO_L1_out_wrapper_172__ap_idle),
    .C_drain_IO_L1_out_wrapper_173__ap_start(C_drain_IO_L1_out_wrapper_173__ap_start),
    .C_drain_IO_L1_out_wrapper_173__ap_ready(C_drain_IO_L1_out_wrapper_173__ap_ready),
    .C_drain_IO_L1_out_wrapper_173__ap_done(C_drain_IO_L1_out_wrapper_173__ap_done),
    .C_drain_IO_L1_out_wrapper_173__ap_idle(C_drain_IO_L1_out_wrapper_173__ap_idle),
    .C_drain_IO_L1_out_wrapper_174__ap_start(C_drain_IO_L1_out_wrapper_174__ap_start),
    .C_drain_IO_L1_out_wrapper_174__ap_ready(C_drain_IO_L1_out_wrapper_174__ap_ready),
    .C_drain_IO_L1_out_wrapper_174__ap_done(C_drain_IO_L1_out_wrapper_174__ap_done),
    .C_drain_IO_L1_out_wrapper_174__ap_idle(C_drain_IO_L1_out_wrapper_174__ap_idle),
    .C_drain_IO_L1_out_wrapper_175__ap_start(C_drain_IO_L1_out_wrapper_175__ap_start),
    .C_drain_IO_L1_out_wrapper_175__ap_ready(C_drain_IO_L1_out_wrapper_175__ap_ready),
    .C_drain_IO_L1_out_wrapper_175__ap_done(C_drain_IO_L1_out_wrapper_175__ap_done),
    .C_drain_IO_L1_out_wrapper_175__ap_idle(C_drain_IO_L1_out_wrapper_175__ap_idle),
    .C_drain_IO_L1_out_wrapper_176__ap_start(C_drain_IO_L1_out_wrapper_176__ap_start),
    .C_drain_IO_L1_out_wrapper_176__ap_ready(C_drain_IO_L1_out_wrapper_176__ap_ready),
    .C_drain_IO_L1_out_wrapper_176__ap_done(C_drain_IO_L1_out_wrapper_176__ap_done),
    .C_drain_IO_L1_out_wrapper_176__ap_idle(C_drain_IO_L1_out_wrapper_176__ap_idle),
    .C_drain_IO_L1_out_wrapper_177__ap_start(C_drain_IO_L1_out_wrapper_177__ap_start),
    .C_drain_IO_L1_out_wrapper_177__ap_ready(C_drain_IO_L1_out_wrapper_177__ap_ready),
    .C_drain_IO_L1_out_wrapper_177__ap_done(C_drain_IO_L1_out_wrapper_177__ap_done),
    .C_drain_IO_L1_out_wrapper_177__ap_idle(C_drain_IO_L1_out_wrapper_177__ap_idle),
    .C_drain_IO_L1_out_wrapper_178__ap_start(C_drain_IO_L1_out_wrapper_178__ap_start),
    .C_drain_IO_L1_out_wrapper_178__ap_ready(C_drain_IO_L1_out_wrapper_178__ap_ready),
    .C_drain_IO_L1_out_wrapper_178__ap_done(C_drain_IO_L1_out_wrapper_178__ap_done),
    .C_drain_IO_L1_out_wrapper_178__ap_idle(C_drain_IO_L1_out_wrapper_178__ap_idle),
    .C_drain_IO_L1_out_wrapper_179__ap_start(C_drain_IO_L1_out_wrapper_179__ap_start),
    .C_drain_IO_L1_out_wrapper_179__ap_ready(C_drain_IO_L1_out_wrapper_179__ap_ready),
    .C_drain_IO_L1_out_wrapper_179__ap_done(C_drain_IO_L1_out_wrapper_179__ap_done),
    .C_drain_IO_L1_out_wrapper_179__ap_idle(C_drain_IO_L1_out_wrapper_179__ap_idle),
    .C_drain_IO_L1_out_wrapper_180__ap_start(C_drain_IO_L1_out_wrapper_180__ap_start),
    .C_drain_IO_L1_out_wrapper_180__ap_ready(C_drain_IO_L1_out_wrapper_180__ap_ready),
    .C_drain_IO_L1_out_wrapper_180__ap_done(C_drain_IO_L1_out_wrapper_180__ap_done),
    .C_drain_IO_L1_out_wrapper_180__ap_idle(C_drain_IO_L1_out_wrapper_180__ap_idle),
    .C_drain_IO_L1_out_wrapper_181__ap_start(C_drain_IO_L1_out_wrapper_181__ap_start),
    .C_drain_IO_L1_out_wrapper_181__ap_ready(C_drain_IO_L1_out_wrapper_181__ap_ready),
    .C_drain_IO_L1_out_wrapper_181__ap_done(C_drain_IO_L1_out_wrapper_181__ap_done),
    .C_drain_IO_L1_out_wrapper_181__ap_idle(C_drain_IO_L1_out_wrapper_181__ap_idle),
    .C_drain_IO_L1_out_wrapper_182__ap_start(C_drain_IO_L1_out_wrapper_182__ap_start),
    .C_drain_IO_L1_out_wrapper_182__ap_ready(C_drain_IO_L1_out_wrapper_182__ap_ready),
    .C_drain_IO_L1_out_wrapper_182__ap_done(C_drain_IO_L1_out_wrapper_182__ap_done),
    .C_drain_IO_L1_out_wrapper_182__ap_idle(C_drain_IO_L1_out_wrapper_182__ap_idle),
    .C_drain_IO_L1_out_wrapper_183__ap_start(C_drain_IO_L1_out_wrapper_183__ap_start),
    .C_drain_IO_L1_out_wrapper_183__ap_ready(C_drain_IO_L1_out_wrapper_183__ap_ready),
    .C_drain_IO_L1_out_wrapper_183__ap_done(C_drain_IO_L1_out_wrapper_183__ap_done),
    .C_drain_IO_L1_out_wrapper_183__ap_idle(C_drain_IO_L1_out_wrapper_183__ap_idle),
    .C_drain_IO_L1_out_wrapper_184__ap_start(C_drain_IO_L1_out_wrapper_184__ap_start),
    .C_drain_IO_L1_out_wrapper_184__ap_ready(C_drain_IO_L1_out_wrapper_184__ap_ready),
    .C_drain_IO_L1_out_wrapper_184__ap_done(C_drain_IO_L1_out_wrapper_184__ap_done),
    .C_drain_IO_L1_out_wrapper_184__ap_idle(C_drain_IO_L1_out_wrapper_184__ap_idle),
    .C_drain_IO_L1_out_wrapper_185__ap_start(C_drain_IO_L1_out_wrapper_185__ap_start),
    .C_drain_IO_L1_out_wrapper_185__ap_ready(C_drain_IO_L1_out_wrapper_185__ap_ready),
    .C_drain_IO_L1_out_wrapper_185__ap_done(C_drain_IO_L1_out_wrapper_185__ap_done),
    .C_drain_IO_L1_out_wrapper_185__ap_idle(C_drain_IO_L1_out_wrapper_185__ap_idle),
    .C_drain_IO_L1_out_wrapper_186__ap_start(C_drain_IO_L1_out_wrapper_186__ap_start),
    .C_drain_IO_L1_out_wrapper_186__ap_ready(C_drain_IO_L1_out_wrapper_186__ap_ready),
    .C_drain_IO_L1_out_wrapper_186__ap_done(C_drain_IO_L1_out_wrapper_186__ap_done),
    .C_drain_IO_L1_out_wrapper_186__ap_idle(C_drain_IO_L1_out_wrapper_186__ap_idle),
    .C_drain_IO_L1_out_wrapper_187__ap_start(C_drain_IO_L1_out_wrapper_187__ap_start),
    .C_drain_IO_L1_out_wrapper_187__ap_ready(C_drain_IO_L1_out_wrapper_187__ap_ready),
    .C_drain_IO_L1_out_wrapper_187__ap_done(C_drain_IO_L1_out_wrapper_187__ap_done),
    .C_drain_IO_L1_out_wrapper_187__ap_idle(C_drain_IO_L1_out_wrapper_187__ap_idle),
    .C_drain_IO_L1_out_wrapper_188__ap_start(C_drain_IO_L1_out_wrapper_188__ap_start),
    .C_drain_IO_L1_out_wrapper_188__ap_ready(C_drain_IO_L1_out_wrapper_188__ap_ready),
    .C_drain_IO_L1_out_wrapper_188__ap_done(C_drain_IO_L1_out_wrapper_188__ap_done),
    .C_drain_IO_L1_out_wrapper_188__ap_idle(C_drain_IO_L1_out_wrapper_188__ap_idle),
    .C_drain_IO_L1_out_wrapper_189__ap_start(C_drain_IO_L1_out_wrapper_189__ap_start),
    .C_drain_IO_L1_out_wrapper_189__ap_ready(C_drain_IO_L1_out_wrapper_189__ap_ready),
    .C_drain_IO_L1_out_wrapper_189__ap_done(C_drain_IO_L1_out_wrapper_189__ap_done),
    .C_drain_IO_L1_out_wrapper_189__ap_idle(C_drain_IO_L1_out_wrapper_189__ap_idle),
    .C_drain_IO_L1_out_wrapper_190__ap_start(C_drain_IO_L1_out_wrapper_190__ap_start),
    .C_drain_IO_L1_out_wrapper_190__ap_ready(C_drain_IO_L1_out_wrapper_190__ap_ready),
    .C_drain_IO_L1_out_wrapper_190__ap_done(C_drain_IO_L1_out_wrapper_190__ap_done),
    .C_drain_IO_L1_out_wrapper_190__ap_idle(C_drain_IO_L1_out_wrapper_190__ap_idle),
    .C_drain_IO_L1_out_wrapper_191__ap_start(C_drain_IO_L1_out_wrapper_191__ap_start),
    .C_drain_IO_L1_out_wrapper_191__ap_ready(C_drain_IO_L1_out_wrapper_191__ap_ready),
    .C_drain_IO_L1_out_wrapper_191__ap_done(C_drain_IO_L1_out_wrapper_191__ap_done),
    .C_drain_IO_L1_out_wrapper_191__ap_idle(C_drain_IO_L1_out_wrapper_191__ap_idle),
    .C_drain_IO_L1_out_wrapper_192__ap_start(C_drain_IO_L1_out_wrapper_192__ap_start),
    .C_drain_IO_L1_out_wrapper_192__ap_ready(C_drain_IO_L1_out_wrapper_192__ap_ready),
    .C_drain_IO_L1_out_wrapper_192__ap_done(C_drain_IO_L1_out_wrapper_192__ap_done),
    .C_drain_IO_L1_out_wrapper_192__ap_idle(C_drain_IO_L1_out_wrapper_192__ap_idle),
    .C_drain_IO_L1_out_wrapper_193__ap_start(C_drain_IO_L1_out_wrapper_193__ap_start),
    .C_drain_IO_L1_out_wrapper_193__ap_ready(C_drain_IO_L1_out_wrapper_193__ap_ready),
    .C_drain_IO_L1_out_wrapper_193__ap_done(C_drain_IO_L1_out_wrapper_193__ap_done),
    .C_drain_IO_L1_out_wrapper_193__ap_idle(C_drain_IO_L1_out_wrapper_193__ap_idle),
    .C_drain_IO_L1_out_wrapper_194__ap_start(C_drain_IO_L1_out_wrapper_194__ap_start),
    .C_drain_IO_L1_out_wrapper_194__ap_ready(C_drain_IO_L1_out_wrapper_194__ap_ready),
    .C_drain_IO_L1_out_wrapper_194__ap_done(C_drain_IO_L1_out_wrapper_194__ap_done),
    .C_drain_IO_L1_out_wrapper_194__ap_idle(C_drain_IO_L1_out_wrapper_194__ap_idle),
    .C_drain_IO_L1_out_wrapper_195__ap_start(C_drain_IO_L1_out_wrapper_195__ap_start),
    .C_drain_IO_L1_out_wrapper_195__ap_ready(C_drain_IO_L1_out_wrapper_195__ap_ready),
    .C_drain_IO_L1_out_wrapper_195__ap_done(C_drain_IO_L1_out_wrapper_195__ap_done),
    .C_drain_IO_L1_out_wrapper_195__ap_idle(C_drain_IO_L1_out_wrapper_195__ap_idle),
    .C_drain_IO_L1_out_wrapper_196__ap_start(C_drain_IO_L1_out_wrapper_196__ap_start),
    .C_drain_IO_L1_out_wrapper_196__ap_ready(C_drain_IO_L1_out_wrapper_196__ap_ready),
    .C_drain_IO_L1_out_wrapper_196__ap_done(C_drain_IO_L1_out_wrapper_196__ap_done),
    .C_drain_IO_L1_out_wrapper_196__ap_idle(C_drain_IO_L1_out_wrapper_196__ap_idle),
    .C_drain_IO_L1_out_wrapper_197__ap_start(C_drain_IO_L1_out_wrapper_197__ap_start),
    .C_drain_IO_L1_out_wrapper_197__ap_ready(C_drain_IO_L1_out_wrapper_197__ap_ready),
    .C_drain_IO_L1_out_wrapper_197__ap_done(C_drain_IO_L1_out_wrapper_197__ap_done),
    .C_drain_IO_L1_out_wrapper_197__ap_idle(C_drain_IO_L1_out_wrapper_197__ap_idle),
    .C_drain_IO_L1_out_wrapper_198__ap_start(C_drain_IO_L1_out_wrapper_198__ap_start),
    .C_drain_IO_L1_out_wrapper_198__ap_ready(C_drain_IO_L1_out_wrapper_198__ap_ready),
    .C_drain_IO_L1_out_wrapper_198__ap_done(C_drain_IO_L1_out_wrapper_198__ap_done),
    .C_drain_IO_L1_out_wrapper_198__ap_idle(C_drain_IO_L1_out_wrapper_198__ap_idle),
    .C_drain_IO_L1_out_wrapper_199__ap_start(C_drain_IO_L1_out_wrapper_199__ap_start),
    .C_drain_IO_L1_out_wrapper_199__ap_ready(C_drain_IO_L1_out_wrapper_199__ap_ready),
    .C_drain_IO_L1_out_wrapper_199__ap_done(C_drain_IO_L1_out_wrapper_199__ap_done),
    .C_drain_IO_L1_out_wrapper_199__ap_idle(C_drain_IO_L1_out_wrapper_199__ap_idle),
    .C_drain_IO_L1_out_wrapper_200__ap_start(C_drain_IO_L1_out_wrapper_200__ap_start),
    .C_drain_IO_L1_out_wrapper_200__ap_ready(C_drain_IO_L1_out_wrapper_200__ap_ready),
    .C_drain_IO_L1_out_wrapper_200__ap_done(C_drain_IO_L1_out_wrapper_200__ap_done),
    .C_drain_IO_L1_out_wrapper_200__ap_idle(C_drain_IO_L1_out_wrapper_200__ap_idle),
    .C_drain_IO_L1_out_wrapper_201__ap_start(C_drain_IO_L1_out_wrapper_201__ap_start),
    .C_drain_IO_L1_out_wrapper_201__ap_ready(C_drain_IO_L1_out_wrapper_201__ap_ready),
    .C_drain_IO_L1_out_wrapper_201__ap_done(C_drain_IO_L1_out_wrapper_201__ap_done),
    .C_drain_IO_L1_out_wrapper_201__ap_idle(C_drain_IO_L1_out_wrapper_201__ap_idle),
    .C_drain_IO_L1_out_wrapper_202__ap_start(C_drain_IO_L1_out_wrapper_202__ap_start),
    .C_drain_IO_L1_out_wrapper_202__ap_ready(C_drain_IO_L1_out_wrapper_202__ap_ready),
    .C_drain_IO_L1_out_wrapper_202__ap_done(C_drain_IO_L1_out_wrapper_202__ap_done),
    .C_drain_IO_L1_out_wrapper_202__ap_idle(C_drain_IO_L1_out_wrapper_202__ap_idle),
    .C_drain_IO_L1_out_wrapper_203__ap_start(C_drain_IO_L1_out_wrapper_203__ap_start),
    .C_drain_IO_L1_out_wrapper_203__ap_ready(C_drain_IO_L1_out_wrapper_203__ap_ready),
    .C_drain_IO_L1_out_wrapper_203__ap_done(C_drain_IO_L1_out_wrapper_203__ap_done),
    .C_drain_IO_L1_out_wrapper_203__ap_idle(C_drain_IO_L1_out_wrapper_203__ap_idle),
    .C_drain_IO_L1_out_wrapper_204__ap_start(C_drain_IO_L1_out_wrapper_204__ap_start),
    .C_drain_IO_L1_out_wrapper_204__ap_ready(C_drain_IO_L1_out_wrapper_204__ap_ready),
    .C_drain_IO_L1_out_wrapper_204__ap_done(C_drain_IO_L1_out_wrapper_204__ap_done),
    .C_drain_IO_L1_out_wrapper_204__ap_idle(C_drain_IO_L1_out_wrapper_204__ap_idle),
    .C_drain_IO_L1_out_wrapper_205__ap_start(C_drain_IO_L1_out_wrapper_205__ap_start),
    .C_drain_IO_L1_out_wrapper_205__ap_ready(C_drain_IO_L1_out_wrapper_205__ap_ready),
    .C_drain_IO_L1_out_wrapper_205__ap_done(C_drain_IO_L1_out_wrapper_205__ap_done),
    .C_drain_IO_L1_out_wrapper_205__ap_idle(C_drain_IO_L1_out_wrapper_205__ap_idle),
    .C_drain_IO_L1_out_wrapper_206__ap_start(C_drain_IO_L1_out_wrapper_206__ap_start),
    .C_drain_IO_L1_out_wrapper_206__ap_ready(C_drain_IO_L1_out_wrapper_206__ap_ready),
    .C_drain_IO_L1_out_wrapper_206__ap_done(C_drain_IO_L1_out_wrapper_206__ap_done),
    .C_drain_IO_L1_out_wrapper_206__ap_idle(C_drain_IO_L1_out_wrapper_206__ap_idle),
    .C_drain_IO_L1_out_wrapper_207__ap_start(C_drain_IO_L1_out_wrapper_207__ap_start),
    .C_drain_IO_L1_out_wrapper_207__ap_ready(C_drain_IO_L1_out_wrapper_207__ap_ready),
    .C_drain_IO_L1_out_wrapper_207__ap_done(C_drain_IO_L1_out_wrapper_207__ap_done),
    .C_drain_IO_L1_out_wrapper_207__ap_idle(C_drain_IO_L1_out_wrapper_207__ap_idle),
    .C_drain_IO_L1_out_wrapper_208__ap_start(C_drain_IO_L1_out_wrapper_208__ap_start),
    .C_drain_IO_L1_out_wrapper_208__ap_ready(C_drain_IO_L1_out_wrapper_208__ap_ready),
    .C_drain_IO_L1_out_wrapper_208__ap_done(C_drain_IO_L1_out_wrapper_208__ap_done),
    .C_drain_IO_L1_out_wrapper_208__ap_idle(C_drain_IO_L1_out_wrapper_208__ap_idle),
    .C_drain_IO_L1_out_wrapper_209__ap_start(C_drain_IO_L1_out_wrapper_209__ap_start),
    .C_drain_IO_L1_out_wrapper_209__ap_ready(C_drain_IO_L1_out_wrapper_209__ap_ready),
    .C_drain_IO_L1_out_wrapper_209__ap_done(C_drain_IO_L1_out_wrapper_209__ap_done),
    .C_drain_IO_L1_out_wrapper_209__ap_idle(C_drain_IO_L1_out_wrapper_209__ap_idle),
    .C_drain_IO_L1_out_wrapper_210__ap_start(C_drain_IO_L1_out_wrapper_210__ap_start),
    .C_drain_IO_L1_out_wrapper_210__ap_ready(C_drain_IO_L1_out_wrapper_210__ap_ready),
    .C_drain_IO_L1_out_wrapper_210__ap_done(C_drain_IO_L1_out_wrapper_210__ap_done),
    .C_drain_IO_L1_out_wrapper_210__ap_idle(C_drain_IO_L1_out_wrapper_210__ap_idle),
    .C_drain_IO_L1_out_wrapper_211__ap_start(C_drain_IO_L1_out_wrapper_211__ap_start),
    .C_drain_IO_L1_out_wrapper_211__ap_ready(C_drain_IO_L1_out_wrapper_211__ap_ready),
    .C_drain_IO_L1_out_wrapper_211__ap_done(C_drain_IO_L1_out_wrapper_211__ap_done),
    .C_drain_IO_L1_out_wrapper_211__ap_idle(C_drain_IO_L1_out_wrapper_211__ap_idle),
    .C_drain_IO_L1_out_wrapper_212__ap_start(C_drain_IO_L1_out_wrapper_212__ap_start),
    .C_drain_IO_L1_out_wrapper_212__ap_ready(C_drain_IO_L1_out_wrapper_212__ap_ready),
    .C_drain_IO_L1_out_wrapper_212__ap_done(C_drain_IO_L1_out_wrapper_212__ap_done),
    .C_drain_IO_L1_out_wrapper_212__ap_idle(C_drain_IO_L1_out_wrapper_212__ap_idle),
    .C_drain_IO_L1_out_wrapper_213__ap_start(C_drain_IO_L1_out_wrapper_213__ap_start),
    .C_drain_IO_L1_out_wrapper_213__ap_ready(C_drain_IO_L1_out_wrapper_213__ap_ready),
    .C_drain_IO_L1_out_wrapper_213__ap_done(C_drain_IO_L1_out_wrapper_213__ap_done),
    .C_drain_IO_L1_out_wrapper_213__ap_idle(C_drain_IO_L1_out_wrapper_213__ap_idle),
    .C_drain_IO_L1_out_wrapper_214__ap_start(C_drain_IO_L1_out_wrapper_214__ap_start),
    .C_drain_IO_L1_out_wrapper_214__ap_ready(C_drain_IO_L1_out_wrapper_214__ap_ready),
    .C_drain_IO_L1_out_wrapper_214__ap_done(C_drain_IO_L1_out_wrapper_214__ap_done),
    .C_drain_IO_L1_out_wrapper_214__ap_idle(C_drain_IO_L1_out_wrapper_214__ap_idle),
    .C_drain_IO_L1_out_wrapper_215__ap_start(C_drain_IO_L1_out_wrapper_215__ap_start),
    .C_drain_IO_L1_out_wrapper_215__ap_ready(C_drain_IO_L1_out_wrapper_215__ap_ready),
    .C_drain_IO_L1_out_wrapper_215__ap_done(C_drain_IO_L1_out_wrapper_215__ap_done),
    .C_drain_IO_L1_out_wrapper_215__ap_idle(C_drain_IO_L1_out_wrapper_215__ap_idle),
    .C_drain_IO_L1_out_wrapper_216__ap_start(C_drain_IO_L1_out_wrapper_216__ap_start),
    .C_drain_IO_L1_out_wrapper_216__ap_ready(C_drain_IO_L1_out_wrapper_216__ap_ready),
    .C_drain_IO_L1_out_wrapper_216__ap_done(C_drain_IO_L1_out_wrapper_216__ap_done),
    .C_drain_IO_L1_out_wrapper_216__ap_idle(C_drain_IO_L1_out_wrapper_216__ap_idle),
    .C_drain_IO_L1_out_wrapper_217__ap_start(C_drain_IO_L1_out_wrapper_217__ap_start),
    .C_drain_IO_L1_out_wrapper_217__ap_ready(C_drain_IO_L1_out_wrapper_217__ap_ready),
    .C_drain_IO_L1_out_wrapper_217__ap_done(C_drain_IO_L1_out_wrapper_217__ap_done),
    .C_drain_IO_L1_out_wrapper_217__ap_idle(C_drain_IO_L1_out_wrapper_217__ap_idle),
    .C_drain_IO_L1_out_wrapper_218__ap_start(C_drain_IO_L1_out_wrapper_218__ap_start),
    .C_drain_IO_L1_out_wrapper_218__ap_ready(C_drain_IO_L1_out_wrapper_218__ap_ready),
    .C_drain_IO_L1_out_wrapper_218__ap_done(C_drain_IO_L1_out_wrapper_218__ap_done),
    .C_drain_IO_L1_out_wrapper_218__ap_idle(C_drain_IO_L1_out_wrapper_218__ap_idle),
    .C_drain_IO_L1_out_wrapper_219__ap_start(C_drain_IO_L1_out_wrapper_219__ap_start),
    .C_drain_IO_L1_out_wrapper_219__ap_ready(C_drain_IO_L1_out_wrapper_219__ap_ready),
    .C_drain_IO_L1_out_wrapper_219__ap_done(C_drain_IO_L1_out_wrapper_219__ap_done),
    .C_drain_IO_L1_out_wrapper_219__ap_idle(C_drain_IO_L1_out_wrapper_219__ap_idle),
    .C_drain_IO_L1_out_wrapper_220__ap_start(C_drain_IO_L1_out_wrapper_220__ap_start),
    .C_drain_IO_L1_out_wrapper_220__ap_ready(C_drain_IO_L1_out_wrapper_220__ap_ready),
    .C_drain_IO_L1_out_wrapper_220__ap_done(C_drain_IO_L1_out_wrapper_220__ap_done),
    .C_drain_IO_L1_out_wrapper_220__ap_idle(C_drain_IO_L1_out_wrapper_220__ap_idle),
    .C_drain_IO_L1_out_wrapper_221__ap_start(C_drain_IO_L1_out_wrapper_221__ap_start),
    .C_drain_IO_L1_out_wrapper_221__ap_ready(C_drain_IO_L1_out_wrapper_221__ap_ready),
    .C_drain_IO_L1_out_wrapper_221__ap_done(C_drain_IO_L1_out_wrapper_221__ap_done),
    .C_drain_IO_L1_out_wrapper_221__ap_idle(C_drain_IO_L1_out_wrapper_221__ap_idle),
    .C_drain_IO_L1_out_wrapper_222__ap_start(C_drain_IO_L1_out_wrapper_222__ap_start),
    .C_drain_IO_L1_out_wrapper_222__ap_ready(C_drain_IO_L1_out_wrapper_222__ap_ready),
    .C_drain_IO_L1_out_wrapper_222__ap_done(C_drain_IO_L1_out_wrapper_222__ap_done),
    .C_drain_IO_L1_out_wrapper_222__ap_idle(C_drain_IO_L1_out_wrapper_222__ap_idle),
    .C_drain_IO_L1_out_wrapper_223__ap_start(C_drain_IO_L1_out_wrapper_223__ap_start),
    .C_drain_IO_L1_out_wrapper_223__ap_ready(C_drain_IO_L1_out_wrapper_223__ap_ready),
    .C_drain_IO_L1_out_wrapper_223__ap_done(C_drain_IO_L1_out_wrapper_223__ap_done),
    .C_drain_IO_L1_out_wrapper_223__ap_idle(C_drain_IO_L1_out_wrapper_223__ap_idle),
    .C_drain_IO_L1_out_wrapper_224__ap_start(C_drain_IO_L1_out_wrapper_224__ap_start),
    .C_drain_IO_L1_out_wrapper_224__ap_ready(C_drain_IO_L1_out_wrapper_224__ap_ready),
    .C_drain_IO_L1_out_wrapper_224__ap_done(C_drain_IO_L1_out_wrapper_224__ap_done),
    .C_drain_IO_L1_out_wrapper_224__ap_idle(C_drain_IO_L1_out_wrapper_224__ap_idle),
    .C_drain_IO_L1_out_wrapper_225__ap_start(C_drain_IO_L1_out_wrapper_225__ap_start),
    .C_drain_IO_L1_out_wrapper_225__ap_ready(C_drain_IO_L1_out_wrapper_225__ap_ready),
    .C_drain_IO_L1_out_wrapper_225__ap_done(C_drain_IO_L1_out_wrapper_225__ap_done),
    .C_drain_IO_L1_out_wrapper_225__ap_idle(C_drain_IO_L1_out_wrapper_225__ap_idle),
    .C_drain_IO_L1_out_wrapper_226__ap_start(C_drain_IO_L1_out_wrapper_226__ap_start),
    .C_drain_IO_L1_out_wrapper_226__ap_ready(C_drain_IO_L1_out_wrapper_226__ap_ready),
    .C_drain_IO_L1_out_wrapper_226__ap_done(C_drain_IO_L1_out_wrapper_226__ap_done),
    .C_drain_IO_L1_out_wrapper_226__ap_idle(C_drain_IO_L1_out_wrapper_226__ap_idle),
    .C_drain_IO_L1_out_wrapper_227__ap_start(C_drain_IO_L1_out_wrapper_227__ap_start),
    .C_drain_IO_L1_out_wrapper_227__ap_ready(C_drain_IO_L1_out_wrapper_227__ap_ready),
    .C_drain_IO_L1_out_wrapper_227__ap_done(C_drain_IO_L1_out_wrapper_227__ap_done),
    .C_drain_IO_L1_out_wrapper_227__ap_idle(C_drain_IO_L1_out_wrapper_227__ap_idle),
    .C_drain_IO_L1_out_wrapper_228__ap_start(C_drain_IO_L1_out_wrapper_228__ap_start),
    .C_drain_IO_L1_out_wrapper_228__ap_ready(C_drain_IO_L1_out_wrapper_228__ap_ready),
    .C_drain_IO_L1_out_wrapper_228__ap_done(C_drain_IO_L1_out_wrapper_228__ap_done),
    .C_drain_IO_L1_out_wrapper_228__ap_idle(C_drain_IO_L1_out_wrapper_228__ap_idle),
    .C_drain_IO_L1_out_wrapper_229__ap_start(C_drain_IO_L1_out_wrapper_229__ap_start),
    .C_drain_IO_L1_out_wrapper_229__ap_ready(C_drain_IO_L1_out_wrapper_229__ap_ready),
    .C_drain_IO_L1_out_wrapper_229__ap_done(C_drain_IO_L1_out_wrapper_229__ap_done),
    .C_drain_IO_L1_out_wrapper_229__ap_idle(C_drain_IO_L1_out_wrapper_229__ap_idle),
    .C_drain_IO_L1_out_wrapper_230__ap_start(C_drain_IO_L1_out_wrapper_230__ap_start),
    .C_drain_IO_L1_out_wrapper_230__ap_ready(C_drain_IO_L1_out_wrapper_230__ap_ready),
    .C_drain_IO_L1_out_wrapper_230__ap_done(C_drain_IO_L1_out_wrapper_230__ap_done),
    .C_drain_IO_L1_out_wrapper_230__ap_idle(C_drain_IO_L1_out_wrapper_230__ap_idle),
    .C_drain_IO_L1_out_wrapper_231__ap_start(C_drain_IO_L1_out_wrapper_231__ap_start),
    .C_drain_IO_L1_out_wrapper_231__ap_ready(C_drain_IO_L1_out_wrapper_231__ap_ready),
    .C_drain_IO_L1_out_wrapper_231__ap_done(C_drain_IO_L1_out_wrapper_231__ap_done),
    .C_drain_IO_L1_out_wrapper_231__ap_idle(C_drain_IO_L1_out_wrapper_231__ap_idle),
    .C_drain_IO_L1_out_wrapper_232__ap_start(C_drain_IO_L1_out_wrapper_232__ap_start),
    .C_drain_IO_L1_out_wrapper_232__ap_ready(C_drain_IO_L1_out_wrapper_232__ap_ready),
    .C_drain_IO_L1_out_wrapper_232__ap_done(C_drain_IO_L1_out_wrapper_232__ap_done),
    .C_drain_IO_L1_out_wrapper_232__ap_idle(C_drain_IO_L1_out_wrapper_232__ap_idle),
    .C_drain_IO_L1_out_wrapper_233__ap_start(C_drain_IO_L1_out_wrapper_233__ap_start),
    .C_drain_IO_L1_out_wrapper_233__ap_ready(C_drain_IO_L1_out_wrapper_233__ap_ready),
    .C_drain_IO_L1_out_wrapper_233__ap_done(C_drain_IO_L1_out_wrapper_233__ap_done),
    .C_drain_IO_L1_out_wrapper_233__ap_idle(C_drain_IO_L1_out_wrapper_233__ap_idle),
    .C_drain_IO_L1_out_wrapper_234__ap_start(C_drain_IO_L1_out_wrapper_234__ap_start),
    .C_drain_IO_L1_out_wrapper_234__ap_ready(C_drain_IO_L1_out_wrapper_234__ap_ready),
    .C_drain_IO_L1_out_wrapper_234__ap_done(C_drain_IO_L1_out_wrapper_234__ap_done),
    .C_drain_IO_L1_out_wrapper_234__ap_idle(C_drain_IO_L1_out_wrapper_234__ap_idle),
    .C_drain_IO_L1_out_wrapper_235__ap_start(C_drain_IO_L1_out_wrapper_235__ap_start),
    .C_drain_IO_L1_out_wrapper_235__ap_ready(C_drain_IO_L1_out_wrapper_235__ap_ready),
    .C_drain_IO_L1_out_wrapper_235__ap_done(C_drain_IO_L1_out_wrapper_235__ap_done),
    .C_drain_IO_L1_out_wrapper_235__ap_idle(C_drain_IO_L1_out_wrapper_235__ap_idle),
    .C_drain_IO_L1_out_wrapper_236__ap_start(C_drain_IO_L1_out_wrapper_236__ap_start),
    .C_drain_IO_L1_out_wrapper_236__ap_ready(C_drain_IO_L1_out_wrapper_236__ap_ready),
    .C_drain_IO_L1_out_wrapper_236__ap_done(C_drain_IO_L1_out_wrapper_236__ap_done),
    .C_drain_IO_L1_out_wrapper_236__ap_idle(C_drain_IO_L1_out_wrapper_236__ap_idle),
    .C_drain_IO_L1_out_wrapper_237__ap_start(C_drain_IO_L1_out_wrapper_237__ap_start),
    .C_drain_IO_L1_out_wrapper_237__ap_ready(C_drain_IO_L1_out_wrapper_237__ap_ready),
    .C_drain_IO_L1_out_wrapper_237__ap_done(C_drain_IO_L1_out_wrapper_237__ap_done),
    .C_drain_IO_L1_out_wrapper_237__ap_idle(C_drain_IO_L1_out_wrapper_237__ap_idle),
    .C_drain_IO_L1_out_wrapper_238__ap_start(C_drain_IO_L1_out_wrapper_238__ap_start),
    .C_drain_IO_L1_out_wrapper_238__ap_ready(C_drain_IO_L1_out_wrapper_238__ap_ready),
    .C_drain_IO_L1_out_wrapper_238__ap_done(C_drain_IO_L1_out_wrapper_238__ap_done),
    .C_drain_IO_L1_out_wrapper_238__ap_idle(C_drain_IO_L1_out_wrapper_238__ap_idle),
    .C_drain_IO_L1_out_wrapper_239__ap_start(C_drain_IO_L1_out_wrapper_239__ap_start),
    .C_drain_IO_L1_out_wrapper_239__ap_ready(C_drain_IO_L1_out_wrapper_239__ap_ready),
    .C_drain_IO_L1_out_wrapper_239__ap_done(C_drain_IO_L1_out_wrapper_239__ap_done),
    .C_drain_IO_L1_out_wrapper_239__ap_idle(C_drain_IO_L1_out_wrapper_239__ap_idle),
    .C_drain_IO_L1_out_wrapper_240__ap_start(C_drain_IO_L1_out_wrapper_240__ap_start),
    .C_drain_IO_L1_out_wrapper_240__ap_ready(C_drain_IO_L1_out_wrapper_240__ap_ready),
    .C_drain_IO_L1_out_wrapper_240__ap_done(C_drain_IO_L1_out_wrapper_240__ap_done),
    .C_drain_IO_L1_out_wrapper_240__ap_idle(C_drain_IO_L1_out_wrapper_240__ap_idle),
    .C_drain_IO_L1_out_wrapper_241__ap_start(C_drain_IO_L1_out_wrapper_241__ap_start),
    .C_drain_IO_L1_out_wrapper_241__ap_ready(C_drain_IO_L1_out_wrapper_241__ap_ready),
    .C_drain_IO_L1_out_wrapper_241__ap_done(C_drain_IO_L1_out_wrapper_241__ap_done),
    .C_drain_IO_L1_out_wrapper_241__ap_idle(C_drain_IO_L1_out_wrapper_241__ap_idle),
    .C_drain_IO_L1_out_wrapper_242__ap_start(C_drain_IO_L1_out_wrapper_242__ap_start),
    .C_drain_IO_L1_out_wrapper_242__ap_ready(C_drain_IO_L1_out_wrapper_242__ap_ready),
    .C_drain_IO_L1_out_wrapper_242__ap_done(C_drain_IO_L1_out_wrapper_242__ap_done),
    .C_drain_IO_L1_out_wrapper_242__ap_idle(C_drain_IO_L1_out_wrapper_242__ap_idle),
    .C_drain_IO_L1_out_wrapper_243__ap_start(C_drain_IO_L1_out_wrapper_243__ap_start),
    .C_drain_IO_L1_out_wrapper_243__ap_ready(C_drain_IO_L1_out_wrapper_243__ap_ready),
    .C_drain_IO_L1_out_wrapper_243__ap_done(C_drain_IO_L1_out_wrapper_243__ap_done),
    .C_drain_IO_L1_out_wrapper_243__ap_idle(C_drain_IO_L1_out_wrapper_243__ap_idle),
    .C_drain_IO_L1_out_wrapper_244__ap_start(C_drain_IO_L1_out_wrapper_244__ap_start),
    .C_drain_IO_L1_out_wrapper_244__ap_ready(C_drain_IO_L1_out_wrapper_244__ap_ready),
    .C_drain_IO_L1_out_wrapper_244__ap_done(C_drain_IO_L1_out_wrapper_244__ap_done),
    .C_drain_IO_L1_out_wrapper_244__ap_idle(C_drain_IO_L1_out_wrapper_244__ap_idle),
    .C_drain_IO_L1_out_wrapper_245__ap_start(C_drain_IO_L1_out_wrapper_245__ap_start),
    .C_drain_IO_L1_out_wrapper_245__ap_ready(C_drain_IO_L1_out_wrapper_245__ap_ready),
    .C_drain_IO_L1_out_wrapper_245__ap_done(C_drain_IO_L1_out_wrapper_245__ap_done),
    .C_drain_IO_L1_out_wrapper_245__ap_idle(C_drain_IO_L1_out_wrapper_245__ap_idle),
    .C_drain_IO_L1_out_wrapper_246__ap_start(C_drain_IO_L1_out_wrapper_246__ap_start),
    .C_drain_IO_L1_out_wrapper_246__ap_ready(C_drain_IO_L1_out_wrapper_246__ap_ready),
    .C_drain_IO_L1_out_wrapper_246__ap_done(C_drain_IO_L1_out_wrapper_246__ap_done),
    .C_drain_IO_L1_out_wrapper_246__ap_idle(C_drain_IO_L1_out_wrapper_246__ap_idle),
    .C_drain_IO_L1_out_wrapper_247__ap_start(C_drain_IO_L1_out_wrapper_247__ap_start),
    .C_drain_IO_L1_out_wrapper_247__ap_ready(C_drain_IO_L1_out_wrapper_247__ap_ready),
    .C_drain_IO_L1_out_wrapper_247__ap_done(C_drain_IO_L1_out_wrapper_247__ap_done),
    .C_drain_IO_L1_out_wrapper_247__ap_idle(C_drain_IO_L1_out_wrapper_247__ap_idle),
    .C_drain_IO_L1_out_wrapper_248__ap_start(C_drain_IO_L1_out_wrapper_248__ap_start),
    .C_drain_IO_L1_out_wrapper_248__ap_ready(C_drain_IO_L1_out_wrapper_248__ap_ready),
    .C_drain_IO_L1_out_wrapper_248__ap_done(C_drain_IO_L1_out_wrapper_248__ap_done),
    .C_drain_IO_L1_out_wrapper_248__ap_idle(C_drain_IO_L1_out_wrapper_248__ap_idle),
    .C_drain_IO_L1_out_wrapper_249__ap_start(C_drain_IO_L1_out_wrapper_249__ap_start),
    .C_drain_IO_L1_out_wrapper_249__ap_ready(C_drain_IO_L1_out_wrapper_249__ap_ready),
    .C_drain_IO_L1_out_wrapper_249__ap_done(C_drain_IO_L1_out_wrapper_249__ap_done),
    .C_drain_IO_L1_out_wrapper_249__ap_idle(C_drain_IO_L1_out_wrapper_249__ap_idle),
    .C_drain_IO_L1_out_wrapper_250__ap_start(C_drain_IO_L1_out_wrapper_250__ap_start),
    .C_drain_IO_L1_out_wrapper_250__ap_ready(C_drain_IO_L1_out_wrapper_250__ap_ready),
    .C_drain_IO_L1_out_wrapper_250__ap_done(C_drain_IO_L1_out_wrapper_250__ap_done),
    .C_drain_IO_L1_out_wrapper_250__ap_idle(C_drain_IO_L1_out_wrapper_250__ap_idle),
    .C_drain_IO_L1_out_wrapper_251__ap_start(C_drain_IO_L1_out_wrapper_251__ap_start),
    .C_drain_IO_L1_out_wrapper_251__ap_ready(C_drain_IO_L1_out_wrapper_251__ap_ready),
    .C_drain_IO_L1_out_wrapper_251__ap_done(C_drain_IO_L1_out_wrapper_251__ap_done),
    .C_drain_IO_L1_out_wrapper_251__ap_idle(C_drain_IO_L1_out_wrapper_251__ap_idle),
    .C_drain_IO_L1_out_wrapper_252__ap_start(C_drain_IO_L1_out_wrapper_252__ap_start),
    .C_drain_IO_L1_out_wrapper_252__ap_ready(C_drain_IO_L1_out_wrapper_252__ap_ready),
    .C_drain_IO_L1_out_wrapper_252__ap_done(C_drain_IO_L1_out_wrapper_252__ap_done),
    .C_drain_IO_L1_out_wrapper_252__ap_idle(C_drain_IO_L1_out_wrapper_252__ap_idle),
    .C_drain_IO_L1_out_wrapper_253__ap_start(C_drain_IO_L1_out_wrapper_253__ap_start),
    .C_drain_IO_L1_out_wrapper_253__ap_ready(C_drain_IO_L1_out_wrapper_253__ap_ready),
    .C_drain_IO_L1_out_wrapper_253__ap_done(C_drain_IO_L1_out_wrapper_253__ap_done),
    .C_drain_IO_L1_out_wrapper_253__ap_idle(C_drain_IO_L1_out_wrapper_253__ap_idle),
    .C_drain_IO_L1_out_wrapper_254__ap_start(C_drain_IO_L1_out_wrapper_254__ap_start),
    .C_drain_IO_L1_out_wrapper_254__ap_ready(C_drain_IO_L1_out_wrapper_254__ap_ready),
    .C_drain_IO_L1_out_wrapper_254__ap_done(C_drain_IO_L1_out_wrapper_254__ap_done),
    .C_drain_IO_L1_out_wrapper_254__ap_idle(C_drain_IO_L1_out_wrapper_254__ap_idle),
    .C_drain_IO_L1_out_wrapper_255__ap_start(C_drain_IO_L1_out_wrapper_255__ap_start),
    .C_drain_IO_L1_out_wrapper_255__ap_ready(C_drain_IO_L1_out_wrapper_255__ap_ready),
    .C_drain_IO_L1_out_wrapper_255__ap_done(C_drain_IO_L1_out_wrapper_255__ap_done),
    .C_drain_IO_L1_out_wrapper_255__ap_idle(C_drain_IO_L1_out_wrapper_255__ap_idle),
    .C_drain_IO_L1_out_wrapper_256__ap_start(C_drain_IO_L1_out_wrapper_256__ap_start),
    .C_drain_IO_L1_out_wrapper_256__ap_ready(C_drain_IO_L1_out_wrapper_256__ap_ready),
    .C_drain_IO_L1_out_wrapper_256__ap_done(C_drain_IO_L1_out_wrapper_256__ap_done),
    .C_drain_IO_L1_out_wrapper_256__ap_idle(C_drain_IO_L1_out_wrapper_256__ap_idle),
    .C_drain_IO_L1_out_wrapper_257__ap_start(C_drain_IO_L1_out_wrapper_257__ap_start),
    .C_drain_IO_L1_out_wrapper_257__ap_ready(C_drain_IO_L1_out_wrapper_257__ap_ready),
    .C_drain_IO_L1_out_wrapper_257__ap_done(C_drain_IO_L1_out_wrapper_257__ap_done),
    .C_drain_IO_L1_out_wrapper_257__ap_idle(C_drain_IO_L1_out_wrapper_257__ap_idle),
    .C_drain_IO_L1_out_wrapper_258__ap_start(C_drain_IO_L1_out_wrapper_258__ap_start),
    .C_drain_IO_L1_out_wrapper_258__ap_ready(C_drain_IO_L1_out_wrapper_258__ap_ready),
    .C_drain_IO_L1_out_wrapper_258__ap_done(C_drain_IO_L1_out_wrapper_258__ap_done),
    .C_drain_IO_L1_out_wrapper_258__ap_idle(C_drain_IO_L1_out_wrapper_258__ap_idle),
    .C_drain_IO_L1_out_wrapper_259__ap_start(C_drain_IO_L1_out_wrapper_259__ap_start),
    .C_drain_IO_L1_out_wrapper_259__ap_ready(C_drain_IO_L1_out_wrapper_259__ap_ready),
    .C_drain_IO_L1_out_wrapper_259__ap_done(C_drain_IO_L1_out_wrapper_259__ap_done),
    .C_drain_IO_L1_out_wrapper_259__ap_idle(C_drain_IO_L1_out_wrapper_259__ap_idle),
    .C_drain_IO_L1_out_wrapper_260__ap_start(C_drain_IO_L1_out_wrapper_260__ap_start),
    .C_drain_IO_L1_out_wrapper_260__ap_ready(C_drain_IO_L1_out_wrapper_260__ap_ready),
    .C_drain_IO_L1_out_wrapper_260__ap_done(C_drain_IO_L1_out_wrapper_260__ap_done),
    .C_drain_IO_L1_out_wrapper_260__ap_idle(C_drain_IO_L1_out_wrapper_260__ap_idle),
    .C_drain_IO_L1_out_wrapper_261__ap_start(C_drain_IO_L1_out_wrapper_261__ap_start),
    .C_drain_IO_L1_out_wrapper_261__ap_ready(C_drain_IO_L1_out_wrapper_261__ap_ready),
    .C_drain_IO_L1_out_wrapper_261__ap_done(C_drain_IO_L1_out_wrapper_261__ap_done),
    .C_drain_IO_L1_out_wrapper_261__ap_idle(C_drain_IO_L1_out_wrapper_261__ap_idle),
    .C_drain_IO_L1_out_wrapper_262__ap_start(C_drain_IO_L1_out_wrapper_262__ap_start),
    .C_drain_IO_L1_out_wrapper_262__ap_ready(C_drain_IO_L1_out_wrapper_262__ap_ready),
    .C_drain_IO_L1_out_wrapper_262__ap_done(C_drain_IO_L1_out_wrapper_262__ap_done),
    .C_drain_IO_L1_out_wrapper_262__ap_idle(C_drain_IO_L1_out_wrapper_262__ap_idle),
    .C_drain_IO_L1_out_wrapper_263__ap_start(C_drain_IO_L1_out_wrapper_263__ap_start),
    .C_drain_IO_L1_out_wrapper_263__ap_ready(C_drain_IO_L1_out_wrapper_263__ap_ready),
    .C_drain_IO_L1_out_wrapper_263__ap_done(C_drain_IO_L1_out_wrapper_263__ap_done),
    .C_drain_IO_L1_out_wrapper_263__ap_idle(C_drain_IO_L1_out_wrapper_263__ap_idle),
    .C_drain_IO_L1_out_wrapper_264__ap_start(C_drain_IO_L1_out_wrapper_264__ap_start),
    .C_drain_IO_L1_out_wrapper_264__ap_ready(C_drain_IO_L1_out_wrapper_264__ap_ready),
    .C_drain_IO_L1_out_wrapper_264__ap_done(C_drain_IO_L1_out_wrapper_264__ap_done),
    .C_drain_IO_L1_out_wrapper_264__ap_idle(C_drain_IO_L1_out_wrapper_264__ap_idle),
    .C_drain_IO_L1_out_wrapper_265__ap_start(C_drain_IO_L1_out_wrapper_265__ap_start),
    .C_drain_IO_L1_out_wrapper_265__ap_ready(C_drain_IO_L1_out_wrapper_265__ap_ready),
    .C_drain_IO_L1_out_wrapper_265__ap_done(C_drain_IO_L1_out_wrapper_265__ap_done),
    .C_drain_IO_L1_out_wrapper_265__ap_idle(C_drain_IO_L1_out_wrapper_265__ap_idle),
    .C_drain_IO_L1_out_wrapper_266__ap_start(C_drain_IO_L1_out_wrapper_266__ap_start),
    .C_drain_IO_L1_out_wrapper_266__ap_ready(C_drain_IO_L1_out_wrapper_266__ap_ready),
    .C_drain_IO_L1_out_wrapper_266__ap_done(C_drain_IO_L1_out_wrapper_266__ap_done),
    .C_drain_IO_L1_out_wrapper_266__ap_idle(C_drain_IO_L1_out_wrapper_266__ap_idle),
    .C_drain_IO_L1_out_wrapper_267__ap_start(C_drain_IO_L1_out_wrapper_267__ap_start),
    .C_drain_IO_L1_out_wrapper_267__ap_ready(C_drain_IO_L1_out_wrapper_267__ap_ready),
    .C_drain_IO_L1_out_wrapper_267__ap_done(C_drain_IO_L1_out_wrapper_267__ap_done),
    .C_drain_IO_L1_out_wrapper_267__ap_idle(C_drain_IO_L1_out_wrapper_267__ap_idle),
    .C_drain_IO_L1_out_wrapper_268__ap_start(C_drain_IO_L1_out_wrapper_268__ap_start),
    .C_drain_IO_L1_out_wrapper_268__ap_ready(C_drain_IO_L1_out_wrapper_268__ap_ready),
    .C_drain_IO_L1_out_wrapper_268__ap_done(C_drain_IO_L1_out_wrapper_268__ap_done),
    .C_drain_IO_L1_out_wrapper_268__ap_idle(C_drain_IO_L1_out_wrapper_268__ap_idle),
    .C_drain_IO_L1_out_wrapper_269__ap_start(C_drain_IO_L1_out_wrapper_269__ap_start),
    .C_drain_IO_L1_out_wrapper_269__ap_ready(C_drain_IO_L1_out_wrapper_269__ap_ready),
    .C_drain_IO_L1_out_wrapper_269__ap_done(C_drain_IO_L1_out_wrapper_269__ap_done),
    .C_drain_IO_L1_out_wrapper_269__ap_idle(C_drain_IO_L1_out_wrapper_269__ap_idle),
    .C_drain_IO_L1_out_wrapper_270__ap_start(C_drain_IO_L1_out_wrapper_270__ap_start),
    .C_drain_IO_L1_out_wrapper_270__ap_ready(C_drain_IO_L1_out_wrapper_270__ap_ready),
    .C_drain_IO_L1_out_wrapper_270__ap_done(C_drain_IO_L1_out_wrapper_270__ap_done),
    .C_drain_IO_L1_out_wrapper_270__ap_idle(C_drain_IO_L1_out_wrapper_270__ap_idle),
    .C_drain_IO_L1_out_wrapper_271__ap_start(C_drain_IO_L1_out_wrapper_271__ap_start),
    .C_drain_IO_L1_out_wrapper_271__ap_ready(C_drain_IO_L1_out_wrapper_271__ap_ready),
    .C_drain_IO_L1_out_wrapper_271__ap_done(C_drain_IO_L1_out_wrapper_271__ap_done),
    .C_drain_IO_L1_out_wrapper_271__ap_idle(C_drain_IO_L1_out_wrapper_271__ap_idle),
    .C_drain_IO_L1_out_wrapper_272__ap_start(C_drain_IO_L1_out_wrapper_272__ap_start),
    .C_drain_IO_L1_out_wrapper_272__ap_ready(C_drain_IO_L1_out_wrapper_272__ap_ready),
    .C_drain_IO_L1_out_wrapper_272__ap_done(C_drain_IO_L1_out_wrapper_272__ap_done),
    .C_drain_IO_L1_out_wrapper_272__ap_idle(C_drain_IO_L1_out_wrapper_272__ap_idle),
    .C_drain_IO_L1_out_wrapper_273__ap_start(C_drain_IO_L1_out_wrapper_273__ap_start),
    .C_drain_IO_L1_out_wrapper_273__ap_ready(C_drain_IO_L1_out_wrapper_273__ap_ready),
    .C_drain_IO_L1_out_wrapper_273__ap_done(C_drain_IO_L1_out_wrapper_273__ap_done),
    .C_drain_IO_L1_out_wrapper_273__ap_idle(C_drain_IO_L1_out_wrapper_273__ap_idle),
    .C_drain_IO_L1_out_wrapper_274__ap_start(C_drain_IO_L1_out_wrapper_274__ap_start),
    .C_drain_IO_L1_out_wrapper_274__ap_ready(C_drain_IO_L1_out_wrapper_274__ap_ready),
    .C_drain_IO_L1_out_wrapper_274__ap_done(C_drain_IO_L1_out_wrapper_274__ap_done),
    .C_drain_IO_L1_out_wrapper_274__ap_idle(C_drain_IO_L1_out_wrapper_274__ap_idle),
    .C_drain_IO_L1_out_wrapper_275__ap_start(C_drain_IO_L1_out_wrapper_275__ap_start),
    .C_drain_IO_L1_out_wrapper_275__ap_ready(C_drain_IO_L1_out_wrapper_275__ap_ready),
    .C_drain_IO_L1_out_wrapper_275__ap_done(C_drain_IO_L1_out_wrapper_275__ap_done),
    .C_drain_IO_L1_out_wrapper_275__ap_idle(C_drain_IO_L1_out_wrapper_275__ap_idle),
    .C_drain_IO_L1_out_wrapper_276__ap_start(C_drain_IO_L1_out_wrapper_276__ap_start),
    .C_drain_IO_L1_out_wrapper_276__ap_ready(C_drain_IO_L1_out_wrapper_276__ap_ready),
    .C_drain_IO_L1_out_wrapper_276__ap_done(C_drain_IO_L1_out_wrapper_276__ap_done),
    .C_drain_IO_L1_out_wrapper_276__ap_idle(C_drain_IO_L1_out_wrapper_276__ap_idle),
    .C_drain_IO_L1_out_wrapper_277__ap_start(C_drain_IO_L1_out_wrapper_277__ap_start),
    .C_drain_IO_L1_out_wrapper_277__ap_ready(C_drain_IO_L1_out_wrapper_277__ap_ready),
    .C_drain_IO_L1_out_wrapper_277__ap_done(C_drain_IO_L1_out_wrapper_277__ap_done),
    .C_drain_IO_L1_out_wrapper_277__ap_idle(C_drain_IO_L1_out_wrapper_277__ap_idle),
    .C_drain_IO_L1_out_wrapper_278__ap_start(C_drain_IO_L1_out_wrapper_278__ap_start),
    .C_drain_IO_L1_out_wrapper_278__ap_ready(C_drain_IO_L1_out_wrapper_278__ap_ready),
    .C_drain_IO_L1_out_wrapper_278__ap_done(C_drain_IO_L1_out_wrapper_278__ap_done),
    .C_drain_IO_L1_out_wrapper_278__ap_idle(C_drain_IO_L1_out_wrapper_278__ap_idle),
    .C_drain_IO_L1_out_wrapper_279__ap_start(C_drain_IO_L1_out_wrapper_279__ap_start),
    .C_drain_IO_L1_out_wrapper_279__ap_ready(C_drain_IO_L1_out_wrapper_279__ap_ready),
    .C_drain_IO_L1_out_wrapper_279__ap_done(C_drain_IO_L1_out_wrapper_279__ap_done),
    .C_drain_IO_L1_out_wrapper_279__ap_idle(C_drain_IO_L1_out_wrapper_279__ap_idle),
    .C_drain_IO_L1_out_wrapper_280__ap_start(C_drain_IO_L1_out_wrapper_280__ap_start),
    .C_drain_IO_L1_out_wrapper_280__ap_ready(C_drain_IO_L1_out_wrapper_280__ap_ready),
    .C_drain_IO_L1_out_wrapper_280__ap_done(C_drain_IO_L1_out_wrapper_280__ap_done),
    .C_drain_IO_L1_out_wrapper_280__ap_idle(C_drain_IO_L1_out_wrapper_280__ap_idle),
    .C_drain_IO_L1_out_wrapper_281__ap_start(C_drain_IO_L1_out_wrapper_281__ap_start),
    .C_drain_IO_L1_out_wrapper_281__ap_ready(C_drain_IO_L1_out_wrapper_281__ap_ready),
    .C_drain_IO_L1_out_wrapper_281__ap_done(C_drain_IO_L1_out_wrapper_281__ap_done),
    .C_drain_IO_L1_out_wrapper_281__ap_idle(C_drain_IO_L1_out_wrapper_281__ap_idle),
    .C_drain_IO_L1_out_wrapper_282__ap_start(C_drain_IO_L1_out_wrapper_282__ap_start),
    .C_drain_IO_L1_out_wrapper_282__ap_ready(C_drain_IO_L1_out_wrapper_282__ap_ready),
    .C_drain_IO_L1_out_wrapper_282__ap_done(C_drain_IO_L1_out_wrapper_282__ap_done),
    .C_drain_IO_L1_out_wrapper_282__ap_idle(C_drain_IO_L1_out_wrapper_282__ap_idle),
    .C_drain_IO_L1_out_wrapper_283__ap_start(C_drain_IO_L1_out_wrapper_283__ap_start),
    .C_drain_IO_L1_out_wrapper_283__ap_ready(C_drain_IO_L1_out_wrapper_283__ap_ready),
    .C_drain_IO_L1_out_wrapper_283__ap_done(C_drain_IO_L1_out_wrapper_283__ap_done),
    .C_drain_IO_L1_out_wrapper_283__ap_idle(C_drain_IO_L1_out_wrapper_283__ap_idle),
    .C_drain_IO_L1_out_wrapper_284__ap_start(C_drain_IO_L1_out_wrapper_284__ap_start),
    .C_drain_IO_L1_out_wrapper_284__ap_ready(C_drain_IO_L1_out_wrapper_284__ap_ready),
    .C_drain_IO_L1_out_wrapper_284__ap_done(C_drain_IO_L1_out_wrapper_284__ap_done),
    .C_drain_IO_L1_out_wrapper_284__ap_idle(C_drain_IO_L1_out_wrapper_284__ap_idle),
    .C_drain_IO_L1_out_wrapper_285__ap_start(C_drain_IO_L1_out_wrapper_285__ap_start),
    .C_drain_IO_L1_out_wrapper_285__ap_ready(C_drain_IO_L1_out_wrapper_285__ap_ready),
    .C_drain_IO_L1_out_wrapper_285__ap_done(C_drain_IO_L1_out_wrapper_285__ap_done),
    .C_drain_IO_L1_out_wrapper_285__ap_idle(C_drain_IO_L1_out_wrapper_285__ap_idle),
    .C_drain_IO_L1_out_wrapper_286__ap_start(C_drain_IO_L1_out_wrapper_286__ap_start),
    .C_drain_IO_L1_out_wrapper_286__ap_ready(C_drain_IO_L1_out_wrapper_286__ap_ready),
    .C_drain_IO_L1_out_wrapper_286__ap_done(C_drain_IO_L1_out_wrapper_286__ap_done),
    .C_drain_IO_L1_out_wrapper_286__ap_idle(C_drain_IO_L1_out_wrapper_286__ap_idle),
    .C_drain_IO_L1_out_wrapper_287__ap_start(C_drain_IO_L1_out_wrapper_287__ap_start),
    .C_drain_IO_L1_out_wrapper_287__ap_ready(C_drain_IO_L1_out_wrapper_287__ap_ready),
    .C_drain_IO_L1_out_wrapper_287__ap_done(C_drain_IO_L1_out_wrapper_287__ap_done),
    .C_drain_IO_L1_out_wrapper_287__ap_idle(C_drain_IO_L1_out_wrapper_287__ap_idle),
    .C_drain_IO_L1_out_wrapper_288__ap_start(C_drain_IO_L1_out_wrapper_288__ap_start),
    .C_drain_IO_L1_out_wrapper_288__ap_ready(C_drain_IO_L1_out_wrapper_288__ap_ready),
    .C_drain_IO_L1_out_wrapper_288__ap_done(C_drain_IO_L1_out_wrapper_288__ap_done),
    .C_drain_IO_L1_out_wrapper_288__ap_idle(C_drain_IO_L1_out_wrapper_288__ap_idle),
    .C_drain_IO_L2_out_0__ap_start(C_drain_IO_L2_out_0__ap_start),
    .C_drain_IO_L2_out_0__ap_ready(C_drain_IO_L2_out_0__ap_ready),
    .C_drain_IO_L2_out_0__ap_done(C_drain_IO_L2_out_0__ap_done),
    .C_drain_IO_L2_out_0__ap_idle(C_drain_IO_L2_out_0__ap_idle),
    .C_drain_IO_L2_out_1__ap_start(C_drain_IO_L2_out_1__ap_start),
    .C_drain_IO_L2_out_1__ap_ready(C_drain_IO_L2_out_1__ap_ready),
    .C_drain_IO_L2_out_1__ap_done(C_drain_IO_L2_out_1__ap_done),
    .C_drain_IO_L2_out_1__ap_idle(C_drain_IO_L2_out_1__ap_idle),
    .C_drain_IO_L2_out_2__ap_start(C_drain_IO_L2_out_2__ap_start),
    .C_drain_IO_L2_out_2__ap_ready(C_drain_IO_L2_out_2__ap_ready),
    .C_drain_IO_L2_out_2__ap_done(C_drain_IO_L2_out_2__ap_done),
    .C_drain_IO_L2_out_2__ap_idle(C_drain_IO_L2_out_2__ap_idle),
    .C_drain_IO_L2_out_3__ap_start(C_drain_IO_L2_out_3__ap_start),
    .C_drain_IO_L2_out_3__ap_ready(C_drain_IO_L2_out_3__ap_ready),
    .C_drain_IO_L2_out_3__ap_done(C_drain_IO_L2_out_3__ap_done),
    .C_drain_IO_L2_out_3__ap_idle(C_drain_IO_L2_out_3__ap_idle),
    .C_drain_IO_L2_out_4__ap_start(C_drain_IO_L2_out_4__ap_start),
    .C_drain_IO_L2_out_4__ap_ready(C_drain_IO_L2_out_4__ap_ready),
    .C_drain_IO_L2_out_4__ap_done(C_drain_IO_L2_out_4__ap_done),
    .C_drain_IO_L2_out_4__ap_idle(C_drain_IO_L2_out_4__ap_idle),
    .C_drain_IO_L2_out_5__ap_start(C_drain_IO_L2_out_5__ap_start),
    .C_drain_IO_L2_out_5__ap_ready(C_drain_IO_L2_out_5__ap_ready),
    .C_drain_IO_L2_out_5__ap_done(C_drain_IO_L2_out_5__ap_done),
    .C_drain_IO_L2_out_5__ap_idle(C_drain_IO_L2_out_5__ap_idle),
    .C_drain_IO_L2_out_6__ap_start(C_drain_IO_L2_out_6__ap_start),
    .C_drain_IO_L2_out_6__ap_ready(C_drain_IO_L2_out_6__ap_ready),
    .C_drain_IO_L2_out_6__ap_done(C_drain_IO_L2_out_6__ap_done),
    .C_drain_IO_L2_out_6__ap_idle(C_drain_IO_L2_out_6__ap_idle),
    .C_drain_IO_L2_out_7__ap_start(C_drain_IO_L2_out_7__ap_start),
    .C_drain_IO_L2_out_7__ap_ready(C_drain_IO_L2_out_7__ap_ready),
    .C_drain_IO_L2_out_7__ap_done(C_drain_IO_L2_out_7__ap_done),
    .C_drain_IO_L2_out_7__ap_idle(C_drain_IO_L2_out_7__ap_idle),
    .C_drain_IO_L2_out_8__ap_start(C_drain_IO_L2_out_8__ap_start),
    .C_drain_IO_L2_out_8__ap_ready(C_drain_IO_L2_out_8__ap_ready),
    .C_drain_IO_L2_out_8__ap_done(C_drain_IO_L2_out_8__ap_done),
    .C_drain_IO_L2_out_8__ap_idle(C_drain_IO_L2_out_8__ap_idle),
    .C_drain_IO_L2_out_9__ap_start(C_drain_IO_L2_out_9__ap_start),
    .C_drain_IO_L2_out_9__ap_ready(C_drain_IO_L2_out_9__ap_ready),
    .C_drain_IO_L2_out_9__ap_done(C_drain_IO_L2_out_9__ap_done),
    .C_drain_IO_L2_out_9__ap_idle(C_drain_IO_L2_out_9__ap_idle),
    .C_drain_IO_L2_out_10__ap_start(C_drain_IO_L2_out_10__ap_start),
    .C_drain_IO_L2_out_10__ap_ready(C_drain_IO_L2_out_10__ap_ready),
    .C_drain_IO_L2_out_10__ap_done(C_drain_IO_L2_out_10__ap_done),
    .C_drain_IO_L2_out_10__ap_idle(C_drain_IO_L2_out_10__ap_idle),
    .C_drain_IO_L2_out_11__ap_start(C_drain_IO_L2_out_11__ap_start),
    .C_drain_IO_L2_out_11__ap_ready(C_drain_IO_L2_out_11__ap_ready),
    .C_drain_IO_L2_out_11__ap_done(C_drain_IO_L2_out_11__ap_done),
    .C_drain_IO_L2_out_11__ap_idle(C_drain_IO_L2_out_11__ap_idle),
    .C_drain_IO_L2_out_12__ap_start(C_drain_IO_L2_out_12__ap_start),
    .C_drain_IO_L2_out_12__ap_ready(C_drain_IO_L2_out_12__ap_ready),
    .C_drain_IO_L2_out_12__ap_done(C_drain_IO_L2_out_12__ap_done),
    .C_drain_IO_L2_out_12__ap_idle(C_drain_IO_L2_out_12__ap_idle),
    .C_drain_IO_L2_out_13__ap_start(C_drain_IO_L2_out_13__ap_start),
    .C_drain_IO_L2_out_13__ap_ready(C_drain_IO_L2_out_13__ap_ready),
    .C_drain_IO_L2_out_13__ap_done(C_drain_IO_L2_out_13__ap_done),
    .C_drain_IO_L2_out_13__ap_idle(C_drain_IO_L2_out_13__ap_idle),
    .C_drain_IO_L2_out_14__ap_start(C_drain_IO_L2_out_14__ap_start),
    .C_drain_IO_L2_out_14__ap_ready(C_drain_IO_L2_out_14__ap_ready),
    .C_drain_IO_L2_out_14__ap_done(C_drain_IO_L2_out_14__ap_done),
    .C_drain_IO_L2_out_14__ap_idle(C_drain_IO_L2_out_14__ap_idle),
    .C_drain_IO_L2_out_15__ap_start(C_drain_IO_L2_out_15__ap_start),
    .C_drain_IO_L2_out_15__ap_ready(C_drain_IO_L2_out_15__ap_ready),
    .C_drain_IO_L2_out_15__ap_done(C_drain_IO_L2_out_15__ap_done),
    .C_drain_IO_L2_out_15__ap_idle(C_drain_IO_L2_out_15__ap_idle),
    .C_drain_IO_L2_out_boundary_0__ap_start(C_drain_IO_L2_out_boundary_0__ap_start),
    .C_drain_IO_L2_out_boundary_0__ap_ready(C_drain_IO_L2_out_boundary_0__ap_ready),
    .C_drain_IO_L2_out_boundary_0__ap_done(C_drain_IO_L2_out_boundary_0__ap_done),
    .C_drain_IO_L2_out_boundary_0__ap_idle(C_drain_IO_L2_out_boundary_0__ap_idle),
    .C_drain_IO_L3_out_0__ap_start(C_drain_IO_L3_out_0__ap_start),
    .C_drain_IO_L3_out_0__ap_ready(C_drain_IO_L3_out_0__ap_ready),
    .C_drain_IO_L3_out_0__ap_done(C_drain_IO_L3_out_0__ap_done),
    .C_drain_IO_L3_out_0__ap_idle(C_drain_IO_L3_out_0__ap_idle),
    .C_drain_IO_L3_out_serialize_0___C__q0(C_drain_IO_L3_out_serialize_0___C__q0),
    .C_drain_IO_L3_out_serialize_0__ap_start(C_drain_IO_L3_out_serialize_0__ap_start),
    .C_drain_IO_L3_out_serialize_0__ap_ready(C_drain_IO_L3_out_serialize_0__ap_ready),
    .C_drain_IO_L3_out_serialize_0__ap_done(C_drain_IO_L3_out_serialize_0__ap_done),
    .C_drain_IO_L3_out_serialize_0__ap_idle(C_drain_IO_L3_out_serialize_0__ap_idle),
    .PE_wrapper_0__ap_start(PE_wrapper_0__ap_start),
    .PE_wrapper_0__ap_ready(PE_wrapper_0__ap_ready),
    .PE_wrapper_0__ap_done(PE_wrapper_0__ap_done),
    .PE_wrapper_0__ap_idle(PE_wrapper_0__ap_idle),
    .PE_wrapper_1__ap_start(PE_wrapper_1__ap_start),
    .PE_wrapper_1__ap_ready(PE_wrapper_1__ap_ready),
    .PE_wrapper_1__ap_done(PE_wrapper_1__ap_done),
    .PE_wrapper_1__ap_idle(PE_wrapper_1__ap_idle),
    .PE_wrapper_2__ap_start(PE_wrapper_2__ap_start),
    .PE_wrapper_2__ap_ready(PE_wrapper_2__ap_ready),
    .PE_wrapper_2__ap_done(PE_wrapper_2__ap_done),
    .PE_wrapper_2__ap_idle(PE_wrapper_2__ap_idle),
    .PE_wrapper_3__ap_start(PE_wrapper_3__ap_start),
    .PE_wrapper_3__ap_ready(PE_wrapper_3__ap_ready),
    .PE_wrapper_3__ap_done(PE_wrapper_3__ap_done),
    .PE_wrapper_3__ap_idle(PE_wrapper_3__ap_idle),
    .PE_wrapper_4__ap_start(PE_wrapper_4__ap_start),
    .PE_wrapper_4__ap_ready(PE_wrapper_4__ap_ready),
    .PE_wrapper_4__ap_done(PE_wrapper_4__ap_done),
    .PE_wrapper_4__ap_idle(PE_wrapper_4__ap_idle),
    .PE_wrapper_5__ap_start(PE_wrapper_5__ap_start),
    .PE_wrapper_5__ap_ready(PE_wrapper_5__ap_ready),
    .PE_wrapper_5__ap_done(PE_wrapper_5__ap_done),
    .PE_wrapper_5__ap_idle(PE_wrapper_5__ap_idle),
    .PE_wrapper_6__ap_start(PE_wrapper_6__ap_start),
    .PE_wrapper_6__ap_ready(PE_wrapper_6__ap_ready),
    .PE_wrapper_6__ap_done(PE_wrapper_6__ap_done),
    .PE_wrapper_6__ap_idle(PE_wrapper_6__ap_idle),
    .PE_wrapper_7__ap_start(PE_wrapper_7__ap_start),
    .PE_wrapper_7__ap_ready(PE_wrapper_7__ap_ready),
    .PE_wrapper_7__ap_done(PE_wrapper_7__ap_done),
    .PE_wrapper_7__ap_idle(PE_wrapper_7__ap_idle),
    .PE_wrapper_8__ap_start(PE_wrapper_8__ap_start),
    .PE_wrapper_8__ap_ready(PE_wrapper_8__ap_ready),
    .PE_wrapper_8__ap_done(PE_wrapper_8__ap_done),
    .PE_wrapper_8__ap_idle(PE_wrapper_8__ap_idle),
    .PE_wrapper_9__ap_start(PE_wrapper_9__ap_start),
    .PE_wrapper_9__ap_ready(PE_wrapper_9__ap_ready),
    .PE_wrapper_9__ap_done(PE_wrapper_9__ap_done),
    .PE_wrapper_9__ap_idle(PE_wrapper_9__ap_idle),
    .PE_wrapper_10__ap_start(PE_wrapper_10__ap_start),
    .PE_wrapper_10__ap_ready(PE_wrapper_10__ap_ready),
    .PE_wrapper_10__ap_done(PE_wrapper_10__ap_done),
    .PE_wrapper_10__ap_idle(PE_wrapper_10__ap_idle),
    .PE_wrapper_11__ap_start(PE_wrapper_11__ap_start),
    .PE_wrapper_11__ap_ready(PE_wrapper_11__ap_ready),
    .PE_wrapper_11__ap_done(PE_wrapper_11__ap_done),
    .PE_wrapper_11__ap_idle(PE_wrapper_11__ap_idle),
    .PE_wrapper_12__ap_start(PE_wrapper_12__ap_start),
    .PE_wrapper_12__ap_ready(PE_wrapper_12__ap_ready),
    .PE_wrapper_12__ap_done(PE_wrapper_12__ap_done),
    .PE_wrapper_12__ap_idle(PE_wrapper_12__ap_idle),
    .PE_wrapper_13__ap_start(PE_wrapper_13__ap_start),
    .PE_wrapper_13__ap_ready(PE_wrapper_13__ap_ready),
    .PE_wrapper_13__ap_done(PE_wrapper_13__ap_done),
    .PE_wrapper_13__ap_idle(PE_wrapper_13__ap_idle),
    .PE_wrapper_14__ap_start(PE_wrapper_14__ap_start),
    .PE_wrapper_14__ap_ready(PE_wrapper_14__ap_ready),
    .PE_wrapper_14__ap_done(PE_wrapper_14__ap_done),
    .PE_wrapper_14__ap_idle(PE_wrapper_14__ap_idle),
    .PE_wrapper_15__ap_start(PE_wrapper_15__ap_start),
    .PE_wrapper_15__ap_ready(PE_wrapper_15__ap_ready),
    .PE_wrapper_15__ap_done(PE_wrapper_15__ap_done),
    .PE_wrapper_15__ap_idle(PE_wrapper_15__ap_idle),
    .PE_wrapper_16__ap_start(PE_wrapper_16__ap_start),
    .PE_wrapper_16__ap_ready(PE_wrapper_16__ap_ready),
    .PE_wrapper_16__ap_done(PE_wrapper_16__ap_done),
    .PE_wrapper_16__ap_idle(PE_wrapper_16__ap_idle),
    .PE_wrapper_17__ap_start(PE_wrapper_17__ap_start),
    .PE_wrapper_17__ap_ready(PE_wrapper_17__ap_ready),
    .PE_wrapper_17__ap_done(PE_wrapper_17__ap_done),
    .PE_wrapper_17__ap_idle(PE_wrapper_17__ap_idle),
    .PE_wrapper_18__ap_start(PE_wrapper_18__ap_start),
    .PE_wrapper_18__ap_ready(PE_wrapper_18__ap_ready),
    .PE_wrapper_18__ap_done(PE_wrapper_18__ap_done),
    .PE_wrapper_18__ap_idle(PE_wrapper_18__ap_idle),
    .PE_wrapper_19__ap_start(PE_wrapper_19__ap_start),
    .PE_wrapper_19__ap_ready(PE_wrapper_19__ap_ready),
    .PE_wrapper_19__ap_done(PE_wrapper_19__ap_done),
    .PE_wrapper_19__ap_idle(PE_wrapper_19__ap_idle),
    .PE_wrapper_20__ap_start(PE_wrapper_20__ap_start),
    .PE_wrapper_20__ap_ready(PE_wrapper_20__ap_ready),
    .PE_wrapper_20__ap_done(PE_wrapper_20__ap_done),
    .PE_wrapper_20__ap_idle(PE_wrapper_20__ap_idle),
    .PE_wrapper_21__ap_start(PE_wrapper_21__ap_start),
    .PE_wrapper_21__ap_ready(PE_wrapper_21__ap_ready),
    .PE_wrapper_21__ap_done(PE_wrapper_21__ap_done),
    .PE_wrapper_21__ap_idle(PE_wrapper_21__ap_idle),
    .PE_wrapper_22__ap_start(PE_wrapper_22__ap_start),
    .PE_wrapper_22__ap_ready(PE_wrapper_22__ap_ready),
    .PE_wrapper_22__ap_done(PE_wrapper_22__ap_done),
    .PE_wrapper_22__ap_idle(PE_wrapper_22__ap_idle),
    .PE_wrapper_23__ap_start(PE_wrapper_23__ap_start),
    .PE_wrapper_23__ap_ready(PE_wrapper_23__ap_ready),
    .PE_wrapper_23__ap_done(PE_wrapper_23__ap_done),
    .PE_wrapper_23__ap_idle(PE_wrapper_23__ap_idle),
    .PE_wrapper_24__ap_start(PE_wrapper_24__ap_start),
    .PE_wrapper_24__ap_ready(PE_wrapper_24__ap_ready),
    .PE_wrapper_24__ap_done(PE_wrapper_24__ap_done),
    .PE_wrapper_24__ap_idle(PE_wrapper_24__ap_idle),
    .PE_wrapper_25__ap_start(PE_wrapper_25__ap_start),
    .PE_wrapper_25__ap_ready(PE_wrapper_25__ap_ready),
    .PE_wrapper_25__ap_done(PE_wrapper_25__ap_done),
    .PE_wrapper_25__ap_idle(PE_wrapper_25__ap_idle),
    .PE_wrapper_26__ap_start(PE_wrapper_26__ap_start),
    .PE_wrapper_26__ap_ready(PE_wrapper_26__ap_ready),
    .PE_wrapper_26__ap_done(PE_wrapper_26__ap_done),
    .PE_wrapper_26__ap_idle(PE_wrapper_26__ap_idle),
    .PE_wrapper_27__ap_start(PE_wrapper_27__ap_start),
    .PE_wrapper_27__ap_ready(PE_wrapper_27__ap_ready),
    .PE_wrapper_27__ap_done(PE_wrapper_27__ap_done),
    .PE_wrapper_27__ap_idle(PE_wrapper_27__ap_idle),
    .PE_wrapper_28__ap_start(PE_wrapper_28__ap_start),
    .PE_wrapper_28__ap_ready(PE_wrapper_28__ap_ready),
    .PE_wrapper_28__ap_done(PE_wrapper_28__ap_done),
    .PE_wrapper_28__ap_idle(PE_wrapper_28__ap_idle),
    .PE_wrapper_29__ap_start(PE_wrapper_29__ap_start),
    .PE_wrapper_29__ap_ready(PE_wrapper_29__ap_ready),
    .PE_wrapper_29__ap_done(PE_wrapper_29__ap_done),
    .PE_wrapper_29__ap_idle(PE_wrapper_29__ap_idle),
    .PE_wrapper_30__ap_start(PE_wrapper_30__ap_start),
    .PE_wrapper_30__ap_ready(PE_wrapper_30__ap_ready),
    .PE_wrapper_30__ap_done(PE_wrapper_30__ap_done),
    .PE_wrapper_30__ap_idle(PE_wrapper_30__ap_idle),
    .PE_wrapper_31__ap_start(PE_wrapper_31__ap_start),
    .PE_wrapper_31__ap_ready(PE_wrapper_31__ap_ready),
    .PE_wrapper_31__ap_done(PE_wrapper_31__ap_done),
    .PE_wrapper_31__ap_idle(PE_wrapper_31__ap_idle),
    .PE_wrapper_32__ap_start(PE_wrapper_32__ap_start),
    .PE_wrapper_32__ap_ready(PE_wrapper_32__ap_ready),
    .PE_wrapper_32__ap_done(PE_wrapper_32__ap_done),
    .PE_wrapper_32__ap_idle(PE_wrapper_32__ap_idle),
    .PE_wrapper_33__ap_start(PE_wrapper_33__ap_start),
    .PE_wrapper_33__ap_ready(PE_wrapper_33__ap_ready),
    .PE_wrapper_33__ap_done(PE_wrapper_33__ap_done),
    .PE_wrapper_33__ap_idle(PE_wrapper_33__ap_idle),
    .PE_wrapper_34__ap_start(PE_wrapper_34__ap_start),
    .PE_wrapper_34__ap_ready(PE_wrapper_34__ap_ready),
    .PE_wrapper_34__ap_done(PE_wrapper_34__ap_done),
    .PE_wrapper_34__ap_idle(PE_wrapper_34__ap_idle),
    .PE_wrapper_35__ap_start(PE_wrapper_35__ap_start),
    .PE_wrapper_35__ap_ready(PE_wrapper_35__ap_ready),
    .PE_wrapper_35__ap_done(PE_wrapper_35__ap_done),
    .PE_wrapper_35__ap_idle(PE_wrapper_35__ap_idle),
    .PE_wrapper_36__ap_start(PE_wrapper_36__ap_start),
    .PE_wrapper_36__ap_ready(PE_wrapper_36__ap_ready),
    .PE_wrapper_36__ap_done(PE_wrapper_36__ap_done),
    .PE_wrapper_36__ap_idle(PE_wrapper_36__ap_idle),
    .PE_wrapper_37__ap_start(PE_wrapper_37__ap_start),
    .PE_wrapper_37__ap_ready(PE_wrapper_37__ap_ready),
    .PE_wrapper_37__ap_done(PE_wrapper_37__ap_done),
    .PE_wrapper_37__ap_idle(PE_wrapper_37__ap_idle),
    .PE_wrapper_38__ap_start(PE_wrapper_38__ap_start),
    .PE_wrapper_38__ap_ready(PE_wrapper_38__ap_ready),
    .PE_wrapper_38__ap_done(PE_wrapper_38__ap_done),
    .PE_wrapper_38__ap_idle(PE_wrapper_38__ap_idle),
    .PE_wrapper_39__ap_start(PE_wrapper_39__ap_start),
    .PE_wrapper_39__ap_ready(PE_wrapper_39__ap_ready),
    .PE_wrapper_39__ap_done(PE_wrapper_39__ap_done),
    .PE_wrapper_39__ap_idle(PE_wrapper_39__ap_idle),
    .PE_wrapper_40__ap_start(PE_wrapper_40__ap_start),
    .PE_wrapper_40__ap_ready(PE_wrapper_40__ap_ready),
    .PE_wrapper_40__ap_done(PE_wrapper_40__ap_done),
    .PE_wrapper_40__ap_idle(PE_wrapper_40__ap_idle),
    .PE_wrapper_41__ap_start(PE_wrapper_41__ap_start),
    .PE_wrapper_41__ap_ready(PE_wrapper_41__ap_ready),
    .PE_wrapper_41__ap_done(PE_wrapper_41__ap_done),
    .PE_wrapper_41__ap_idle(PE_wrapper_41__ap_idle),
    .PE_wrapper_42__ap_start(PE_wrapper_42__ap_start),
    .PE_wrapper_42__ap_ready(PE_wrapper_42__ap_ready),
    .PE_wrapper_42__ap_done(PE_wrapper_42__ap_done),
    .PE_wrapper_42__ap_idle(PE_wrapper_42__ap_idle),
    .PE_wrapper_43__ap_start(PE_wrapper_43__ap_start),
    .PE_wrapper_43__ap_ready(PE_wrapper_43__ap_ready),
    .PE_wrapper_43__ap_done(PE_wrapper_43__ap_done),
    .PE_wrapper_43__ap_idle(PE_wrapper_43__ap_idle),
    .PE_wrapper_44__ap_start(PE_wrapper_44__ap_start),
    .PE_wrapper_44__ap_ready(PE_wrapper_44__ap_ready),
    .PE_wrapper_44__ap_done(PE_wrapper_44__ap_done),
    .PE_wrapper_44__ap_idle(PE_wrapper_44__ap_idle),
    .PE_wrapper_45__ap_start(PE_wrapper_45__ap_start),
    .PE_wrapper_45__ap_ready(PE_wrapper_45__ap_ready),
    .PE_wrapper_45__ap_done(PE_wrapper_45__ap_done),
    .PE_wrapper_45__ap_idle(PE_wrapper_45__ap_idle),
    .PE_wrapper_46__ap_start(PE_wrapper_46__ap_start),
    .PE_wrapper_46__ap_ready(PE_wrapper_46__ap_ready),
    .PE_wrapper_46__ap_done(PE_wrapper_46__ap_done),
    .PE_wrapper_46__ap_idle(PE_wrapper_46__ap_idle),
    .PE_wrapper_47__ap_start(PE_wrapper_47__ap_start),
    .PE_wrapper_47__ap_ready(PE_wrapper_47__ap_ready),
    .PE_wrapper_47__ap_done(PE_wrapper_47__ap_done),
    .PE_wrapper_47__ap_idle(PE_wrapper_47__ap_idle),
    .PE_wrapper_48__ap_start(PE_wrapper_48__ap_start),
    .PE_wrapper_48__ap_ready(PE_wrapper_48__ap_ready),
    .PE_wrapper_48__ap_done(PE_wrapper_48__ap_done),
    .PE_wrapper_48__ap_idle(PE_wrapper_48__ap_idle),
    .PE_wrapper_49__ap_start(PE_wrapper_49__ap_start),
    .PE_wrapper_49__ap_ready(PE_wrapper_49__ap_ready),
    .PE_wrapper_49__ap_done(PE_wrapper_49__ap_done),
    .PE_wrapper_49__ap_idle(PE_wrapper_49__ap_idle),
    .PE_wrapper_50__ap_start(PE_wrapper_50__ap_start),
    .PE_wrapper_50__ap_ready(PE_wrapper_50__ap_ready),
    .PE_wrapper_50__ap_done(PE_wrapper_50__ap_done),
    .PE_wrapper_50__ap_idle(PE_wrapper_50__ap_idle),
    .PE_wrapper_51__ap_start(PE_wrapper_51__ap_start),
    .PE_wrapper_51__ap_ready(PE_wrapper_51__ap_ready),
    .PE_wrapper_51__ap_done(PE_wrapper_51__ap_done),
    .PE_wrapper_51__ap_idle(PE_wrapper_51__ap_idle),
    .PE_wrapper_52__ap_start(PE_wrapper_52__ap_start),
    .PE_wrapper_52__ap_ready(PE_wrapper_52__ap_ready),
    .PE_wrapper_52__ap_done(PE_wrapper_52__ap_done),
    .PE_wrapper_52__ap_idle(PE_wrapper_52__ap_idle),
    .PE_wrapper_53__ap_start(PE_wrapper_53__ap_start),
    .PE_wrapper_53__ap_ready(PE_wrapper_53__ap_ready),
    .PE_wrapper_53__ap_done(PE_wrapper_53__ap_done),
    .PE_wrapper_53__ap_idle(PE_wrapper_53__ap_idle),
    .PE_wrapper_54__ap_start(PE_wrapper_54__ap_start),
    .PE_wrapper_54__ap_ready(PE_wrapper_54__ap_ready),
    .PE_wrapper_54__ap_done(PE_wrapper_54__ap_done),
    .PE_wrapper_54__ap_idle(PE_wrapper_54__ap_idle),
    .PE_wrapper_55__ap_start(PE_wrapper_55__ap_start),
    .PE_wrapper_55__ap_ready(PE_wrapper_55__ap_ready),
    .PE_wrapper_55__ap_done(PE_wrapper_55__ap_done),
    .PE_wrapper_55__ap_idle(PE_wrapper_55__ap_idle),
    .PE_wrapper_56__ap_start(PE_wrapper_56__ap_start),
    .PE_wrapper_56__ap_ready(PE_wrapper_56__ap_ready),
    .PE_wrapper_56__ap_done(PE_wrapper_56__ap_done),
    .PE_wrapper_56__ap_idle(PE_wrapper_56__ap_idle),
    .PE_wrapper_57__ap_start(PE_wrapper_57__ap_start),
    .PE_wrapper_57__ap_ready(PE_wrapper_57__ap_ready),
    .PE_wrapper_57__ap_done(PE_wrapper_57__ap_done),
    .PE_wrapper_57__ap_idle(PE_wrapper_57__ap_idle),
    .PE_wrapper_58__ap_start(PE_wrapper_58__ap_start),
    .PE_wrapper_58__ap_ready(PE_wrapper_58__ap_ready),
    .PE_wrapper_58__ap_done(PE_wrapper_58__ap_done),
    .PE_wrapper_58__ap_idle(PE_wrapper_58__ap_idle),
    .PE_wrapper_59__ap_start(PE_wrapper_59__ap_start),
    .PE_wrapper_59__ap_ready(PE_wrapper_59__ap_ready),
    .PE_wrapper_59__ap_done(PE_wrapper_59__ap_done),
    .PE_wrapper_59__ap_idle(PE_wrapper_59__ap_idle),
    .PE_wrapper_60__ap_start(PE_wrapper_60__ap_start),
    .PE_wrapper_60__ap_ready(PE_wrapper_60__ap_ready),
    .PE_wrapper_60__ap_done(PE_wrapper_60__ap_done),
    .PE_wrapper_60__ap_idle(PE_wrapper_60__ap_idle),
    .PE_wrapper_61__ap_start(PE_wrapper_61__ap_start),
    .PE_wrapper_61__ap_ready(PE_wrapper_61__ap_ready),
    .PE_wrapper_61__ap_done(PE_wrapper_61__ap_done),
    .PE_wrapper_61__ap_idle(PE_wrapper_61__ap_idle),
    .PE_wrapper_62__ap_start(PE_wrapper_62__ap_start),
    .PE_wrapper_62__ap_ready(PE_wrapper_62__ap_ready),
    .PE_wrapper_62__ap_done(PE_wrapper_62__ap_done),
    .PE_wrapper_62__ap_idle(PE_wrapper_62__ap_idle),
    .PE_wrapper_63__ap_start(PE_wrapper_63__ap_start),
    .PE_wrapper_63__ap_ready(PE_wrapper_63__ap_ready),
    .PE_wrapper_63__ap_done(PE_wrapper_63__ap_done),
    .PE_wrapper_63__ap_idle(PE_wrapper_63__ap_idle),
    .PE_wrapper_64__ap_start(PE_wrapper_64__ap_start),
    .PE_wrapper_64__ap_ready(PE_wrapper_64__ap_ready),
    .PE_wrapper_64__ap_done(PE_wrapper_64__ap_done),
    .PE_wrapper_64__ap_idle(PE_wrapper_64__ap_idle),
    .PE_wrapper_65__ap_start(PE_wrapper_65__ap_start),
    .PE_wrapper_65__ap_ready(PE_wrapper_65__ap_ready),
    .PE_wrapper_65__ap_done(PE_wrapper_65__ap_done),
    .PE_wrapper_65__ap_idle(PE_wrapper_65__ap_idle),
    .PE_wrapper_66__ap_start(PE_wrapper_66__ap_start),
    .PE_wrapper_66__ap_ready(PE_wrapper_66__ap_ready),
    .PE_wrapper_66__ap_done(PE_wrapper_66__ap_done),
    .PE_wrapper_66__ap_idle(PE_wrapper_66__ap_idle),
    .PE_wrapper_67__ap_start(PE_wrapper_67__ap_start),
    .PE_wrapper_67__ap_ready(PE_wrapper_67__ap_ready),
    .PE_wrapper_67__ap_done(PE_wrapper_67__ap_done),
    .PE_wrapper_67__ap_idle(PE_wrapper_67__ap_idle),
    .PE_wrapper_68__ap_start(PE_wrapper_68__ap_start),
    .PE_wrapper_68__ap_ready(PE_wrapper_68__ap_ready),
    .PE_wrapper_68__ap_done(PE_wrapper_68__ap_done),
    .PE_wrapper_68__ap_idle(PE_wrapper_68__ap_idle),
    .PE_wrapper_69__ap_start(PE_wrapper_69__ap_start),
    .PE_wrapper_69__ap_ready(PE_wrapper_69__ap_ready),
    .PE_wrapper_69__ap_done(PE_wrapper_69__ap_done),
    .PE_wrapper_69__ap_idle(PE_wrapper_69__ap_idle),
    .PE_wrapper_70__ap_start(PE_wrapper_70__ap_start),
    .PE_wrapper_70__ap_ready(PE_wrapper_70__ap_ready),
    .PE_wrapper_70__ap_done(PE_wrapper_70__ap_done),
    .PE_wrapper_70__ap_idle(PE_wrapper_70__ap_idle),
    .PE_wrapper_71__ap_start(PE_wrapper_71__ap_start),
    .PE_wrapper_71__ap_ready(PE_wrapper_71__ap_ready),
    .PE_wrapper_71__ap_done(PE_wrapper_71__ap_done),
    .PE_wrapper_71__ap_idle(PE_wrapper_71__ap_idle),
    .PE_wrapper_72__ap_start(PE_wrapper_72__ap_start),
    .PE_wrapper_72__ap_ready(PE_wrapper_72__ap_ready),
    .PE_wrapper_72__ap_done(PE_wrapper_72__ap_done),
    .PE_wrapper_72__ap_idle(PE_wrapper_72__ap_idle),
    .PE_wrapper_73__ap_start(PE_wrapper_73__ap_start),
    .PE_wrapper_73__ap_ready(PE_wrapper_73__ap_ready),
    .PE_wrapper_73__ap_done(PE_wrapper_73__ap_done),
    .PE_wrapper_73__ap_idle(PE_wrapper_73__ap_idle),
    .PE_wrapper_74__ap_start(PE_wrapper_74__ap_start),
    .PE_wrapper_74__ap_ready(PE_wrapper_74__ap_ready),
    .PE_wrapper_74__ap_done(PE_wrapper_74__ap_done),
    .PE_wrapper_74__ap_idle(PE_wrapper_74__ap_idle),
    .PE_wrapper_75__ap_start(PE_wrapper_75__ap_start),
    .PE_wrapper_75__ap_ready(PE_wrapper_75__ap_ready),
    .PE_wrapper_75__ap_done(PE_wrapper_75__ap_done),
    .PE_wrapper_75__ap_idle(PE_wrapper_75__ap_idle),
    .PE_wrapper_76__ap_start(PE_wrapper_76__ap_start),
    .PE_wrapper_76__ap_ready(PE_wrapper_76__ap_ready),
    .PE_wrapper_76__ap_done(PE_wrapper_76__ap_done),
    .PE_wrapper_76__ap_idle(PE_wrapper_76__ap_idle),
    .PE_wrapper_77__ap_start(PE_wrapper_77__ap_start),
    .PE_wrapper_77__ap_ready(PE_wrapper_77__ap_ready),
    .PE_wrapper_77__ap_done(PE_wrapper_77__ap_done),
    .PE_wrapper_77__ap_idle(PE_wrapper_77__ap_idle),
    .PE_wrapper_78__ap_start(PE_wrapper_78__ap_start),
    .PE_wrapper_78__ap_ready(PE_wrapper_78__ap_ready),
    .PE_wrapper_78__ap_done(PE_wrapper_78__ap_done),
    .PE_wrapper_78__ap_idle(PE_wrapper_78__ap_idle),
    .PE_wrapper_79__ap_start(PE_wrapper_79__ap_start),
    .PE_wrapper_79__ap_ready(PE_wrapper_79__ap_ready),
    .PE_wrapper_79__ap_done(PE_wrapper_79__ap_done),
    .PE_wrapper_79__ap_idle(PE_wrapper_79__ap_idle),
    .PE_wrapper_80__ap_start(PE_wrapper_80__ap_start),
    .PE_wrapper_80__ap_ready(PE_wrapper_80__ap_ready),
    .PE_wrapper_80__ap_done(PE_wrapper_80__ap_done),
    .PE_wrapper_80__ap_idle(PE_wrapper_80__ap_idle),
    .PE_wrapper_81__ap_start(PE_wrapper_81__ap_start),
    .PE_wrapper_81__ap_ready(PE_wrapper_81__ap_ready),
    .PE_wrapper_81__ap_done(PE_wrapper_81__ap_done),
    .PE_wrapper_81__ap_idle(PE_wrapper_81__ap_idle),
    .PE_wrapper_82__ap_start(PE_wrapper_82__ap_start),
    .PE_wrapper_82__ap_ready(PE_wrapper_82__ap_ready),
    .PE_wrapper_82__ap_done(PE_wrapper_82__ap_done),
    .PE_wrapper_82__ap_idle(PE_wrapper_82__ap_idle),
    .PE_wrapper_83__ap_start(PE_wrapper_83__ap_start),
    .PE_wrapper_83__ap_ready(PE_wrapper_83__ap_ready),
    .PE_wrapper_83__ap_done(PE_wrapper_83__ap_done),
    .PE_wrapper_83__ap_idle(PE_wrapper_83__ap_idle),
    .PE_wrapper_84__ap_start(PE_wrapper_84__ap_start),
    .PE_wrapper_84__ap_ready(PE_wrapper_84__ap_ready),
    .PE_wrapper_84__ap_done(PE_wrapper_84__ap_done),
    .PE_wrapper_84__ap_idle(PE_wrapper_84__ap_idle),
    .PE_wrapper_85__ap_start(PE_wrapper_85__ap_start),
    .PE_wrapper_85__ap_ready(PE_wrapper_85__ap_ready),
    .PE_wrapper_85__ap_done(PE_wrapper_85__ap_done),
    .PE_wrapper_85__ap_idle(PE_wrapper_85__ap_idle),
    .PE_wrapper_86__ap_start(PE_wrapper_86__ap_start),
    .PE_wrapper_86__ap_ready(PE_wrapper_86__ap_ready),
    .PE_wrapper_86__ap_done(PE_wrapper_86__ap_done),
    .PE_wrapper_86__ap_idle(PE_wrapper_86__ap_idle),
    .PE_wrapper_87__ap_start(PE_wrapper_87__ap_start),
    .PE_wrapper_87__ap_ready(PE_wrapper_87__ap_ready),
    .PE_wrapper_87__ap_done(PE_wrapper_87__ap_done),
    .PE_wrapper_87__ap_idle(PE_wrapper_87__ap_idle),
    .PE_wrapper_88__ap_start(PE_wrapper_88__ap_start),
    .PE_wrapper_88__ap_ready(PE_wrapper_88__ap_ready),
    .PE_wrapper_88__ap_done(PE_wrapper_88__ap_done),
    .PE_wrapper_88__ap_idle(PE_wrapper_88__ap_idle),
    .PE_wrapper_89__ap_start(PE_wrapper_89__ap_start),
    .PE_wrapper_89__ap_ready(PE_wrapper_89__ap_ready),
    .PE_wrapper_89__ap_done(PE_wrapper_89__ap_done),
    .PE_wrapper_89__ap_idle(PE_wrapper_89__ap_idle),
    .PE_wrapper_90__ap_start(PE_wrapper_90__ap_start),
    .PE_wrapper_90__ap_ready(PE_wrapper_90__ap_ready),
    .PE_wrapper_90__ap_done(PE_wrapper_90__ap_done),
    .PE_wrapper_90__ap_idle(PE_wrapper_90__ap_idle),
    .PE_wrapper_91__ap_start(PE_wrapper_91__ap_start),
    .PE_wrapper_91__ap_ready(PE_wrapper_91__ap_ready),
    .PE_wrapper_91__ap_done(PE_wrapper_91__ap_done),
    .PE_wrapper_91__ap_idle(PE_wrapper_91__ap_idle),
    .PE_wrapper_92__ap_start(PE_wrapper_92__ap_start),
    .PE_wrapper_92__ap_ready(PE_wrapper_92__ap_ready),
    .PE_wrapper_92__ap_done(PE_wrapper_92__ap_done),
    .PE_wrapper_92__ap_idle(PE_wrapper_92__ap_idle),
    .PE_wrapper_93__ap_start(PE_wrapper_93__ap_start),
    .PE_wrapper_93__ap_ready(PE_wrapper_93__ap_ready),
    .PE_wrapper_93__ap_done(PE_wrapper_93__ap_done),
    .PE_wrapper_93__ap_idle(PE_wrapper_93__ap_idle),
    .PE_wrapper_94__ap_start(PE_wrapper_94__ap_start),
    .PE_wrapper_94__ap_ready(PE_wrapper_94__ap_ready),
    .PE_wrapper_94__ap_done(PE_wrapper_94__ap_done),
    .PE_wrapper_94__ap_idle(PE_wrapper_94__ap_idle),
    .PE_wrapper_95__ap_start(PE_wrapper_95__ap_start),
    .PE_wrapper_95__ap_ready(PE_wrapper_95__ap_ready),
    .PE_wrapper_95__ap_done(PE_wrapper_95__ap_done),
    .PE_wrapper_95__ap_idle(PE_wrapper_95__ap_idle),
    .PE_wrapper_96__ap_start(PE_wrapper_96__ap_start),
    .PE_wrapper_96__ap_ready(PE_wrapper_96__ap_ready),
    .PE_wrapper_96__ap_done(PE_wrapper_96__ap_done),
    .PE_wrapper_96__ap_idle(PE_wrapper_96__ap_idle),
    .PE_wrapper_97__ap_start(PE_wrapper_97__ap_start),
    .PE_wrapper_97__ap_ready(PE_wrapper_97__ap_ready),
    .PE_wrapper_97__ap_done(PE_wrapper_97__ap_done),
    .PE_wrapper_97__ap_idle(PE_wrapper_97__ap_idle),
    .PE_wrapper_98__ap_start(PE_wrapper_98__ap_start),
    .PE_wrapper_98__ap_ready(PE_wrapper_98__ap_ready),
    .PE_wrapper_98__ap_done(PE_wrapper_98__ap_done),
    .PE_wrapper_98__ap_idle(PE_wrapper_98__ap_idle),
    .PE_wrapper_99__ap_start(PE_wrapper_99__ap_start),
    .PE_wrapper_99__ap_ready(PE_wrapper_99__ap_ready),
    .PE_wrapper_99__ap_done(PE_wrapper_99__ap_done),
    .PE_wrapper_99__ap_idle(PE_wrapper_99__ap_idle),
    .PE_wrapper_100__ap_start(PE_wrapper_100__ap_start),
    .PE_wrapper_100__ap_ready(PE_wrapper_100__ap_ready),
    .PE_wrapper_100__ap_done(PE_wrapper_100__ap_done),
    .PE_wrapper_100__ap_idle(PE_wrapper_100__ap_idle),
    .PE_wrapper_101__ap_start(PE_wrapper_101__ap_start),
    .PE_wrapper_101__ap_ready(PE_wrapper_101__ap_ready),
    .PE_wrapper_101__ap_done(PE_wrapper_101__ap_done),
    .PE_wrapper_101__ap_idle(PE_wrapper_101__ap_idle),
    .PE_wrapper_102__ap_start(PE_wrapper_102__ap_start),
    .PE_wrapper_102__ap_ready(PE_wrapper_102__ap_ready),
    .PE_wrapper_102__ap_done(PE_wrapper_102__ap_done),
    .PE_wrapper_102__ap_idle(PE_wrapper_102__ap_idle),
    .PE_wrapper_103__ap_start(PE_wrapper_103__ap_start),
    .PE_wrapper_103__ap_ready(PE_wrapper_103__ap_ready),
    .PE_wrapper_103__ap_done(PE_wrapper_103__ap_done),
    .PE_wrapper_103__ap_idle(PE_wrapper_103__ap_idle),
    .PE_wrapper_104__ap_start(PE_wrapper_104__ap_start),
    .PE_wrapper_104__ap_ready(PE_wrapper_104__ap_ready),
    .PE_wrapper_104__ap_done(PE_wrapper_104__ap_done),
    .PE_wrapper_104__ap_idle(PE_wrapper_104__ap_idle),
    .PE_wrapper_105__ap_start(PE_wrapper_105__ap_start),
    .PE_wrapper_105__ap_ready(PE_wrapper_105__ap_ready),
    .PE_wrapper_105__ap_done(PE_wrapper_105__ap_done),
    .PE_wrapper_105__ap_idle(PE_wrapper_105__ap_idle),
    .PE_wrapper_106__ap_start(PE_wrapper_106__ap_start),
    .PE_wrapper_106__ap_ready(PE_wrapper_106__ap_ready),
    .PE_wrapper_106__ap_done(PE_wrapper_106__ap_done),
    .PE_wrapper_106__ap_idle(PE_wrapper_106__ap_idle),
    .PE_wrapper_107__ap_start(PE_wrapper_107__ap_start),
    .PE_wrapper_107__ap_ready(PE_wrapper_107__ap_ready),
    .PE_wrapper_107__ap_done(PE_wrapper_107__ap_done),
    .PE_wrapper_107__ap_idle(PE_wrapper_107__ap_idle),
    .PE_wrapper_108__ap_start(PE_wrapper_108__ap_start),
    .PE_wrapper_108__ap_ready(PE_wrapper_108__ap_ready),
    .PE_wrapper_108__ap_done(PE_wrapper_108__ap_done),
    .PE_wrapper_108__ap_idle(PE_wrapper_108__ap_idle),
    .PE_wrapper_109__ap_start(PE_wrapper_109__ap_start),
    .PE_wrapper_109__ap_ready(PE_wrapper_109__ap_ready),
    .PE_wrapper_109__ap_done(PE_wrapper_109__ap_done),
    .PE_wrapper_109__ap_idle(PE_wrapper_109__ap_idle),
    .PE_wrapper_110__ap_start(PE_wrapper_110__ap_start),
    .PE_wrapper_110__ap_ready(PE_wrapper_110__ap_ready),
    .PE_wrapper_110__ap_done(PE_wrapper_110__ap_done),
    .PE_wrapper_110__ap_idle(PE_wrapper_110__ap_idle),
    .PE_wrapper_111__ap_start(PE_wrapper_111__ap_start),
    .PE_wrapper_111__ap_ready(PE_wrapper_111__ap_ready),
    .PE_wrapper_111__ap_done(PE_wrapper_111__ap_done),
    .PE_wrapper_111__ap_idle(PE_wrapper_111__ap_idle),
    .PE_wrapper_112__ap_start(PE_wrapper_112__ap_start),
    .PE_wrapper_112__ap_ready(PE_wrapper_112__ap_ready),
    .PE_wrapper_112__ap_done(PE_wrapper_112__ap_done),
    .PE_wrapper_112__ap_idle(PE_wrapper_112__ap_idle),
    .PE_wrapper_113__ap_start(PE_wrapper_113__ap_start),
    .PE_wrapper_113__ap_ready(PE_wrapper_113__ap_ready),
    .PE_wrapper_113__ap_done(PE_wrapper_113__ap_done),
    .PE_wrapper_113__ap_idle(PE_wrapper_113__ap_idle),
    .PE_wrapper_114__ap_start(PE_wrapper_114__ap_start),
    .PE_wrapper_114__ap_ready(PE_wrapper_114__ap_ready),
    .PE_wrapper_114__ap_done(PE_wrapper_114__ap_done),
    .PE_wrapper_114__ap_idle(PE_wrapper_114__ap_idle),
    .PE_wrapper_115__ap_start(PE_wrapper_115__ap_start),
    .PE_wrapper_115__ap_ready(PE_wrapper_115__ap_ready),
    .PE_wrapper_115__ap_done(PE_wrapper_115__ap_done),
    .PE_wrapper_115__ap_idle(PE_wrapper_115__ap_idle),
    .PE_wrapper_116__ap_start(PE_wrapper_116__ap_start),
    .PE_wrapper_116__ap_ready(PE_wrapper_116__ap_ready),
    .PE_wrapper_116__ap_done(PE_wrapper_116__ap_done),
    .PE_wrapper_116__ap_idle(PE_wrapper_116__ap_idle),
    .PE_wrapper_117__ap_start(PE_wrapper_117__ap_start),
    .PE_wrapper_117__ap_ready(PE_wrapper_117__ap_ready),
    .PE_wrapper_117__ap_done(PE_wrapper_117__ap_done),
    .PE_wrapper_117__ap_idle(PE_wrapper_117__ap_idle),
    .PE_wrapper_118__ap_start(PE_wrapper_118__ap_start),
    .PE_wrapper_118__ap_ready(PE_wrapper_118__ap_ready),
    .PE_wrapper_118__ap_done(PE_wrapper_118__ap_done),
    .PE_wrapper_118__ap_idle(PE_wrapper_118__ap_idle),
    .PE_wrapper_119__ap_start(PE_wrapper_119__ap_start),
    .PE_wrapper_119__ap_ready(PE_wrapper_119__ap_ready),
    .PE_wrapper_119__ap_done(PE_wrapper_119__ap_done),
    .PE_wrapper_119__ap_idle(PE_wrapper_119__ap_idle),
    .PE_wrapper_120__ap_start(PE_wrapper_120__ap_start),
    .PE_wrapper_120__ap_ready(PE_wrapper_120__ap_ready),
    .PE_wrapper_120__ap_done(PE_wrapper_120__ap_done),
    .PE_wrapper_120__ap_idle(PE_wrapper_120__ap_idle),
    .PE_wrapper_121__ap_start(PE_wrapper_121__ap_start),
    .PE_wrapper_121__ap_ready(PE_wrapper_121__ap_ready),
    .PE_wrapper_121__ap_done(PE_wrapper_121__ap_done),
    .PE_wrapper_121__ap_idle(PE_wrapper_121__ap_idle),
    .PE_wrapper_122__ap_start(PE_wrapper_122__ap_start),
    .PE_wrapper_122__ap_ready(PE_wrapper_122__ap_ready),
    .PE_wrapper_122__ap_done(PE_wrapper_122__ap_done),
    .PE_wrapper_122__ap_idle(PE_wrapper_122__ap_idle),
    .PE_wrapper_123__ap_start(PE_wrapper_123__ap_start),
    .PE_wrapper_123__ap_ready(PE_wrapper_123__ap_ready),
    .PE_wrapper_123__ap_done(PE_wrapper_123__ap_done),
    .PE_wrapper_123__ap_idle(PE_wrapper_123__ap_idle),
    .PE_wrapper_124__ap_start(PE_wrapper_124__ap_start),
    .PE_wrapper_124__ap_ready(PE_wrapper_124__ap_ready),
    .PE_wrapper_124__ap_done(PE_wrapper_124__ap_done),
    .PE_wrapper_124__ap_idle(PE_wrapper_124__ap_idle),
    .PE_wrapper_125__ap_start(PE_wrapper_125__ap_start),
    .PE_wrapper_125__ap_ready(PE_wrapper_125__ap_ready),
    .PE_wrapper_125__ap_done(PE_wrapper_125__ap_done),
    .PE_wrapper_125__ap_idle(PE_wrapper_125__ap_idle),
    .PE_wrapper_126__ap_start(PE_wrapper_126__ap_start),
    .PE_wrapper_126__ap_ready(PE_wrapper_126__ap_ready),
    .PE_wrapper_126__ap_done(PE_wrapper_126__ap_done),
    .PE_wrapper_126__ap_idle(PE_wrapper_126__ap_idle),
    .PE_wrapper_127__ap_start(PE_wrapper_127__ap_start),
    .PE_wrapper_127__ap_ready(PE_wrapper_127__ap_ready),
    .PE_wrapper_127__ap_done(PE_wrapper_127__ap_done),
    .PE_wrapper_127__ap_idle(PE_wrapper_127__ap_idle),
    .PE_wrapper_128__ap_start(PE_wrapper_128__ap_start),
    .PE_wrapper_128__ap_ready(PE_wrapper_128__ap_ready),
    .PE_wrapper_128__ap_done(PE_wrapper_128__ap_done),
    .PE_wrapper_128__ap_idle(PE_wrapper_128__ap_idle),
    .PE_wrapper_129__ap_start(PE_wrapper_129__ap_start),
    .PE_wrapper_129__ap_ready(PE_wrapper_129__ap_ready),
    .PE_wrapper_129__ap_done(PE_wrapper_129__ap_done),
    .PE_wrapper_129__ap_idle(PE_wrapper_129__ap_idle),
    .PE_wrapper_130__ap_start(PE_wrapper_130__ap_start),
    .PE_wrapper_130__ap_ready(PE_wrapper_130__ap_ready),
    .PE_wrapper_130__ap_done(PE_wrapper_130__ap_done),
    .PE_wrapper_130__ap_idle(PE_wrapper_130__ap_idle),
    .PE_wrapper_131__ap_start(PE_wrapper_131__ap_start),
    .PE_wrapper_131__ap_ready(PE_wrapper_131__ap_ready),
    .PE_wrapper_131__ap_done(PE_wrapper_131__ap_done),
    .PE_wrapper_131__ap_idle(PE_wrapper_131__ap_idle),
    .PE_wrapper_132__ap_start(PE_wrapper_132__ap_start),
    .PE_wrapper_132__ap_ready(PE_wrapper_132__ap_ready),
    .PE_wrapper_132__ap_done(PE_wrapper_132__ap_done),
    .PE_wrapper_132__ap_idle(PE_wrapper_132__ap_idle),
    .PE_wrapper_133__ap_start(PE_wrapper_133__ap_start),
    .PE_wrapper_133__ap_ready(PE_wrapper_133__ap_ready),
    .PE_wrapper_133__ap_done(PE_wrapper_133__ap_done),
    .PE_wrapper_133__ap_idle(PE_wrapper_133__ap_idle),
    .PE_wrapper_134__ap_start(PE_wrapper_134__ap_start),
    .PE_wrapper_134__ap_ready(PE_wrapper_134__ap_ready),
    .PE_wrapper_134__ap_done(PE_wrapper_134__ap_done),
    .PE_wrapper_134__ap_idle(PE_wrapper_134__ap_idle),
    .PE_wrapper_135__ap_start(PE_wrapper_135__ap_start),
    .PE_wrapper_135__ap_ready(PE_wrapper_135__ap_ready),
    .PE_wrapper_135__ap_done(PE_wrapper_135__ap_done),
    .PE_wrapper_135__ap_idle(PE_wrapper_135__ap_idle),
    .PE_wrapper_136__ap_start(PE_wrapper_136__ap_start),
    .PE_wrapper_136__ap_ready(PE_wrapper_136__ap_ready),
    .PE_wrapper_136__ap_done(PE_wrapper_136__ap_done),
    .PE_wrapper_136__ap_idle(PE_wrapper_136__ap_idle),
    .PE_wrapper_137__ap_start(PE_wrapper_137__ap_start),
    .PE_wrapper_137__ap_ready(PE_wrapper_137__ap_ready),
    .PE_wrapper_137__ap_done(PE_wrapper_137__ap_done),
    .PE_wrapper_137__ap_idle(PE_wrapper_137__ap_idle),
    .PE_wrapper_138__ap_start(PE_wrapper_138__ap_start),
    .PE_wrapper_138__ap_ready(PE_wrapper_138__ap_ready),
    .PE_wrapper_138__ap_done(PE_wrapper_138__ap_done),
    .PE_wrapper_138__ap_idle(PE_wrapper_138__ap_idle),
    .PE_wrapper_139__ap_start(PE_wrapper_139__ap_start),
    .PE_wrapper_139__ap_ready(PE_wrapper_139__ap_ready),
    .PE_wrapper_139__ap_done(PE_wrapper_139__ap_done),
    .PE_wrapper_139__ap_idle(PE_wrapper_139__ap_idle),
    .PE_wrapper_140__ap_start(PE_wrapper_140__ap_start),
    .PE_wrapper_140__ap_ready(PE_wrapper_140__ap_ready),
    .PE_wrapper_140__ap_done(PE_wrapper_140__ap_done),
    .PE_wrapper_140__ap_idle(PE_wrapper_140__ap_idle),
    .PE_wrapper_141__ap_start(PE_wrapper_141__ap_start),
    .PE_wrapper_141__ap_ready(PE_wrapper_141__ap_ready),
    .PE_wrapper_141__ap_done(PE_wrapper_141__ap_done),
    .PE_wrapper_141__ap_idle(PE_wrapper_141__ap_idle),
    .PE_wrapper_142__ap_start(PE_wrapper_142__ap_start),
    .PE_wrapper_142__ap_ready(PE_wrapper_142__ap_ready),
    .PE_wrapper_142__ap_done(PE_wrapper_142__ap_done),
    .PE_wrapper_142__ap_idle(PE_wrapper_142__ap_idle),
    .PE_wrapper_143__ap_start(PE_wrapper_143__ap_start),
    .PE_wrapper_143__ap_ready(PE_wrapper_143__ap_ready),
    .PE_wrapper_143__ap_done(PE_wrapper_143__ap_done),
    .PE_wrapper_143__ap_idle(PE_wrapper_143__ap_idle),
    .PE_wrapper_144__ap_start(PE_wrapper_144__ap_start),
    .PE_wrapper_144__ap_ready(PE_wrapper_144__ap_ready),
    .PE_wrapper_144__ap_done(PE_wrapper_144__ap_done),
    .PE_wrapper_144__ap_idle(PE_wrapper_144__ap_idle),
    .PE_wrapper_145__ap_start(PE_wrapper_145__ap_start),
    .PE_wrapper_145__ap_ready(PE_wrapper_145__ap_ready),
    .PE_wrapper_145__ap_done(PE_wrapper_145__ap_done),
    .PE_wrapper_145__ap_idle(PE_wrapper_145__ap_idle),
    .PE_wrapper_146__ap_start(PE_wrapper_146__ap_start),
    .PE_wrapper_146__ap_ready(PE_wrapper_146__ap_ready),
    .PE_wrapper_146__ap_done(PE_wrapper_146__ap_done),
    .PE_wrapper_146__ap_idle(PE_wrapper_146__ap_idle),
    .PE_wrapper_147__ap_start(PE_wrapper_147__ap_start),
    .PE_wrapper_147__ap_ready(PE_wrapper_147__ap_ready),
    .PE_wrapper_147__ap_done(PE_wrapper_147__ap_done),
    .PE_wrapper_147__ap_idle(PE_wrapper_147__ap_idle),
    .PE_wrapper_148__ap_start(PE_wrapper_148__ap_start),
    .PE_wrapper_148__ap_ready(PE_wrapper_148__ap_ready),
    .PE_wrapper_148__ap_done(PE_wrapper_148__ap_done),
    .PE_wrapper_148__ap_idle(PE_wrapper_148__ap_idle),
    .PE_wrapper_149__ap_start(PE_wrapper_149__ap_start),
    .PE_wrapper_149__ap_ready(PE_wrapper_149__ap_ready),
    .PE_wrapper_149__ap_done(PE_wrapper_149__ap_done),
    .PE_wrapper_149__ap_idle(PE_wrapper_149__ap_idle),
    .PE_wrapper_150__ap_start(PE_wrapper_150__ap_start),
    .PE_wrapper_150__ap_ready(PE_wrapper_150__ap_ready),
    .PE_wrapper_150__ap_done(PE_wrapper_150__ap_done),
    .PE_wrapper_150__ap_idle(PE_wrapper_150__ap_idle),
    .PE_wrapper_151__ap_start(PE_wrapper_151__ap_start),
    .PE_wrapper_151__ap_ready(PE_wrapper_151__ap_ready),
    .PE_wrapper_151__ap_done(PE_wrapper_151__ap_done),
    .PE_wrapper_151__ap_idle(PE_wrapper_151__ap_idle),
    .PE_wrapper_152__ap_start(PE_wrapper_152__ap_start),
    .PE_wrapper_152__ap_ready(PE_wrapper_152__ap_ready),
    .PE_wrapper_152__ap_done(PE_wrapper_152__ap_done),
    .PE_wrapper_152__ap_idle(PE_wrapper_152__ap_idle),
    .PE_wrapper_153__ap_start(PE_wrapper_153__ap_start),
    .PE_wrapper_153__ap_ready(PE_wrapper_153__ap_ready),
    .PE_wrapper_153__ap_done(PE_wrapper_153__ap_done),
    .PE_wrapper_153__ap_idle(PE_wrapper_153__ap_idle),
    .PE_wrapper_154__ap_start(PE_wrapper_154__ap_start),
    .PE_wrapper_154__ap_ready(PE_wrapper_154__ap_ready),
    .PE_wrapper_154__ap_done(PE_wrapper_154__ap_done),
    .PE_wrapper_154__ap_idle(PE_wrapper_154__ap_idle),
    .PE_wrapper_155__ap_start(PE_wrapper_155__ap_start),
    .PE_wrapper_155__ap_ready(PE_wrapper_155__ap_ready),
    .PE_wrapper_155__ap_done(PE_wrapper_155__ap_done),
    .PE_wrapper_155__ap_idle(PE_wrapper_155__ap_idle),
    .PE_wrapper_156__ap_start(PE_wrapper_156__ap_start),
    .PE_wrapper_156__ap_ready(PE_wrapper_156__ap_ready),
    .PE_wrapper_156__ap_done(PE_wrapper_156__ap_done),
    .PE_wrapper_156__ap_idle(PE_wrapper_156__ap_idle),
    .PE_wrapper_157__ap_start(PE_wrapper_157__ap_start),
    .PE_wrapper_157__ap_ready(PE_wrapper_157__ap_ready),
    .PE_wrapper_157__ap_done(PE_wrapper_157__ap_done),
    .PE_wrapper_157__ap_idle(PE_wrapper_157__ap_idle),
    .PE_wrapper_158__ap_start(PE_wrapper_158__ap_start),
    .PE_wrapper_158__ap_ready(PE_wrapper_158__ap_ready),
    .PE_wrapper_158__ap_done(PE_wrapper_158__ap_done),
    .PE_wrapper_158__ap_idle(PE_wrapper_158__ap_idle),
    .PE_wrapper_159__ap_start(PE_wrapper_159__ap_start),
    .PE_wrapper_159__ap_ready(PE_wrapper_159__ap_ready),
    .PE_wrapper_159__ap_done(PE_wrapper_159__ap_done),
    .PE_wrapper_159__ap_idle(PE_wrapper_159__ap_idle),
    .PE_wrapper_160__ap_start(PE_wrapper_160__ap_start),
    .PE_wrapper_160__ap_ready(PE_wrapper_160__ap_ready),
    .PE_wrapper_160__ap_done(PE_wrapper_160__ap_done),
    .PE_wrapper_160__ap_idle(PE_wrapper_160__ap_idle),
    .PE_wrapper_161__ap_start(PE_wrapper_161__ap_start),
    .PE_wrapper_161__ap_ready(PE_wrapper_161__ap_ready),
    .PE_wrapper_161__ap_done(PE_wrapper_161__ap_done),
    .PE_wrapper_161__ap_idle(PE_wrapper_161__ap_idle),
    .PE_wrapper_162__ap_start(PE_wrapper_162__ap_start),
    .PE_wrapper_162__ap_ready(PE_wrapper_162__ap_ready),
    .PE_wrapper_162__ap_done(PE_wrapper_162__ap_done),
    .PE_wrapper_162__ap_idle(PE_wrapper_162__ap_idle),
    .PE_wrapper_163__ap_start(PE_wrapper_163__ap_start),
    .PE_wrapper_163__ap_ready(PE_wrapper_163__ap_ready),
    .PE_wrapper_163__ap_done(PE_wrapper_163__ap_done),
    .PE_wrapper_163__ap_idle(PE_wrapper_163__ap_idle),
    .PE_wrapper_164__ap_start(PE_wrapper_164__ap_start),
    .PE_wrapper_164__ap_ready(PE_wrapper_164__ap_ready),
    .PE_wrapper_164__ap_done(PE_wrapper_164__ap_done),
    .PE_wrapper_164__ap_idle(PE_wrapper_164__ap_idle),
    .PE_wrapper_165__ap_start(PE_wrapper_165__ap_start),
    .PE_wrapper_165__ap_ready(PE_wrapper_165__ap_ready),
    .PE_wrapper_165__ap_done(PE_wrapper_165__ap_done),
    .PE_wrapper_165__ap_idle(PE_wrapper_165__ap_idle),
    .PE_wrapper_166__ap_start(PE_wrapper_166__ap_start),
    .PE_wrapper_166__ap_ready(PE_wrapper_166__ap_ready),
    .PE_wrapper_166__ap_done(PE_wrapper_166__ap_done),
    .PE_wrapper_166__ap_idle(PE_wrapper_166__ap_idle),
    .PE_wrapper_167__ap_start(PE_wrapper_167__ap_start),
    .PE_wrapper_167__ap_ready(PE_wrapper_167__ap_ready),
    .PE_wrapper_167__ap_done(PE_wrapper_167__ap_done),
    .PE_wrapper_167__ap_idle(PE_wrapper_167__ap_idle),
    .PE_wrapper_168__ap_start(PE_wrapper_168__ap_start),
    .PE_wrapper_168__ap_ready(PE_wrapper_168__ap_ready),
    .PE_wrapper_168__ap_done(PE_wrapper_168__ap_done),
    .PE_wrapper_168__ap_idle(PE_wrapper_168__ap_idle),
    .PE_wrapper_169__ap_start(PE_wrapper_169__ap_start),
    .PE_wrapper_169__ap_ready(PE_wrapper_169__ap_ready),
    .PE_wrapper_169__ap_done(PE_wrapper_169__ap_done),
    .PE_wrapper_169__ap_idle(PE_wrapper_169__ap_idle),
    .PE_wrapper_170__ap_start(PE_wrapper_170__ap_start),
    .PE_wrapper_170__ap_ready(PE_wrapper_170__ap_ready),
    .PE_wrapper_170__ap_done(PE_wrapper_170__ap_done),
    .PE_wrapper_170__ap_idle(PE_wrapper_170__ap_idle),
    .PE_wrapper_171__ap_start(PE_wrapper_171__ap_start),
    .PE_wrapper_171__ap_ready(PE_wrapper_171__ap_ready),
    .PE_wrapper_171__ap_done(PE_wrapper_171__ap_done),
    .PE_wrapper_171__ap_idle(PE_wrapper_171__ap_idle),
    .PE_wrapper_172__ap_start(PE_wrapper_172__ap_start),
    .PE_wrapper_172__ap_ready(PE_wrapper_172__ap_ready),
    .PE_wrapper_172__ap_done(PE_wrapper_172__ap_done),
    .PE_wrapper_172__ap_idle(PE_wrapper_172__ap_idle),
    .PE_wrapper_173__ap_start(PE_wrapper_173__ap_start),
    .PE_wrapper_173__ap_ready(PE_wrapper_173__ap_ready),
    .PE_wrapper_173__ap_done(PE_wrapper_173__ap_done),
    .PE_wrapper_173__ap_idle(PE_wrapper_173__ap_idle),
    .PE_wrapper_174__ap_start(PE_wrapper_174__ap_start),
    .PE_wrapper_174__ap_ready(PE_wrapper_174__ap_ready),
    .PE_wrapper_174__ap_done(PE_wrapper_174__ap_done),
    .PE_wrapper_174__ap_idle(PE_wrapper_174__ap_idle),
    .PE_wrapper_175__ap_start(PE_wrapper_175__ap_start),
    .PE_wrapper_175__ap_ready(PE_wrapper_175__ap_ready),
    .PE_wrapper_175__ap_done(PE_wrapper_175__ap_done),
    .PE_wrapper_175__ap_idle(PE_wrapper_175__ap_idle),
    .PE_wrapper_176__ap_start(PE_wrapper_176__ap_start),
    .PE_wrapper_176__ap_ready(PE_wrapper_176__ap_ready),
    .PE_wrapper_176__ap_done(PE_wrapper_176__ap_done),
    .PE_wrapper_176__ap_idle(PE_wrapper_176__ap_idle),
    .PE_wrapper_177__ap_start(PE_wrapper_177__ap_start),
    .PE_wrapper_177__ap_ready(PE_wrapper_177__ap_ready),
    .PE_wrapper_177__ap_done(PE_wrapper_177__ap_done),
    .PE_wrapper_177__ap_idle(PE_wrapper_177__ap_idle),
    .PE_wrapper_178__ap_start(PE_wrapper_178__ap_start),
    .PE_wrapper_178__ap_ready(PE_wrapper_178__ap_ready),
    .PE_wrapper_178__ap_done(PE_wrapper_178__ap_done),
    .PE_wrapper_178__ap_idle(PE_wrapper_178__ap_idle),
    .PE_wrapper_179__ap_start(PE_wrapper_179__ap_start),
    .PE_wrapper_179__ap_ready(PE_wrapper_179__ap_ready),
    .PE_wrapper_179__ap_done(PE_wrapper_179__ap_done),
    .PE_wrapper_179__ap_idle(PE_wrapper_179__ap_idle),
    .PE_wrapper_180__ap_start(PE_wrapper_180__ap_start),
    .PE_wrapper_180__ap_ready(PE_wrapper_180__ap_ready),
    .PE_wrapper_180__ap_done(PE_wrapper_180__ap_done),
    .PE_wrapper_180__ap_idle(PE_wrapper_180__ap_idle),
    .PE_wrapper_181__ap_start(PE_wrapper_181__ap_start),
    .PE_wrapper_181__ap_ready(PE_wrapper_181__ap_ready),
    .PE_wrapper_181__ap_done(PE_wrapper_181__ap_done),
    .PE_wrapper_181__ap_idle(PE_wrapper_181__ap_idle),
    .PE_wrapper_182__ap_start(PE_wrapper_182__ap_start),
    .PE_wrapper_182__ap_ready(PE_wrapper_182__ap_ready),
    .PE_wrapper_182__ap_done(PE_wrapper_182__ap_done),
    .PE_wrapper_182__ap_idle(PE_wrapper_182__ap_idle),
    .PE_wrapper_183__ap_start(PE_wrapper_183__ap_start),
    .PE_wrapper_183__ap_ready(PE_wrapper_183__ap_ready),
    .PE_wrapper_183__ap_done(PE_wrapper_183__ap_done),
    .PE_wrapper_183__ap_idle(PE_wrapper_183__ap_idle),
    .PE_wrapper_184__ap_start(PE_wrapper_184__ap_start),
    .PE_wrapper_184__ap_ready(PE_wrapper_184__ap_ready),
    .PE_wrapper_184__ap_done(PE_wrapper_184__ap_done),
    .PE_wrapper_184__ap_idle(PE_wrapper_184__ap_idle),
    .PE_wrapper_185__ap_start(PE_wrapper_185__ap_start),
    .PE_wrapper_185__ap_ready(PE_wrapper_185__ap_ready),
    .PE_wrapper_185__ap_done(PE_wrapper_185__ap_done),
    .PE_wrapper_185__ap_idle(PE_wrapper_185__ap_idle),
    .PE_wrapper_186__ap_start(PE_wrapper_186__ap_start),
    .PE_wrapper_186__ap_ready(PE_wrapper_186__ap_ready),
    .PE_wrapper_186__ap_done(PE_wrapper_186__ap_done),
    .PE_wrapper_186__ap_idle(PE_wrapper_186__ap_idle),
    .PE_wrapper_187__ap_start(PE_wrapper_187__ap_start),
    .PE_wrapper_187__ap_ready(PE_wrapper_187__ap_ready),
    .PE_wrapper_187__ap_done(PE_wrapper_187__ap_done),
    .PE_wrapper_187__ap_idle(PE_wrapper_187__ap_idle),
    .PE_wrapper_188__ap_start(PE_wrapper_188__ap_start),
    .PE_wrapper_188__ap_ready(PE_wrapper_188__ap_ready),
    .PE_wrapper_188__ap_done(PE_wrapper_188__ap_done),
    .PE_wrapper_188__ap_idle(PE_wrapper_188__ap_idle),
    .PE_wrapper_189__ap_start(PE_wrapper_189__ap_start),
    .PE_wrapper_189__ap_ready(PE_wrapper_189__ap_ready),
    .PE_wrapper_189__ap_done(PE_wrapper_189__ap_done),
    .PE_wrapper_189__ap_idle(PE_wrapper_189__ap_idle),
    .PE_wrapper_190__ap_start(PE_wrapper_190__ap_start),
    .PE_wrapper_190__ap_ready(PE_wrapper_190__ap_ready),
    .PE_wrapper_190__ap_done(PE_wrapper_190__ap_done),
    .PE_wrapper_190__ap_idle(PE_wrapper_190__ap_idle),
    .PE_wrapper_191__ap_start(PE_wrapper_191__ap_start),
    .PE_wrapper_191__ap_ready(PE_wrapper_191__ap_ready),
    .PE_wrapper_191__ap_done(PE_wrapper_191__ap_done),
    .PE_wrapper_191__ap_idle(PE_wrapper_191__ap_idle),
    .PE_wrapper_192__ap_start(PE_wrapper_192__ap_start),
    .PE_wrapper_192__ap_ready(PE_wrapper_192__ap_ready),
    .PE_wrapper_192__ap_done(PE_wrapper_192__ap_done),
    .PE_wrapper_192__ap_idle(PE_wrapper_192__ap_idle),
    .PE_wrapper_193__ap_start(PE_wrapper_193__ap_start),
    .PE_wrapper_193__ap_ready(PE_wrapper_193__ap_ready),
    .PE_wrapper_193__ap_done(PE_wrapper_193__ap_done),
    .PE_wrapper_193__ap_idle(PE_wrapper_193__ap_idle),
    .PE_wrapper_194__ap_start(PE_wrapper_194__ap_start),
    .PE_wrapper_194__ap_ready(PE_wrapper_194__ap_ready),
    .PE_wrapper_194__ap_done(PE_wrapper_194__ap_done),
    .PE_wrapper_194__ap_idle(PE_wrapper_194__ap_idle),
    .PE_wrapper_195__ap_start(PE_wrapper_195__ap_start),
    .PE_wrapper_195__ap_ready(PE_wrapper_195__ap_ready),
    .PE_wrapper_195__ap_done(PE_wrapper_195__ap_done),
    .PE_wrapper_195__ap_idle(PE_wrapper_195__ap_idle),
    .PE_wrapper_196__ap_start(PE_wrapper_196__ap_start),
    .PE_wrapper_196__ap_ready(PE_wrapper_196__ap_ready),
    .PE_wrapper_196__ap_done(PE_wrapper_196__ap_done),
    .PE_wrapper_196__ap_idle(PE_wrapper_196__ap_idle),
    .PE_wrapper_197__ap_start(PE_wrapper_197__ap_start),
    .PE_wrapper_197__ap_ready(PE_wrapper_197__ap_ready),
    .PE_wrapper_197__ap_done(PE_wrapper_197__ap_done),
    .PE_wrapper_197__ap_idle(PE_wrapper_197__ap_idle),
    .PE_wrapper_198__ap_start(PE_wrapper_198__ap_start),
    .PE_wrapper_198__ap_ready(PE_wrapper_198__ap_ready),
    .PE_wrapper_198__ap_done(PE_wrapper_198__ap_done),
    .PE_wrapper_198__ap_idle(PE_wrapper_198__ap_idle),
    .PE_wrapper_199__ap_start(PE_wrapper_199__ap_start),
    .PE_wrapper_199__ap_ready(PE_wrapper_199__ap_ready),
    .PE_wrapper_199__ap_done(PE_wrapper_199__ap_done),
    .PE_wrapper_199__ap_idle(PE_wrapper_199__ap_idle),
    .PE_wrapper_200__ap_start(PE_wrapper_200__ap_start),
    .PE_wrapper_200__ap_ready(PE_wrapper_200__ap_ready),
    .PE_wrapper_200__ap_done(PE_wrapper_200__ap_done),
    .PE_wrapper_200__ap_idle(PE_wrapper_200__ap_idle),
    .PE_wrapper_201__ap_start(PE_wrapper_201__ap_start),
    .PE_wrapper_201__ap_ready(PE_wrapper_201__ap_ready),
    .PE_wrapper_201__ap_done(PE_wrapper_201__ap_done),
    .PE_wrapper_201__ap_idle(PE_wrapper_201__ap_idle),
    .PE_wrapper_202__ap_start(PE_wrapper_202__ap_start),
    .PE_wrapper_202__ap_ready(PE_wrapper_202__ap_ready),
    .PE_wrapper_202__ap_done(PE_wrapper_202__ap_done),
    .PE_wrapper_202__ap_idle(PE_wrapper_202__ap_idle),
    .PE_wrapper_203__ap_start(PE_wrapper_203__ap_start),
    .PE_wrapper_203__ap_ready(PE_wrapper_203__ap_ready),
    .PE_wrapper_203__ap_done(PE_wrapper_203__ap_done),
    .PE_wrapper_203__ap_idle(PE_wrapper_203__ap_idle),
    .PE_wrapper_204__ap_start(PE_wrapper_204__ap_start),
    .PE_wrapper_204__ap_ready(PE_wrapper_204__ap_ready),
    .PE_wrapper_204__ap_done(PE_wrapper_204__ap_done),
    .PE_wrapper_204__ap_idle(PE_wrapper_204__ap_idle),
    .PE_wrapper_205__ap_start(PE_wrapper_205__ap_start),
    .PE_wrapper_205__ap_ready(PE_wrapper_205__ap_ready),
    .PE_wrapper_205__ap_done(PE_wrapper_205__ap_done),
    .PE_wrapper_205__ap_idle(PE_wrapper_205__ap_idle),
    .PE_wrapper_206__ap_start(PE_wrapper_206__ap_start),
    .PE_wrapper_206__ap_ready(PE_wrapper_206__ap_ready),
    .PE_wrapper_206__ap_done(PE_wrapper_206__ap_done),
    .PE_wrapper_206__ap_idle(PE_wrapper_206__ap_idle),
    .PE_wrapper_207__ap_start(PE_wrapper_207__ap_start),
    .PE_wrapper_207__ap_ready(PE_wrapper_207__ap_ready),
    .PE_wrapper_207__ap_done(PE_wrapper_207__ap_done),
    .PE_wrapper_207__ap_idle(PE_wrapper_207__ap_idle),
    .PE_wrapper_208__ap_start(PE_wrapper_208__ap_start),
    .PE_wrapper_208__ap_ready(PE_wrapper_208__ap_ready),
    .PE_wrapper_208__ap_done(PE_wrapper_208__ap_done),
    .PE_wrapper_208__ap_idle(PE_wrapper_208__ap_idle),
    .PE_wrapper_209__ap_start(PE_wrapper_209__ap_start),
    .PE_wrapper_209__ap_ready(PE_wrapper_209__ap_ready),
    .PE_wrapper_209__ap_done(PE_wrapper_209__ap_done),
    .PE_wrapper_209__ap_idle(PE_wrapper_209__ap_idle),
    .PE_wrapper_210__ap_start(PE_wrapper_210__ap_start),
    .PE_wrapper_210__ap_ready(PE_wrapper_210__ap_ready),
    .PE_wrapper_210__ap_done(PE_wrapper_210__ap_done),
    .PE_wrapper_210__ap_idle(PE_wrapper_210__ap_idle),
    .PE_wrapper_211__ap_start(PE_wrapper_211__ap_start),
    .PE_wrapper_211__ap_ready(PE_wrapper_211__ap_ready),
    .PE_wrapper_211__ap_done(PE_wrapper_211__ap_done),
    .PE_wrapper_211__ap_idle(PE_wrapper_211__ap_idle),
    .PE_wrapper_212__ap_start(PE_wrapper_212__ap_start),
    .PE_wrapper_212__ap_ready(PE_wrapper_212__ap_ready),
    .PE_wrapper_212__ap_done(PE_wrapper_212__ap_done),
    .PE_wrapper_212__ap_idle(PE_wrapper_212__ap_idle),
    .PE_wrapper_213__ap_start(PE_wrapper_213__ap_start),
    .PE_wrapper_213__ap_ready(PE_wrapper_213__ap_ready),
    .PE_wrapper_213__ap_done(PE_wrapper_213__ap_done),
    .PE_wrapper_213__ap_idle(PE_wrapper_213__ap_idle),
    .PE_wrapper_214__ap_start(PE_wrapper_214__ap_start),
    .PE_wrapper_214__ap_ready(PE_wrapper_214__ap_ready),
    .PE_wrapper_214__ap_done(PE_wrapper_214__ap_done),
    .PE_wrapper_214__ap_idle(PE_wrapper_214__ap_idle),
    .PE_wrapper_215__ap_start(PE_wrapper_215__ap_start),
    .PE_wrapper_215__ap_ready(PE_wrapper_215__ap_ready),
    .PE_wrapper_215__ap_done(PE_wrapper_215__ap_done),
    .PE_wrapper_215__ap_idle(PE_wrapper_215__ap_idle),
    .PE_wrapper_216__ap_start(PE_wrapper_216__ap_start),
    .PE_wrapper_216__ap_ready(PE_wrapper_216__ap_ready),
    .PE_wrapper_216__ap_done(PE_wrapper_216__ap_done),
    .PE_wrapper_216__ap_idle(PE_wrapper_216__ap_idle),
    .PE_wrapper_217__ap_start(PE_wrapper_217__ap_start),
    .PE_wrapper_217__ap_ready(PE_wrapper_217__ap_ready),
    .PE_wrapper_217__ap_done(PE_wrapper_217__ap_done),
    .PE_wrapper_217__ap_idle(PE_wrapper_217__ap_idle),
    .PE_wrapper_218__ap_start(PE_wrapper_218__ap_start),
    .PE_wrapper_218__ap_ready(PE_wrapper_218__ap_ready),
    .PE_wrapper_218__ap_done(PE_wrapper_218__ap_done),
    .PE_wrapper_218__ap_idle(PE_wrapper_218__ap_idle),
    .PE_wrapper_219__ap_start(PE_wrapper_219__ap_start),
    .PE_wrapper_219__ap_ready(PE_wrapper_219__ap_ready),
    .PE_wrapper_219__ap_done(PE_wrapper_219__ap_done),
    .PE_wrapper_219__ap_idle(PE_wrapper_219__ap_idle),
    .PE_wrapper_220__ap_start(PE_wrapper_220__ap_start),
    .PE_wrapper_220__ap_ready(PE_wrapper_220__ap_ready),
    .PE_wrapper_220__ap_done(PE_wrapper_220__ap_done),
    .PE_wrapper_220__ap_idle(PE_wrapper_220__ap_idle),
    .PE_wrapper_221__ap_start(PE_wrapper_221__ap_start),
    .PE_wrapper_221__ap_ready(PE_wrapper_221__ap_ready),
    .PE_wrapper_221__ap_done(PE_wrapper_221__ap_done),
    .PE_wrapper_221__ap_idle(PE_wrapper_221__ap_idle),
    .PE_wrapper_222__ap_start(PE_wrapper_222__ap_start),
    .PE_wrapper_222__ap_ready(PE_wrapper_222__ap_ready),
    .PE_wrapper_222__ap_done(PE_wrapper_222__ap_done),
    .PE_wrapper_222__ap_idle(PE_wrapper_222__ap_idle),
    .PE_wrapper_223__ap_start(PE_wrapper_223__ap_start),
    .PE_wrapper_223__ap_ready(PE_wrapper_223__ap_ready),
    .PE_wrapper_223__ap_done(PE_wrapper_223__ap_done),
    .PE_wrapper_223__ap_idle(PE_wrapper_223__ap_idle),
    .PE_wrapper_224__ap_start(PE_wrapper_224__ap_start),
    .PE_wrapper_224__ap_ready(PE_wrapper_224__ap_ready),
    .PE_wrapper_224__ap_done(PE_wrapper_224__ap_done),
    .PE_wrapper_224__ap_idle(PE_wrapper_224__ap_idle),
    .PE_wrapper_225__ap_start(PE_wrapper_225__ap_start),
    .PE_wrapper_225__ap_ready(PE_wrapper_225__ap_ready),
    .PE_wrapper_225__ap_done(PE_wrapper_225__ap_done),
    .PE_wrapper_225__ap_idle(PE_wrapper_225__ap_idle),
    .PE_wrapper_226__ap_start(PE_wrapper_226__ap_start),
    .PE_wrapper_226__ap_ready(PE_wrapper_226__ap_ready),
    .PE_wrapper_226__ap_done(PE_wrapper_226__ap_done),
    .PE_wrapper_226__ap_idle(PE_wrapper_226__ap_idle),
    .PE_wrapper_227__ap_start(PE_wrapper_227__ap_start),
    .PE_wrapper_227__ap_ready(PE_wrapper_227__ap_ready),
    .PE_wrapper_227__ap_done(PE_wrapper_227__ap_done),
    .PE_wrapper_227__ap_idle(PE_wrapper_227__ap_idle),
    .PE_wrapper_228__ap_start(PE_wrapper_228__ap_start),
    .PE_wrapper_228__ap_ready(PE_wrapper_228__ap_ready),
    .PE_wrapper_228__ap_done(PE_wrapper_228__ap_done),
    .PE_wrapper_228__ap_idle(PE_wrapper_228__ap_idle),
    .PE_wrapper_229__ap_start(PE_wrapper_229__ap_start),
    .PE_wrapper_229__ap_ready(PE_wrapper_229__ap_ready),
    .PE_wrapper_229__ap_done(PE_wrapper_229__ap_done),
    .PE_wrapper_229__ap_idle(PE_wrapper_229__ap_idle),
    .PE_wrapper_230__ap_start(PE_wrapper_230__ap_start),
    .PE_wrapper_230__ap_ready(PE_wrapper_230__ap_ready),
    .PE_wrapper_230__ap_done(PE_wrapper_230__ap_done),
    .PE_wrapper_230__ap_idle(PE_wrapper_230__ap_idle),
    .PE_wrapper_231__ap_start(PE_wrapper_231__ap_start),
    .PE_wrapper_231__ap_ready(PE_wrapper_231__ap_ready),
    .PE_wrapper_231__ap_done(PE_wrapper_231__ap_done),
    .PE_wrapper_231__ap_idle(PE_wrapper_231__ap_idle),
    .PE_wrapper_232__ap_start(PE_wrapper_232__ap_start),
    .PE_wrapper_232__ap_ready(PE_wrapper_232__ap_ready),
    .PE_wrapper_232__ap_done(PE_wrapper_232__ap_done),
    .PE_wrapper_232__ap_idle(PE_wrapper_232__ap_idle),
    .PE_wrapper_233__ap_start(PE_wrapper_233__ap_start),
    .PE_wrapper_233__ap_ready(PE_wrapper_233__ap_ready),
    .PE_wrapper_233__ap_done(PE_wrapper_233__ap_done),
    .PE_wrapper_233__ap_idle(PE_wrapper_233__ap_idle),
    .PE_wrapper_234__ap_start(PE_wrapper_234__ap_start),
    .PE_wrapper_234__ap_ready(PE_wrapper_234__ap_ready),
    .PE_wrapper_234__ap_done(PE_wrapper_234__ap_done),
    .PE_wrapper_234__ap_idle(PE_wrapper_234__ap_idle),
    .PE_wrapper_235__ap_start(PE_wrapper_235__ap_start),
    .PE_wrapper_235__ap_ready(PE_wrapper_235__ap_ready),
    .PE_wrapper_235__ap_done(PE_wrapper_235__ap_done),
    .PE_wrapper_235__ap_idle(PE_wrapper_235__ap_idle),
    .PE_wrapper_236__ap_start(PE_wrapper_236__ap_start),
    .PE_wrapper_236__ap_ready(PE_wrapper_236__ap_ready),
    .PE_wrapper_236__ap_done(PE_wrapper_236__ap_done),
    .PE_wrapper_236__ap_idle(PE_wrapper_236__ap_idle),
    .PE_wrapper_237__ap_start(PE_wrapper_237__ap_start),
    .PE_wrapper_237__ap_ready(PE_wrapper_237__ap_ready),
    .PE_wrapper_237__ap_done(PE_wrapper_237__ap_done),
    .PE_wrapper_237__ap_idle(PE_wrapper_237__ap_idle),
    .PE_wrapper_238__ap_start(PE_wrapper_238__ap_start),
    .PE_wrapper_238__ap_ready(PE_wrapper_238__ap_ready),
    .PE_wrapper_238__ap_done(PE_wrapper_238__ap_done),
    .PE_wrapper_238__ap_idle(PE_wrapper_238__ap_idle),
    .PE_wrapper_239__ap_start(PE_wrapper_239__ap_start),
    .PE_wrapper_239__ap_ready(PE_wrapper_239__ap_ready),
    .PE_wrapper_239__ap_done(PE_wrapper_239__ap_done),
    .PE_wrapper_239__ap_idle(PE_wrapper_239__ap_idle),
    .PE_wrapper_240__ap_start(PE_wrapper_240__ap_start),
    .PE_wrapper_240__ap_ready(PE_wrapper_240__ap_ready),
    .PE_wrapper_240__ap_done(PE_wrapper_240__ap_done),
    .PE_wrapper_240__ap_idle(PE_wrapper_240__ap_idle),
    .PE_wrapper_241__ap_start(PE_wrapper_241__ap_start),
    .PE_wrapper_241__ap_ready(PE_wrapper_241__ap_ready),
    .PE_wrapper_241__ap_done(PE_wrapper_241__ap_done),
    .PE_wrapper_241__ap_idle(PE_wrapper_241__ap_idle),
    .PE_wrapper_242__ap_start(PE_wrapper_242__ap_start),
    .PE_wrapper_242__ap_ready(PE_wrapper_242__ap_ready),
    .PE_wrapper_242__ap_done(PE_wrapper_242__ap_done),
    .PE_wrapper_242__ap_idle(PE_wrapper_242__ap_idle),
    .PE_wrapper_243__ap_start(PE_wrapper_243__ap_start),
    .PE_wrapper_243__ap_ready(PE_wrapper_243__ap_ready),
    .PE_wrapper_243__ap_done(PE_wrapper_243__ap_done),
    .PE_wrapper_243__ap_idle(PE_wrapper_243__ap_idle),
    .PE_wrapper_244__ap_start(PE_wrapper_244__ap_start),
    .PE_wrapper_244__ap_ready(PE_wrapper_244__ap_ready),
    .PE_wrapper_244__ap_done(PE_wrapper_244__ap_done),
    .PE_wrapper_244__ap_idle(PE_wrapper_244__ap_idle),
    .PE_wrapper_245__ap_start(PE_wrapper_245__ap_start),
    .PE_wrapper_245__ap_ready(PE_wrapper_245__ap_ready),
    .PE_wrapper_245__ap_done(PE_wrapper_245__ap_done),
    .PE_wrapper_245__ap_idle(PE_wrapper_245__ap_idle),
    .PE_wrapper_246__ap_start(PE_wrapper_246__ap_start),
    .PE_wrapper_246__ap_ready(PE_wrapper_246__ap_ready),
    .PE_wrapper_246__ap_done(PE_wrapper_246__ap_done),
    .PE_wrapper_246__ap_idle(PE_wrapper_246__ap_idle),
    .PE_wrapper_247__ap_start(PE_wrapper_247__ap_start),
    .PE_wrapper_247__ap_ready(PE_wrapper_247__ap_ready),
    .PE_wrapper_247__ap_done(PE_wrapper_247__ap_done),
    .PE_wrapper_247__ap_idle(PE_wrapper_247__ap_idle),
    .PE_wrapper_248__ap_start(PE_wrapper_248__ap_start),
    .PE_wrapper_248__ap_ready(PE_wrapper_248__ap_ready),
    .PE_wrapper_248__ap_done(PE_wrapper_248__ap_done),
    .PE_wrapper_248__ap_idle(PE_wrapper_248__ap_idle),
    .PE_wrapper_249__ap_start(PE_wrapper_249__ap_start),
    .PE_wrapper_249__ap_ready(PE_wrapper_249__ap_ready),
    .PE_wrapper_249__ap_done(PE_wrapper_249__ap_done),
    .PE_wrapper_249__ap_idle(PE_wrapper_249__ap_idle),
    .PE_wrapper_250__ap_start(PE_wrapper_250__ap_start),
    .PE_wrapper_250__ap_ready(PE_wrapper_250__ap_ready),
    .PE_wrapper_250__ap_done(PE_wrapper_250__ap_done),
    .PE_wrapper_250__ap_idle(PE_wrapper_250__ap_idle),
    .PE_wrapper_251__ap_start(PE_wrapper_251__ap_start),
    .PE_wrapper_251__ap_ready(PE_wrapper_251__ap_ready),
    .PE_wrapper_251__ap_done(PE_wrapper_251__ap_done),
    .PE_wrapper_251__ap_idle(PE_wrapper_251__ap_idle),
    .PE_wrapper_252__ap_start(PE_wrapper_252__ap_start),
    .PE_wrapper_252__ap_ready(PE_wrapper_252__ap_ready),
    .PE_wrapper_252__ap_done(PE_wrapper_252__ap_done),
    .PE_wrapper_252__ap_idle(PE_wrapper_252__ap_idle),
    .PE_wrapper_253__ap_start(PE_wrapper_253__ap_start),
    .PE_wrapper_253__ap_ready(PE_wrapper_253__ap_ready),
    .PE_wrapper_253__ap_done(PE_wrapper_253__ap_done),
    .PE_wrapper_253__ap_idle(PE_wrapper_253__ap_idle),
    .PE_wrapper_254__ap_start(PE_wrapper_254__ap_start),
    .PE_wrapper_254__ap_ready(PE_wrapper_254__ap_ready),
    .PE_wrapper_254__ap_done(PE_wrapper_254__ap_done),
    .PE_wrapper_254__ap_idle(PE_wrapper_254__ap_idle),
    .PE_wrapper_255__ap_start(PE_wrapper_255__ap_start),
    .PE_wrapper_255__ap_ready(PE_wrapper_255__ap_ready),
    .PE_wrapper_255__ap_done(PE_wrapper_255__ap_done),
    .PE_wrapper_255__ap_idle(PE_wrapper_255__ap_idle),
    .PE_wrapper_256__ap_start(PE_wrapper_256__ap_start),
    .PE_wrapper_256__ap_ready(PE_wrapper_256__ap_ready),
    .PE_wrapper_256__ap_done(PE_wrapper_256__ap_done),
    .PE_wrapper_256__ap_idle(PE_wrapper_256__ap_idle),
    .PE_wrapper_257__ap_start(PE_wrapper_257__ap_start),
    .PE_wrapper_257__ap_ready(PE_wrapper_257__ap_ready),
    .PE_wrapper_257__ap_done(PE_wrapper_257__ap_done),
    .PE_wrapper_257__ap_idle(PE_wrapper_257__ap_idle),
    .PE_wrapper_258__ap_start(PE_wrapper_258__ap_start),
    .PE_wrapper_258__ap_ready(PE_wrapper_258__ap_ready),
    .PE_wrapper_258__ap_done(PE_wrapper_258__ap_done),
    .PE_wrapper_258__ap_idle(PE_wrapper_258__ap_idle),
    .PE_wrapper_259__ap_start(PE_wrapper_259__ap_start),
    .PE_wrapper_259__ap_ready(PE_wrapper_259__ap_ready),
    .PE_wrapper_259__ap_done(PE_wrapper_259__ap_done),
    .PE_wrapper_259__ap_idle(PE_wrapper_259__ap_idle),
    .PE_wrapper_260__ap_start(PE_wrapper_260__ap_start),
    .PE_wrapper_260__ap_ready(PE_wrapper_260__ap_ready),
    .PE_wrapper_260__ap_done(PE_wrapper_260__ap_done),
    .PE_wrapper_260__ap_idle(PE_wrapper_260__ap_idle),
    .PE_wrapper_261__ap_start(PE_wrapper_261__ap_start),
    .PE_wrapper_261__ap_ready(PE_wrapper_261__ap_ready),
    .PE_wrapper_261__ap_done(PE_wrapper_261__ap_done),
    .PE_wrapper_261__ap_idle(PE_wrapper_261__ap_idle),
    .PE_wrapper_262__ap_start(PE_wrapper_262__ap_start),
    .PE_wrapper_262__ap_ready(PE_wrapper_262__ap_ready),
    .PE_wrapper_262__ap_done(PE_wrapper_262__ap_done),
    .PE_wrapper_262__ap_idle(PE_wrapper_262__ap_idle),
    .PE_wrapper_263__ap_start(PE_wrapper_263__ap_start),
    .PE_wrapper_263__ap_ready(PE_wrapper_263__ap_ready),
    .PE_wrapper_263__ap_done(PE_wrapper_263__ap_done),
    .PE_wrapper_263__ap_idle(PE_wrapper_263__ap_idle),
    .PE_wrapper_264__ap_start(PE_wrapper_264__ap_start),
    .PE_wrapper_264__ap_ready(PE_wrapper_264__ap_ready),
    .PE_wrapper_264__ap_done(PE_wrapper_264__ap_done),
    .PE_wrapper_264__ap_idle(PE_wrapper_264__ap_idle),
    .PE_wrapper_265__ap_start(PE_wrapper_265__ap_start),
    .PE_wrapper_265__ap_ready(PE_wrapper_265__ap_ready),
    .PE_wrapper_265__ap_done(PE_wrapper_265__ap_done),
    .PE_wrapper_265__ap_idle(PE_wrapper_265__ap_idle),
    .PE_wrapper_266__ap_start(PE_wrapper_266__ap_start),
    .PE_wrapper_266__ap_ready(PE_wrapper_266__ap_ready),
    .PE_wrapper_266__ap_done(PE_wrapper_266__ap_done),
    .PE_wrapper_266__ap_idle(PE_wrapper_266__ap_idle),
    .PE_wrapper_267__ap_start(PE_wrapper_267__ap_start),
    .PE_wrapper_267__ap_ready(PE_wrapper_267__ap_ready),
    .PE_wrapper_267__ap_done(PE_wrapper_267__ap_done),
    .PE_wrapper_267__ap_idle(PE_wrapper_267__ap_idle),
    .PE_wrapper_268__ap_start(PE_wrapper_268__ap_start),
    .PE_wrapper_268__ap_ready(PE_wrapper_268__ap_ready),
    .PE_wrapper_268__ap_done(PE_wrapper_268__ap_done),
    .PE_wrapper_268__ap_idle(PE_wrapper_268__ap_idle),
    .PE_wrapper_269__ap_start(PE_wrapper_269__ap_start),
    .PE_wrapper_269__ap_ready(PE_wrapper_269__ap_ready),
    .PE_wrapper_269__ap_done(PE_wrapper_269__ap_done),
    .PE_wrapper_269__ap_idle(PE_wrapper_269__ap_idle),
    .PE_wrapper_270__ap_start(PE_wrapper_270__ap_start),
    .PE_wrapper_270__ap_ready(PE_wrapper_270__ap_ready),
    .PE_wrapper_270__ap_done(PE_wrapper_270__ap_done),
    .PE_wrapper_270__ap_idle(PE_wrapper_270__ap_idle),
    .PE_wrapper_271__ap_start(PE_wrapper_271__ap_start),
    .PE_wrapper_271__ap_ready(PE_wrapper_271__ap_ready),
    .PE_wrapper_271__ap_done(PE_wrapper_271__ap_done),
    .PE_wrapper_271__ap_idle(PE_wrapper_271__ap_idle),
    .PE_wrapper_272__ap_start(PE_wrapper_272__ap_start),
    .PE_wrapper_272__ap_ready(PE_wrapper_272__ap_ready),
    .PE_wrapper_272__ap_done(PE_wrapper_272__ap_done),
    .PE_wrapper_272__ap_idle(PE_wrapper_272__ap_idle),
    .PE_wrapper_273__ap_start(PE_wrapper_273__ap_start),
    .PE_wrapper_273__ap_ready(PE_wrapper_273__ap_ready),
    .PE_wrapper_273__ap_done(PE_wrapper_273__ap_done),
    .PE_wrapper_273__ap_idle(PE_wrapper_273__ap_idle),
    .PE_wrapper_274__ap_start(PE_wrapper_274__ap_start),
    .PE_wrapper_274__ap_ready(PE_wrapper_274__ap_ready),
    .PE_wrapper_274__ap_done(PE_wrapper_274__ap_done),
    .PE_wrapper_274__ap_idle(PE_wrapper_274__ap_idle),
    .PE_wrapper_275__ap_start(PE_wrapper_275__ap_start),
    .PE_wrapper_275__ap_ready(PE_wrapper_275__ap_ready),
    .PE_wrapper_275__ap_done(PE_wrapper_275__ap_done),
    .PE_wrapper_275__ap_idle(PE_wrapper_275__ap_idle),
    .PE_wrapper_276__ap_start(PE_wrapper_276__ap_start),
    .PE_wrapper_276__ap_ready(PE_wrapper_276__ap_ready),
    .PE_wrapper_276__ap_done(PE_wrapper_276__ap_done),
    .PE_wrapper_276__ap_idle(PE_wrapper_276__ap_idle),
    .PE_wrapper_277__ap_start(PE_wrapper_277__ap_start),
    .PE_wrapper_277__ap_ready(PE_wrapper_277__ap_ready),
    .PE_wrapper_277__ap_done(PE_wrapper_277__ap_done),
    .PE_wrapper_277__ap_idle(PE_wrapper_277__ap_idle),
    .PE_wrapper_278__ap_start(PE_wrapper_278__ap_start),
    .PE_wrapper_278__ap_ready(PE_wrapper_278__ap_ready),
    .PE_wrapper_278__ap_done(PE_wrapper_278__ap_done),
    .PE_wrapper_278__ap_idle(PE_wrapper_278__ap_idle),
    .PE_wrapper_279__ap_start(PE_wrapper_279__ap_start),
    .PE_wrapper_279__ap_ready(PE_wrapper_279__ap_ready),
    .PE_wrapper_279__ap_done(PE_wrapper_279__ap_done),
    .PE_wrapper_279__ap_idle(PE_wrapper_279__ap_idle),
    .PE_wrapper_280__ap_start(PE_wrapper_280__ap_start),
    .PE_wrapper_280__ap_ready(PE_wrapper_280__ap_ready),
    .PE_wrapper_280__ap_done(PE_wrapper_280__ap_done),
    .PE_wrapper_280__ap_idle(PE_wrapper_280__ap_idle),
    .PE_wrapper_281__ap_start(PE_wrapper_281__ap_start),
    .PE_wrapper_281__ap_ready(PE_wrapper_281__ap_ready),
    .PE_wrapper_281__ap_done(PE_wrapper_281__ap_done),
    .PE_wrapper_281__ap_idle(PE_wrapper_281__ap_idle),
    .PE_wrapper_282__ap_start(PE_wrapper_282__ap_start),
    .PE_wrapper_282__ap_ready(PE_wrapper_282__ap_ready),
    .PE_wrapper_282__ap_done(PE_wrapper_282__ap_done),
    .PE_wrapper_282__ap_idle(PE_wrapper_282__ap_idle),
    .PE_wrapper_283__ap_start(PE_wrapper_283__ap_start),
    .PE_wrapper_283__ap_ready(PE_wrapper_283__ap_ready),
    .PE_wrapper_283__ap_done(PE_wrapper_283__ap_done),
    .PE_wrapper_283__ap_idle(PE_wrapper_283__ap_idle),
    .PE_wrapper_284__ap_start(PE_wrapper_284__ap_start),
    .PE_wrapper_284__ap_ready(PE_wrapper_284__ap_ready),
    .PE_wrapper_284__ap_done(PE_wrapper_284__ap_done),
    .PE_wrapper_284__ap_idle(PE_wrapper_284__ap_idle),
    .PE_wrapper_285__ap_start(PE_wrapper_285__ap_start),
    .PE_wrapper_285__ap_ready(PE_wrapper_285__ap_ready),
    .PE_wrapper_285__ap_done(PE_wrapper_285__ap_done),
    .PE_wrapper_285__ap_idle(PE_wrapper_285__ap_idle),
    .PE_wrapper_286__ap_start(PE_wrapper_286__ap_start),
    .PE_wrapper_286__ap_ready(PE_wrapper_286__ap_ready),
    .PE_wrapper_286__ap_done(PE_wrapper_286__ap_done),
    .PE_wrapper_286__ap_idle(PE_wrapper_286__ap_idle),
    .PE_wrapper_287__ap_start(PE_wrapper_287__ap_start),
    .PE_wrapper_287__ap_ready(PE_wrapper_287__ap_ready),
    .PE_wrapper_287__ap_done(PE_wrapper_287__ap_done),
    .PE_wrapper_287__ap_idle(PE_wrapper_287__ap_idle),
    .PE_wrapper_288__ap_start(PE_wrapper_288__ap_start),
    .PE_wrapper_288__ap_ready(PE_wrapper_288__ap_ready),
    .PE_wrapper_288__ap_done(PE_wrapper_288__ap_done),
    .PE_wrapper_288__ap_idle(PE_wrapper_288__ap_idle),
    .PE_wrapper_289__ap_start(PE_wrapper_289__ap_start),
    .PE_wrapper_289__ap_ready(PE_wrapper_289__ap_ready),
    .PE_wrapper_289__ap_done(PE_wrapper_289__ap_done),
    .PE_wrapper_289__ap_idle(PE_wrapper_289__ap_idle),
    .PE_wrapper_290__ap_start(PE_wrapper_290__ap_start),
    .PE_wrapper_290__ap_ready(PE_wrapper_290__ap_ready),
    .PE_wrapper_290__ap_done(PE_wrapper_290__ap_done),
    .PE_wrapper_290__ap_idle(PE_wrapper_290__ap_idle),
    .PE_wrapper_291__ap_start(PE_wrapper_291__ap_start),
    .PE_wrapper_291__ap_ready(PE_wrapper_291__ap_ready),
    .PE_wrapper_291__ap_done(PE_wrapper_291__ap_done),
    .PE_wrapper_291__ap_idle(PE_wrapper_291__ap_idle),
    .PE_wrapper_292__ap_start(PE_wrapper_292__ap_start),
    .PE_wrapper_292__ap_ready(PE_wrapper_292__ap_ready),
    .PE_wrapper_292__ap_done(PE_wrapper_292__ap_done),
    .PE_wrapper_292__ap_idle(PE_wrapper_292__ap_idle),
    .PE_wrapper_293__ap_start(PE_wrapper_293__ap_start),
    .PE_wrapper_293__ap_ready(PE_wrapper_293__ap_ready),
    .PE_wrapper_293__ap_done(PE_wrapper_293__ap_done),
    .PE_wrapper_293__ap_idle(PE_wrapper_293__ap_idle),
    .PE_wrapper_294__ap_start(PE_wrapper_294__ap_start),
    .PE_wrapper_294__ap_ready(PE_wrapper_294__ap_ready),
    .PE_wrapper_294__ap_done(PE_wrapper_294__ap_done),
    .PE_wrapper_294__ap_idle(PE_wrapper_294__ap_idle),
    .PE_wrapper_295__ap_start(PE_wrapper_295__ap_start),
    .PE_wrapper_295__ap_ready(PE_wrapper_295__ap_ready),
    .PE_wrapper_295__ap_done(PE_wrapper_295__ap_done),
    .PE_wrapper_295__ap_idle(PE_wrapper_295__ap_idle),
    .PE_wrapper_296__ap_start(PE_wrapper_296__ap_start),
    .PE_wrapper_296__ap_ready(PE_wrapper_296__ap_ready),
    .PE_wrapper_296__ap_done(PE_wrapper_296__ap_done),
    .PE_wrapper_296__ap_idle(PE_wrapper_296__ap_idle),
    .PE_wrapper_297__ap_start(PE_wrapper_297__ap_start),
    .PE_wrapper_297__ap_ready(PE_wrapper_297__ap_ready),
    .PE_wrapper_297__ap_done(PE_wrapper_297__ap_done),
    .PE_wrapper_297__ap_idle(PE_wrapper_297__ap_idle),
    .PE_wrapper_298__ap_start(PE_wrapper_298__ap_start),
    .PE_wrapper_298__ap_ready(PE_wrapper_298__ap_ready),
    .PE_wrapper_298__ap_done(PE_wrapper_298__ap_done),
    .PE_wrapper_298__ap_idle(PE_wrapper_298__ap_idle),
    .PE_wrapper_299__ap_start(PE_wrapper_299__ap_start),
    .PE_wrapper_299__ap_ready(PE_wrapper_299__ap_ready),
    .PE_wrapper_299__ap_done(PE_wrapper_299__ap_done),
    .PE_wrapper_299__ap_idle(PE_wrapper_299__ap_idle),
    .PE_wrapper_300__ap_start(PE_wrapper_300__ap_start),
    .PE_wrapper_300__ap_ready(PE_wrapper_300__ap_ready),
    .PE_wrapper_300__ap_done(PE_wrapper_300__ap_done),
    .PE_wrapper_300__ap_idle(PE_wrapper_300__ap_idle),
    .PE_wrapper_301__ap_start(PE_wrapper_301__ap_start),
    .PE_wrapper_301__ap_ready(PE_wrapper_301__ap_ready),
    .PE_wrapper_301__ap_done(PE_wrapper_301__ap_done),
    .PE_wrapper_301__ap_idle(PE_wrapper_301__ap_idle),
    .PE_wrapper_302__ap_start(PE_wrapper_302__ap_start),
    .PE_wrapper_302__ap_ready(PE_wrapper_302__ap_ready),
    .PE_wrapper_302__ap_done(PE_wrapper_302__ap_done),
    .PE_wrapper_302__ap_idle(PE_wrapper_302__ap_idle),
    .PE_wrapper_303__ap_start(PE_wrapper_303__ap_start),
    .PE_wrapper_303__ap_ready(PE_wrapper_303__ap_ready),
    .PE_wrapper_303__ap_done(PE_wrapper_303__ap_done),
    .PE_wrapper_303__ap_idle(PE_wrapper_303__ap_idle),
    .PE_wrapper_304__ap_start(PE_wrapper_304__ap_start),
    .PE_wrapper_304__ap_ready(PE_wrapper_304__ap_ready),
    .PE_wrapper_304__ap_done(PE_wrapper_304__ap_done),
    .PE_wrapper_304__ap_idle(PE_wrapper_304__ap_idle),
    .PE_wrapper_305__ap_start(PE_wrapper_305__ap_start),
    .PE_wrapper_305__ap_ready(PE_wrapper_305__ap_ready),
    .PE_wrapper_305__ap_done(PE_wrapper_305__ap_done),
    .PE_wrapper_305__ap_idle(PE_wrapper_305__ap_idle)
  );

  assign ap_rst_n_inv = (~ap_rst_n);

endmodule

