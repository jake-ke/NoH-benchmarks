`timescale 1 ns / 1 ps
 
(* CORE_GENERATION_INFO = "Knn_Knn,hls_ip_2023_2_2,{HLS_INPUT_TYPE=cxx,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=0,HLS_INPUT_PART=xcvh1582-vsva3697-2MP-e-S,HLS_INPUT_CLOCK=3.330000,HLS_INPUT_ARCH=others,HLS_SYN_CLOCK=1.000000,HLS_SYN_LAT=0,HLS_SYN_TPT=none,HLS_SYN_MEM=0,HLS_SYN_DSP=0,HLS_SYN_FF=3956,HLS_SYN_LUT=7208,HLS_VERSION=2023_2_2}" *)module __rs_Knn_aux #(
    parameter C_S_AXI_CONTROL_DATA_WIDTH  = 32,
    parameter C_S_AXI_CONTROL_ADDR_WIDTH  = 10,
    parameter C_S_AXI_DATA_WIDTH          = 32,
    parameter C_S_AXI_CONTROL_WSTRB_WIDTH = 4,
    parameter C_S_AXI_WSTRB_WIDTH         = 4
) (
    input wire                                           s_axi_control_AWVALID,
    output wire                                          s_axi_control_AWREADY,
    input wire  [    (C_S_AXI_CONTROL_ADDR_WIDTH - 1):0] s_axi_control_AWADDR,
    input wire                                           s_axi_control_WVALID,
    output wire                                          s_axi_control_WREADY,
    input wire  [    (C_S_AXI_CONTROL_DATA_WIDTH - 1):0] s_axi_control_WDATA,
    input wire  [   (C_S_AXI_CONTROL_WSTRB_WIDTH - 1):0] s_axi_control_WSTRB,
    input wire                                           s_axi_control_ARVALID,
    output wire                                          s_axi_control_ARREADY,
    input wire  [    (C_S_AXI_CONTROL_ADDR_WIDTH - 1):0] s_axi_control_ARADDR,
    output wire                                          s_axi_control_RVALID,
    input wire                                           s_axi_control_RREADY,
    output wire [    (C_S_AXI_CONTROL_DATA_WIDTH - 1):0] s_axi_control_RDATA,
    output wire [                                   1:0] s_axi_control_RRESP,
    output wire                                          s_axi_control_BVALID,
    input wire                                           s_axi_control_BREADY,
    output wire [                                   1:0] s_axi_control_BRESP,
    input wire                                           ap_clk,
    input wire                                           ap_rst_n,
    output wire                                          interrupt,
    output wire [                                  63:0] m_axi_L4_out_dist_ARADDR,
    output wire [                                   1:0] m_axi_L4_out_dist_ARBURST,
    output wire [                                   3:0] m_axi_L4_out_dist_ARCACHE,
    output wire [                                   0:0] m_axi_L4_out_dist_ARID,
    output wire [                                   7:0] m_axi_L4_out_dist_ARLEN,
    output wire                                          m_axi_L4_out_dist_ARLOCK,
    output wire [                                   2:0] m_axi_L4_out_dist_ARPROT,
    output wire [                                   3:0] m_axi_L4_out_dist_ARQOS,
    input wire                                           m_axi_L4_out_dist_ARREADY,
    output wire [                                   2:0] m_axi_L4_out_dist_ARSIZE,
    output wire                                          m_axi_L4_out_dist_ARVALID,
    output wire [                                  63:0] m_axi_L4_out_dist_AWADDR,
    output wire [                                   1:0] m_axi_L4_out_dist_AWBURST,
    output wire [                                   3:0] m_axi_L4_out_dist_AWCACHE,
    output wire [                                   0:0] m_axi_L4_out_dist_AWID,
    output wire [                                   7:0] m_axi_L4_out_dist_AWLEN,
    output wire                                          m_axi_L4_out_dist_AWLOCK,
    output wire [                                   2:0] m_axi_L4_out_dist_AWPROT,
    output wire [                                   3:0] m_axi_L4_out_dist_AWQOS,
    input wire                                           m_axi_L4_out_dist_AWREADY,
    output wire [                                   2:0] m_axi_L4_out_dist_AWSIZE,
    output wire                                          m_axi_L4_out_dist_AWVALID,
    input wire  [                                   0:0] m_axi_L4_out_dist_BID,
    output wire                                          m_axi_L4_out_dist_BREADY,
    input wire  [                                   1:0] m_axi_L4_out_dist_BRESP,
    input wire                                           m_axi_L4_out_dist_BVALID,
    input wire  [                                  31:0] m_axi_L4_out_dist_RDATA,
    input wire  [                                   0:0] m_axi_L4_out_dist_RID,
    input wire                                           m_axi_L4_out_dist_RLAST,
    output wire                                          m_axi_L4_out_dist_RREADY,
    input wire  [                                   1:0] m_axi_L4_out_dist_RRESP,
    input wire                                           m_axi_L4_out_dist_RVALID,
    output wire [                                  31:0] m_axi_L4_out_dist_WDATA,
    output wire                                          m_axi_L4_out_dist_WLAST,
    input wire                                           m_axi_L4_out_dist_WREADY,
    output wire [                                   3:0] m_axi_L4_out_dist_WSTRB,
    output wire                                          m_axi_L4_out_dist_WVALID,
    output wire [                                  63:0] m_axi_L4_out_id_ARADDR,
    output wire [                                   1:0] m_axi_L4_out_id_ARBURST,
    output wire [                                   3:0] m_axi_L4_out_id_ARCACHE,
    output wire [                                   0:0] m_axi_L4_out_id_ARID,
    output wire [                                   7:0] m_axi_L4_out_id_ARLEN,
    output wire                                          m_axi_L4_out_id_ARLOCK,
    output wire [                                   2:0] m_axi_L4_out_id_ARPROT,
    output wire [                                   3:0] m_axi_L4_out_id_ARQOS,
    input wire                                           m_axi_L4_out_id_ARREADY,
    output wire [                                   2:0] m_axi_L4_out_id_ARSIZE,
    output wire                                          m_axi_L4_out_id_ARVALID,
    output wire [                                  63:0] m_axi_L4_out_id_AWADDR,
    output wire [                                   1:0] m_axi_L4_out_id_AWBURST,
    output wire [                                   3:0] m_axi_L4_out_id_AWCACHE,
    output wire [                                   0:0] m_axi_L4_out_id_AWID,
    output wire [                                   7:0] m_axi_L4_out_id_AWLEN,
    output wire                                          m_axi_L4_out_id_AWLOCK,
    output wire [                                   2:0] m_axi_L4_out_id_AWPROT,
    output wire [                                   3:0] m_axi_L4_out_id_AWQOS,
    input wire                                           m_axi_L4_out_id_AWREADY,
    output wire [                                   2:0] m_axi_L4_out_id_AWSIZE,
    output wire                                          m_axi_L4_out_id_AWVALID,
    input wire  [                                   0:0] m_axi_L4_out_id_BID,
    output wire                                          m_axi_L4_out_id_BREADY,
    input wire  [                                   1:0] m_axi_L4_out_id_BRESP,
    input wire                                           m_axi_L4_out_id_BVALID,
    input wire  [                                  31:0] m_axi_L4_out_id_RDATA,
    input wire  [                                   0:0] m_axi_L4_out_id_RID,
    input wire                                           m_axi_L4_out_id_RLAST,
    output wire                                          m_axi_L4_out_id_RREADY,
    input wire  [                                   1:0] m_axi_L4_out_id_RRESP,
    input wire                                           m_axi_L4_out_id_RVALID,
    output wire [                                  31:0] m_axi_L4_out_id_WDATA,
    output wire                                          m_axi_L4_out_id_WLAST,
    input wire                                           m_axi_L4_out_id_WREADY,
    output wire [                                   3:0] m_axi_L4_out_id_WSTRB,
    output wire                                          m_axi_L4_out_id_WVALID,
    output wire [                                  63:0] m_axi_in_0_ARADDR,
    output wire [                                   1:0] m_axi_in_0_ARBURST,
    output wire [                                   3:0] m_axi_in_0_ARCACHE,
    output wire [                                   0:0] m_axi_in_0_ARID,
    output wire [                                   7:0] m_axi_in_0_ARLEN,
    output wire                                          m_axi_in_0_ARLOCK,
    output wire [                                   2:0] m_axi_in_0_ARPROT,
    output wire [                                   3:0] m_axi_in_0_ARQOS,
    input wire                                           m_axi_in_0_ARREADY,
    output wire [                                   2:0] m_axi_in_0_ARSIZE,
    output wire                                          m_axi_in_0_ARVALID,
    output wire [                                  63:0] m_axi_in_0_AWADDR,
    output wire [                                   1:0] m_axi_in_0_AWBURST,
    output wire [                                   3:0] m_axi_in_0_AWCACHE,
    output wire [                                   0:0] m_axi_in_0_AWID,
    output wire [                                   7:0] m_axi_in_0_AWLEN,
    output wire                                          m_axi_in_0_AWLOCK,
    output wire [                                   2:0] m_axi_in_0_AWPROT,
    output wire [                                   3:0] m_axi_in_0_AWQOS,
    input wire                                           m_axi_in_0_AWREADY,
    output wire [                                   2:0] m_axi_in_0_AWSIZE,
    output wire                                          m_axi_in_0_AWVALID,
    input wire  [                                   0:0] m_axi_in_0_BID,
    output wire                                          m_axi_in_0_BREADY,
    input wire  [                                   1:0] m_axi_in_0_BRESP,
    input wire                                           m_axi_in_0_BVALID,
    input wire  [                                 255:0] m_axi_in_0_RDATA,
    input wire  [                                   0:0] m_axi_in_0_RID,
    input wire                                           m_axi_in_0_RLAST,
    output wire                                          m_axi_in_0_RREADY,
    input wire  [                                   1:0] m_axi_in_0_RRESP,
    input wire                                           m_axi_in_0_RVALID,
    output wire [                                 255:0] m_axi_in_0_WDATA,
    output wire                                          m_axi_in_0_WLAST,
    input wire                                           m_axi_in_0_WREADY,
    output wire [                                  31:0] m_axi_in_0_WSTRB,
    output wire                                          m_axi_in_0_WVALID,
    output wire [                                  63:0] m_axi_in_1_ARADDR,
    output wire [                                   1:0] m_axi_in_1_ARBURST,
    output wire [                                   3:0] m_axi_in_1_ARCACHE,
    output wire [                                   0:0] m_axi_in_1_ARID,
    output wire [                                   7:0] m_axi_in_1_ARLEN,
    output wire                                          m_axi_in_1_ARLOCK,
    output wire [                                   2:0] m_axi_in_1_ARPROT,
    output wire [                                   3:0] m_axi_in_1_ARQOS,
    input wire                                           m_axi_in_1_ARREADY,
    output wire [                                   2:0] m_axi_in_1_ARSIZE,
    output wire                                          m_axi_in_1_ARVALID,
    output wire [                                  63:0] m_axi_in_1_AWADDR,
    output wire [                                   1:0] m_axi_in_1_AWBURST,
    output wire [                                   3:0] m_axi_in_1_AWCACHE,
    output wire [                                   0:0] m_axi_in_1_AWID,
    output wire [                                   7:0] m_axi_in_1_AWLEN,
    output wire                                          m_axi_in_1_AWLOCK,
    output wire [                                   2:0] m_axi_in_1_AWPROT,
    output wire [                                   3:0] m_axi_in_1_AWQOS,
    input wire                                           m_axi_in_1_AWREADY,
    output wire [                                   2:0] m_axi_in_1_AWSIZE,
    output wire                                          m_axi_in_1_AWVALID,
    input wire  [                                   0:0] m_axi_in_1_BID,
    output wire                                          m_axi_in_1_BREADY,
    input wire  [                                   1:0] m_axi_in_1_BRESP,
    input wire                                           m_axi_in_1_BVALID,
    input wire  [                                 255:0] m_axi_in_1_RDATA,
    input wire  [                                   0:0] m_axi_in_1_RID,
    input wire                                           m_axi_in_1_RLAST,
    output wire                                          m_axi_in_1_RREADY,
    input wire  [                                   1:0] m_axi_in_1_RRESP,
    input wire                                           m_axi_in_1_RVALID,
    output wire [                                 255:0] m_axi_in_1_WDATA,
    output wire                                          m_axi_in_1_WLAST,
    input wire                                           m_axi_in_1_WREADY,
    output wire [                                  31:0] m_axi_in_1_WSTRB,
    output wire                                          m_axi_in_1_WVALID,
    output wire [                                  63:0] m_axi_in_10_ARADDR,
    output wire [                                   1:0] m_axi_in_10_ARBURST,
    output wire [                                   3:0] m_axi_in_10_ARCACHE,
    output wire [                                   0:0] m_axi_in_10_ARID,
    output wire [                                   7:0] m_axi_in_10_ARLEN,
    output wire                                          m_axi_in_10_ARLOCK,
    output wire [                                   2:0] m_axi_in_10_ARPROT,
    output wire [                                   3:0] m_axi_in_10_ARQOS,
    input wire                                           m_axi_in_10_ARREADY,
    output wire [                                   2:0] m_axi_in_10_ARSIZE,
    output wire                                          m_axi_in_10_ARVALID,
    output wire [                                  63:0] m_axi_in_10_AWADDR,
    output wire [                                   1:0] m_axi_in_10_AWBURST,
    output wire [                                   3:0] m_axi_in_10_AWCACHE,
    output wire [                                   0:0] m_axi_in_10_AWID,
    output wire [                                   7:0] m_axi_in_10_AWLEN,
    output wire                                          m_axi_in_10_AWLOCK,
    output wire [                                   2:0] m_axi_in_10_AWPROT,
    output wire [                                   3:0] m_axi_in_10_AWQOS,
    input wire                                           m_axi_in_10_AWREADY,
    output wire [                                   2:0] m_axi_in_10_AWSIZE,
    output wire                                          m_axi_in_10_AWVALID,
    input wire  [                                   0:0] m_axi_in_10_BID,
    output wire                                          m_axi_in_10_BREADY,
    input wire  [                                   1:0] m_axi_in_10_BRESP,
    input wire                                           m_axi_in_10_BVALID,
    input wire  [                                 255:0] m_axi_in_10_RDATA,
    input wire  [                                   0:0] m_axi_in_10_RID,
    input wire                                           m_axi_in_10_RLAST,
    output wire                                          m_axi_in_10_RREADY,
    input wire  [                                   1:0] m_axi_in_10_RRESP,
    input wire                                           m_axi_in_10_RVALID,
    output wire [                                 255:0] m_axi_in_10_WDATA,
    output wire                                          m_axi_in_10_WLAST,
    input wire                                           m_axi_in_10_WREADY,
    output wire [                                  31:0] m_axi_in_10_WSTRB,
    output wire                                          m_axi_in_10_WVALID,
    output wire [                                  63:0] m_axi_in_11_ARADDR,
    output wire [                                   1:0] m_axi_in_11_ARBURST,
    output wire [                                   3:0] m_axi_in_11_ARCACHE,
    output wire [                                   0:0] m_axi_in_11_ARID,
    output wire [                                   7:0] m_axi_in_11_ARLEN,
    output wire                                          m_axi_in_11_ARLOCK,
    output wire [                                   2:0] m_axi_in_11_ARPROT,
    output wire [                                   3:0] m_axi_in_11_ARQOS,
    input wire                                           m_axi_in_11_ARREADY,
    output wire [                                   2:0] m_axi_in_11_ARSIZE,
    output wire                                          m_axi_in_11_ARVALID,
    output wire [                                  63:0] m_axi_in_11_AWADDR,
    output wire [                                   1:0] m_axi_in_11_AWBURST,
    output wire [                                   3:0] m_axi_in_11_AWCACHE,
    output wire [                                   0:0] m_axi_in_11_AWID,
    output wire [                                   7:0] m_axi_in_11_AWLEN,
    output wire                                          m_axi_in_11_AWLOCK,
    output wire [                                   2:0] m_axi_in_11_AWPROT,
    output wire [                                   3:0] m_axi_in_11_AWQOS,
    input wire                                           m_axi_in_11_AWREADY,
    output wire [                                   2:0] m_axi_in_11_AWSIZE,
    output wire                                          m_axi_in_11_AWVALID,
    input wire  [                                   0:0] m_axi_in_11_BID,
    output wire                                          m_axi_in_11_BREADY,
    input wire  [                                   1:0] m_axi_in_11_BRESP,
    input wire                                           m_axi_in_11_BVALID,
    input wire  [                                 255:0] m_axi_in_11_RDATA,
    input wire  [                                   0:0] m_axi_in_11_RID,
    input wire                                           m_axi_in_11_RLAST,
    output wire                                          m_axi_in_11_RREADY,
    input wire  [                                   1:0] m_axi_in_11_RRESP,
    input wire                                           m_axi_in_11_RVALID,
    output wire [                                 255:0] m_axi_in_11_WDATA,
    output wire                                          m_axi_in_11_WLAST,
    input wire                                           m_axi_in_11_WREADY,
    output wire [                                  31:0] m_axi_in_11_WSTRB,
    output wire                                          m_axi_in_11_WVALID,
    output wire [                                  63:0] m_axi_in_12_ARADDR,
    output wire [                                   1:0] m_axi_in_12_ARBURST,
    output wire [                                   3:0] m_axi_in_12_ARCACHE,
    output wire [                                   0:0] m_axi_in_12_ARID,
    output wire [                                   7:0] m_axi_in_12_ARLEN,
    output wire                                          m_axi_in_12_ARLOCK,
    output wire [                                   2:0] m_axi_in_12_ARPROT,
    output wire [                                   3:0] m_axi_in_12_ARQOS,
    input wire                                           m_axi_in_12_ARREADY,
    output wire [                                   2:0] m_axi_in_12_ARSIZE,
    output wire                                          m_axi_in_12_ARVALID,
    output wire [                                  63:0] m_axi_in_12_AWADDR,
    output wire [                                   1:0] m_axi_in_12_AWBURST,
    output wire [                                   3:0] m_axi_in_12_AWCACHE,
    output wire [                                   0:0] m_axi_in_12_AWID,
    output wire [                                   7:0] m_axi_in_12_AWLEN,
    output wire                                          m_axi_in_12_AWLOCK,
    output wire [                                   2:0] m_axi_in_12_AWPROT,
    output wire [                                   3:0] m_axi_in_12_AWQOS,
    input wire                                           m_axi_in_12_AWREADY,
    output wire [                                   2:0] m_axi_in_12_AWSIZE,
    output wire                                          m_axi_in_12_AWVALID,
    input wire  [                                   0:0] m_axi_in_12_BID,
    output wire                                          m_axi_in_12_BREADY,
    input wire  [                                   1:0] m_axi_in_12_BRESP,
    input wire                                           m_axi_in_12_BVALID,
    input wire  [                                 255:0] m_axi_in_12_RDATA,
    input wire  [                                   0:0] m_axi_in_12_RID,
    input wire                                           m_axi_in_12_RLAST,
    output wire                                          m_axi_in_12_RREADY,
    input wire  [                                   1:0] m_axi_in_12_RRESP,
    input wire                                           m_axi_in_12_RVALID,
    output wire [                                 255:0] m_axi_in_12_WDATA,
    output wire                                          m_axi_in_12_WLAST,
    input wire                                           m_axi_in_12_WREADY,
    output wire [                                  31:0] m_axi_in_12_WSTRB,
    output wire                                          m_axi_in_12_WVALID,
    output wire [                                  63:0] m_axi_in_13_ARADDR,
    output wire [                                   1:0] m_axi_in_13_ARBURST,
    output wire [                                   3:0] m_axi_in_13_ARCACHE,
    output wire [                                   0:0] m_axi_in_13_ARID,
    output wire [                                   7:0] m_axi_in_13_ARLEN,
    output wire                                          m_axi_in_13_ARLOCK,
    output wire [                                   2:0] m_axi_in_13_ARPROT,
    output wire [                                   3:0] m_axi_in_13_ARQOS,
    input wire                                           m_axi_in_13_ARREADY,
    output wire [                                   2:0] m_axi_in_13_ARSIZE,
    output wire                                          m_axi_in_13_ARVALID,
    output wire [                                  63:0] m_axi_in_13_AWADDR,
    output wire [                                   1:0] m_axi_in_13_AWBURST,
    output wire [                                   3:0] m_axi_in_13_AWCACHE,
    output wire [                                   0:0] m_axi_in_13_AWID,
    output wire [                                   7:0] m_axi_in_13_AWLEN,
    output wire                                          m_axi_in_13_AWLOCK,
    output wire [                                   2:0] m_axi_in_13_AWPROT,
    output wire [                                   3:0] m_axi_in_13_AWQOS,
    input wire                                           m_axi_in_13_AWREADY,
    output wire [                                   2:0] m_axi_in_13_AWSIZE,
    output wire                                          m_axi_in_13_AWVALID,
    input wire  [                                   0:0] m_axi_in_13_BID,
    output wire                                          m_axi_in_13_BREADY,
    input wire  [                                   1:0] m_axi_in_13_BRESP,
    input wire                                           m_axi_in_13_BVALID,
    input wire  [                                 255:0] m_axi_in_13_RDATA,
    input wire  [                                   0:0] m_axi_in_13_RID,
    input wire                                           m_axi_in_13_RLAST,
    output wire                                          m_axi_in_13_RREADY,
    input wire  [                                   1:0] m_axi_in_13_RRESP,
    input wire                                           m_axi_in_13_RVALID,
    output wire [                                 255:0] m_axi_in_13_WDATA,
    output wire                                          m_axi_in_13_WLAST,
    input wire                                           m_axi_in_13_WREADY,
    output wire [                                  31:0] m_axi_in_13_WSTRB,
    output wire                                          m_axi_in_13_WVALID,
    output wire [                                  63:0] m_axi_in_14_ARADDR,
    output wire [                                   1:0] m_axi_in_14_ARBURST,
    output wire [                                   3:0] m_axi_in_14_ARCACHE,
    output wire [                                   0:0] m_axi_in_14_ARID,
    output wire [                                   7:0] m_axi_in_14_ARLEN,
    output wire                                          m_axi_in_14_ARLOCK,
    output wire [                                   2:0] m_axi_in_14_ARPROT,
    output wire [                                   3:0] m_axi_in_14_ARQOS,
    input wire                                           m_axi_in_14_ARREADY,
    output wire [                                   2:0] m_axi_in_14_ARSIZE,
    output wire                                          m_axi_in_14_ARVALID,
    output wire [                                  63:0] m_axi_in_14_AWADDR,
    output wire [                                   1:0] m_axi_in_14_AWBURST,
    output wire [                                   3:0] m_axi_in_14_AWCACHE,
    output wire [                                   0:0] m_axi_in_14_AWID,
    output wire [                                   7:0] m_axi_in_14_AWLEN,
    output wire                                          m_axi_in_14_AWLOCK,
    output wire [                                   2:0] m_axi_in_14_AWPROT,
    output wire [                                   3:0] m_axi_in_14_AWQOS,
    input wire                                           m_axi_in_14_AWREADY,
    output wire [                                   2:0] m_axi_in_14_AWSIZE,
    output wire                                          m_axi_in_14_AWVALID,
    input wire  [                                   0:0] m_axi_in_14_BID,
    output wire                                          m_axi_in_14_BREADY,
    input wire  [                                   1:0] m_axi_in_14_BRESP,
    input wire                                           m_axi_in_14_BVALID,
    input wire  [                                 255:0] m_axi_in_14_RDATA,
    input wire  [                                   0:0] m_axi_in_14_RID,
    input wire                                           m_axi_in_14_RLAST,
    output wire                                          m_axi_in_14_RREADY,
    input wire  [                                   1:0] m_axi_in_14_RRESP,
    input wire                                           m_axi_in_14_RVALID,
    output wire [                                 255:0] m_axi_in_14_WDATA,
    output wire                                          m_axi_in_14_WLAST,
    input wire                                           m_axi_in_14_WREADY,
    output wire [                                  31:0] m_axi_in_14_WSTRB,
    output wire                                          m_axi_in_14_WVALID,
    output wire [                                  63:0] m_axi_in_15_ARADDR,
    output wire [                                   1:0] m_axi_in_15_ARBURST,
    output wire [                                   3:0] m_axi_in_15_ARCACHE,
    output wire [                                   0:0] m_axi_in_15_ARID,
    output wire [                                   7:0] m_axi_in_15_ARLEN,
    output wire                                          m_axi_in_15_ARLOCK,
    output wire [                                   2:0] m_axi_in_15_ARPROT,
    output wire [                                   3:0] m_axi_in_15_ARQOS,
    input wire                                           m_axi_in_15_ARREADY,
    output wire [                                   2:0] m_axi_in_15_ARSIZE,
    output wire                                          m_axi_in_15_ARVALID,
    output wire [                                  63:0] m_axi_in_15_AWADDR,
    output wire [                                   1:0] m_axi_in_15_AWBURST,
    output wire [                                   3:0] m_axi_in_15_AWCACHE,
    output wire [                                   0:0] m_axi_in_15_AWID,
    output wire [                                   7:0] m_axi_in_15_AWLEN,
    output wire                                          m_axi_in_15_AWLOCK,
    output wire [                                   2:0] m_axi_in_15_AWPROT,
    output wire [                                   3:0] m_axi_in_15_AWQOS,
    input wire                                           m_axi_in_15_AWREADY,
    output wire [                                   2:0] m_axi_in_15_AWSIZE,
    output wire                                          m_axi_in_15_AWVALID,
    input wire  [                                   0:0] m_axi_in_15_BID,
    output wire                                          m_axi_in_15_BREADY,
    input wire  [                                   1:0] m_axi_in_15_BRESP,
    input wire                                           m_axi_in_15_BVALID,
    input wire  [                                 255:0] m_axi_in_15_RDATA,
    input wire  [                                   0:0] m_axi_in_15_RID,
    input wire                                           m_axi_in_15_RLAST,
    output wire                                          m_axi_in_15_RREADY,
    input wire  [                                   1:0] m_axi_in_15_RRESP,
    input wire                                           m_axi_in_15_RVALID,
    output wire [                                 255:0] m_axi_in_15_WDATA,
    output wire                                          m_axi_in_15_WLAST,
    input wire                                           m_axi_in_15_WREADY,
    output wire [                                  31:0] m_axi_in_15_WSTRB,
    output wire                                          m_axi_in_15_WVALID,
    output wire [                                  63:0] m_axi_in_16_ARADDR,
    output wire [                                   1:0] m_axi_in_16_ARBURST,
    output wire [                                   3:0] m_axi_in_16_ARCACHE,
    output wire [                                   0:0] m_axi_in_16_ARID,
    output wire [                                   7:0] m_axi_in_16_ARLEN,
    output wire                                          m_axi_in_16_ARLOCK,
    output wire [                                   2:0] m_axi_in_16_ARPROT,
    output wire [                                   3:0] m_axi_in_16_ARQOS,
    input wire                                           m_axi_in_16_ARREADY,
    output wire [                                   2:0] m_axi_in_16_ARSIZE,
    output wire                                          m_axi_in_16_ARVALID,
    output wire [                                  63:0] m_axi_in_16_AWADDR,
    output wire [                                   1:0] m_axi_in_16_AWBURST,
    output wire [                                   3:0] m_axi_in_16_AWCACHE,
    output wire [                                   0:0] m_axi_in_16_AWID,
    output wire [                                   7:0] m_axi_in_16_AWLEN,
    output wire                                          m_axi_in_16_AWLOCK,
    output wire [                                   2:0] m_axi_in_16_AWPROT,
    output wire [                                   3:0] m_axi_in_16_AWQOS,
    input wire                                           m_axi_in_16_AWREADY,
    output wire [                                   2:0] m_axi_in_16_AWSIZE,
    output wire                                          m_axi_in_16_AWVALID,
    input wire  [                                   0:0] m_axi_in_16_BID,
    output wire                                          m_axi_in_16_BREADY,
    input wire  [                                   1:0] m_axi_in_16_BRESP,
    input wire                                           m_axi_in_16_BVALID,
    input wire  [                                 255:0] m_axi_in_16_RDATA,
    input wire  [                                   0:0] m_axi_in_16_RID,
    input wire                                           m_axi_in_16_RLAST,
    output wire                                          m_axi_in_16_RREADY,
    input wire  [                                   1:0] m_axi_in_16_RRESP,
    input wire                                           m_axi_in_16_RVALID,
    output wire [                                 255:0] m_axi_in_16_WDATA,
    output wire                                          m_axi_in_16_WLAST,
    input wire                                           m_axi_in_16_WREADY,
    output wire [                                  31:0] m_axi_in_16_WSTRB,
    output wire                                          m_axi_in_16_WVALID,
    output wire [                                  63:0] m_axi_in_17_ARADDR,
    output wire [                                   1:0] m_axi_in_17_ARBURST,
    output wire [                                   3:0] m_axi_in_17_ARCACHE,
    output wire [                                   0:0] m_axi_in_17_ARID,
    output wire [                                   7:0] m_axi_in_17_ARLEN,
    output wire                                          m_axi_in_17_ARLOCK,
    output wire [                                   2:0] m_axi_in_17_ARPROT,
    output wire [                                   3:0] m_axi_in_17_ARQOS,
    input wire                                           m_axi_in_17_ARREADY,
    output wire [                                   2:0] m_axi_in_17_ARSIZE,
    output wire                                          m_axi_in_17_ARVALID,
    output wire [                                  63:0] m_axi_in_17_AWADDR,
    output wire [                                   1:0] m_axi_in_17_AWBURST,
    output wire [                                   3:0] m_axi_in_17_AWCACHE,
    output wire [                                   0:0] m_axi_in_17_AWID,
    output wire [                                   7:0] m_axi_in_17_AWLEN,
    output wire                                          m_axi_in_17_AWLOCK,
    output wire [                                   2:0] m_axi_in_17_AWPROT,
    output wire [                                   3:0] m_axi_in_17_AWQOS,
    input wire                                           m_axi_in_17_AWREADY,
    output wire [                                   2:0] m_axi_in_17_AWSIZE,
    output wire                                          m_axi_in_17_AWVALID,
    input wire  [                                   0:0] m_axi_in_17_BID,
    output wire                                          m_axi_in_17_BREADY,
    input wire  [                                   1:0] m_axi_in_17_BRESP,
    input wire                                           m_axi_in_17_BVALID,
    input wire  [                                 255:0] m_axi_in_17_RDATA,
    input wire  [                                   0:0] m_axi_in_17_RID,
    input wire                                           m_axi_in_17_RLAST,
    output wire                                          m_axi_in_17_RREADY,
    input wire  [                                   1:0] m_axi_in_17_RRESP,
    input wire                                           m_axi_in_17_RVALID,
    output wire [                                 255:0] m_axi_in_17_WDATA,
    output wire                                          m_axi_in_17_WLAST,
    input wire                                           m_axi_in_17_WREADY,
    output wire [                                  31:0] m_axi_in_17_WSTRB,
    output wire                                          m_axi_in_17_WVALID,
    output wire [                                  63:0] m_axi_in_18_ARADDR,
    output wire [                                   1:0] m_axi_in_18_ARBURST,
    output wire [                                   3:0] m_axi_in_18_ARCACHE,
    output wire [                                   0:0] m_axi_in_18_ARID,
    output wire [                                   7:0] m_axi_in_18_ARLEN,
    output wire                                          m_axi_in_18_ARLOCK,
    output wire [                                   2:0] m_axi_in_18_ARPROT,
    output wire [                                   3:0] m_axi_in_18_ARQOS,
    input wire                                           m_axi_in_18_ARREADY,
    output wire [                                   2:0] m_axi_in_18_ARSIZE,
    output wire                                          m_axi_in_18_ARVALID,
    output wire [                                  63:0] m_axi_in_18_AWADDR,
    output wire [                                   1:0] m_axi_in_18_AWBURST,
    output wire [                                   3:0] m_axi_in_18_AWCACHE,
    output wire [                                   0:0] m_axi_in_18_AWID,
    output wire [                                   7:0] m_axi_in_18_AWLEN,
    output wire                                          m_axi_in_18_AWLOCK,
    output wire [                                   2:0] m_axi_in_18_AWPROT,
    output wire [                                   3:0] m_axi_in_18_AWQOS,
    input wire                                           m_axi_in_18_AWREADY,
    output wire [                                   2:0] m_axi_in_18_AWSIZE,
    output wire                                          m_axi_in_18_AWVALID,
    input wire  [                                   0:0] m_axi_in_18_BID,
    output wire                                          m_axi_in_18_BREADY,
    input wire  [                                   1:0] m_axi_in_18_BRESP,
    input wire                                           m_axi_in_18_BVALID,
    input wire  [                                 255:0] m_axi_in_18_RDATA,
    input wire  [                                   0:0] m_axi_in_18_RID,
    input wire                                           m_axi_in_18_RLAST,
    output wire                                          m_axi_in_18_RREADY,
    input wire  [                                   1:0] m_axi_in_18_RRESP,
    input wire                                           m_axi_in_18_RVALID,
    output wire [                                 255:0] m_axi_in_18_WDATA,
    output wire                                          m_axi_in_18_WLAST,
    input wire                                           m_axi_in_18_WREADY,
    output wire [                                  31:0] m_axi_in_18_WSTRB,
    output wire                                          m_axi_in_18_WVALID,
    output wire [                                  63:0] m_axi_in_19_ARADDR,
    output wire [                                   1:0] m_axi_in_19_ARBURST,
    output wire [                                   3:0] m_axi_in_19_ARCACHE,
    output wire [                                   0:0] m_axi_in_19_ARID,
    output wire [                                   7:0] m_axi_in_19_ARLEN,
    output wire                                          m_axi_in_19_ARLOCK,
    output wire [                                   2:0] m_axi_in_19_ARPROT,
    output wire [                                   3:0] m_axi_in_19_ARQOS,
    input wire                                           m_axi_in_19_ARREADY,
    output wire [                                   2:0] m_axi_in_19_ARSIZE,
    output wire                                          m_axi_in_19_ARVALID,
    output wire [                                  63:0] m_axi_in_19_AWADDR,
    output wire [                                   1:0] m_axi_in_19_AWBURST,
    output wire [                                   3:0] m_axi_in_19_AWCACHE,
    output wire [                                   0:0] m_axi_in_19_AWID,
    output wire [                                   7:0] m_axi_in_19_AWLEN,
    output wire                                          m_axi_in_19_AWLOCK,
    output wire [                                   2:0] m_axi_in_19_AWPROT,
    output wire [                                   3:0] m_axi_in_19_AWQOS,
    input wire                                           m_axi_in_19_AWREADY,
    output wire [                                   2:0] m_axi_in_19_AWSIZE,
    output wire                                          m_axi_in_19_AWVALID,
    input wire  [                                   0:0] m_axi_in_19_BID,
    output wire                                          m_axi_in_19_BREADY,
    input wire  [                                   1:0] m_axi_in_19_BRESP,
    input wire                                           m_axi_in_19_BVALID,
    input wire  [                                 255:0] m_axi_in_19_RDATA,
    input wire  [                                   0:0] m_axi_in_19_RID,
    input wire                                           m_axi_in_19_RLAST,
    output wire                                          m_axi_in_19_RREADY,
    input wire  [                                   1:0] m_axi_in_19_RRESP,
    input wire                                           m_axi_in_19_RVALID,
    output wire [                                 255:0] m_axi_in_19_WDATA,
    output wire                                          m_axi_in_19_WLAST,
    input wire                                           m_axi_in_19_WREADY,
    output wire [                                  31:0] m_axi_in_19_WSTRB,
    output wire                                          m_axi_in_19_WVALID,
    output wire [                                  63:0] m_axi_in_2_ARADDR,
    output wire [                                   1:0] m_axi_in_2_ARBURST,
    output wire [                                   3:0] m_axi_in_2_ARCACHE,
    output wire [                                   0:0] m_axi_in_2_ARID,
    output wire [                                   7:0] m_axi_in_2_ARLEN,
    output wire                                          m_axi_in_2_ARLOCK,
    output wire [                                   2:0] m_axi_in_2_ARPROT,
    output wire [                                   3:0] m_axi_in_2_ARQOS,
    input wire                                           m_axi_in_2_ARREADY,
    output wire [                                   2:0] m_axi_in_2_ARSIZE,
    output wire                                          m_axi_in_2_ARVALID,
    output wire [                                  63:0] m_axi_in_2_AWADDR,
    output wire [                                   1:0] m_axi_in_2_AWBURST,
    output wire [                                   3:0] m_axi_in_2_AWCACHE,
    output wire [                                   0:0] m_axi_in_2_AWID,
    output wire [                                   7:0] m_axi_in_2_AWLEN,
    output wire                                          m_axi_in_2_AWLOCK,
    output wire [                                   2:0] m_axi_in_2_AWPROT,
    output wire [                                   3:0] m_axi_in_2_AWQOS,
    input wire                                           m_axi_in_2_AWREADY,
    output wire [                                   2:0] m_axi_in_2_AWSIZE,
    output wire                                          m_axi_in_2_AWVALID,
    input wire  [                                   0:0] m_axi_in_2_BID,
    output wire                                          m_axi_in_2_BREADY,
    input wire  [                                   1:0] m_axi_in_2_BRESP,
    input wire                                           m_axi_in_2_BVALID,
    input wire  [                                 255:0] m_axi_in_2_RDATA,
    input wire  [                                   0:0] m_axi_in_2_RID,
    input wire                                           m_axi_in_2_RLAST,
    output wire                                          m_axi_in_2_RREADY,
    input wire  [                                   1:0] m_axi_in_2_RRESP,
    input wire                                           m_axi_in_2_RVALID,
    output wire [                                 255:0] m_axi_in_2_WDATA,
    output wire                                          m_axi_in_2_WLAST,
    input wire                                           m_axi_in_2_WREADY,
    output wire [                                  31:0] m_axi_in_2_WSTRB,
    output wire                                          m_axi_in_2_WVALID,
    output wire [                                  63:0] m_axi_in_20_ARADDR,
    output wire [                                   1:0] m_axi_in_20_ARBURST,
    output wire [                                   3:0] m_axi_in_20_ARCACHE,
    output wire [                                   0:0] m_axi_in_20_ARID,
    output wire [                                   7:0] m_axi_in_20_ARLEN,
    output wire                                          m_axi_in_20_ARLOCK,
    output wire [                                   2:0] m_axi_in_20_ARPROT,
    output wire [                                   3:0] m_axi_in_20_ARQOS,
    input wire                                           m_axi_in_20_ARREADY,
    output wire [                                   2:0] m_axi_in_20_ARSIZE,
    output wire                                          m_axi_in_20_ARVALID,
    output wire [                                  63:0] m_axi_in_20_AWADDR,
    output wire [                                   1:0] m_axi_in_20_AWBURST,
    output wire [                                   3:0] m_axi_in_20_AWCACHE,
    output wire [                                   0:0] m_axi_in_20_AWID,
    output wire [                                   7:0] m_axi_in_20_AWLEN,
    output wire                                          m_axi_in_20_AWLOCK,
    output wire [                                   2:0] m_axi_in_20_AWPROT,
    output wire [                                   3:0] m_axi_in_20_AWQOS,
    input wire                                           m_axi_in_20_AWREADY,
    output wire [                                   2:0] m_axi_in_20_AWSIZE,
    output wire                                          m_axi_in_20_AWVALID,
    input wire  [                                   0:0] m_axi_in_20_BID,
    output wire                                          m_axi_in_20_BREADY,
    input wire  [                                   1:0] m_axi_in_20_BRESP,
    input wire                                           m_axi_in_20_BVALID,
    input wire  [                                 255:0] m_axi_in_20_RDATA,
    input wire  [                                   0:0] m_axi_in_20_RID,
    input wire                                           m_axi_in_20_RLAST,
    output wire                                          m_axi_in_20_RREADY,
    input wire  [                                   1:0] m_axi_in_20_RRESP,
    input wire                                           m_axi_in_20_RVALID,
    output wire [                                 255:0] m_axi_in_20_WDATA,
    output wire                                          m_axi_in_20_WLAST,
    input wire                                           m_axi_in_20_WREADY,
    output wire [                                  31:0] m_axi_in_20_WSTRB,
    output wire                                          m_axi_in_20_WVALID,
    output wire [                                  63:0] m_axi_in_21_ARADDR,
    output wire [                                   1:0] m_axi_in_21_ARBURST,
    output wire [                                   3:0] m_axi_in_21_ARCACHE,
    output wire [                                   0:0] m_axi_in_21_ARID,
    output wire [                                   7:0] m_axi_in_21_ARLEN,
    output wire                                          m_axi_in_21_ARLOCK,
    output wire [                                   2:0] m_axi_in_21_ARPROT,
    output wire [                                   3:0] m_axi_in_21_ARQOS,
    input wire                                           m_axi_in_21_ARREADY,
    output wire [                                   2:0] m_axi_in_21_ARSIZE,
    output wire                                          m_axi_in_21_ARVALID,
    output wire [                                  63:0] m_axi_in_21_AWADDR,
    output wire [                                   1:0] m_axi_in_21_AWBURST,
    output wire [                                   3:0] m_axi_in_21_AWCACHE,
    output wire [                                   0:0] m_axi_in_21_AWID,
    output wire [                                   7:0] m_axi_in_21_AWLEN,
    output wire                                          m_axi_in_21_AWLOCK,
    output wire [                                   2:0] m_axi_in_21_AWPROT,
    output wire [                                   3:0] m_axi_in_21_AWQOS,
    input wire                                           m_axi_in_21_AWREADY,
    output wire [                                   2:0] m_axi_in_21_AWSIZE,
    output wire                                          m_axi_in_21_AWVALID,
    input wire  [                                   0:0] m_axi_in_21_BID,
    output wire                                          m_axi_in_21_BREADY,
    input wire  [                                   1:0] m_axi_in_21_BRESP,
    input wire                                           m_axi_in_21_BVALID,
    input wire  [                                 255:0] m_axi_in_21_RDATA,
    input wire  [                                   0:0] m_axi_in_21_RID,
    input wire                                           m_axi_in_21_RLAST,
    output wire                                          m_axi_in_21_RREADY,
    input wire  [                                   1:0] m_axi_in_21_RRESP,
    input wire                                           m_axi_in_21_RVALID,
    output wire [                                 255:0] m_axi_in_21_WDATA,
    output wire                                          m_axi_in_21_WLAST,
    input wire                                           m_axi_in_21_WREADY,
    output wire [                                  31:0] m_axi_in_21_WSTRB,
    output wire                                          m_axi_in_21_WVALID,
    output wire [                                  63:0] m_axi_in_22_ARADDR,
    output wire [                                   1:0] m_axi_in_22_ARBURST,
    output wire [                                   3:0] m_axi_in_22_ARCACHE,
    output wire [                                   0:0] m_axi_in_22_ARID,
    output wire [                                   7:0] m_axi_in_22_ARLEN,
    output wire                                          m_axi_in_22_ARLOCK,
    output wire [                                   2:0] m_axi_in_22_ARPROT,
    output wire [                                   3:0] m_axi_in_22_ARQOS,
    input wire                                           m_axi_in_22_ARREADY,
    output wire [                                   2:0] m_axi_in_22_ARSIZE,
    output wire                                          m_axi_in_22_ARVALID,
    output wire [                                  63:0] m_axi_in_22_AWADDR,
    output wire [                                   1:0] m_axi_in_22_AWBURST,
    output wire [                                   3:0] m_axi_in_22_AWCACHE,
    output wire [                                   0:0] m_axi_in_22_AWID,
    output wire [                                   7:0] m_axi_in_22_AWLEN,
    output wire                                          m_axi_in_22_AWLOCK,
    output wire [                                   2:0] m_axi_in_22_AWPROT,
    output wire [                                   3:0] m_axi_in_22_AWQOS,
    input wire                                           m_axi_in_22_AWREADY,
    output wire [                                   2:0] m_axi_in_22_AWSIZE,
    output wire                                          m_axi_in_22_AWVALID,
    input wire  [                                   0:0] m_axi_in_22_BID,
    output wire                                          m_axi_in_22_BREADY,
    input wire  [                                   1:0] m_axi_in_22_BRESP,
    input wire                                           m_axi_in_22_BVALID,
    input wire  [                                 255:0] m_axi_in_22_RDATA,
    input wire  [                                   0:0] m_axi_in_22_RID,
    input wire                                           m_axi_in_22_RLAST,
    output wire                                          m_axi_in_22_RREADY,
    input wire  [                                   1:0] m_axi_in_22_RRESP,
    input wire                                           m_axi_in_22_RVALID,
    output wire [                                 255:0] m_axi_in_22_WDATA,
    output wire                                          m_axi_in_22_WLAST,
    input wire                                           m_axi_in_22_WREADY,
    output wire [                                  31:0] m_axi_in_22_WSTRB,
    output wire                                          m_axi_in_22_WVALID,
    output wire [                                  63:0] m_axi_in_23_ARADDR,
    output wire [                                   1:0] m_axi_in_23_ARBURST,
    output wire [                                   3:0] m_axi_in_23_ARCACHE,
    output wire [                                   0:0] m_axi_in_23_ARID,
    output wire [                                   7:0] m_axi_in_23_ARLEN,
    output wire                                          m_axi_in_23_ARLOCK,
    output wire [                                   2:0] m_axi_in_23_ARPROT,
    output wire [                                   3:0] m_axi_in_23_ARQOS,
    input wire                                           m_axi_in_23_ARREADY,
    output wire [                                   2:0] m_axi_in_23_ARSIZE,
    output wire                                          m_axi_in_23_ARVALID,
    output wire [                                  63:0] m_axi_in_23_AWADDR,
    output wire [                                   1:0] m_axi_in_23_AWBURST,
    output wire [                                   3:0] m_axi_in_23_AWCACHE,
    output wire [                                   0:0] m_axi_in_23_AWID,
    output wire [                                   7:0] m_axi_in_23_AWLEN,
    output wire                                          m_axi_in_23_AWLOCK,
    output wire [                                   2:0] m_axi_in_23_AWPROT,
    output wire [                                   3:0] m_axi_in_23_AWQOS,
    input wire                                           m_axi_in_23_AWREADY,
    output wire [                                   2:0] m_axi_in_23_AWSIZE,
    output wire                                          m_axi_in_23_AWVALID,
    input wire  [                                   0:0] m_axi_in_23_BID,
    output wire                                          m_axi_in_23_BREADY,
    input wire  [                                   1:0] m_axi_in_23_BRESP,
    input wire                                           m_axi_in_23_BVALID,
    input wire  [                                 255:0] m_axi_in_23_RDATA,
    input wire  [                                   0:0] m_axi_in_23_RID,
    input wire                                           m_axi_in_23_RLAST,
    output wire                                          m_axi_in_23_RREADY,
    input wire  [                                   1:0] m_axi_in_23_RRESP,
    input wire                                           m_axi_in_23_RVALID,
    output wire [                                 255:0] m_axi_in_23_WDATA,
    output wire                                          m_axi_in_23_WLAST,
    input wire                                           m_axi_in_23_WREADY,
    output wire [                                  31:0] m_axi_in_23_WSTRB,
    output wire                                          m_axi_in_23_WVALID,
    output wire [                                  63:0] m_axi_in_24_ARADDR,
    output wire [                                   1:0] m_axi_in_24_ARBURST,
    output wire [                                   3:0] m_axi_in_24_ARCACHE,
    output wire [                                   0:0] m_axi_in_24_ARID,
    output wire [                                   7:0] m_axi_in_24_ARLEN,
    output wire                                          m_axi_in_24_ARLOCK,
    output wire [                                   2:0] m_axi_in_24_ARPROT,
    output wire [                                   3:0] m_axi_in_24_ARQOS,
    input wire                                           m_axi_in_24_ARREADY,
    output wire [                                   2:0] m_axi_in_24_ARSIZE,
    output wire                                          m_axi_in_24_ARVALID,
    output wire [                                  63:0] m_axi_in_24_AWADDR,
    output wire [                                   1:0] m_axi_in_24_AWBURST,
    output wire [                                   3:0] m_axi_in_24_AWCACHE,
    output wire [                                   0:0] m_axi_in_24_AWID,
    output wire [                                   7:0] m_axi_in_24_AWLEN,
    output wire                                          m_axi_in_24_AWLOCK,
    output wire [                                   2:0] m_axi_in_24_AWPROT,
    output wire [                                   3:0] m_axi_in_24_AWQOS,
    input wire                                           m_axi_in_24_AWREADY,
    output wire [                                   2:0] m_axi_in_24_AWSIZE,
    output wire                                          m_axi_in_24_AWVALID,
    input wire  [                                   0:0] m_axi_in_24_BID,
    output wire                                          m_axi_in_24_BREADY,
    input wire  [                                   1:0] m_axi_in_24_BRESP,
    input wire                                           m_axi_in_24_BVALID,
    input wire  [                                 255:0] m_axi_in_24_RDATA,
    input wire  [                                   0:0] m_axi_in_24_RID,
    input wire                                           m_axi_in_24_RLAST,
    output wire                                          m_axi_in_24_RREADY,
    input wire  [                                   1:0] m_axi_in_24_RRESP,
    input wire                                           m_axi_in_24_RVALID,
    output wire [                                 255:0] m_axi_in_24_WDATA,
    output wire                                          m_axi_in_24_WLAST,
    input wire                                           m_axi_in_24_WREADY,
    output wire [                                  31:0] m_axi_in_24_WSTRB,
    output wire                                          m_axi_in_24_WVALID,
    output wire [                                  63:0] m_axi_in_25_ARADDR,
    output wire [                                   1:0] m_axi_in_25_ARBURST,
    output wire [                                   3:0] m_axi_in_25_ARCACHE,
    output wire [                                   0:0] m_axi_in_25_ARID,
    output wire [                                   7:0] m_axi_in_25_ARLEN,
    output wire                                          m_axi_in_25_ARLOCK,
    output wire [                                   2:0] m_axi_in_25_ARPROT,
    output wire [                                   3:0] m_axi_in_25_ARQOS,
    input wire                                           m_axi_in_25_ARREADY,
    output wire [                                   2:0] m_axi_in_25_ARSIZE,
    output wire                                          m_axi_in_25_ARVALID,
    output wire [                                  63:0] m_axi_in_25_AWADDR,
    output wire [                                   1:0] m_axi_in_25_AWBURST,
    output wire [                                   3:0] m_axi_in_25_AWCACHE,
    output wire [                                   0:0] m_axi_in_25_AWID,
    output wire [                                   7:0] m_axi_in_25_AWLEN,
    output wire                                          m_axi_in_25_AWLOCK,
    output wire [                                   2:0] m_axi_in_25_AWPROT,
    output wire [                                   3:0] m_axi_in_25_AWQOS,
    input wire                                           m_axi_in_25_AWREADY,
    output wire [                                   2:0] m_axi_in_25_AWSIZE,
    output wire                                          m_axi_in_25_AWVALID,
    input wire  [                                   0:0] m_axi_in_25_BID,
    output wire                                          m_axi_in_25_BREADY,
    input wire  [                                   1:0] m_axi_in_25_BRESP,
    input wire                                           m_axi_in_25_BVALID,
    input wire  [                                 255:0] m_axi_in_25_RDATA,
    input wire  [                                   0:0] m_axi_in_25_RID,
    input wire                                           m_axi_in_25_RLAST,
    output wire                                          m_axi_in_25_RREADY,
    input wire  [                                   1:0] m_axi_in_25_RRESP,
    input wire                                           m_axi_in_25_RVALID,
    output wire [                                 255:0] m_axi_in_25_WDATA,
    output wire                                          m_axi_in_25_WLAST,
    input wire                                           m_axi_in_25_WREADY,
    output wire [                                  31:0] m_axi_in_25_WSTRB,
    output wire                                          m_axi_in_25_WVALID,
    output wire [                                  63:0] m_axi_in_26_ARADDR,
    output wire [                                   1:0] m_axi_in_26_ARBURST,
    output wire [                                   3:0] m_axi_in_26_ARCACHE,
    output wire [                                   0:0] m_axi_in_26_ARID,
    output wire [                                   7:0] m_axi_in_26_ARLEN,
    output wire                                          m_axi_in_26_ARLOCK,
    output wire [                                   2:0] m_axi_in_26_ARPROT,
    output wire [                                   3:0] m_axi_in_26_ARQOS,
    input wire                                           m_axi_in_26_ARREADY,
    output wire [                                   2:0] m_axi_in_26_ARSIZE,
    output wire                                          m_axi_in_26_ARVALID,
    output wire [                                  63:0] m_axi_in_26_AWADDR,
    output wire [                                   1:0] m_axi_in_26_AWBURST,
    output wire [                                   3:0] m_axi_in_26_AWCACHE,
    output wire [                                   0:0] m_axi_in_26_AWID,
    output wire [                                   7:0] m_axi_in_26_AWLEN,
    output wire                                          m_axi_in_26_AWLOCK,
    output wire [                                   2:0] m_axi_in_26_AWPROT,
    output wire [                                   3:0] m_axi_in_26_AWQOS,
    input wire                                           m_axi_in_26_AWREADY,
    output wire [                                   2:0] m_axi_in_26_AWSIZE,
    output wire                                          m_axi_in_26_AWVALID,
    input wire  [                                   0:0] m_axi_in_26_BID,
    output wire                                          m_axi_in_26_BREADY,
    input wire  [                                   1:0] m_axi_in_26_BRESP,
    input wire                                           m_axi_in_26_BVALID,
    input wire  [                                 255:0] m_axi_in_26_RDATA,
    input wire  [                                   0:0] m_axi_in_26_RID,
    input wire                                           m_axi_in_26_RLAST,
    output wire                                          m_axi_in_26_RREADY,
    input wire  [                                   1:0] m_axi_in_26_RRESP,
    input wire                                           m_axi_in_26_RVALID,
    output wire [                                 255:0] m_axi_in_26_WDATA,
    output wire                                          m_axi_in_26_WLAST,
    input wire                                           m_axi_in_26_WREADY,
    output wire [                                  31:0] m_axi_in_26_WSTRB,
    output wire                                          m_axi_in_26_WVALID,
    output wire [                                  63:0] m_axi_in_27_ARADDR,
    output wire [                                   1:0] m_axi_in_27_ARBURST,
    output wire [                                   3:0] m_axi_in_27_ARCACHE,
    output wire [                                   0:0] m_axi_in_27_ARID,
    output wire [                                   7:0] m_axi_in_27_ARLEN,
    output wire                                          m_axi_in_27_ARLOCK,
    output wire [                                   2:0] m_axi_in_27_ARPROT,
    output wire [                                   3:0] m_axi_in_27_ARQOS,
    input wire                                           m_axi_in_27_ARREADY,
    output wire [                                   2:0] m_axi_in_27_ARSIZE,
    output wire                                          m_axi_in_27_ARVALID,
    output wire [                                  63:0] m_axi_in_27_AWADDR,
    output wire [                                   1:0] m_axi_in_27_AWBURST,
    output wire [                                   3:0] m_axi_in_27_AWCACHE,
    output wire [                                   0:0] m_axi_in_27_AWID,
    output wire [                                   7:0] m_axi_in_27_AWLEN,
    output wire                                          m_axi_in_27_AWLOCK,
    output wire [                                   2:0] m_axi_in_27_AWPROT,
    output wire [                                   3:0] m_axi_in_27_AWQOS,
    input wire                                           m_axi_in_27_AWREADY,
    output wire [                                   2:0] m_axi_in_27_AWSIZE,
    output wire                                          m_axi_in_27_AWVALID,
    input wire  [                                   0:0] m_axi_in_27_BID,
    output wire                                          m_axi_in_27_BREADY,
    input wire  [                                   1:0] m_axi_in_27_BRESP,
    input wire                                           m_axi_in_27_BVALID,
    input wire  [                                 255:0] m_axi_in_27_RDATA,
    input wire  [                                   0:0] m_axi_in_27_RID,
    input wire                                           m_axi_in_27_RLAST,
    output wire                                          m_axi_in_27_RREADY,
    input wire  [                                   1:0] m_axi_in_27_RRESP,
    input wire                                           m_axi_in_27_RVALID,
    output wire [                                 255:0] m_axi_in_27_WDATA,
    output wire                                          m_axi_in_27_WLAST,
    input wire                                           m_axi_in_27_WREADY,
    output wire [                                  31:0] m_axi_in_27_WSTRB,
    output wire                                          m_axi_in_27_WVALID,
    output wire [                                  63:0] m_axi_in_28_ARADDR,
    output wire [                                   1:0] m_axi_in_28_ARBURST,
    output wire [                                   3:0] m_axi_in_28_ARCACHE,
    output wire [                                   0:0] m_axi_in_28_ARID,
    output wire [                                   7:0] m_axi_in_28_ARLEN,
    output wire                                          m_axi_in_28_ARLOCK,
    output wire [                                   2:0] m_axi_in_28_ARPROT,
    output wire [                                   3:0] m_axi_in_28_ARQOS,
    input wire                                           m_axi_in_28_ARREADY,
    output wire [                                   2:0] m_axi_in_28_ARSIZE,
    output wire                                          m_axi_in_28_ARVALID,
    output wire [                                  63:0] m_axi_in_28_AWADDR,
    output wire [                                   1:0] m_axi_in_28_AWBURST,
    output wire [                                   3:0] m_axi_in_28_AWCACHE,
    output wire [                                   0:0] m_axi_in_28_AWID,
    output wire [                                   7:0] m_axi_in_28_AWLEN,
    output wire                                          m_axi_in_28_AWLOCK,
    output wire [                                   2:0] m_axi_in_28_AWPROT,
    output wire [                                   3:0] m_axi_in_28_AWQOS,
    input wire                                           m_axi_in_28_AWREADY,
    output wire [                                   2:0] m_axi_in_28_AWSIZE,
    output wire                                          m_axi_in_28_AWVALID,
    input wire  [                                   0:0] m_axi_in_28_BID,
    output wire                                          m_axi_in_28_BREADY,
    input wire  [                                   1:0] m_axi_in_28_BRESP,
    input wire                                           m_axi_in_28_BVALID,
    input wire  [                                 255:0] m_axi_in_28_RDATA,
    input wire  [                                   0:0] m_axi_in_28_RID,
    input wire                                           m_axi_in_28_RLAST,
    output wire                                          m_axi_in_28_RREADY,
    input wire  [                                   1:0] m_axi_in_28_RRESP,
    input wire                                           m_axi_in_28_RVALID,
    output wire [                                 255:0] m_axi_in_28_WDATA,
    output wire                                          m_axi_in_28_WLAST,
    input wire                                           m_axi_in_28_WREADY,
    output wire [                                  31:0] m_axi_in_28_WSTRB,
    output wire                                          m_axi_in_28_WVALID,
    output wire [                                  63:0] m_axi_in_29_ARADDR,
    output wire [                                   1:0] m_axi_in_29_ARBURST,
    output wire [                                   3:0] m_axi_in_29_ARCACHE,
    output wire [                                   0:0] m_axi_in_29_ARID,
    output wire [                                   7:0] m_axi_in_29_ARLEN,
    output wire                                          m_axi_in_29_ARLOCK,
    output wire [                                   2:0] m_axi_in_29_ARPROT,
    output wire [                                   3:0] m_axi_in_29_ARQOS,
    input wire                                           m_axi_in_29_ARREADY,
    output wire [                                   2:0] m_axi_in_29_ARSIZE,
    output wire                                          m_axi_in_29_ARVALID,
    output wire [                                  63:0] m_axi_in_29_AWADDR,
    output wire [                                   1:0] m_axi_in_29_AWBURST,
    output wire [                                   3:0] m_axi_in_29_AWCACHE,
    output wire [                                   0:0] m_axi_in_29_AWID,
    output wire [                                   7:0] m_axi_in_29_AWLEN,
    output wire                                          m_axi_in_29_AWLOCK,
    output wire [                                   2:0] m_axi_in_29_AWPROT,
    output wire [                                   3:0] m_axi_in_29_AWQOS,
    input wire                                           m_axi_in_29_AWREADY,
    output wire [                                   2:0] m_axi_in_29_AWSIZE,
    output wire                                          m_axi_in_29_AWVALID,
    input wire  [                                   0:0] m_axi_in_29_BID,
    output wire                                          m_axi_in_29_BREADY,
    input wire  [                                   1:0] m_axi_in_29_BRESP,
    input wire                                           m_axi_in_29_BVALID,
    input wire  [                                 255:0] m_axi_in_29_RDATA,
    input wire  [                                   0:0] m_axi_in_29_RID,
    input wire                                           m_axi_in_29_RLAST,
    output wire                                          m_axi_in_29_RREADY,
    input wire  [                                   1:0] m_axi_in_29_RRESP,
    input wire                                           m_axi_in_29_RVALID,
    output wire [                                 255:0] m_axi_in_29_WDATA,
    output wire                                          m_axi_in_29_WLAST,
    input wire                                           m_axi_in_29_WREADY,
    output wire [                                  31:0] m_axi_in_29_WSTRB,
    output wire                                          m_axi_in_29_WVALID,
    output wire [                                  63:0] m_axi_in_3_ARADDR,
    output wire [                                   1:0] m_axi_in_3_ARBURST,
    output wire [                                   3:0] m_axi_in_3_ARCACHE,
    output wire [                                   0:0] m_axi_in_3_ARID,
    output wire [                                   7:0] m_axi_in_3_ARLEN,
    output wire                                          m_axi_in_3_ARLOCK,
    output wire [                                   2:0] m_axi_in_3_ARPROT,
    output wire [                                   3:0] m_axi_in_3_ARQOS,
    input wire                                           m_axi_in_3_ARREADY,
    output wire [                                   2:0] m_axi_in_3_ARSIZE,
    output wire                                          m_axi_in_3_ARVALID,
    output wire [                                  63:0] m_axi_in_3_AWADDR,
    output wire [                                   1:0] m_axi_in_3_AWBURST,
    output wire [                                   3:0] m_axi_in_3_AWCACHE,
    output wire [                                   0:0] m_axi_in_3_AWID,
    output wire [                                   7:0] m_axi_in_3_AWLEN,
    output wire                                          m_axi_in_3_AWLOCK,
    output wire [                                   2:0] m_axi_in_3_AWPROT,
    output wire [                                   3:0] m_axi_in_3_AWQOS,
    input wire                                           m_axi_in_3_AWREADY,
    output wire [                                   2:0] m_axi_in_3_AWSIZE,
    output wire                                          m_axi_in_3_AWVALID,
    input wire  [                                   0:0] m_axi_in_3_BID,
    output wire                                          m_axi_in_3_BREADY,
    input wire  [                                   1:0] m_axi_in_3_BRESP,
    input wire                                           m_axi_in_3_BVALID,
    input wire  [                                 255:0] m_axi_in_3_RDATA,
    input wire  [                                   0:0] m_axi_in_3_RID,
    input wire                                           m_axi_in_3_RLAST,
    output wire                                          m_axi_in_3_RREADY,
    input wire  [                                   1:0] m_axi_in_3_RRESP,
    input wire                                           m_axi_in_3_RVALID,
    output wire [                                 255:0] m_axi_in_3_WDATA,
    output wire                                          m_axi_in_3_WLAST,
    input wire                                           m_axi_in_3_WREADY,
    output wire [                                  31:0] m_axi_in_3_WSTRB,
    output wire                                          m_axi_in_3_WVALID,
    output wire [                                  63:0] m_axi_in_30_ARADDR,
    output wire [                                   1:0] m_axi_in_30_ARBURST,
    output wire [                                   3:0] m_axi_in_30_ARCACHE,
    output wire [                                   0:0] m_axi_in_30_ARID,
    output wire [                                   7:0] m_axi_in_30_ARLEN,
    output wire                                          m_axi_in_30_ARLOCK,
    output wire [                                   2:0] m_axi_in_30_ARPROT,
    output wire [                                   3:0] m_axi_in_30_ARQOS,
    input wire                                           m_axi_in_30_ARREADY,
    output wire [                                   2:0] m_axi_in_30_ARSIZE,
    output wire                                          m_axi_in_30_ARVALID,
    output wire [                                  63:0] m_axi_in_30_AWADDR,
    output wire [                                   1:0] m_axi_in_30_AWBURST,
    output wire [                                   3:0] m_axi_in_30_AWCACHE,
    output wire [                                   0:0] m_axi_in_30_AWID,
    output wire [                                   7:0] m_axi_in_30_AWLEN,
    output wire                                          m_axi_in_30_AWLOCK,
    output wire [                                   2:0] m_axi_in_30_AWPROT,
    output wire [                                   3:0] m_axi_in_30_AWQOS,
    input wire                                           m_axi_in_30_AWREADY,
    output wire [                                   2:0] m_axi_in_30_AWSIZE,
    output wire                                          m_axi_in_30_AWVALID,
    input wire  [                                   0:0] m_axi_in_30_BID,
    output wire                                          m_axi_in_30_BREADY,
    input wire  [                                   1:0] m_axi_in_30_BRESP,
    input wire                                           m_axi_in_30_BVALID,
    input wire  [                                 255:0] m_axi_in_30_RDATA,
    input wire  [                                   0:0] m_axi_in_30_RID,
    input wire                                           m_axi_in_30_RLAST,
    output wire                                          m_axi_in_30_RREADY,
    input wire  [                                   1:0] m_axi_in_30_RRESP,
    input wire                                           m_axi_in_30_RVALID,
    output wire [                                 255:0] m_axi_in_30_WDATA,
    output wire                                          m_axi_in_30_WLAST,
    input wire                                           m_axi_in_30_WREADY,
    output wire [                                  31:0] m_axi_in_30_WSTRB,
    output wire                                          m_axi_in_30_WVALID,
    output wire [                                  63:0] m_axi_in_31_ARADDR,
    output wire [                                   1:0] m_axi_in_31_ARBURST,
    output wire [                                   3:0] m_axi_in_31_ARCACHE,
    output wire [                                   0:0] m_axi_in_31_ARID,
    output wire [                                   7:0] m_axi_in_31_ARLEN,
    output wire                                          m_axi_in_31_ARLOCK,
    output wire [                                   2:0] m_axi_in_31_ARPROT,
    output wire [                                   3:0] m_axi_in_31_ARQOS,
    input wire                                           m_axi_in_31_ARREADY,
    output wire [                                   2:0] m_axi_in_31_ARSIZE,
    output wire                                          m_axi_in_31_ARVALID,
    output wire [                                  63:0] m_axi_in_31_AWADDR,
    output wire [                                   1:0] m_axi_in_31_AWBURST,
    output wire [                                   3:0] m_axi_in_31_AWCACHE,
    output wire [                                   0:0] m_axi_in_31_AWID,
    output wire [                                   7:0] m_axi_in_31_AWLEN,
    output wire                                          m_axi_in_31_AWLOCK,
    output wire [                                   2:0] m_axi_in_31_AWPROT,
    output wire [                                   3:0] m_axi_in_31_AWQOS,
    input wire                                           m_axi_in_31_AWREADY,
    output wire [                                   2:0] m_axi_in_31_AWSIZE,
    output wire                                          m_axi_in_31_AWVALID,
    input wire  [                                   0:0] m_axi_in_31_BID,
    output wire                                          m_axi_in_31_BREADY,
    input wire  [                                   1:0] m_axi_in_31_BRESP,
    input wire                                           m_axi_in_31_BVALID,
    input wire  [                                 255:0] m_axi_in_31_RDATA,
    input wire  [                                   0:0] m_axi_in_31_RID,
    input wire                                           m_axi_in_31_RLAST,
    output wire                                          m_axi_in_31_RREADY,
    input wire  [                                   1:0] m_axi_in_31_RRESP,
    input wire                                           m_axi_in_31_RVALID,
    output wire [                                 255:0] m_axi_in_31_WDATA,
    output wire                                          m_axi_in_31_WLAST,
    input wire                                           m_axi_in_31_WREADY,
    output wire [                                  31:0] m_axi_in_31_WSTRB,
    output wire                                          m_axi_in_31_WVALID,
    output wire [                                  63:0] m_axi_in_32_ARADDR,
    output wire [                                   1:0] m_axi_in_32_ARBURST,
    output wire [                                   3:0] m_axi_in_32_ARCACHE,
    output wire [                                   0:0] m_axi_in_32_ARID,
    output wire [                                   7:0] m_axi_in_32_ARLEN,
    output wire                                          m_axi_in_32_ARLOCK,
    output wire [                                   2:0] m_axi_in_32_ARPROT,
    output wire [                                   3:0] m_axi_in_32_ARQOS,
    input wire                                           m_axi_in_32_ARREADY,
    output wire [                                   2:0] m_axi_in_32_ARSIZE,
    output wire                                          m_axi_in_32_ARVALID,
    output wire [                                  63:0] m_axi_in_32_AWADDR,
    output wire [                                   1:0] m_axi_in_32_AWBURST,
    output wire [                                   3:0] m_axi_in_32_AWCACHE,
    output wire [                                   0:0] m_axi_in_32_AWID,
    output wire [                                   7:0] m_axi_in_32_AWLEN,
    output wire                                          m_axi_in_32_AWLOCK,
    output wire [                                   2:0] m_axi_in_32_AWPROT,
    output wire [                                   3:0] m_axi_in_32_AWQOS,
    input wire                                           m_axi_in_32_AWREADY,
    output wire [                                   2:0] m_axi_in_32_AWSIZE,
    output wire                                          m_axi_in_32_AWVALID,
    input wire  [                                   0:0] m_axi_in_32_BID,
    output wire                                          m_axi_in_32_BREADY,
    input wire  [                                   1:0] m_axi_in_32_BRESP,
    input wire                                           m_axi_in_32_BVALID,
    input wire  [                                 255:0] m_axi_in_32_RDATA,
    input wire  [                                   0:0] m_axi_in_32_RID,
    input wire                                           m_axi_in_32_RLAST,
    output wire                                          m_axi_in_32_RREADY,
    input wire  [                                   1:0] m_axi_in_32_RRESP,
    input wire                                           m_axi_in_32_RVALID,
    output wire [                                 255:0] m_axi_in_32_WDATA,
    output wire                                          m_axi_in_32_WLAST,
    input wire                                           m_axi_in_32_WREADY,
    output wire [                                  31:0] m_axi_in_32_WSTRB,
    output wire                                          m_axi_in_32_WVALID,
    output wire [                                  63:0] m_axi_in_33_ARADDR,
    output wire [                                   1:0] m_axi_in_33_ARBURST,
    output wire [                                   3:0] m_axi_in_33_ARCACHE,
    output wire [                                   0:0] m_axi_in_33_ARID,
    output wire [                                   7:0] m_axi_in_33_ARLEN,
    output wire                                          m_axi_in_33_ARLOCK,
    output wire [                                   2:0] m_axi_in_33_ARPROT,
    output wire [                                   3:0] m_axi_in_33_ARQOS,
    input wire                                           m_axi_in_33_ARREADY,
    output wire [                                   2:0] m_axi_in_33_ARSIZE,
    output wire                                          m_axi_in_33_ARVALID,
    output wire [                                  63:0] m_axi_in_33_AWADDR,
    output wire [                                   1:0] m_axi_in_33_AWBURST,
    output wire [                                   3:0] m_axi_in_33_AWCACHE,
    output wire [                                   0:0] m_axi_in_33_AWID,
    output wire [                                   7:0] m_axi_in_33_AWLEN,
    output wire                                          m_axi_in_33_AWLOCK,
    output wire [                                   2:0] m_axi_in_33_AWPROT,
    output wire [                                   3:0] m_axi_in_33_AWQOS,
    input wire                                           m_axi_in_33_AWREADY,
    output wire [                                   2:0] m_axi_in_33_AWSIZE,
    output wire                                          m_axi_in_33_AWVALID,
    input wire  [                                   0:0] m_axi_in_33_BID,
    output wire                                          m_axi_in_33_BREADY,
    input wire  [                                   1:0] m_axi_in_33_BRESP,
    input wire                                           m_axi_in_33_BVALID,
    input wire  [                                 255:0] m_axi_in_33_RDATA,
    input wire  [                                   0:0] m_axi_in_33_RID,
    input wire                                           m_axi_in_33_RLAST,
    output wire                                          m_axi_in_33_RREADY,
    input wire  [                                   1:0] m_axi_in_33_RRESP,
    input wire                                           m_axi_in_33_RVALID,
    output wire [                                 255:0] m_axi_in_33_WDATA,
    output wire                                          m_axi_in_33_WLAST,
    input wire                                           m_axi_in_33_WREADY,
    output wire [                                  31:0] m_axi_in_33_WSTRB,
    output wire                                          m_axi_in_33_WVALID,
    output wire [                                  63:0] m_axi_in_34_ARADDR,
    output wire [                                   1:0] m_axi_in_34_ARBURST,
    output wire [                                   3:0] m_axi_in_34_ARCACHE,
    output wire [                                   0:0] m_axi_in_34_ARID,
    output wire [                                   7:0] m_axi_in_34_ARLEN,
    output wire                                          m_axi_in_34_ARLOCK,
    output wire [                                   2:0] m_axi_in_34_ARPROT,
    output wire [                                   3:0] m_axi_in_34_ARQOS,
    input wire                                           m_axi_in_34_ARREADY,
    output wire [                                   2:0] m_axi_in_34_ARSIZE,
    output wire                                          m_axi_in_34_ARVALID,
    output wire [                                  63:0] m_axi_in_34_AWADDR,
    output wire [                                   1:0] m_axi_in_34_AWBURST,
    output wire [                                   3:0] m_axi_in_34_AWCACHE,
    output wire [                                   0:0] m_axi_in_34_AWID,
    output wire [                                   7:0] m_axi_in_34_AWLEN,
    output wire                                          m_axi_in_34_AWLOCK,
    output wire [                                   2:0] m_axi_in_34_AWPROT,
    output wire [                                   3:0] m_axi_in_34_AWQOS,
    input wire                                           m_axi_in_34_AWREADY,
    output wire [                                   2:0] m_axi_in_34_AWSIZE,
    output wire                                          m_axi_in_34_AWVALID,
    input wire  [                                   0:0] m_axi_in_34_BID,
    output wire                                          m_axi_in_34_BREADY,
    input wire  [                                   1:0] m_axi_in_34_BRESP,
    input wire                                           m_axi_in_34_BVALID,
    input wire  [                                 255:0] m_axi_in_34_RDATA,
    input wire  [                                   0:0] m_axi_in_34_RID,
    input wire                                           m_axi_in_34_RLAST,
    output wire                                          m_axi_in_34_RREADY,
    input wire  [                                   1:0] m_axi_in_34_RRESP,
    input wire                                           m_axi_in_34_RVALID,
    output wire [                                 255:0] m_axi_in_34_WDATA,
    output wire                                          m_axi_in_34_WLAST,
    input wire                                           m_axi_in_34_WREADY,
    output wire [                                  31:0] m_axi_in_34_WSTRB,
    output wire                                          m_axi_in_34_WVALID,
    output wire [                                  63:0] m_axi_in_35_ARADDR,
    output wire [                                   1:0] m_axi_in_35_ARBURST,
    output wire [                                   3:0] m_axi_in_35_ARCACHE,
    output wire [                                   0:0] m_axi_in_35_ARID,
    output wire [                                   7:0] m_axi_in_35_ARLEN,
    output wire                                          m_axi_in_35_ARLOCK,
    output wire [                                   2:0] m_axi_in_35_ARPROT,
    output wire [                                   3:0] m_axi_in_35_ARQOS,
    input wire                                           m_axi_in_35_ARREADY,
    output wire [                                   2:0] m_axi_in_35_ARSIZE,
    output wire                                          m_axi_in_35_ARVALID,
    output wire [                                  63:0] m_axi_in_35_AWADDR,
    output wire [                                   1:0] m_axi_in_35_AWBURST,
    output wire [                                   3:0] m_axi_in_35_AWCACHE,
    output wire [                                   0:0] m_axi_in_35_AWID,
    output wire [                                   7:0] m_axi_in_35_AWLEN,
    output wire                                          m_axi_in_35_AWLOCK,
    output wire [                                   2:0] m_axi_in_35_AWPROT,
    output wire [                                   3:0] m_axi_in_35_AWQOS,
    input wire                                           m_axi_in_35_AWREADY,
    output wire [                                   2:0] m_axi_in_35_AWSIZE,
    output wire                                          m_axi_in_35_AWVALID,
    input wire  [                                   0:0] m_axi_in_35_BID,
    output wire                                          m_axi_in_35_BREADY,
    input wire  [                                   1:0] m_axi_in_35_BRESP,
    input wire                                           m_axi_in_35_BVALID,
    input wire  [                                 255:0] m_axi_in_35_RDATA,
    input wire  [                                   0:0] m_axi_in_35_RID,
    input wire                                           m_axi_in_35_RLAST,
    output wire                                          m_axi_in_35_RREADY,
    input wire  [                                   1:0] m_axi_in_35_RRESP,
    input wire                                           m_axi_in_35_RVALID,
    output wire [                                 255:0] m_axi_in_35_WDATA,
    output wire                                          m_axi_in_35_WLAST,
    input wire                                           m_axi_in_35_WREADY,
    output wire [                                  31:0] m_axi_in_35_WSTRB,
    output wire                                          m_axi_in_35_WVALID,
    output wire [                                  63:0] m_axi_in_36_ARADDR,
    output wire [                                   1:0] m_axi_in_36_ARBURST,
    output wire [                                   3:0] m_axi_in_36_ARCACHE,
    output wire [                                   0:0] m_axi_in_36_ARID,
    output wire [                                   7:0] m_axi_in_36_ARLEN,
    output wire                                          m_axi_in_36_ARLOCK,
    output wire [                                   2:0] m_axi_in_36_ARPROT,
    output wire [                                   3:0] m_axi_in_36_ARQOS,
    input wire                                           m_axi_in_36_ARREADY,
    output wire [                                   2:0] m_axi_in_36_ARSIZE,
    output wire                                          m_axi_in_36_ARVALID,
    output wire [                                  63:0] m_axi_in_36_AWADDR,
    output wire [                                   1:0] m_axi_in_36_AWBURST,
    output wire [                                   3:0] m_axi_in_36_AWCACHE,
    output wire [                                   0:0] m_axi_in_36_AWID,
    output wire [                                   7:0] m_axi_in_36_AWLEN,
    output wire                                          m_axi_in_36_AWLOCK,
    output wire [                                   2:0] m_axi_in_36_AWPROT,
    output wire [                                   3:0] m_axi_in_36_AWQOS,
    input wire                                           m_axi_in_36_AWREADY,
    output wire [                                   2:0] m_axi_in_36_AWSIZE,
    output wire                                          m_axi_in_36_AWVALID,
    input wire  [                                   0:0] m_axi_in_36_BID,
    output wire                                          m_axi_in_36_BREADY,
    input wire  [                                   1:0] m_axi_in_36_BRESP,
    input wire                                           m_axi_in_36_BVALID,
    input wire  [                                 255:0] m_axi_in_36_RDATA,
    input wire  [                                   0:0] m_axi_in_36_RID,
    input wire                                           m_axi_in_36_RLAST,
    output wire                                          m_axi_in_36_RREADY,
    input wire  [                                   1:0] m_axi_in_36_RRESP,
    input wire                                           m_axi_in_36_RVALID,
    output wire [                                 255:0] m_axi_in_36_WDATA,
    output wire                                          m_axi_in_36_WLAST,
    input wire                                           m_axi_in_36_WREADY,
    output wire [                                  31:0] m_axi_in_36_WSTRB,
    output wire                                          m_axi_in_36_WVALID,
    output wire [                                  63:0] m_axi_in_37_ARADDR,
    output wire [                                   1:0] m_axi_in_37_ARBURST,
    output wire [                                   3:0] m_axi_in_37_ARCACHE,
    output wire [                                   0:0] m_axi_in_37_ARID,
    output wire [                                   7:0] m_axi_in_37_ARLEN,
    output wire                                          m_axi_in_37_ARLOCK,
    output wire [                                   2:0] m_axi_in_37_ARPROT,
    output wire [                                   3:0] m_axi_in_37_ARQOS,
    input wire                                           m_axi_in_37_ARREADY,
    output wire [                                   2:0] m_axi_in_37_ARSIZE,
    output wire                                          m_axi_in_37_ARVALID,
    output wire [                                  63:0] m_axi_in_37_AWADDR,
    output wire [                                   1:0] m_axi_in_37_AWBURST,
    output wire [                                   3:0] m_axi_in_37_AWCACHE,
    output wire [                                   0:0] m_axi_in_37_AWID,
    output wire [                                   7:0] m_axi_in_37_AWLEN,
    output wire                                          m_axi_in_37_AWLOCK,
    output wire [                                   2:0] m_axi_in_37_AWPROT,
    output wire [                                   3:0] m_axi_in_37_AWQOS,
    input wire                                           m_axi_in_37_AWREADY,
    output wire [                                   2:0] m_axi_in_37_AWSIZE,
    output wire                                          m_axi_in_37_AWVALID,
    input wire  [                                   0:0] m_axi_in_37_BID,
    output wire                                          m_axi_in_37_BREADY,
    input wire  [                                   1:0] m_axi_in_37_BRESP,
    input wire                                           m_axi_in_37_BVALID,
    input wire  [                                 255:0] m_axi_in_37_RDATA,
    input wire  [                                   0:0] m_axi_in_37_RID,
    input wire                                           m_axi_in_37_RLAST,
    output wire                                          m_axi_in_37_RREADY,
    input wire  [                                   1:0] m_axi_in_37_RRESP,
    input wire                                           m_axi_in_37_RVALID,
    output wire [                                 255:0] m_axi_in_37_WDATA,
    output wire                                          m_axi_in_37_WLAST,
    input wire                                           m_axi_in_37_WREADY,
    output wire [                                  31:0] m_axi_in_37_WSTRB,
    output wire                                          m_axi_in_37_WVALID,
    output wire [                                  63:0] m_axi_in_38_ARADDR,
    output wire [                                   1:0] m_axi_in_38_ARBURST,
    output wire [                                   3:0] m_axi_in_38_ARCACHE,
    output wire [                                   0:0] m_axi_in_38_ARID,
    output wire [                                   7:0] m_axi_in_38_ARLEN,
    output wire                                          m_axi_in_38_ARLOCK,
    output wire [                                   2:0] m_axi_in_38_ARPROT,
    output wire [                                   3:0] m_axi_in_38_ARQOS,
    input wire                                           m_axi_in_38_ARREADY,
    output wire [                                   2:0] m_axi_in_38_ARSIZE,
    output wire                                          m_axi_in_38_ARVALID,
    output wire [                                  63:0] m_axi_in_38_AWADDR,
    output wire [                                   1:0] m_axi_in_38_AWBURST,
    output wire [                                   3:0] m_axi_in_38_AWCACHE,
    output wire [                                   0:0] m_axi_in_38_AWID,
    output wire [                                   7:0] m_axi_in_38_AWLEN,
    output wire                                          m_axi_in_38_AWLOCK,
    output wire [                                   2:0] m_axi_in_38_AWPROT,
    output wire [                                   3:0] m_axi_in_38_AWQOS,
    input wire                                           m_axi_in_38_AWREADY,
    output wire [                                   2:0] m_axi_in_38_AWSIZE,
    output wire                                          m_axi_in_38_AWVALID,
    input wire  [                                   0:0] m_axi_in_38_BID,
    output wire                                          m_axi_in_38_BREADY,
    input wire  [                                   1:0] m_axi_in_38_BRESP,
    input wire                                           m_axi_in_38_BVALID,
    input wire  [                                 255:0] m_axi_in_38_RDATA,
    input wire  [                                   0:0] m_axi_in_38_RID,
    input wire                                           m_axi_in_38_RLAST,
    output wire                                          m_axi_in_38_RREADY,
    input wire  [                                   1:0] m_axi_in_38_RRESP,
    input wire                                           m_axi_in_38_RVALID,
    output wire [                                 255:0] m_axi_in_38_WDATA,
    output wire                                          m_axi_in_38_WLAST,
    input wire                                           m_axi_in_38_WREADY,
    output wire [                                  31:0] m_axi_in_38_WSTRB,
    output wire                                          m_axi_in_38_WVALID,
    output wire [                                  63:0] m_axi_in_39_ARADDR,
    output wire [                                   1:0] m_axi_in_39_ARBURST,
    output wire [                                   3:0] m_axi_in_39_ARCACHE,
    output wire [                                   0:0] m_axi_in_39_ARID,
    output wire [                                   7:0] m_axi_in_39_ARLEN,
    output wire                                          m_axi_in_39_ARLOCK,
    output wire [                                   2:0] m_axi_in_39_ARPROT,
    output wire [                                   3:0] m_axi_in_39_ARQOS,
    input wire                                           m_axi_in_39_ARREADY,
    output wire [                                   2:0] m_axi_in_39_ARSIZE,
    output wire                                          m_axi_in_39_ARVALID,
    output wire [                                  63:0] m_axi_in_39_AWADDR,
    output wire [                                   1:0] m_axi_in_39_AWBURST,
    output wire [                                   3:0] m_axi_in_39_AWCACHE,
    output wire [                                   0:0] m_axi_in_39_AWID,
    output wire [                                   7:0] m_axi_in_39_AWLEN,
    output wire                                          m_axi_in_39_AWLOCK,
    output wire [                                   2:0] m_axi_in_39_AWPROT,
    output wire [                                   3:0] m_axi_in_39_AWQOS,
    input wire                                           m_axi_in_39_AWREADY,
    output wire [                                   2:0] m_axi_in_39_AWSIZE,
    output wire                                          m_axi_in_39_AWVALID,
    input wire  [                                   0:0] m_axi_in_39_BID,
    output wire                                          m_axi_in_39_BREADY,
    input wire  [                                   1:0] m_axi_in_39_BRESP,
    input wire                                           m_axi_in_39_BVALID,
    input wire  [                                 255:0] m_axi_in_39_RDATA,
    input wire  [                                   0:0] m_axi_in_39_RID,
    input wire                                           m_axi_in_39_RLAST,
    output wire                                          m_axi_in_39_RREADY,
    input wire  [                                   1:0] m_axi_in_39_RRESP,
    input wire                                           m_axi_in_39_RVALID,
    output wire [                                 255:0] m_axi_in_39_WDATA,
    output wire                                          m_axi_in_39_WLAST,
    input wire                                           m_axi_in_39_WREADY,
    output wire [                                  31:0] m_axi_in_39_WSTRB,
    output wire                                          m_axi_in_39_WVALID,
    output wire [                                  63:0] m_axi_in_4_ARADDR,
    output wire [                                   1:0] m_axi_in_4_ARBURST,
    output wire [                                   3:0] m_axi_in_4_ARCACHE,
    output wire [                                   0:0] m_axi_in_4_ARID,
    output wire [                                   7:0] m_axi_in_4_ARLEN,
    output wire                                          m_axi_in_4_ARLOCK,
    output wire [                                   2:0] m_axi_in_4_ARPROT,
    output wire [                                   3:0] m_axi_in_4_ARQOS,
    input wire                                           m_axi_in_4_ARREADY,
    output wire [                                   2:0] m_axi_in_4_ARSIZE,
    output wire                                          m_axi_in_4_ARVALID,
    output wire [                                  63:0] m_axi_in_4_AWADDR,
    output wire [                                   1:0] m_axi_in_4_AWBURST,
    output wire [                                   3:0] m_axi_in_4_AWCACHE,
    output wire [                                   0:0] m_axi_in_4_AWID,
    output wire [                                   7:0] m_axi_in_4_AWLEN,
    output wire                                          m_axi_in_4_AWLOCK,
    output wire [                                   2:0] m_axi_in_4_AWPROT,
    output wire [                                   3:0] m_axi_in_4_AWQOS,
    input wire                                           m_axi_in_4_AWREADY,
    output wire [                                   2:0] m_axi_in_4_AWSIZE,
    output wire                                          m_axi_in_4_AWVALID,
    input wire  [                                   0:0] m_axi_in_4_BID,
    output wire                                          m_axi_in_4_BREADY,
    input wire  [                                   1:0] m_axi_in_4_BRESP,
    input wire                                           m_axi_in_4_BVALID,
    input wire  [                                 255:0] m_axi_in_4_RDATA,
    input wire  [                                   0:0] m_axi_in_4_RID,
    input wire                                           m_axi_in_4_RLAST,
    output wire                                          m_axi_in_4_RREADY,
    input wire  [                                   1:0] m_axi_in_4_RRESP,
    input wire                                           m_axi_in_4_RVALID,
    output wire [                                 255:0] m_axi_in_4_WDATA,
    output wire                                          m_axi_in_4_WLAST,
    input wire                                           m_axi_in_4_WREADY,
    output wire [                                  31:0] m_axi_in_4_WSTRB,
    output wire                                          m_axi_in_4_WVALID,
    output wire [                                  63:0] m_axi_in_40_ARADDR,
    output wire [                                   1:0] m_axi_in_40_ARBURST,
    output wire [                                   3:0] m_axi_in_40_ARCACHE,
    output wire [                                   0:0] m_axi_in_40_ARID,
    output wire [                                   7:0] m_axi_in_40_ARLEN,
    output wire                                          m_axi_in_40_ARLOCK,
    output wire [                                   2:0] m_axi_in_40_ARPROT,
    output wire [                                   3:0] m_axi_in_40_ARQOS,
    input wire                                           m_axi_in_40_ARREADY,
    output wire [                                   2:0] m_axi_in_40_ARSIZE,
    output wire                                          m_axi_in_40_ARVALID,
    output wire [                                  63:0] m_axi_in_40_AWADDR,
    output wire [                                   1:0] m_axi_in_40_AWBURST,
    output wire [                                   3:0] m_axi_in_40_AWCACHE,
    output wire [                                   0:0] m_axi_in_40_AWID,
    output wire [                                   7:0] m_axi_in_40_AWLEN,
    output wire                                          m_axi_in_40_AWLOCK,
    output wire [                                   2:0] m_axi_in_40_AWPROT,
    output wire [                                   3:0] m_axi_in_40_AWQOS,
    input wire                                           m_axi_in_40_AWREADY,
    output wire [                                   2:0] m_axi_in_40_AWSIZE,
    output wire                                          m_axi_in_40_AWVALID,
    input wire  [                                   0:0] m_axi_in_40_BID,
    output wire                                          m_axi_in_40_BREADY,
    input wire  [                                   1:0] m_axi_in_40_BRESP,
    input wire                                           m_axi_in_40_BVALID,
    input wire  [                                 255:0] m_axi_in_40_RDATA,
    input wire  [                                   0:0] m_axi_in_40_RID,
    input wire                                           m_axi_in_40_RLAST,
    output wire                                          m_axi_in_40_RREADY,
    input wire  [                                   1:0] m_axi_in_40_RRESP,
    input wire                                           m_axi_in_40_RVALID,
    output wire [                                 255:0] m_axi_in_40_WDATA,
    output wire                                          m_axi_in_40_WLAST,
    input wire                                           m_axi_in_40_WREADY,
    output wire [                                  31:0] m_axi_in_40_WSTRB,
    output wire                                          m_axi_in_40_WVALID,
    output wire [                                  63:0] m_axi_in_41_ARADDR,
    output wire [                                   1:0] m_axi_in_41_ARBURST,
    output wire [                                   3:0] m_axi_in_41_ARCACHE,
    output wire [                                   0:0] m_axi_in_41_ARID,
    output wire [                                   7:0] m_axi_in_41_ARLEN,
    output wire                                          m_axi_in_41_ARLOCK,
    output wire [                                   2:0] m_axi_in_41_ARPROT,
    output wire [                                   3:0] m_axi_in_41_ARQOS,
    input wire                                           m_axi_in_41_ARREADY,
    output wire [                                   2:0] m_axi_in_41_ARSIZE,
    output wire                                          m_axi_in_41_ARVALID,
    output wire [                                  63:0] m_axi_in_41_AWADDR,
    output wire [                                   1:0] m_axi_in_41_AWBURST,
    output wire [                                   3:0] m_axi_in_41_AWCACHE,
    output wire [                                   0:0] m_axi_in_41_AWID,
    output wire [                                   7:0] m_axi_in_41_AWLEN,
    output wire                                          m_axi_in_41_AWLOCK,
    output wire [                                   2:0] m_axi_in_41_AWPROT,
    output wire [                                   3:0] m_axi_in_41_AWQOS,
    input wire                                           m_axi_in_41_AWREADY,
    output wire [                                   2:0] m_axi_in_41_AWSIZE,
    output wire                                          m_axi_in_41_AWVALID,
    input wire  [                                   0:0] m_axi_in_41_BID,
    output wire                                          m_axi_in_41_BREADY,
    input wire  [                                   1:0] m_axi_in_41_BRESP,
    input wire                                           m_axi_in_41_BVALID,
    input wire  [                                 255:0] m_axi_in_41_RDATA,
    input wire  [                                   0:0] m_axi_in_41_RID,
    input wire                                           m_axi_in_41_RLAST,
    output wire                                          m_axi_in_41_RREADY,
    input wire  [                                   1:0] m_axi_in_41_RRESP,
    input wire                                           m_axi_in_41_RVALID,
    output wire [                                 255:0] m_axi_in_41_WDATA,
    output wire                                          m_axi_in_41_WLAST,
    input wire                                           m_axi_in_41_WREADY,
    output wire [                                  31:0] m_axi_in_41_WSTRB,
    output wire                                          m_axi_in_41_WVALID,
    output wire [                                  63:0] m_axi_in_42_ARADDR,
    output wire [                                   1:0] m_axi_in_42_ARBURST,
    output wire [                                   3:0] m_axi_in_42_ARCACHE,
    output wire [                                   0:0] m_axi_in_42_ARID,
    output wire [                                   7:0] m_axi_in_42_ARLEN,
    output wire                                          m_axi_in_42_ARLOCK,
    output wire [                                   2:0] m_axi_in_42_ARPROT,
    output wire [                                   3:0] m_axi_in_42_ARQOS,
    input wire                                           m_axi_in_42_ARREADY,
    output wire [                                   2:0] m_axi_in_42_ARSIZE,
    output wire                                          m_axi_in_42_ARVALID,
    output wire [                                  63:0] m_axi_in_42_AWADDR,
    output wire [                                   1:0] m_axi_in_42_AWBURST,
    output wire [                                   3:0] m_axi_in_42_AWCACHE,
    output wire [                                   0:0] m_axi_in_42_AWID,
    output wire [                                   7:0] m_axi_in_42_AWLEN,
    output wire                                          m_axi_in_42_AWLOCK,
    output wire [                                   2:0] m_axi_in_42_AWPROT,
    output wire [                                   3:0] m_axi_in_42_AWQOS,
    input wire                                           m_axi_in_42_AWREADY,
    output wire [                                   2:0] m_axi_in_42_AWSIZE,
    output wire                                          m_axi_in_42_AWVALID,
    input wire  [                                   0:0] m_axi_in_42_BID,
    output wire                                          m_axi_in_42_BREADY,
    input wire  [                                   1:0] m_axi_in_42_BRESP,
    input wire                                           m_axi_in_42_BVALID,
    input wire  [                                 255:0] m_axi_in_42_RDATA,
    input wire  [                                   0:0] m_axi_in_42_RID,
    input wire                                           m_axi_in_42_RLAST,
    output wire                                          m_axi_in_42_RREADY,
    input wire  [                                   1:0] m_axi_in_42_RRESP,
    input wire                                           m_axi_in_42_RVALID,
    output wire [                                 255:0] m_axi_in_42_WDATA,
    output wire                                          m_axi_in_42_WLAST,
    input wire                                           m_axi_in_42_WREADY,
    output wire [                                  31:0] m_axi_in_42_WSTRB,
    output wire                                          m_axi_in_42_WVALID,
    output wire [                                  63:0] m_axi_in_43_ARADDR,
    output wire [                                   1:0] m_axi_in_43_ARBURST,
    output wire [                                   3:0] m_axi_in_43_ARCACHE,
    output wire [                                   0:0] m_axi_in_43_ARID,
    output wire [                                   7:0] m_axi_in_43_ARLEN,
    output wire                                          m_axi_in_43_ARLOCK,
    output wire [                                   2:0] m_axi_in_43_ARPROT,
    output wire [                                   3:0] m_axi_in_43_ARQOS,
    input wire                                           m_axi_in_43_ARREADY,
    output wire [                                   2:0] m_axi_in_43_ARSIZE,
    output wire                                          m_axi_in_43_ARVALID,
    output wire [                                  63:0] m_axi_in_43_AWADDR,
    output wire [                                   1:0] m_axi_in_43_AWBURST,
    output wire [                                   3:0] m_axi_in_43_AWCACHE,
    output wire [                                   0:0] m_axi_in_43_AWID,
    output wire [                                   7:0] m_axi_in_43_AWLEN,
    output wire                                          m_axi_in_43_AWLOCK,
    output wire [                                   2:0] m_axi_in_43_AWPROT,
    output wire [                                   3:0] m_axi_in_43_AWQOS,
    input wire                                           m_axi_in_43_AWREADY,
    output wire [                                   2:0] m_axi_in_43_AWSIZE,
    output wire                                          m_axi_in_43_AWVALID,
    input wire  [                                   0:0] m_axi_in_43_BID,
    output wire                                          m_axi_in_43_BREADY,
    input wire  [                                   1:0] m_axi_in_43_BRESP,
    input wire                                           m_axi_in_43_BVALID,
    input wire  [                                 255:0] m_axi_in_43_RDATA,
    input wire  [                                   0:0] m_axi_in_43_RID,
    input wire                                           m_axi_in_43_RLAST,
    output wire                                          m_axi_in_43_RREADY,
    input wire  [                                   1:0] m_axi_in_43_RRESP,
    input wire                                           m_axi_in_43_RVALID,
    output wire [                                 255:0] m_axi_in_43_WDATA,
    output wire                                          m_axi_in_43_WLAST,
    input wire                                           m_axi_in_43_WREADY,
    output wire [                                  31:0] m_axi_in_43_WSTRB,
    output wire                                          m_axi_in_43_WVALID,
    output wire [                                  63:0] m_axi_in_44_ARADDR,
    output wire [                                   1:0] m_axi_in_44_ARBURST,
    output wire [                                   3:0] m_axi_in_44_ARCACHE,
    output wire [                                   0:0] m_axi_in_44_ARID,
    output wire [                                   7:0] m_axi_in_44_ARLEN,
    output wire                                          m_axi_in_44_ARLOCK,
    output wire [                                   2:0] m_axi_in_44_ARPROT,
    output wire [                                   3:0] m_axi_in_44_ARQOS,
    input wire                                           m_axi_in_44_ARREADY,
    output wire [                                   2:0] m_axi_in_44_ARSIZE,
    output wire                                          m_axi_in_44_ARVALID,
    output wire [                                  63:0] m_axi_in_44_AWADDR,
    output wire [                                   1:0] m_axi_in_44_AWBURST,
    output wire [                                   3:0] m_axi_in_44_AWCACHE,
    output wire [                                   0:0] m_axi_in_44_AWID,
    output wire [                                   7:0] m_axi_in_44_AWLEN,
    output wire                                          m_axi_in_44_AWLOCK,
    output wire [                                   2:0] m_axi_in_44_AWPROT,
    output wire [                                   3:0] m_axi_in_44_AWQOS,
    input wire                                           m_axi_in_44_AWREADY,
    output wire [                                   2:0] m_axi_in_44_AWSIZE,
    output wire                                          m_axi_in_44_AWVALID,
    input wire  [                                   0:0] m_axi_in_44_BID,
    output wire                                          m_axi_in_44_BREADY,
    input wire  [                                   1:0] m_axi_in_44_BRESP,
    input wire                                           m_axi_in_44_BVALID,
    input wire  [                                 255:0] m_axi_in_44_RDATA,
    input wire  [                                   0:0] m_axi_in_44_RID,
    input wire                                           m_axi_in_44_RLAST,
    output wire                                          m_axi_in_44_RREADY,
    input wire  [                                   1:0] m_axi_in_44_RRESP,
    input wire                                           m_axi_in_44_RVALID,
    output wire [                                 255:0] m_axi_in_44_WDATA,
    output wire                                          m_axi_in_44_WLAST,
    input wire                                           m_axi_in_44_WREADY,
    output wire [                                  31:0] m_axi_in_44_WSTRB,
    output wire                                          m_axi_in_44_WVALID,
    output wire [                                  63:0] m_axi_in_45_ARADDR,
    output wire [                                   1:0] m_axi_in_45_ARBURST,
    output wire [                                   3:0] m_axi_in_45_ARCACHE,
    output wire [                                   0:0] m_axi_in_45_ARID,
    output wire [                                   7:0] m_axi_in_45_ARLEN,
    output wire                                          m_axi_in_45_ARLOCK,
    output wire [                                   2:0] m_axi_in_45_ARPROT,
    output wire [                                   3:0] m_axi_in_45_ARQOS,
    input wire                                           m_axi_in_45_ARREADY,
    output wire [                                   2:0] m_axi_in_45_ARSIZE,
    output wire                                          m_axi_in_45_ARVALID,
    output wire [                                  63:0] m_axi_in_45_AWADDR,
    output wire [                                   1:0] m_axi_in_45_AWBURST,
    output wire [                                   3:0] m_axi_in_45_AWCACHE,
    output wire [                                   0:0] m_axi_in_45_AWID,
    output wire [                                   7:0] m_axi_in_45_AWLEN,
    output wire                                          m_axi_in_45_AWLOCK,
    output wire [                                   2:0] m_axi_in_45_AWPROT,
    output wire [                                   3:0] m_axi_in_45_AWQOS,
    input wire                                           m_axi_in_45_AWREADY,
    output wire [                                   2:0] m_axi_in_45_AWSIZE,
    output wire                                          m_axi_in_45_AWVALID,
    input wire  [                                   0:0] m_axi_in_45_BID,
    output wire                                          m_axi_in_45_BREADY,
    input wire  [                                   1:0] m_axi_in_45_BRESP,
    input wire                                           m_axi_in_45_BVALID,
    input wire  [                                 255:0] m_axi_in_45_RDATA,
    input wire  [                                   0:0] m_axi_in_45_RID,
    input wire                                           m_axi_in_45_RLAST,
    output wire                                          m_axi_in_45_RREADY,
    input wire  [                                   1:0] m_axi_in_45_RRESP,
    input wire                                           m_axi_in_45_RVALID,
    output wire [                                 255:0] m_axi_in_45_WDATA,
    output wire                                          m_axi_in_45_WLAST,
    input wire                                           m_axi_in_45_WREADY,
    output wire [                                  31:0] m_axi_in_45_WSTRB,
    output wire                                          m_axi_in_45_WVALID,
    output wire [                                  63:0] m_axi_in_46_ARADDR,
    output wire [                                   1:0] m_axi_in_46_ARBURST,
    output wire [                                   3:0] m_axi_in_46_ARCACHE,
    output wire [                                   0:0] m_axi_in_46_ARID,
    output wire [                                   7:0] m_axi_in_46_ARLEN,
    output wire                                          m_axi_in_46_ARLOCK,
    output wire [                                   2:0] m_axi_in_46_ARPROT,
    output wire [                                   3:0] m_axi_in_46_ARQOS,
    input wire                                           m_axi_in_46_ARREADY,
    output wire [                                   2:0] m_axi_in_46_ARSIZE,
    output wire                                          m_axi_in_46_ARVALID,
    output wire [                                  63:0] m_axi_in_46_AWADDR,
    output wire [                                   1:0] m_axi_in_46_AWBURST,
    output wire [                                   3:0] m_axi_in_46_AWCACHE,
    output wire [                                   0:0] m_axi_in_46_AWID,
    output wire [                                   7:0] m_axi_in_46_AWLEN,
    output wire                                          m_axi_in_46_AWLOCK,
    output wire [                                   2:0] m_axi_in_46_AWPROT,
    output wire [                                   3:0] m_axi_in_46_AWQOS,
    input wire                                           m_axi_in_46_AWREADY,
    output wire [                                   2:0] m_axi_in_46_AWSIZE,
    output wire                                          m_axi_in_46_AWVALID,
    input wire  [                                   0:0] m_axi_in_46_BID,
    output wire                                          m_axi_in_46_BREADY,
    input wire  [                                   1:0] m_axi_in_46_BRESP,
    input wire                                           m_axi_in_46_BVALID,
    input wire  [                                 255:0] m_axi_in_46_RDATA,
    input wire  [                                   0:0] m_axi_in_46_RID,
    input wire                                           m_axi_in_46_RLAST,
    output wire                                          m_axi_in_46_RREADY,
    input wire  [                                   1:0] m_axi_in_46_RRESP,
    input wire                                           m_axi_in_46_RVALID,
    output wire [                                 255:0] m_axi_in_46_WDATA,
    output wire                                          m_axi_in_46_WLAST,
    input wire                                           m_axi_in_46_WREADY,
    output wire [                                  31:0] m_axi_in_46_WSTRB,
    output wire                                          m_axi_in_46_WVALID,
    output wire [                                  63:0] m_axi_in_47_ARADDR,
    output wire [                                   1:0] m_axi_in_47_ARBURST,
    output wire [                                   3:0] m_axi_in_47_ARCACHE,
    output wire [                                   0:0] m_axi_in_47_ARID,
    output wire [                                   7:0] m_axi_in_47_ARLEN,
    output wire                                          m_axi_in_47_ARLOCK,
    output wire [                                   2:0] m_axi_in_47_ARPROT,
    output wire [                                   3:0] m_axi_in_47_ARQOS,
    input wire                                           m_axi_in_47_ARREADY,
    output wire [                                   2:0] m_axi_in_47_ARSIZE,
    output wire                                          m_axi_in_47_ARVALID,
    output wire [                                  63:0] m_axi_in_47_AWADDR,
    output wire [                                   1:0] m_axi_in_47_AWBURST,
    output wire [                                   3:0] m_axi_in_47_AWCACHE,
    output wire [                                   0:0] m_axi_in_47_AWID,
    output wire [                                   7:0] m_axi_in_47_AWLEN,
    output wire                                          m_axi_in_47_AWLOCK,
    output wire [                                   2:0] m_axi_in_47_AWPROT,
    output wire [                                   3:0] m_axi_in_47_AWQOS,
    input wire                                           m_axi_in_47_AWREADY,
    output wire [                                   2:0] m_axi_in_47_AWSIZE,
    output wire                                          m_axi_in_47_AWVALID,
    input wire  [                                   0:0] m_axi_in_47_BID,
    output wire                                          m_axi_in_47_BREADY,
    input wire  [                                   1:0] m_axi_in_47_BRESP,
    input wire                                           m_axi_in_47_BVALID,
    input wire  [                                 255:0] m_axi_in_47_RDATA,
    input wire  [                                   0:0] m_axi_in_47_RID,
    input wire                                           m_axi_in_47_RLAST,
    output wire                                          m_axi_in_47_RREADY,
    input wire  [                                   1:0] m_axi_in_47_RRESP,
    input wire                                           m_axi_in_47_RVALID,
    output wire [                                 255:0] m_axi_in_47_WDATA,
    output wire                                          m_axi_in_47_WLAST,
    input wire                                           m_axi_in_47_WREADY,
    output wire [                                  31:0] m_axi_in_47_WSTRB,
    output wire                                          m_axi_in_47_WVALID,
    output wire [                                  63:0] m_axi_in_48_ARADDR,
    output wire [                                   1:0] m_axi_in_48_ARBURST,
    output wire [                                   3:0] m_axi_in_48_ARCACHE,
    output wire [                                   0:0] m_axi_in_48_ARID,
    output wire [                                   7:0] m_axi_in_48_ARLEN,
    output wire                                          m_axi_in_48_ARLOCK,
    output wire [                                   2:0] m_axi_in_48_ARPROT,
    output wire [                                   3:0] m_axi_in_48_ARQOS,
    input wire                                           m_axi_in_48_ARREADY,
    output wire [                                   2:0] m_axi_in_48_ARSIZE,
    output wire                                          m_axi_in_48_ARVALID,
    output wire [                                  63:0] m_axi_in_48_AWADDR,
    output wire [                                   1:0] m_axi_in_48_AWBURST,
    output wire [                                   3:0] m_axi_in_48_AWCACHE,
    output wire [                                   0:0] m_axi_in_48_AWID,
    output wire [                                   7:0] m_axi_in_48_AWLEN,
    output wire                                          m_axi_in_48_AWLOCK,
    output wire [                                   2:0] m_axi_in_48_AWPROT,
    output wire [                                   3:0] m_axi_in_48_AWQOS,
    input wire                                           m_axi_in_48_AWREADY,
    output wire [                                   2:0] m_axi_in_48_AWSIZE,
    output wire                                          m_axi_in_48_AWVALID,
    input wire  [                                   0:0] m_axi_in_48_BID,
    output wire                                          m_axi_in_48_BREADY,
    input wire  [                                   1:0] m_axi_in_48_BRESP,
    input wire                                           m_axi_in_48_BVALID,
    input wire  [                                 255:0] m_axi_in_48_RDATA,
    input wire  [                                   0:0] m_axi_in_48_RID,
    input wire                                           m_axi_in_48_RLAST,
    output wire                                          m_axi_in_48_RREADY,
    input wire  [                                   1:0] m_axi_in_48_RRESP,
    input wire                                           m_axi_in_48_RVALID,
    output wire [                                 255:0] m_axi_in_48_WDATA,
    output wire                                          m_axi_in_48_WLAST,
    input wire                                           m_axi_in_48_WREADY,
    output wire [                                  31:0] m_axi_in_48_WSTRB,
    output wire                                          m_axi_in_48_WVALID,
    output wire [                                  63:0] m_axi_in_49_ARADDR,
    output wire [                                   1:0] m_axi_in_49_ARBURST,
    output wire [                                   3:0] m_axi_in_49_ARCACHE,
    output wire [                                   0:0] m_axi_in_49_ARID,
    output wire [                                   7:0] m_axi_in_49_ARLEN,
    output wire                                          m_axi_in_49_ARLOCK,
    output wire [                                   2:0] m_axi_in_49_ARPROT,
    output wire [                                   3:0] m_axi_in_49_ARQOS,
    input wire                                           m_axi_in_49_ARREADY,
    output wire [                                   2:0] m_axi_in_49_ARSIZE,
    output wire                                          m_axi_in_49_ARVALID,
    output wire [                                  63:0] m_axi_in_49_AWADDR,
    output wire [                                   1:0] m_axi_in_49_AWBURST,
    output wire [                                   3:0] m_axi_in_49_AWCACHE,
    output wire [                                   0:0] m_axi_in_49_AWID,
    output wire [                                   7:0] m_axi_in_49_AWLEN,
    output wire                                          m_axi_in_49_AWLOCK,
    output wire [                                   2:0] m_axi_in_49_AWPROT,
    output wire [                                   3:0] m_axi_in_49_AWQOS,
    input wire                                           m_axi_in_49_AWREADY,
    output wire [                                   2:0] m_axi_in_49_AWSIZE,
    output wire                                          m_axi_in_49_AWVALID,
    input wire  [                                   0:0] m_axi_in_49_BID,
    output wire                                          m_axi_in_49_BREADY,
    input wire  [                                   1:0] m_axi_in_49_BRESP,
    input wire                                           m_axi_in_49_BVALID,
    input wire  [                                 255:0] m_axi_in_49_RDATA,
    input wire  [                                   0:0] m_axi_in_49_RID,
    input wire                                           m_axi_in_49_RLAST,
    output wire                                          m_axi_in_49_RREADY,
    input wire  [                                   1:0] m_axi_in_49_RRESP,
    input wire                                           m_axi_in_49_RVALID,
    output wire [                                 255:0] m_axi_in_49_WDATA,
    output wire                                          m_axi_in_49_WLAST,
    input wire                                           m_axi_in_49_WREADY,
    output wire [                                  31:0] m_axi_in_49_WSTRB,
    output wire                                          m_axi_in_49_WVALID,
    output wire [                                  63:0] m_axi_in_5_ARADDR,
    output wire [                                   1:0] m_axi_in_5_ARBURST,
    output wire [                                   3:0] m_axi_in_5_ARCACHE,
    output wire [                                   0:0] m_axi_in_5_ARID,
    output wire [                                   7:0] m_axi_in_5_ARLEN,
    output wire                                          m_axi_in_5_ARLOCK,
    output wire [                                   2:0] m_axi_in_5_ARPROT,
    output wire [                                   3:0] m_axi_in_5_ARQOS,
    input wire                                           m_axi_in_5_ARREADY,
    output wire [                                   2:0] m_axi_in_5_ARSIZE,
    output wire                                          m_axi_in_5_ARVALID,
    output wire [                                  63:0] m_axi_in_5_AWADDR,
    output wire [                                   1:0] m_axi_in_5_AWBURST,
    output wire [                                   3:0] m_axi_in_5_AWCACHE,
    output wire [                                   0:0] m_axi_in_5_AWID,
    output wire [                                   7:0] m_axi_in_5_AWLEN,
    output wire                                          m_axi_in_5_AWLOCK,
    output wire [                                   2:0] m_axi_in_5_AWPROT,
    output wire [                                   3:0] m_axi_in_5_AWQOS,
    input wire                                           m_axi_in_5_AWREADY,
    output wire [                                   2:0] m_axi_in_5_AWSIZE,
    output wire                                          m_axi_in_5_AWVALID,
    input wire  [                                   0:0] m_axi_in_5_BID,
    output wire                                          m_axi_in_5_BREADY,
    input wire  [                                   1:0] m_axi_in_5_BRESP,
    input wire                                           m_axi_in_5_BVALID,
    input wire  [                                 255:0] m_axi_in_5_RDATA,
    input wire  [                                   0:0] m_axi_in_5_RID,
    input wire                                           m_axi_in_5_RLAST,
    output wire                                          m_axi_in_5_RREADY,
    input wire  [                                   1:0] m_axi_in_5_RRESP,
    input wire                                           m_axi_in_5_RVALID,
    output wire [                                 255:0] m_axi_in_5_WDATA,
    output wire                                          m_axi_in_5_WLAST,
    input wire                                           m_axi_in_5_WREADY,
    output wire [                                  31:0] m_axi_in_5_WSTRB,
    output wire                                          m_axi_in_5_WVALID,
    output wire [                                  63:0] m_axi_in_50_ARADDR,
    output wire [                                   1:0] m_axi_in_50_ARBURST,
    output wire [                                   3:0] m_axi_in_50_ARCACHE,
    output wire [                                   0:0] m_axi_in_50_ARID,
    output wire [                                   7:0] m_axi_in_50_ARLEN,
    output wire                                          m_axi_in_50_ARLOCK,
    output wire [                                   2:0] m_axi_in_50_ARPROT,
    output wire [                                   3:0] m_axi_in_50_ARQOS,
    input wire                                           m_axi_in_50_ARREADY,
    output wire [                                   2:0] m_axi_in_50_ARSIZE,
    output wire                                          m_axi_in_50_ARVALID,
    output wire [                                  63:0] m_axi_in_50_AWADDR,
    output wire [                                   1:0] m_axi_in_50_AWBURST,
    output wire [                                   3:0] m_axi_in_50_AWCACHE,
    output wire [                                   0:0] m_axi_in_50_AWID,
    output wire [                                   7:0] m_axi_in_50_AWLEN,
    output wire                                          m_axi_in_50_AWLOCK,
    output wire [                                   2:0] m_axi_in_50_AWPROT,
    output wire [                                   3:0] m_axi_in_50_AWQOS,
    input wire                                           m_axi_in_50_AWREADY,
    output wire [                                   2:0] m_axi_in_50_AWSIZE,
    output wire                                          m_axi_in_50_AWVALID,
    input wire  [                                   0:0] m_axi_in_50_BID,
    output wire                                          m_axi_in_50_BREADY,
    input wire  [                                   1:0] m_axi_in_50_BRESP,
    input wire                                           m_axi_in_50_BVALID,
    input wire  [                                 255:0] m_axi_in_50_RDATA,
    input wire  [                                   0:0] m_axi_in_50_RID,
    input wire                                           m_axi_in_50_RLAST,
    output wire                                          m_axi_in_50_RREADY,
    input wire  [                                   1:0] m_axi_in_50_RRESP,
    input wire                                           m_axi_in_50_RVALID,
    output wire [                                 255:0] m_axi_in_50_WDATA,
    output wire                                          m_axi_in_50_WLAST,
    input wire                                           m_axi_in_50_WREADY,
    output wire [                                  31:0] m_axi_in_50_WSTRB,
    output wire                                          m_axi_in_50_WVALID,
    output wire [                                  63:0] m_axi_in_51_ARADDR,
    output wire [                                   1:0] m_axi_in_51_ARBURST,
    output wire [                                   3:0] m_axi_in_51_ARCACHE,
    output wire [                                   0:0] m_axi_in_51_ARID,
    output wire [                                   7:0] m_axi_in_51_ARLEN,
    output wire                                          m_axi_in_51_ARLOCK,
    output wire [                                   2:0] m_axi_in_51_ARPROT,
    output wire [                                   3:0] m_axi_in_51_ARQOS,
    input wire                                           m_axi_in_51_ARREADY,
    output wire [                                   2:0] m_axi_in_51_ARSIZE,
    output wire                                          m_axi_in_51_ARVALID,
    output wire [                                  63:0] m_axi_in_51_AWADDR,
    output wire [                                   1:0] m_axi_in_51_AWBURST,
    output wire [                                   3:0] m_axi_in_51_AWCACHE,
    output wire [                                   0:0] m_axi_in_51_AWID,
    output wire [                                   7:0] m_axi_in_51_AWLEN,
    output wire                                          m_axi_in_51_AWLOCK,
    output wire [                                   2:0] m_axi_in_51_AWPROT,
    output wire [                                   3:0] m_axi_in_51_AWQOS,
    input wire                                           m_axi_in_51_AWREADY,
    output wire [                                   2:0] m_axi_in_51_AWSIZE,
    output wire                                          m_axi_in_51_AWVALID,
    input wire  [                                   0:0] m_axi_in_51_BID,
    output wire                                          m_axi_in_51_BREADY,
    input wire  [                                   1:0] m_axi_in_51_BRESP,
    input wire                                           m_axi_in_51_BVALID,
    input wire  [                                 255:0] m_axi_in_51_RDATA,
    input wire  [                                   0:0] m_axi_in_51_RID,
    input wire                                           m_axi_in_51_RLAST,
    output wire                                          m_axi_in_51_RREADY,
    input wire  [                                   1:0] m_axi_in_51_RRESP,
    input wire                                           m_axi_in_51_RVALID,
    output wire [                                 255:0] m_axi_in_51_WDATA,
    output wire                                          m_axi_in_51_WLAST,
    input wire                                           m_axi_in_51_WREADY,
    output wire [                                  31:0] m_axi_in_51_WSTRB,
    output wire                                          m_axi_in_51_WVALID,
    output wire [                                  63:0] m_axi_in_52_ARADDR,
    output wire [                                   1:0] m_axi_in_52_ARBURST,
    output wire [                                   3:0] m_axi_in_52_ARCACHE,
    output wire [                                   0:0] m_axi_in_52_ARID,
    output wire [                                   7:0] m_axi_in_52_ARLEN,
    output wire                                          m_axi_in_52_ARLOCK,
    output wire [                                   2:0] m_axi_in_52_ARPROT,
    output wire [                                   3:0] m_axi_in_52_ARQOS,
    input wire                                           m_axi_in_52_ARREADY,
    output wire [                                   2:0] m_axi_in_52_ARSIZE,
    output wire                                          m_axi_in_52_ARVALID,
    output wire [                                  63:0] m_axi_in_52_AWADDR,
    output wire [                                   1:0] m_axi_in_52_AWBURST,
    output wire [                                   3:0] m_axi_in_52_AWCACHE,
    output wire [                                   0:0] m_axi_in_52_AWID,
    output wire [                                   7:0] m_axi_in_52_AWLEN,
    output wire                                          m_axi_in_52_AWLOCK,
    output wire [                                   2:0] m_axi_in_52_AWPROT,
    output wire [                                   3:0] m_axi_in_52_AWQOS,
    input wire                                           m_axi_in_52_AWREADY,
    output wire [                                   2:0] m_axi_in_52_AWSIZE,
    output wire                                          m_axi_in_52_AWVALID,
    input wire  [                                   0:0] m_axi_in_52_BID,
    output wire                                          m_axi_in_52_BREADY,
    input wire  [                                   1:0] m_axi_in_52_BRESP,
    input wire                                           m_axi_in_52_BVALID,
    input wire  [                                 255:0] m_axi_in_52_RDATA,
    input wire  [                                   0:0] m_axi_in_52_RID,
    input wire                                           m_axi_in_52_RLAST,
    output wire                                          m_axi_in_52_RREADY,
    input wire  [                                   1:0] m_axi_in_52_RRESP,
    input wire                                           m_axi_in_52_RVALID,
    output wire [                                 255:0] m_axi_in_52_WDATA,
    output wire                                          m_axi_in_52_WLAST,
    input wire                                           m_axi_in_52_WREADY,
    output wire [                                  31:0] m_axi_in_52_WSTRB,
    output wire                                          m_axi_in_52_WVALID,
    output wire [                                  63:0] m_axi_in_53_ARADDR,
    output wire [                                   1:0] m_axi_in_53_ARBURST,
    output wire [                                   3:0] m_axi_in_53_ARCACHE,
    output wire [                                   0:0] m_axi_in_53_ARID,
    output wire [                                   7:0] m_axi_in_53_ARLEN,
    output wire                                          m_axi_in_53_ARLOCK,
    output wire [                                   2:0] m_axi_in_53_ARPROT,
    output wire [                                   3:0] m_axi_in_53_ARQOS,
    input wire                                           m_axi_in_53_ARREADY,
    output wire [                                   2:0] m_axi_in_53_ARSIZE,
    output wire                                          m_axi_in_53_ARVALID,
    output wire [                                  63:0] m_axi_in_53_AWADDR,
    output wire [                                   1:0] m_axi_in_53_AWBURST,
    output wire [                                   3:0] m_axi_in_53_AWCACHE,
    output wire [                                   0:0] m_axi_in_53_AWID,
    output wire [                                   7:0] m_axi_in_53_AWLEN,
    output wire                                          m_axi_in_53_AWLOCK,
    output wire [                                   2:0] m_axi_in_53_AWPROT,
    output wire [                                   3:0] m_axi_in_53_AWQOS,
    input wire                                           m_axi_in_53_AWREADY,
    output wire [                                   2:0] m_axi_in_53_AWSIZE,
    output wire                                          m_axi_in_53_AWVALID,
    input wire  [                                   0:0] m_axi_in_53_BID,
    output wire                                          m_axi_in_53_BREADY,
    input wire  [                                   1:0] m_axi_in_53_BRESP,
    input wire                                           m_axi_in_53_BVALID,
    input wire  [                                 255:0] m_axi_in_53_RDATA,
    input wire  [                                   0:0] m_axi_in_53_RID,
    input wire                                           m_axi_in_53_RLAST,
    output wire                                          m_axi_in_53_RREADY,
    input wire  [                                   1:0] m_axi_in_53_RRESP,
    input wire                                           m_axi_in_53_RVALID,
    output wire [                                 255:0] m_axi_in_53_WDATA,
    output wire                                          m_axi_in_53_WLAST,
    input wire                                           m_axi_in_53_WREADY,
    output wire [                                  31:0] m_axi_in_53_WSTRB,
    output wire                                          m_axi_in_53_WVALID,
    output wire [                                  63:0] m_axi_in_6_ARADDR,
    output wire [                                   1:0] m_axi_in_6_ARBURST,
    output wire [                                   3:0] m_axi_in_6_ARCACHE,
    output wire [                                   0:0] m_axi_in_6_ARID,
    output wire [                                   7:0] m_axi_in_6_ARLEN,
    output wire                                          m_axi_in_6_ARLOCK,
    output wire [                                   2:0] m_axi_in_6_ARPROT,
    output wire [                                   3:0] m_axi_in_6_ARQOS,
    input wire                                           m_axi_in_6_ARREADY,
    output wire [                                   2:0] m_axi_in_6_ARSIZE,
    output wire                                          m_axi_in_6_ARVALID,
    output wire [                                  63:0] m_axi_in_6_AWADDR,
    output wire [                                   1:0] m_axi_in_6_AWBURST,
    output wire [                                   3:0] m_axi_in_6_AWCACHE,
    output wire [                                   0:0] m_axi_in_6_AWID,
    output wire [                                   7:0] m_axi_in_6_AWLEN,
    output wire                                          m_axi_in_6_AWLOCK,
    output wire [                                   2:0] m_axi_in_6_AWPROT,
    output wire [                                   3:0] m_axi_in_6_AWQOS,
    input wire                                           m_axi_in_6_AWREADY,
    output wire [                                   2:0] m_axi_in_6_AWSIZE,
    output wire                                          m_axi_in_6_AWVALID,
    input wire  [                                   0:0] m_axi_in_6_BID,
    output wire                                          m_axi_in_6_BREADY,
    input wire  [                                   1:0] m_axi_in_6_BRESP,
    input wire                                           m_axi_in_6_BVALID,
    input wire  [                                 255:0] m_axi_in_6_RDATA,
    input wire  [                                   0:0] m_axi_in_6_RID,
    input wire                                           m_axi_in_6_RLAST,
    output wire                                          m_axi_in_6_RREADY,
    input wire  [                                   1:0] m_axi_in_6_RRESP,
    input wire                                           m_axi_in_6_RVALID,
    output wire [                                 255:0] m_axi_in_6_WDATA,
    output wire                                          m_axi_in_6_WLAST,
    input wire                                           m_axi_in_6_WREADY,
    output wire [                                  31:0] m_axi_in_6_WSTRB,
    output wire                                          m_axi_in_6_WVALID,
    output wire [                                  63:0] m_axi_in_7_ARADDR,
    output wire [                                   1:0] m_axi_in_7_ARBURST,
    output wire [                                   3:0] m_axi_in_7_ARCACHE,
    output wire [                                   0:0] m_axi_in_7_ARID,
    output wire [                                   7:0] m_axi_in_7_ARLEN,
    output wire                                          m_axi_in_7_ARLOCK,
    output wire [                                   2:0] m_axi_in_7_ARPROT,
    output wire [                                   3:0] m_axi_in_7_ARQOS,
    input wire                                           m_axi_in_7_ARREADY,
    output wire [                                   2:0] m_axi_in_7_ARSIZE,
    output wire                                          m_axi_in_7_ARVALID,
    output wire [                                  63:0] m_axi_in_7_AWADDR,
    output wire [                                   1:0] m_axi_in_7_AWBURST,
    output wire [                                   3:0] m_axi_in_7_AWCACHE,
    output wire [                                   0:0] m_axi_in_7_AWID,
    output wire [                                   7:0] m_axi_in_7_AWLEN,
    output wire                                          m_axi_in_7_AWLOCK,
    output wire [                                   2:0] m_axi_in_7_AWPROT,
    output wire [                                   3:0] m_axi_in_7_AWQOS,
    input wire                                           m_axi_in_7_AWREADY,
    output wire [                                   2:0] m_axi_in_7_AWSIZE,
    output wire                                          m_axi_in_7_AWVALID,
    input wire  [                                   0:0] m_axi_in_7_BID,
    output wire                                          m_axi_in_7_BREADY,
    input wire  [                                   1:0] m_axi_in_7_BRESP,
    input wire                                           m_axi_in_7_BVALID,
    input wire  [                                 255:0] m_axi_in_7_RDATA,
    input wire  [                                   0:0] m_axi_in_7_RID,
    input wire                                           m_axi_in_7_RLAST,
    output wire                                          m_axi_in_7_RREADY,
    input wire  [                                   1:0] m_axi_in_7_RRESP,
    input wire                                           m_axi_in_7_RVALID,
    output wire [                                 255:0] m_axi_in_7_WDATA,
    output wire                                          m_axi_in_7_WLAST,
    input wire                                           m_axi_in_7_WREADY,
    output wire [                                  31:0] m_axi_in_7_WSTRB,
    output wire                                          m_axi_in_7_WVALID,
    output wire [                                  63:0] m_axi_in_8_ARADDR,
    output wire [                                   1:0] m_axi_in_8_ARBURST,
    output wire [                                   3:0] m_axi_in_8_ARCACHE,
    output wire [                                   0:0] m_axi_in_8_ARID,
    output wire [                                   7:0] m_axi_in_8_ARLEN,
    output wire                                          m_axi_in_8_ARLOCK,
    output wire [                                   2:0] m_axi_in_8_ARPROT,
    output wire [                                   3:0] m_axi_in_8_ARQOS,
    input wire                                           m_axi_in_8_ARREADY,
    output wire [                                   2:0] m_axi_in_8_ARSIZE,
    output wire                                          m_axi_in_8_ARVALID,
    output wire [                                  63:0] m_axi_in_8_AWADDR,
    output wire [                                   1:0] m_axi_in_8_AWBURST,
    output wire [                                   3:0] m_axi_in_8_AWCACHE,
    output wire [                                   0:0] m_axi_in_8_AWID,
    output wire [                                   7:0] m_axi_in_8_AWLEN,
    output wire                                          m_axi_in_8_AWLOCK,
    output wire [                                   2:0] m_axi_in_8_AWPROT,
    output wire [                                   3:0] m_axi_in_8_AWQOS,
    input wire                                           m_axi_in_8_AWREADY,
    output wire [                                   2:0] m_axi_in_8_AWSIZE,
    output wire                                          m_axi_in_8_AWVALID,
    input wire  [                                   0:0] m_axi_in_8_BID,
    output wire                                          m_axi_in_8_BREADY,
    input wire  [                                   1:0] m_axi_in_8_BRESP,
    input wire                                           m_axi_in_8_BVALID,
    input wire  [                                 255:0] m_axi_in_8_RDATA,
    input wire  [                                   0:0] m_axi_in_8_RID,
    input wire                                           m_axi_in_8_RLAST,
    output wire                                          m_axi_in_8_RREADY,
    input wire  [                                   1:0] m_axi_in_8_RRESP,
    input wire                                           m_axi_in_8_RVALID,
    output wire [                                 255:0] m_axi_in_8_WDATA,
    output wire                                          m_axi_in_8_WLAST,
    input wire                                           m_axi_in_8_WREADY,
    output wire [                                  31:0] m_axi_in_8_WSTRB,
    output wire                                          m_axi_in_8_WVALID,
    output wire [                                  63:0] m_axi_in_9_ARADDR,
    output wire [                                   1:0] m_axi_in_9_ARBURST,
    output wire [                                   3:0] m_axi_in_9_ARCACHE,
    output wire [                                   0:0] m_axi_in_9_ARID,
    output wire [                                   7:0] m_axi_in_9_ARLEN,
    output wire                                          m_axi_in_9_ARLOCK,
    output wire [                                   2:0] m_axi_in_9_ARPROT,
    output wire [                                   3:0] m_axi_in_9_ARQOS,
    input wire                                           m_axi_in_9_ARREADY,
    output wire [                                   2:0] m_axi_in_9_ARSIZE,
    output wire                                          m_axi_in_9_ARVALID,
    output wire [                                  63:0] m_axi_in_9_AWADDR,
    output wire [                                   1:0] m_axi_in_9_AWBURST,
    output wire [                                   3:0] m_axi_in_9_AWCACHE,
    output wire [                                   0:0] m_axi_in_9_AWID,
    output wire [                                   7:0] m_axi_in_9_AWLEN,
    output wire                                          m_axi_in_9_AWLOCK,
    output wire [                                   2:0] m_axi_in_9_AWPROT,
    output wire [                                   3:0] m_axi_in_9_AWQOS,
    input wire                                           m_axi_in_9_AWREADY,
    output wire [                                   2:0] m_axi_in_9_AWSIZE,
    output wire                                          m_axi_in_9_AWVALID,
    input wire  [                                   0:0] m_axi_in_9_BID,
    output wire                                          m_axi_in_9_BREADY,
    input wire  [                                   1:0] m_axi_in_9_BRESP,
    input wire                                           m_axi_in_9_BVALID,
    input wire  [                                 255:0] m_axi_in_9_RDATA,
    input wire  [                                   0:0] m_axi_in_9_RID,
    input wire                                           m_axi_in_9_RLAST,
    output wire                                          m_axi_in_9_RREADY,
    input wire  [                                   1:0] m_axi_in_9_RRESP,
    input wire                                           m_axi_in_9_RVALID,
    output wire [                                 255:0] m_axi_in_9_WDATA,
    output wire                                          m_axi_in_9_WLAST,
    input wire                                           m_axi_in_9_WREADY,
    output wire [                                  31:0] m_axi_in_9_WSTRB,
    output wire                                          m_axi_in_9_WVALID,
    output wire                                          control_s_axi_U_ACLK,
    output wire                                          control_s_axi_U_ACLK_EN,
    output wire [    (C_S_AXI_CONTROL_ADDR_WIDTH - 1):0] control_s_axi_U_ARADDR,
    output wire                                          control_s_axi_U_ARESET,
    input wire                                           control_s_axi_U_ARREADY,
    output wire                                          control_s_axi_U_ARVALID,
    output wire [    (C_S_AXI_CONTROL_ADDR_WIDTH - 1):0] control_s_axi_U_AWADDR,
    input wire                                           control_s_axi_U_AWREADY,
    output wire                                          control_s_axi_U_AWVALID,
    output wire                                          control_s_axi_U_BREADY,
    input wire  [                                   1:0] control_s_axi_U_BRESP,
    input wire                                           control_s_axi_U_BVALID,
    input wire  [                                  63:0] control_s_axi_U_L4_out_dist,
    input wire  [                                  63:0] control_s_axi_U_L4_out_id,
    input wire  [    (C_S_AXI_CONTROL_DATA_WIDTH - 1):0] control_s_axi_U_RDATA,
    output wire                                          control_s_axi_U_RREADY,
    input wire  [                                   1:0] control_s_axi_U_RRESP,
    input wire                                           control_s_axi_U_RVALID,
    output wire [    (C_S_AXI_CONTROL_DATA_WIDTH - 1):0] control_s_axi_U_WDATA,
    input wire                                           control_s_axi_U_WREADY,
    output wire [(C_S_AXI_CONTROL_DATA_WIDTH / 8 - 1):0] control_s_axi_U_WSTRB,
    output wire                                          control_s_axi_U_WVALID,
    output wire                                          control_s_axi_U_ap_done,
    output wire                                          control_s_axi_U_ap_idle,
    output wire                                          control_s_axi_U_ap_ready,
    input wire                                           control_s_axi_U_ap_start,
    input wire  [                                  63:0] control_s_axi_U_in_0,
    input wire  [                                  63:0] control_s_axi_U_in_1,
    input wire  [                                  63:0] control_s_axi_U_in_10,
    input wire  [                                  63:0] control_s_axi_U_in_11,
    input wire  [                                  63:0] control_s_axi_U_in_12,
    input wire  [                                  63:0] control_s_axi_U_in_13,
    input wire  [                                  63:0] control_s_axi_U_in_14,
    input wire  [                                  63:0] control_s_axi_U_in_15,
    input wire  [                                  63:0] control_s_axi_U_in_16,
    input wire  [                                  63:0] control_s_axi_U_in_17,
    input wire  [                                  63:0] control_s_axi_U_in_18,
    input wire  [                                  63:0] control_s_axi_U_in_19,
    input wire  [                                  63:0] control_s_axi_U_in_2,
    input wire  [                                  63:0] control_s_axi_U_in_20,
    input wire  [                                  63:0] control_s_axi_U_in_21,
    input wire  [                                  63:0] control_s_axi_U_in_22,
    input wire  [                                  63:0] control_s_axi_U_in_23,
    input wire  [                                  63:0] control_s_axi_U_in_24,
    input wire  [                                  63:0] control_s_axi_U_in_25,
    input wire  [                                  63:0] control_s_axi_U_in_26,
    input wire  [                                  63:0] control_s_axi_U_in_27,
    input wire  [                                  63:0] control_s_axi_U_in_28,
    input wire  [                                  63:0] control_s_axi_U_in_29,
    input wire  [                                  63:0] control_s_axi_U_in_3,
    input wire  [                                  63:0] control_s_axi_U_in_30,
    input wire  [                                  63:0] control_s_axi_U_in_31,
    input wire  [                                  63:0] control_s_axi_U_in_32,
    input wire  [                                  63:0] control_s_axi_U_in_33,
    input wire  [                                  63:0] control_s_axi_U_in_34,
    input wire  [                                  63:0] control_s_axi_U_in_35,
    input wire  [                                  63:0] control_s_axi_U_in_36,
    input wire  [                                  63:0] control_s_axi_U_in_37,
    input wire  [                                  63:0] control_s_axi_U_in_38,
    input wire  [                                  63:0] control_s_axi_U_in_39,
    input wire  [                                  63:0] control_s_axi_U_in_4,
    input wire  [                                  63:0] control_s_axi_U_in_40,
    input wire  [                                  63:0] control_s_axi_U_in_41,
    input wire  [                                  63:0] control_s_axi_U_in_42,
    input wire  [                                  63:0] control_s_axi_U_in_43,
    input wire  [                                  63:0] control_s_axi_U_in_44,
    input wire  [                                  63:0] control_s_axi_U_in_45,
    input wire  [                                  63:0] control_s_axi_U_in_46,
    input wire  [                                  63:0] control_s_axi_U_in_47,
    input wire  [                                  63:0] control_s_axi_U_in_48,
    input wire  [                                  63:0] control_s_axi_U_in_49,
    input wire  [                                  63:0] control_s_axi_U_in_5,
    input wire  [                                  63:0] control_s_axi_U_in_50,
    input wire  [                                  63:0] control_s_axi_U_in_51,
    input wire  [                                  63:0] control_s_axi_U_in_52,
    input wire  [                                  63:0] control_s_axi_U_in_53,
    input wire  [                                  63:0] control_s_axi_U_in_6,
    input wire  [                                  63:0] control_s_axi_U_in_7,
    input wire  [                                  63:0] control_s_axi_U_in_8,
    input wire  [                                  63:0] control_s_axi_U_in_9,
    input wire                                           control_s_axi_U_interrupt,
    output wire                                          L1_out_dist_0_clk,
    output wire [                                  65:0] L1_out_dist_0_if_din,
    input wire  [                                  65:0] L1_out_dist_0_if_dout,
    input wire                                           L1_out_dist_0_if_empty_n,
    input wire                                           L1_out_dist_0_if_full_n,
    output wire                                          L1_out_dist_0_if_read,
    output wire                                          L1_out_dist_0_if_read_ce,
    output wire                                          L1_out_dist_0_if_write,
    output wire                                          L1_out_dist_0_if_write_ce,
    output wire                                          L1_out_dist_0_reset,
    output wire                                          L1_out_dist_10_clk,
    output wire [                                  65:0] L1_out_dist_10_if_din,
    input wire  [                                  65:0] L1_out_dist_10_if_dout,
    input wire                                           L1_out_dist_10_if_empty_n,
    input wire                                           L1_out_dist_10_if_full_n,
    output wire                                          L1_out_dist_10_if_read,
    output wire                                          L1_out_dist_10_if_read_ce,
    output wire                                          L1_out_dist_10_if_write,
    output wire                                          L1_out_dist_10_if_write_ce,
    output wire                                          L1_out_dist_10_reset,
    output wire                                          L1_out_dist_11_clk,
    output wire [                                  65:0] L1_out_dist_11_if_din,
    input wire  [                                  65:0] L1_out_dist_11_if_dout,
    input wire                                           L1_out_dist_11_if_empty_n,
    input wire                                           L1_out_dist_11_if_full_n,
    output wire                                          L1_out_dist_11_if_read,
    output wire                                          L1_out_dist_11_if_read_ce,
    output wire                                          L1_out_dist_11_if_write,
    output wire                                          L1_out_dist_11_if_write_ce,
    output wire                                          L1_out_dist_11_reset,
    output wire                                          L1_out_dist_12_clk,
    output wire [                                  65:0] L1_out_dist_12_if_din,
    input wire  [                                  65:0] L1_out_dist_12_if_dout,
    input wire                                           L1_out_dist_12_if_empty_n,
    input wire                                           L1_out_dist_12_if_full_n,
    output wire                                          L1_out_dist_12_if_read,
    output wire                                          L1_out_dist_12_if_read_ce,
    output wire                                          L1_out_dist_12_if_write,
    output wire                                          L1_out_dist_12_if_write_ce,
    output wire                                          L1_out_dist_12_reset,
    output wire                                          L1_out_dist_13_clk,
    output wire [                                  65:0] L1_out_dist_13_if_din,
    input wire  [                                  65:0] L1_out_dist_13_if_dout,
    input wire                                           L1_out_dist_13_if_empty_n,
    input wire                                           L1_out_dist_13_if_full_n,
    output wire                                          L1_out_dist_13_if_read,
    output wire                                          L1_out_dist_13_if_read_ce,
    output wire                                          L1_out_dist_13_if_write,
    output wire                                          L1_out_dist_13_if_write_ce,
    output wire                                          L1_out_dist_13_reset,
    output wire                                          L1_out_dist_14_clk,
    output wire [                                  65:0] L1_out_dist_14_if_din,
    input wire  [                                  65:0] L1_out_dist_14_if_dout,
    input wire                                           L1_out_dist_14_if_empty_n,
    input wire                                           L1_out_dist_14_if_full_n,
    output wire                                          L1_out_dist_14_if_read,
    output wire                                          L1_out_dist_14_if_read_ce,
    output wire                                          L1_out_dist_14_if_write,
    output wire                                          L1_out_dist_14_if_write_ce,
    output wire                                          L1_out_dist_14_reset,
    output wire                                          L1_out_dist_15_clk,
    output wire [                                  65:0] L1_out_dist_15_if_din,
    input wire  [                                  65:0] L1_out_dist_15_if_dout,
    input wire                                           L1_out_dist_15_if_empty_n,
    input wire                                           L1_out_dist_15_if_full_n,
    output wire                                          L1_out_dist_15_if_read,
    output wire                                          L1_out_dist_15_if_read_ce,
    output wire                                          L1_out_dist_15_if_write,
    output wire                                          L1_out_dist_15_if_write_ce,
    output wire                                          L1_out_dist_15_reset,
    output wire                                          L1_out_dist_16_clk,
    output wire [                                  65:0] L1_out_dist_16_if_din,
    input wire  [                                  65:0] L1_out_dist_16_if_dout,
    input wire                                           L1_out_dist_16_if_empty_n,
    input wire                                           L1_out_dist_16_if_full_n,
    output wire                                          L1_out_dist_16_if_read,
    output wire                                          L1_out_dist_16_if_read_ce,
    output wire                                          L1_out_dist_16_if_write,
    output wire                                          L1_out_dist_16_if_write_ce,
    output wire                                          L1_out_dist_16_reset,
    output wire                                          L1_out_dist_17_clk,
    output wire [                                  65:0] L1_out_dist_17_if_din,
    input wire  [                                  65:0] L1_out_dist_17_if_dout,
    input wire                                           L1_out_dist_17_if_empty_n,
    input wire                                           L1_out_dist_17_if_full_n,
    output wire                                          L1_out_dist_17_if_read,
    output wire                                          L1_out_dist_17_if_read_ce,
    output wire                                          L1_out_dist_17_if_write,
    output wire                                          L1_out_dist_17_if_write_ce,
    output wire                                          L1_out_dist_17_reset,
    output wire                                          L1_out_dist_1_clk,
    output wire [                                  65:0] L1_out_dist_1_if_din,
    input wire  [                                  65:0] L1_out_dist_1_if_dout,
    input wire                                           L1_out_dist_1_if_empty_n,
    input wire                                           L1_out_dist_1_if_full_n,
    output wire                                          L1_out_dist_1_if_read,
    output wire                                          L1_out_dist_1_if_read_ce,
    output wire                                          L1_out_dist_1_if_write,
    output wire                                          L1_out_dist_1_if_write_ce,
    output wire                                          L1_out_dist_1_reset,
    output wire                                          L1_out_dist_2_clk,
    output wire [                                  65:0] L1_out_dist_2_if_din,
    input wire  [                                  65:0] L1_out_dist_2_if_dout,
    input wire                                           L1_out_dist_2_if_empty_n,
    input wire                                           L1_out_dist_2_if_full_n,
    output wire                                          L1_out_dist_2_if_read,
    output wire                                          L1_out_dist_2_if_read_ce,
    output wire                                          L1_out_dist_2_if_write,
    output wire                                          L1_out_dist_2_if_write_ce,
    output wire                                          L1_out_dist_2_reset,
    output wire                                          L1_out_dist_3_clk,
    output wire [                                  65:0] L1_out_dist_3_if_din,
    input wire  [                                  65:0] L1_out_dist_3_if_dout,
    input wire                                           L1_out_dist_3_if_empty_n,
    input wire                                           L1_out_dist_3_if_full_n,
    output wire                                          L1_out_dist_3_if_read,
    output wire                                          L1_out_dist_3_if_read_ce,
    output wire                                          L1_out_dist_3_if_write,
    output wire                                          L1_out_dist_3_if_write_ce,
    output wire                                          L1_out_dist_3_reset,
    output wire                                          L1_out_dist_4_clk,
    output wire [                                  65:0] L1_out_dist_4_if_din,
    input wire  [                                  65:0] L1_out_dist_4_if_dout,
    input wire                                           L1_out_dist_4_if_empty_n,
    input wire                                           L1_out_dist_4_if_full_n,
    output wire                                          L1_out_dist_4_if_read,
    output wire                                          L1_out_dist_4_if_read_ce,
    output wire                                          L1_out_dist_4_if_write,
    output wire                                          L1_out_dist_4_if_write_ce,
    output wire                                          L1_out_dist_4_reset,
    output wire                                          L1_out_dist_5_clk,
    output wire [                                  65:0] L1_out_dist_5_if_din,
    input wire  [                                  65:0] L1_out_dist_5_if_dout,
    input wire                                           L1_out_dist_5_if_empty_n,
    input wire                                           L1_out_dist_5_if_full_n,
    output wire                                          L1_out_dist_5_if_read,
    output wire                                          L1_out_dist_5_if_read_ce,
    output wire                                          L1_out_dist_5_if_write,
    output wire                                          L1_out_dist_5_if_write_ce,
    output wire                                          L1_out_dist_5_reset,
    output wire                                          L1_out_dist_6_clk,
    output wire [                                  65:0] L1_out_dist_6_if_din,
    input wire  [                                  65:0] L1_out_dist_6_if_dout,
    input wire                                           L1_out_dist_6_if_empty_n,
    input wire                                           L1_out_dist_6_if_full_n,
    output wire                                          L1_out_dist_6_if_read,
    output wire                                          L1_out_dist_6_if_read_ce,
    output wire                                          L1_out_dist_6_if_write,
    output wire                                          L1_out_dist_6_if_write_ce,
    output wire                                          L1_out_dist_6_reset,
    output wire                                          L1_out_dist_7_clk,
    output wire [                                  65:0] L1_out_dist_7_if_din,
    input wire  [                                  65:0] L1_out_dist_7_if_dout,
    input wire                                           L1_out_dist_7_if_empty_n,
    input wire                                           L1_out_dist_7_if_full_n,
    output wire                                          L1_out_dist_7_if_read,
    output wire                                          L1_out_dist_7_if_read_ce,
    output wire                                          L1_out_dist_7_if_write,
    output wire                                          L1_out_dist_7_if_write_ce,
    output wire                                          L1_out_dist_7_reset,
    output wire                                          L1_out_dist_8_clk,
    output wire [                                  65:0] L1_out_dist_8_if_din,
    input wire  [                                  65:0] L1_out_dist_8_if_dout,
    input wire                                           L1_out_dist_8_if_empty_n,
    input wire                                           L1_out_dist_8_if_full_n,
    output wire                                          L1_out_dist_8_if_read,
    output wire                                          L1_out_dist_8_if_read_ce,
    output wire                                          L1_out_dist_8_if_write,
    output wire                                          L1_out_dist_8_if_write_ce,
    output wire                                          L1_out_dist_8_reset,
    output wire                                          L1_out_dist_9_clk,
    output wire [                                  65:0] L1_out_dist_9_if_din,
    input wire  [                                  65:0] L1_out_dist_9_if_dout,
    input wire                                           L1_out_dist_9_if_empty_n,
    input wire                                           L1_out_dist_9_if_full_n,
    output wire                                          L1_out_dist_9_if_read,
    output wire                                          L1_out_dist_9_if_read_ce,
    output wire                                          L1_out_dist_9_if_write,
    output wire                                          L1_out_dist_9_if_write_ce,
    output wire                                          L1_out_dist_9_reset,
    output wire                                          L1_out_id_0_clk,
    output wire [                                  65:0] L1_out_id_0_if_din,
    input wire  [                                  65:0] L1_out_id_0_if_dout,
    input wire                                           L1_out_id_0_if_empty_n,
    input wire                                           L1_out_id_0_if_full_n,
    output wire                                          L1_out_id_0_if_read,
    output wire                                          L1_out_id_0_if_read_ce,
    output wire                                          L1_out_id_0_if_write,
    output wire                                          L1_out_id_0_if_write_ce,
    output wire                                          L1_out_id_0_reset,
    output wire                                          L1_out_id_10_clk,
    output wire [                                  65:0] L1_out_id_10_if_din,
    input wire  [                                  65:0] L1_out_id_10_if_dout,
    input wire                                           L1_out_id_10_if_empty_n,
    input wire                                           L1_out_id_10_if_full_n,
    output wire                                          L1_out_id_10_if_read,
    output wire                                          L1_out_id_10_if_read_ce,
    output wire                                          L1_out_id_10_if_write,
    output wire                                          L1_out_id_10_if_write_ce,
    output wire                                          L1_out_id_10_reset,
    output wire                                          L1_out_id_11_clk,
    output wire [                                  65:0] L1_out_id_11_if_din,
    input wire  [                                  65:0] L1_out_id_11_if_dout,
    input wire                                           L1_out_id_11_if_empty_n,
    input wire                                           L1_out_id_11_if_full_n,
    output wire                                          L1_out_id_11_if_read,
    output wire                                          L1_out_id_11_if_read_ce,
    output wire                                          L1_out_id_11_if_write,
    output wire                                          L1_out_id_11_if_write_ce,
    output wire                                          L1_out_id_11_reset,
    output wire                                          L1_out_id_12_clk,
    output wire [                                  65:0] L1_out_id_12_if_din,
    input wire  [                                  65:0] L1_out_id_12_if_dout,
    input wire                                           L1_out_id_12_if_empty_n,
    input wire                                           L1_out_id_12_if_full_n,
    output wire                                          L1_out_id_12_if_read,
    output wire                                          L1_out_id_12_if_read_ce,
    output wire                                          L1_out_id_12_if_write,
    output wire                                          L1_out_id_12_if_write_ce,
    output wire                                          L1_out_id_12_reset,
    output wire                                          L1_out_id_13_clk,
    output wire [                                  65:0] L1_out_id_13_if_din,
    input wire  [                                  65:0] L1_out_id_13_if_dout,
    input wire                                           L1_out_id_13_if_empty_n,
    input wire                                           L1_out_id_13_if_full_n,
    output wire                                          L1_out_id_13_if_read,
    output wire                                          L1_out_id_13_if_read_ce,
    output wire                                          L1_out_id_13_if_write,
    output wire                                          L1_out_id_13_if_write_ce,
    output wire                                          L1_out_id_13_reset,
    output wire                                          L1_out_id_14_clk,
    output wire [                                  65:0] L1_out_id_14_if_din,
    input wire  [                                  65:0] L1_out_id_14_if_dout,
    input wire                                           L1_out_id_14_if_empty_n,
    input wire                                           L1_out_id_14_if_full_n,
    output wire                                          L1_out_id_14_if_read,
    output wire                                          L1_out_id_14_if_read_ce,
    output wire                                          L1_out_id_14_if_write,
    output wire                                          L1_out_id_14_if_write_ce,
    output wire                                          L1_out_id_14_reset,
    output wire                                          L1_out_id_15_clk,
    output wire [                                  65:0] L1_out_id_15_if_din,
    input wire  [                                  65:0] L1_out_id_15_if_dout,
    input wire                                           L1_out_id_15_if_empty_n,
    input wire                                           L1_out_id_15_if_full_n,
    output wire                                          L1_out_id_15_if_read,
    output wire                                          L1_out_id_15_if_read_ce,
    output wire                                          L1_out_id_15_if_write,
    output wire                                          L1_out_id_15_if_write_ce,
    output wire                                          L1_out_id_15_reset,
    output wire                                          L1_out_id_16_clk,
    output wire [                                  65:0] L1_out_id_16_if_din,
    input wire  [                                  65:0] L1_out_id_16_if_dout,
    input wire                                           L1_out_id_16_if_empty_n,
    input wire                                           L1_out_id_16_if_full_n,
    output wire                                          L1_out_id_16_if_read,
    output wire                                          L1_out_id_16_if_read_ce,
    output wire                                          L1_out_id_16_if_write,
    output wire                                          L1_out_id_16_if_write_ce,
    output wire                                          L1_out_id_16_reset,
    output wire                                          L1_out_id_17_clk,
    output wire [                                  65:0] L1_out_id_17_if_din,
    input wire  [                                  65:0] L1_out_id_17_if_dout,
    input wire                                           L1_out_id_17_if_empty_n,
    input wire                                           L1_out_id_17_if_full_n,
    output wire                                          L1_out_id_17_if_read,
    output wire                                          L1_out_id_17_if_read_ce,
    output wire                                          L1_out_id_17_if_write,
    output wire                                          L1_out_id_17_if_write_ce,
    output wire                                          L1_out_id_17_reset,
    output wire                                          L1_out_id_1_clk,
    output wire [                                  65:0] L1_out_id_1_if_din,
    input wire  [                                  65:0] L1_out_id_1_if_dout,
    input wire                                           L1_out_id_1_if_empty_n,
    input wire                                           L1_out_id_1_if_full_n,
    output wire                                          L1_out_id_1_if_read,
    output wire                                          L1_out_id_1_if_read_ce,
    output wire                                          L1_out_id_1_if_write,
    output wire                                          L1_out_id_1_if_write_ce,
    output wire                                          L1_out_id_1_reset,
    output wire                                          L1_out_id_2_clk,
    output wire [                                  65:0] L1_out_id_2_if_din,
    input wire  [                                  65:0] L1_out_id_2_if_dout,
    input wire                                           L1_out_id_2_if_empty_n,
    input wire                                           L1_out_id_2_if_full_n,
    output wire                                          L1_out_id_2_if_read,
    output wire                                          L1_out_id_2_if_read_ce,
    output wire                                          L1_out_id_2_if_write,
    output wire                                          L1_out_id_2_if_write_ce,
    output wire                                          L1_out_id_2_reset,
    output wire                                          L1_out_id_3_clk,
    output wire [                                  65:0] L1_out_id_3_if_din,
    input wire  [                                  65:0] L1_out_id_3_if_dout,
    input wire                                           L1_out_id_3_if_empty_n,
    input wire                                           L1_out_id_3_if_full_n,
    output wire                                          L1_out_id_3_if_read,
    output wire                                          L1_out_id_3_if_read_ce,
    output wire                                          L1_out_id_3_if_write,
    output wire                                          L1_out_id_3_if_write_ce,
    output wire                                          L1_out_id_3_reset,
    output wire                                          L1_out_id_4_clk,
    output wire [                                  65:0] L1_out_id_4_if_din,
    input wire  [                                  65:0] L1_out_id_4_if_dout,
    input wire                                           L1_out_id_4_if_empty_n,
    input wire                                           L1_out_id_4_if_full_n,
    output wire                                          L1_out_id_4_if_read,
    output wire                                          L1_out_id_4_if_read_ce,
    output wire                                          L1_out_id_4_if_write,
    output wire                                          L1_out_id_4_if_write_ce,
    output wire                                          L1_out_id_4_reset,
    output wire                                          L1_out_id_5_clk,
    output wire [                                  65:0] L1_out_id_5_if_din,
    input wire  [                                  65:0] L1_out_id_5_if_dout,
    input wire                                           L1_out_id_5_if_empty_n,
    input wire                                           L1_out_id_5_if_full_n,
    output wire                                          L1_out_id_5_if_read,
    output wire                                          L1_out_id_5_if_read_ce,
    output wire                                          L1_out_id_5_if_write,
    output wire                                          L1_out_id_5_if_write_ce,
    output wire                                          L1_out_id_5_reset,
    output wire                                          L1_out_id_6_clk,
    output wire [                                  65:0] L1_out_id_6_if_din,
    input wire  [                                  65:0] L1_out_id_6_if_dout,
    input wire                                           L1_out_id_6_if_empty_n,
    input wire                                           L1_out_id_6_if_full_n,
    output wire                                          L1_out_id_6_if_read,
    output wire                                          L1_out_id_6_if_read_ce,
    output wire                                          L1_out_id_6_if_write,
    output wire                                          L1_out_id_6_if_write_ce,
    output wire                                          L1_out_id_6_reset,
    output wire                                          L1_out_id_7_clk,
    output wire [                                  65:0] L1_out_id_7_if_din,
    input wire  [                                  65:0] L1_out_id_7_if_dout,
    input wire                                           L1_out_id_7_if_empty_n,
    input wire                                           L1_out_id_7_if_full_n,
    output wire                                          L1_out_id_7_if_read,
    output wire                                          L1_out_id_7_if_read_ce,
    output wire                                          L1_out_id_7_if_write,
    output wire                                          L1_out_id_7_if_write_ce,
    output wire                                          L1_out_id_7_reset,
    output wire                                          L1_out_id_8_clk,
    output wire [                                  65:0] L1_out_id_8_if_din,
    input wire  [                                  65:0] L1_out_id_8_if_dout,
    input wire                                           L1_out_id_8_if_empty_n,
    input wire                                           L1_out_id_8_if_full_n,
    output wire                                          L1_out_id_8_if_read,
    output wire                                          L1_out_id_8_if_read_ce,
    output wire                                          L1_out_id_8_if_write,
    output wire                                          L1_out_id_8_if_write_ce,
    output wire                                          L1_out_id_8_reset,
    output wire                                          L1_out_id_9_clk,
    output wire [                                  65:0] L1_out_id_9_if_din,
    input wire  [                                  65:0] L1_out_id_9_if_dout,
    input wire                                           L1_out_id_9_if_empty_n,
    input wire                                           L1_out_id_9_if_full_n,
    output wire                                          L1_out_id_9_if_read,
    output wire                                          L1_out_id_9_if_read_ce,
    output wire                                          L1_out_id_9_if_write,
    output wire                                          L1_out_id_9_if_write_ce,
    output wire                                          L1_out_id_9_reset,
    output wire                                          L2_out_dist0_clk,
    output wire [                                  65:0] L2_out_dist0_if_din,
    input wire  [                                  65:0] L2_out_dist0_if_dout,
    input wire                                           L2_out_dist0_if_empty_n,
    input wire                                           L2_out_dist0_if_full_n,
    output wire                                          L2_out_dist0_if_read,
    output wire                                          L2_out_dist0_if_read_ce,
    output wire                                          L2_out_dist0_if_write,
    output wire                                          L2_out_dist0_if_write_ce,
    output wire                                          L2_out_dist0_reset,
    output wire                                          L2_out_dist1_clk,
    output wire [                                  65:0] L2_out_dist1_if_din,
    input wire  [                                  65:0] L2_out_dist1_if_dout,
    input wire                                           L2_out_dist1_if_empty_n,
    input wire                                           L2_out_dist1_if_full_n,
    output wire                                          L2_out_dist1_if_read,
    output wire                                          L2_out_dist1_if_read_ce,
    output wire                                          L2_out_dist1_if_write,
    output wire                                          L2_out_dist1_if_write_ce,
    output wire                                          L2_out_dist1_reset,
    output wire                                          L2_out_dist2_clk,
    output wire [                                  65:0] L2_out_dist2_if_din,
    input wire  [                                  65:0] L2_out_dist2_if_dout,
    input wire                                           L2_out_dist2_if_empty_n,
    input wire                                           L2_out_dist2_if_full_n,
    output wire                                          L2_out_dist2_if_read,
    output wire                                          L2_out_dist2_if_read_ce,
    output wire                                          L2_out_dist2_if_write,
    output wire                                          L2_out_dist2_if_write_ce,
    output wire                                          L2_out_dist2_reset,
    output wire                                          L2_out_dist3_clk,
    output wire [                                  65:0] L2_out_dist3_if_din,
    input wire  [                                  65:0] L2_out_dist3_if_dout,
    input wire                                           L2_out_dist3_if_empty_n,
    input wire                                           L2_out_dist3_if_full_n,
    output wire                                          L2_out_dist3_if_read,
    output wire                                          L2_out_dist3_if_read_ce,
    output wire                                          L2_out_dist3_if_write,
    output wire                                          L2_out_dist3_if_write_ce,
    output wire                                          L2_out_dist3_reset,
    output wire                                          L2_out_dist4_clk,
    output wire [                                  65:0] L2_out_dist4_if_din,
    input wire  [                                  65:0] L2_out_dist4_if_dout,
    input wire                                           L2_out_dist4_if_empty_n,
    input wire                                           L2_out_dist4_if_full_n,
    output wire                                          L2_out_dist4_if_read,
    output wire                                          L2_out_dist4_if_read_ce,
    output wire                                          L2_out_dist4_if_write,
    output wire                                          L2_out_dist4_if_write_ce,
    output wire                                          L2_out_dist4_reset,
    output wire                                          L2_out_dist5_clk,
    output wire [                                  65:0] L2_out_dist5_if_din,
    input wire  [                                  65:0] L2_out_dist5_if_dout,
    input wire                                           L2_out_dist5_if_empty_n,
    input wire                                           L2_out_dist5_if_full_n,
    output wire                                          L2_out_dist5_if_read,
    output wire                                          L2_out_dist5_if_read_ce,
    output wire                                          L2_out_dist5_if_write,
    output wire                                          L2_out_dist5_if_write_ce,
    output wire                                          L2_out_dist5_reset,
    output wire                                          L2_out_id0_clk,
    output wire [                                  65:0] L2_out_id0_if_din,
    input wire  [                                  65:0] L2_out_id0_if_dout,
    input wire                                           L2_out_id0_if_empty_n,
    input wire                                           L2_out_id0_if_full_n,
    output wire                                          L2_out_id0_if_read,
    output wire                                          L2_out_id0_if_read_ce,
    output wire                                          L2_out_id0_if_write,
    output wire                                          L2_out_id0_if_write_ce,
    output wire                                          L2_out_id0_reset,
    output wire                                          L2_out_id1_clk,
    output wire [                                  65:0] L2_out_id1_if_din,
    input wire  [                                  65:0] L2_out_id1_if_dout,
    input wire                                           L2_out_id1_if_empty_n,
    input wire                                           L2_out_id1_if_full_n,
    output wire                                          L2_out_id1_if_read,
    output wire                                          L2_out_id1_if_read_ce,
    output wire                                          L2_out_id1_if_write,
    output wire                                          L2_out_id1_if_write_ce,
    output wire                                          L2_out_id1_reset,
    output wire                                          L2_out_id2_clk,
    output wire [                                  65:0] L2_out_id2_if_din,
    input wire  [                                  65:0] L2_out_id2_if_dout,
    input wire                                           L2_out_id2_if_empty_n,
    input wire                                           L2_out_id2_if_full_n,
    output wire                                          L2_out_id2_if_read,
    output wire                                          L2_out_id2_if_read_ce,
    output wire                                          L2_out_id2_if_write,
    output wire                                          L2_out_id2_if_write_ce,
    output wire                                          L2_out_id2_reset,
    output wire                                          L2_out_id3_clk,
    output wire [                                  65:0] L2_out_id3_if_din,
    input wire  [                                  65:0] L2_out_id3_if_dout,
    input wire                                           L2_out_id3_if_empty_n,
    input wire                                           L2_out_id3_if_full_n,
    output wire                                          L2_out_id3_if_read,
    output wire                                          L2_out_id3_if_read_ce,
    output wire                                          L2_out_id3_if_write,
    output wire                                          L2_out_id3_if_write_ce,
    output wire                                          L2_out_id3_reset,
    output wire                                          L2_out_id4_clk,
    output wire [                                  65:0] L2_out_id4_if_din,
    input wire  [                                  65:0] L2_out_id4_if_dout,
    input wire                                           L2_out_id4_if_empty_n,
    input wire                                           L2_out_id4_if_full_n,
    output wire                                          L2_out_id4_if_read,
    output wire                                          L2_out_id4_if_read_ce,
    output wire                                          L2_out_id4_if_write,
    output wire                                          L2_out_id4_if_write_ce,
    output wire                                          L2_out_id4_reset,
    output wire                                          L2_out_id5_clk,
    output wire [                                  65:0] L2_out_id5_if_din,
    input wire  [                                  65:0] L2_out_id5_if_dout,
    input wire                                           L2_out_id5_if_empty_n,
    input wire                                           L2_out_id5_if_full_n,
    output wire                                          L2_out_id5_if_read,
    output wire                                          L2_out_id5_if_read_ce,
    output wire                                          L2_out_id5_if_write,
    output wire                                          L2_out_id5_if_write_ce,
    output wire                                          L2_out_id5_reset,
    output wire                                          L3_out_dist0_clk,
    output wire [                                  65:0] L3_out_dist0_if_din,
    input wire  [                                  65:0] L3_out_dist0_if_dout,
    input wire                                           L3_out_dist0_if_empty_n,
    input wire                                           L3_out_dist0_if_full_n,
    output wire                                          L3_out_dist0_if_read,
    output wire                                          L3_out_dist0_if_read_ce,
    output wire                                          L3_out_dist0_if_write,
    output wire                                          L3_out_dist0_if_write_ce,
    output wire                                          L3_out_dist0_reset,
    output wire                                          L3_out_dist1_clk,
    output wire [                                  65:0] L3_out_dist1_if_din,
    input wire  [                                  65:0] L3_out_dist1_if_dout,
    input wire                                           L3_out_dist1_if_empty_n,
    input wire                                           L3_out_dist1_if_full_n,
    output wire                                          L3_out_dist1_if_read,
    output wire                                          L3_out_dist1_if_read_ce,
    output wire                                          L3_out_dist1_if_write,
    output wire                                          L3_out_dist1_if_write_ce,
    output wire                                          L3_out_dist1_reset,
    output wire                                          L3_out_id0_clk,
    output wire [                                  65:0] L3_out_id0_if_din,
    input wire  [                                  65:0] L3_out_id0_if_dout,
    input wire                                           L3_out_id0_if_empty_n,
    input wire                                           L3_out_id0_if_full_n,
    output wire                                          L3_out_id0_if_read,
    output wire                                          L3_out_id0_if_read_ce,
    output wire                                          L3_out_id0_if_write,
    output wire                                          L3_out_id0_if_write_ce,
    output wire                                          L3_out_id0_reset,
    output wire                                          L3_out_id1_clk,
    output wire [                                  65:0] L3_out_id1_if_din,
    input wire  [                                  65:0] L3_out_id1_if_dout,
    input wire                                           L3_out_id1_if_empty_n,
    input wire                                           L3_out_id1_if_full_n,
    output wire                                          L3_out_id1_if_read,
    output wire                                          L3_out_id1_if_read_ce,
    output wire                                          L3_out_id1_if_write,
    output wire                                          L3_out_id1_if_write_ce,
    output wire                                          L3_out_id1_reset,
    output wire                                          out_dist_0_clk,
    output wire [                                  65:0] out_dist_0_if_din,
    input wire  [                                  65:0] out_dist_0_if_dout,
    input wire                                           out_dist_0_if_empty_n,
    input wire                                           out_dist_0_if_full_n,
    output wire                                          out_dist_0_if_read,
    output wire                                          out_dist_0_if_read_ce,
    output wire                                          out_dist_0_if_write,
    output wire                                          out_dist_0_if_write_ce,
    output wire                                          out_dist_0_reset,
    output wire                                          out_dist_10_clk,
    output wire [                                  65:0] out_dist_10_if_din,
    input wire  [                                  65:0] out_dist_10_if_dout,
    input wire                                           out_dist_10_if_empty_n,
    input wire                                           out_dist_10_if_full_n,
    output wire                                          out_dist_10_if_read,
    output wire                                          out_dist_10_if_read_ce,
    output wire                                          out_dist_10_if_write,
    output wire                                          out_dist_10_if_write_ce,
    output wire                                          out_dist_10_reset,
    output wire                                          out_dist_11_clk,
    output wire [                                  65:0] out_dist_11_if_din,
    input wire  [                                  65:0] out_dist_11_if_dout,
    input wire                                           out_dist_11_if_empty_n,
    input wire                                           out_dist_11_if_full_n,
    output wire                                          out_dist_11_if_read,
    output wire                                          out_dist_11_if_read_ce,
    output wire                                          out_dist_11_if_write,
    output wire                                          out_dist_11_if_write_ce,
    output wire                                          out_dist_11_reset,
    output wire                                          out_dist_12_clk,
    output wire [                                  65:0] out_dist_12_if_din,
    input wire  [                                  65:0] out_dist_12_if_dout,
    input wire                                           out_dist_12_if_empty_n,
    input wire                                           out_dist_12_if_full_n,
    output wire                                          out_dist_12_if_read,
    output wire                                          out_dist_12_if_read_ce,
    output wire                                          out_dist_12_if_write,
    output wire                                          out_dist_12_if_write_ce,
    output wire                                          out_dist_12_reset,
    output wire                                          out_dist_13_clk,
    output wire [                                  65:0] out_dist_13_if_din,
    input wire  [                                  65:0] out_dist_13_if_dout,
    input wire                                           out_dist_13_if_empty_n,
    input wire                                           out_dist_13_if_full_n,
    output wire                                          out_dist_13_if_read,
    output wire                                          out_dist_13_if_read_ce,
    output wire                                          out_dist_13_if_write,
    output wire                                          out_dist_13_if_write_ce,
    output wire                                          out_dist_13_reset,
    output wire                                          out_dist_14_clk,
    output wire [                                  65:0] out_dist_14_if_din,
    input wire  [                                  65:0] out_dist_14_if_dout,
    input wire                                           out_dist_14_if_empty_n,
    input wire                                           out_dist_14_if_full_n,
    output wire                                          out_dist_14_if_read,
    output wire                                          out_dist_14_if_read_ce,
    output wire                                          out_dist_14_if_write,
    output wire                                          out_dist_14_if_write_ce,
    output wire                                          out_dist_14_reset,
    output wire                                          out_dist_15_clk,
    output wire [                                  65:0] out_dist_15_if_din,
    input wire  [                                  65:0] out_dist_15_if_dout,
    input wire                                           out_dist_15_if_empty_n,
    input wire                                           out_dist_15_if_full_n,
    output wire                                          out_dist_15_if_read,
    output wire                                          out_dist_15_if_read_ce,
    output wire                                          out_dist_15_if_write,
    output wire                                          out_dist_15_if_write_ce,
    output wire                                          out_dist_15_reset,
    output wire                                          out_dist_16_clk,
    output wire [                                  65:0] out_dist_16_if_din,
    input wire  [                                  65:0] out_dist_16_if_dout,
    input wire                                           out_dist_16_if_empty_n,
    input wire                                           out_dist_16_if_full_n,
    output wire                                          out_dist_16_if_read,
    output wire                                          out_dist_16_if_read_ce,
    output wire                                          out_dist_16_if_write,
    output wire                                          out_dist_16_if_write_ce,
    output wire                                          out_dist_16_reset,
    output wire                                          out_dist_17_clk,
    output wire [                                  65:0] out_dist_17_if_din,
    input wire  [                                  65:0] out_dist_17_if_dout,
    input wire                                           out_dist_17_if_empty_n,
    input wire                                           out_dist_17_if_full_n,
    output wire                                          out_dist_17_if_read,
    output wire                                          out_dist_17_if_read_ce,
    output wire                                          out_dist_17_if_write,
    output wire                                          out_dist_17_if_write_ce,
    output wire                                          out_dist_17_reset,
    output wire                                          out_dist_18_clk,
    output wire [                                  65:0] out_dist_18_if_din,
    input wire  [                                  65:0] out_dist_18_if_dout,
    input wire                                           out_dist_18_if_empty_n,
    input wire                                           out_dist_18_if_full_n,
    output wire                                          out_dist_18_if_read,
    output wire                                          out_dist_18_if_read_ce,
    output wire                                          out_dist_18_if_write,
    output wire                                          out_dist_18_if_write_ce,
    output wire                                          out_dist_18_reset,
    output wire                                          out_dist_19_clk,
    output wire [                                  65:0] out_dist_19_if_din,
    input wire  [                                  65:0] out_dist_19_if_dout,
    input wire                                           out_dist_19_if_empty_n,
    input wire                                           out_dist_19_if_full_n,
    output wire                                          out_dist_19_if_read,
    output wire                                          out_dist_19_if_read_ce,
    output wire                                          out_dist_19_if_write,
    output wire                                          out_dist_19_if_write_ce,
    output wire                                          out_dist_19_reset,
    output wire                                          out_dist_1_clk,
    output wire [                                  65:0] out_dist_1_if_din,
    input wire  [                                  65:0] out_dist_1_if_dout,
    input wire                                           out_dist_1_if_empty_n,
    input wire                                           out_dist_1_if_full_n,
    output wire                                          out_dist_1_if_read,
    output wire                                          out_dist_1_if_read_ce,
    output wire                                          out_dist_1_if_write,
    output wire                                          out_dist_1_if_write_ce,
    output wire                                          out_dist_1_reset,
    output wire                                          out_dist_20_clk,
    output wire [                                  65:0] out_dist_20_if_din,
    input wire  [                                  65:0] out_dist_20_if_dout,
    input wire                                           out_dist_20_if_empty_n,
    input wire                                           out_dist_20_if_full_n,
    output wire                                          out_dist_20_if_read,
    output wire                                          out_dist_20_if_read_ce,
    output wire                                          out_dist_20_if_write,
    output wire                                          out_dist_20_if_write_ce,
    output wire                                          out_dist_20_reset,
    output wire                                          out_dist_21_clk,
    output wire [                                  65:0] out_dist_21_if_din,
    input wire  [                                  65:0] out_dist_21_if_dout,
    input wire                                           out_dist_21_if_empty_n,
    input wire                                           out_dist_21_if_full_n,
    output wire                                          out_dist_21_if_read,
    output wire                                          out_dist_21_if_read_ce,
    output wire                                          out_dist_21_if_write,
    output wire                                          out_dist_21_if_write_ce,
    output wire                                          out_dist_21_reset,
    output wire                                          out_dist_22_clk,
    output wire [                                  65:0] out_dist_22_if_din,
    input wire  [                                  65:0] out_dist_22_if_dout,
    input wire                                           out_dist_22_if_empty_n,
    input wire                                           out_dist_22_if_full_n,
    output wire                                          out_dist_22_if_read,
    output wire                                          out_dist_22_if_read_ce,
    output wire                                          out_dist_22_if_write,
    output wire                                          out_dist_22_if_write_ce,
    output wire                                          out_dist_22_reset,
    output wire                                          out_dist_23_clk,
    output wire [                                  65:0] out_dist_23_if_din,
    input wire  [                                  65:0] out_dist_23_if_dout,
    input wire                                           out_dist_23_if_empty_n,
    input wire                                           out_dist_23_if_full_n,
    output wire                                          out_dist_23_if_read,
    output wire                                          out_dist_23_if_read_ce,
    output wire                                          out_dist_23_if_write,
    output wire                                          out_dist_23_if_write_ce,
    output wire                                          out_dist_23_reset,
    output wire                                          out_dist_24_clk,
    output wire [                                  65:0] out_dist_24_if_din,
    input wire  [                                  65:0] out_dist_24_if_dout,
    input wire                                           out_dist_24_if_empty_n,
    input wire                                           out_dist_24_if_full_n,
    output wire                                          out_dist_24_if_read,
    output wire                                          out_dist_24_if_read_ce,
    output wire                                          out_dist_24_if_write,
    output wire                                          out_dist_24_if_write_ce,
    output wire                                          out_dist_24_reset,
    output wire                                          out_dist_25_clk,
    output wire [                                  65:0] out_dist_25_if_din,
    input wire  [                                  65:0] out_dist_25_if_dout,
    input wire                                           out_dist_25_if_empty_n,
    input wire                                           out_dist_25_if_full_n,
    output wire                                          out_dist_25_if_read,
    output wire                                          out_dist_25_if_read_ce,
    output wire                                          out_dist_25_if_write,
    output wire                                          out_dist_25_if_write_ce,
    output wire                                          out_dist_25_reset,
    output wire                                          out_dist_26_clk,
    output wire [                                  65:0] out_dist_26_if_din,
    input wire  [                                  65:0] out_dist_26_if_dout,
    input wire                                           out_dist_26_if_empty_n,
    input wire                                           out_dist_26_if_full_n,
    output wire                                          out_dist_26_if_read,
    output wire                                          out_dist_26_if_read_ce,
    output wire                                          out_dist_26_if_write,
    output wire                                          out_dist_26_if_write_ce,
    output wire                                          out_dist_26_reset,
    output wire                                          out_dist_27_clk,
    output wire [                                  65:0] out_dist_27_if_din,
    input wire  [                                  65:0] out_dist_27_if_dout,
    input wire                                           out_dist_27_if_empty_n,
    input wire                                           out_dist_27_if_full_n,
    output wire                                          out_dist_27_if_read,
    output wire                                          out_dist_27_if_read_ce,
    output wire                                          out_dist_27_if_write,
    output wire                                          out_dist_27_if_write_ce,
    output wire                                          out_dist_27_reset,
    output wire                                          out_dist_28_clk,
    output wire [                                  65:0] out_dist_28_if_din,
    input wire  [                                  65:0] out_dist_28_if_dout,
    input wire                                           out_dist_28_if_empty_n,
    input wire                                           out_dist_28_if_full_n,
    output wire                                          out_dist_28_if_read,
    output wire                                          out_dist_28_if_read_ce,
    output wire                                          out_dist_28_if_write,
    output wire                                          out_dist_28_if_write_ce,
    output wire                                          out_dist_28_reset,
    output wire                                          out_dist_29_clk,
    output wire [                                  65:0] out_dist_29_if_din,
    input wire  [                                  65:0] out_dist_29_if_dout,
    input wire                                           out_dist_29_if_empty_n,
    input wire                                           out_dist_29_if_full_n,
    output wire                                          out_dist_29_if_read,
    output wire                                          out_dist_29_if_read_ce,
    output wire                                          out_dist_29_if_write,
    output wire                                          out_dist_29_if_write_ce,
    output wire                                          out_dist_29_reset,
    output wire                                          out_dist_2_clk,
    output wire [                                  65:0] out_dist_2_if_din,
    input wire  [                                  65:0] out_dist_2_if_dout,
    input wire                                           out_dist_2_if_empty_n,
    input wire                                           out_dist_2_if_full_n,
    output wire                                          out_dist_2_if_read,
    output wire                                          out_dist_2_if_read_ce,
    output wire                                          out_dist_2_if_write,
    output wire                                          out_dist_2_if_write_ce,
    output wire                                          out_dist_2_reset,
    output wire                                          out_dist_30_clk,
    output wire [                                  65:0] out_dist_30_if_din,
    input wire  [                                  65:0] out_dist_30_if_dout,
    input wire                                           out_dist_30_if_empty_n,
    input wire                                           out_dist_30_if_full_n,
    output wire                                          out_dist_30_if_read,
    output wire                                          out_dist_30_if_read_ce,
    output wire                                          out_dist_30_if_write,
    output wire                                          out_dist_30_if_write_ce,
    output wire                                          out_dist_30_reset,
    output wire                                          out_dist_31_clk,
    output wire [                                  65:0] out_dist_31_if_din,
    input wire  [                                  65:0] out_dist_31_if_dout,
    input wire                                           out_dist_31_if_empty_n,
    input wire                                           out_dist_31_if_full_n,
    output wire                                          out_dist_31_if_read,
    output wire                                          out_dist_31_if_read_ce,
    output wire                                          out_dist_31_if_write,
    output wire                                          out_dist_31_if_write_ce,
    output wire                                          out_dist_31_reset,
    output wire                                          out_dist_32_clk,
    output wire [                                  65:0] out_dist_32_if_din,
    input wire  [                                  65:0] out_dist_32_if_dout,
    input wire                                           out_dist_32_if_empty_n,
    input wire                                           out_dist_32_if_full_n,
    output wire                                          out_dist_32_if_read,
    output wire                                          out_dist_32_if_read_ce,
    output wire                                          out_dist_32_if_write,
    output wire                                          out_dist_32_if_write_ce,
    output wire                                          out_dist_32_reset,
    output wire                                          out_dist_33_clk,
    output wire [                                  65:0] out_dist_33_if_din,
    input wire  [                                  65:0] out_dist_33_if_dout,
    input wire                                           out_dist_33_if_empty_n,
    input wire                                           out_dist_33_if_full_n,
    output wire                                          out_dist_33_if_read,
    output wire                                          out_dist_33_if_read_ce,
    output wire                                          out_dist_33_if_write,
    output wire                                          out_dist_33_if_write_ce,
    output wire                                          out_dist_33_reset,
    output wire                                          out_dist_34_clk,
    output wire [                                  65:0] out_dist_34_if_din,
    input wire  [                                  65:0] out_dist_34_if_dout,
    input wire                                           out_dist_34_if_empty_n,
    input wire                                           out_dist_34_if_full_n,
    output wire                                          out_dist_34_if_read,
    output wire                                          out_dist_34_if_read_ce,
    output wire                                          out_dist_34_if_write,
    output wire                                          out_dist_34_if_write_ce,
    output wire                                          out_dist_34_reset,
    output wire                                          out_dist_35_clk,
    output wire [                                  65:0] out_dist_35_if_din,
    input wire  [                                  65:0] out_dist_35_if_dout,
    input wire                                           out_dist_35_if_empty_n,
    input wire                                           out_dist_35_if_full_n,
    output wire                                          out_dist_35_if_read,
    output wire                                          out_dist_35_if_read_ce,
    output wire                                          out_dist_35_if_write,
    output wire                                          out_dist_35_if_write_ce,
    output wire                                          out_dist_35_reset,
    output wire                                          out_dist_36_clk,
    output wire [                                  65:0] out_dist_36_if_din,
    input wire  [                                  65:0] out_dist_36_if_dout,
    input wire                                           out_dist_36_if_empty_n,
    input wire                                           out_dist_36_if_full_n,
    output wire                                          out_dist_36_if_read,
    output wire                                          out_dist_36_if_read_ce,
    output wire                                          out_dist_36_if_write,
    output wire                                          out_dist_36_if_write_ce,
    output wire                                          out_dist_36_reset,
    output wire                                          out_dist_37_clk,
    output wire [                                  65:0] out_dist_37_if_din,
    input wire  [                                  65:0] out_dist_37_if_dout,
    input wire                                           out_dist_37_if_empty_n,
    input wire                                           out_dist_37_if_full_n,
    output wire                                          out_dist_37_if_read,
    output wire                                          out_dist_37_if_read_ce,
    output wire                                          out_dist_37_if_write,
    output wire                                          out_dist_37_if_write_ce,
    output wire                                          out_dist_37_reset,
    output wire                                          out_dist_38_clk,
    output wire [                                  65:0] out_dist_38_if_din,
    input wire  [                                  65:0] out_dist_38_if_dout,
    input wire                                           out_dist_38_if_empty_n,
    input wire                                           out_dist_38_if_full_n,
    output wire                                          out_dist_38_if_read,
    output wire                                          out_dist_38_if_read_ce,
    output wire                                          out_dist_38_if_write,
    output wire                                          out_dist_38_if_write_ce,
    output wire                                          out_dist_38_reset,
    output wire                                          out_dist_39_clk,
    output wire [                                  65:0] out_dist_39_if_din,
    input wire  [                                  65:0] out_dist_39_if_dout,
    input wire                                           out_dist_39_if_empty_n,
    input wire                                           out_dist_39_if_full_n,
    output wire                                          out_dist_39_if_read,
    output wire                                          out_dist_39_if_read_ce,
    output wire                                          out_dist_39_if_write,
    output wire                                          out_dist_39_if_write_ce,
    output wire                                          out_dist_39_reset,
    output wire                                          out_dist_3_clk,
    output wire [                                  65:0] out_dist_3_if_din,
    input wire  [                                  65:0] out_dist_3_if_dout,
    input wire                                           out_dist_3_if_empty_n,
    input wire                                           out_dist_3_if_full_n,
    output wire                                          out_dist_3_if_read,
    output wire                                          out_dist_3_if_read_ce,
    output wire                                          out_dist_3_if_write,
    output wire                                          out_dist_3_if_write_ce,
    output wire                                          out_dist_3_reset,
    output wire                                          out_dist_40_clk,
    output wire [                                  65:0] out_dist_40_if_din,
    input wire  [                                  65:0] out_dist_40_if_dout,
    input wire                                           out_dist_40_if_empty_n,
    input wire                                           out_dist_40_if_full_n,
    output wire                                          out_dist_40_if_read,
    output wire                                          out_dist_40_if_read_ce,
    output wire                                          out_dist_40_if_write,
    output wire                                          out_dist_40_if_write_ce,
    output wire                                          out_dist_40_reset,
    output wire                                          out_dist_41_clk,
    output wire [                                  65:0] out_dist_41_if_din,
    input wire  [                                  65:0] out_dist_41_if_dout,
    input wire                                           out_dist_41_if_empty_n,
    input wire                                           out_dist_41_if_full_n,
    output wire                                          out_dist_41_if_read,
    output wire                                          out_dist_41_if_read_ce,
    output wire                                          out_dist_41_if_write,
    output wire                                          out_dist_41_if_write_ce,
    output wire                                          out_dist_41_reset,
    output wire                                          out_dist_42_clk,
    output wire [                                  65:0] out_dist_42_if_din,
    input wire  [                                  65:0] out_dist_42_if_dout,
    input wire                                           out_dist_42_if_empty_n,
    input wire                                           out_dist_42_if_full_n,
    output wire                                          out_dist_42_if_read,
    output wire                                          out_dist_42_if_read_ce,
    output wire                                          out_dist_42_if_write,
    output wire                                          out_dist_42_if_write_ce,
    output wire                                          out_dist_42_reset,
    output wire                                          out_dist_43_clk,
    output wire [                                  65:0] out_dist_43_if_din,
    input wire  [                                  65:0] out_dist_43_if_dout,
    input wire                                           out_dist_43_if_empty_n,
    input wire                                           out_dist_43_if_full_n,
    output wire                                          out_dist_43_if_read,
    output wire                                          out_dist_43_if_read_ce,
    output wire                                          out_dist_43_if_write,
    output wire                                          out_dist_43_if_write_ce,
    output wire                                          out_dist_43_reset,
    output wire                                          out_dist_44_clk,
    output wire [                                  65:0] out_dist_44_if_din,
    input wire  [                                  65:0] out_dist_44_if_dout,
    input wire                                           out_dist_44_if_empty_n,
    input wire                                           out_dist_44_if_full_n,
    output wire                                          out_dist_44_if_read,
    output wire                                          out_dist_44_if_read_ce,
    output wire                                          out_dist_44_if_write,
    output wire                                          out_dist_44_if_write_ce,
    output wire                                          out_dist_44_reset,
    output wire                                          out_dist_45_clk,
    output wire [                                  65:0] out_dist_45_if_din,
    input wire  [                                  65:0] out_dist_45_if_dout,
    input wire                                           out_dist_45_if_empty_n,
    input wire                                           out_dist_45_if_full_n,
    output wire                                          out_dist_45_if_read,
    output wire                                          out_dist_45_if_read_ce,
    output wire                                          out_dist_45_if_write,
    output wire                                          out_dist_45_if_write_ce,
    output wire                                          out_dist_45_reset,
    output wire                                          out_dist_46_clk,
    output wire [                                  65:0] out_dist_46_if_din,
    input wire  [                                  65:0] out_dist_46_if_dout,
    input wire                                           out_dist_46_if_empty_n,
    input wire                                           out_dist_46_if_full_n,
    output wire                                          out_dist_46_if_read,
    output wire                                          out_dist_46_if_read_ce,
    output wire                                          out_dist_46_if_write,
    output wire                                          out_dist_46_if_write_ce,
    output wire                                          out_dist_46_reset,
    output wire                                          out_dist_47_clk,
    output wire [                                  65:0] out_dist_47_if_din,
    input wire  [                                  65:0] out_dist_47_if_dout,
    input wire                                           out_dist_47_if_empty_n,
    input wire                                           out_dist_47_if_full_n,
    output wire                                          out_dist_47_if_read,
    output wire                                          out_dist_47_if_read_ce,
    output wire                                          out_dist_47_if_write,
    output wire                                          out_dist_47_if_write_ce,
    output wire                                          out_dist_47_reset,
    output wire                                          out_dist_48_clk,
    output wire [                                  65:0] out_dist_48_if_din,
    input wire  [                                  65:0] out_dist_48_if_dout,
    input wire                                           out_dist_48_if_empty_n,
    input wire                                           out_dist_48_if_full_n,
    output wire                                          out_dist_48_if_read,
    output wire                                          out_dist_48_if_read_ce,
    output wire                                          out_dist_48_if_write,
    output wire                                          out_dist_48_if_write_ce,
    output wire                                          out_dist_48_reset,
    output wire                                          out_dist_49_clk,
    output wire [                                  65:0] out_dist_49_if_din,
    input wire  [                                  65:0] out_dist_49_if_dout,
    input wire                                           out_dist_49_if_empty_n,
    input wire                                           out_dist_49_if_full_n,
    output wire                                          out_dist_49_if_read,
    output wire                                          out_dist_49_if_read_ce,
    output wire                                          out_dist_49_if_write,
    output wire                                          out_dist_49_if_write_ce,
    output wire                                          out_dist_49_reset,
    output wire                                          out_dist_4_clk,
    output wire [                                  65:0] out_dist_4_if_din,
    input wire  [                                  65:0] out_dist_4_if_dout,
    input wire                                           out_dist_4_if_empty_n,
    input wire                                           out_dist_4_if_full_n,
    output wire                                          out_dist_4_if_read,
    output wire                                          out_dist_4_if_read_ce,
    output wire                                          out_dist_4_if_write,
    output wire                                          out_dist_4_if_write_ce,
    output wire                                          out_dist_4_reset,
    output wire                                          out_dist_50_clk,
    output wire [                                  65:0] out_dist_50_if_din,
    input wire  [                                  65:0] out_dist_50_if_dout,
    input wire                                           out_dist_50_if_empty_n,
    input wire                                           out_dist_50_if_full_n,
    output wire                                          out_dist_50_if_read,
    output wire                                          out_dist_50_if_read_ce,
    output wire                                          out_dist_50_if_write,
    output wire                                          out_dist_50_if_write_ce,
    output wire                                          out_dist_50_reset,
    output wire                                          out_dist_51_clk,
    output wire [                                  65:0] out_dist_51_if_din,
    input wire  [                                  65:0] out_dist_51_if_dout,
    input wire                                           out_dist_51_if_empty_n,
    input wire                                           out_dist_51_if_full_n,
    output wire                                          out_dist_51_if_read,
    output wire                                          out_dist_51_if_read_ce,
    output wire                                          out_dist_51_if_write,
    output wire                                          out_dist_51_if_write_ce,
    output wire                                          out_dist_51_reset,
    output wire                                          out_dist_52_clk,
    output wire [                                  65:0] out_dist_52_if_din,
    input wire  [                                  65:0] out_dist_52_if_dout,
    input wire                                           out_dist_52_if_empty_n,
    input wire                                           out_dist_52_if_full_n,
    output wire                                          out_dist_52_if_read,
    output wire                                          out_dist_52_if_read_ce,
    output wire                                          out_dist_52_if_write,
    output wire                                          out_dist_52_if_write_ce,
    output wire                                          out_dist_52_reset,
    output wire                                          out_dist_53_clk,
    output wire [                                  65:0] out_dist_53_if_din,
    input wire  [                                  65:0] out_dist_53_if_dout,
    input wire                                           out_dist_53_if_empty_n,
    input wire                                           out_dist_53_if_full_n,
    output wire                                          out_dist_53_if_read,
    output wire                                          out_dist_53_if_read_ce,
    output wire                                          out_dist_53_if_write,
    output wire                                          out_dist_53_if_write_ce,
    output wire                                          out_dist_53_reset,
    output wire                                          out_dist_5_clk,
    output wire [                                  65:0] out_dist_5_if_din,
    input wire  [                                  65:0] out_dist_5_if_dout,
    input wire                                           out_dist_5_if_empty_n,
    input wire                                           out_dist_5_if_full_n,
    output wire                                          out_dist_5_if_read,
    output wire                                          out_dist_5_if_read_ce,
    output wire                                          out_dist_5_if_write,
    output wire                                          out_dist_5_if_write_ce,
    output wire                                          out_dist_5_reset,
    output wire                                          out_dist_6_clk,
    output wire [                                  65:0] out_dist_6_if_din,
    input wire  [                                  65:0] out_dist_6_if_dout,
    input wire                                           out_dist_6_if_empty_n,
    input wire                                           out_dist_6_if_full_n,
    output wire                                          out_dist_6_if_read,
    output wire                                          out_dist_6_if_read_ce,
    output wire                                          out_dist_6_if_write,
    output wire                                          out_dist_6_if_write_ce,
    output wire                                          out_dist_6_reset,
    output wire                                          out_dist_7_clk,
    output wire [                                  65:0] out_dist_7_if_din,
    input wire  [                                  65:0] out_dist_7_if_dout,
    input wire                                           out_dist_7_if_empty_n,
    input wire                                           out_dist_7_if_full_n,
    output wire                                          out_dist_7_if_read,
    output wire                                          out_dist_7_if_read_ce,
    output wire                                          out_dist_7_if_write,
    output wire                                          out_dist_7_if_write_ce,
    output wire                                          out_dist_7_reset,
    output wire                                          out_dist_8_clk,
    output wire [                                  65:0] out_dist_8_if_din,
    input wire  [                                  65:0] out_dist_8_if_dout,
    input wire                                           out_dist_8_if_empty_n,
    input wire                                           out_dist_8_if_full_n,
    output wire                                          out_dist_8_if_read,
    output wire                                          out_dist_8_if_read_ce,
    output wire                                          out_dist_8_if_write,
    output wire                                          out_dist_8_if_write_ce,
    output wire                                          out_dist_8_reset,
    output wire                                          out_dist_9_clk,
    output wire [                                  65:0] out_dist_9_if_din,
    input wire  [                                  65:0] out_dist_9_if_dout,
    input wire                                           out_dist_9_if_empty_n,
    input wire                                           out_dist_9_if_full_n,
    output wire                                          out_dist_9_if_read,
    output wire                                          out_dist_9_if_read_ce,
    output wire                                          out_dist_9_if_write,
    output wire                                          out_dist_9_if_write_ce,
    output wire                                          out_dist_9_reset,
    output wire                                          out_id_0_clk,
    output wire [                                  65:0] out_id_0_if_din,
    input wire  [                                  65:0] out_id_0_if_dout,
    input wire                                           out_id_0_if_empty_n,
    input wire                                           out_id_0_if_full_n,
    output wire                                          out_id_0_if_read,
    output wire                                          out_id_0_if_read_ce,
    output wire                                          out_id_0_if_write,
    output wire                                          out_id_0_if_write_ce,
    output wire                                          out_id_0_reset,
    output wire                                          out_id_10_clk,
    output wire [                                  65:0] out_id_10_if_din,
    input wire  [                                  65:0] out_id_10_if_dout,
    input wire                                           out_id_10_if_empty_n,
    input wire                                           out_id_10_if_full_n,
    output wire                                          out_id_10_if_read,
    output wire                                          out_id_10_if_read_ce,
    output wire                                          out_id_10_if_write,
    output wire                                          out_id_10_if_write_ce,
    output wire                                          out_id_10_reset,
    output wire                                          out_id_11_clk,
    output wire [                                  65:0] out_id_11_if_din,
    input wire  [                                  65:0] out_id_11_if_dout,
    input wire                                           out_id_11_if_empty_n,
    input wire                                           out_id_11_if_full_n,
    output wire                                          out_id_11_if_read,
    output wire                                          out_id_11_if_read_ce,
    output wire                                          out_id_11_if_write,
    output wire                                          out_id_11_if_write_ce,
    output wire                                          out_id_11_reset,
    output wire                                          out_id_12_clk,
    output wire [                                  65:0] out_id_12_if_din,
    input wire  [                                  65:0] out_id_12_if_dout,
    input wire                                           out_id_12_if_empty_n,
    input wire                                           out_id_12_if_full_n,
    output wire                                          out_id_12_if_read,
    output wire                                          out_id_12_if_read_ce,
    output wire                                          out_id_12_if_write,
    output wire                                          out_id_12_if_write_ce,
    output wire                                          out_id_12_reset,
    output wire                                          out_id_13_clk,
    output wire [                                  65:0] out_id_13_if_din,
    input wire  [                                  65:0] out_id_13_if_dout,
    input wire                                           out_id_13_if_empty_n,
    input wire                                           out_id_13_if_full_n,
    output wire                                          out_id_13_if_read,
    output wire                                          out_id_13_if_read_ce,
    output wire                                          out_id_13_if_write,
    output wire                                          out_id_13_if_write_ce,
    output wire                                          out_id_13_reset,
    output wire                                          out_id_14_clk,
    output wire [                                  65:0] out_id_14_if_din,
    input wire  [                                  65:0] out_id_14_if_dout,
    input wire                                           out_id_14_if_empty_n,
    input wire                                           out_id_14_if_full_n,
    output wire                                          out_id_14_if_read,
    output wire                                          out_id_14_if_read_ce,
    output wire                                          out_id_14_if_write,
    output wire                                          out_id_14_if_write_ce,
    output wire                                          out_id_14_reset,
    output wire                                          out_id_15_clk,
    output wire [                                  65:0] out_id_15_if_din,
    input wire  [                                  65:0] out_id_15_if_dout,
    input wire                                           out_id_15_if_empty_n,
    input wire                                           out_id_15_if_full_n,
    output wire                                          out_id_15_if_read,
    output wire                                          out_id_15_if_read_ce,
    output wire                                          out_id_15_if_write,
    output wire                                          out_id_15_if_write_ce,
    output wire                                          out_id_15_reset,
    output wire                                          out_id_16_clk,
    output wire [                                  65:0] out_id_16_if_din,
    input wire  [                                  65:0] out_id_16_if_dout,
    input wire                                           out_id_16_if_empty_n,
    input wire                                           out_id_16_if_full_n,
    output wire                                          out_id_16_if_read,
    output wire                                          out_id_16_if_read_ce,
    output wire                                          out_id_16_if_write,
    output wire                                          out_id_16_if_write_ce,
    output wire                                          out_id_16_reset,
    output wire                                          out_id_17_clk,
    output wire [                                  65:0] out_id_17_if_din,
    input wire  [                                  65:0] out_id_17_if_dout,
    input wire                                           out_id_17_if_empty_n,
    input wire                                           out_id_17_if_full_n,
    output wire                                          out_id_17_if_read,
    output wire                                          out_id_17_if_read_ce,
    output wire                                          out_id_17_if_write,
    output wire                                          out_id_17_if_write_ce,
    output wire                                          out_id_17_reset,
    output wire                                          out_id_18_clk,
    output wire [                                  65:0] out_id_18_if_din,
    input wire  [                                  65:0] out_id_18_if_dout,
    input wire                                           out_id_18_if_empty_n,
    input wire                                           out_id_18_if_full_n,
    output wire                                          out_id_18_if_read,
    output wire                                          out_id_18_if_read_ce,
    output wire                                          out_id_18_if_write,
    output wire                                          out_id_18_if_write_ce,
    output wire                                          out_id_18_reset,
    output wire                                          out_id_19_clk,
    output wire [                                  65:0] out_id_19_if_din,
    input wire  [                                  65:0] out_id_19_if_dout,
    input wire                                           out_id_19_if_empty_n,
    input wire                                           out_id_19_if_full_n,
    output wire                                          out_id_19_if_read,
    output wire                                          out_id_19_if_read_ce,
    output wire                                          out_id_19_if_write,
    output wire                                          out_id_19_if_write_ce,
    output wire                                          out_id_19_reset,
    output wire                                          out_id_1_clk,
    output wire [                                  65:0] out_id_1_if_din,
    input wire  [                                  65:0] out_id_1_if_dout,
    input wire                                           out_id_1_if_empty_n,
    input wire                                           out_id_1_if_full_n,
    output wire                                          out_id_1_if_read,
    output wire                                          out_id_1_if_read_ce,
    output wire                                          out_id_1_if_write,
    output wire                                          out_id_1_if_write_ce,
    output wire                                          out_id_1_reset,
    output wire                                          out_id_20_clk,
    output wire [                                  65:0] out_id_20_if_din,
    input wire  [                                  65:0] out_id_20_if_dout,
    input wire                                           out_id_20_if_empty_n,
    input wire                                           out_id_20_if_full_n,
    output wire                                          out_id_20_if_read,
    output wire                                          out_id_20_if_read_ce,
    output wire                                          out_id_20_if_write,
    output wire                                          out_id_20_if_write_ce,
    output wire                                          out_id_20_reset,
    output wire                                          out_id_21_clk,
    output wire [                                  65:0] out_id_21_if_din,
    input wire  [                                  65:0] out_id_21_if_dout,
    input wire                                           out_id_21_if_empty_n,
    input wire                                           out_id_21_if_full_n,
    output wire                                          out_id_21_if_read,
    output wire                                          out_id_21_if_read_ce,
    output wire                                          out_id_21_if_write,
    output wire                                          out_id_21_if_write_ce,
    output wire                                          out_id_21_reset,
    output wire                                          out_id_22_clk,
    output wire [                                  65:0] out_id_22_if_din,
    input wire  [                                  65:0] out_id_22_if_dout,
    input wire                                           out_id_22_if_empty_n,
    input wire                                           out_id_22_if_full_n,
    output wire                                          out_id_22_if_read,
    output wire                                          out_id_22_if_read_ce,
    output wire                                          out_id_22_if_write,
    output wire                                          out_id_22_if_write_ce,
    output wire                                          out_id_22_reset,
    output wire                                          out_id_23_clk,
    output wire [                                  65:0] out_id_23_if_din,
    input wire  [                                  65:0] out_id_23_if_dout,
    input wire                                           out_id_23_if_empty_n,
    input wire                                           out_id_23_if_full_n,
    output wire                                          out_id_23_if_read,
    output wire                                          out_id_23_if_read_ce,
    output wire                                          out_id_23_if_write,
    output wire                                          out_id_23_if_write_ce,
    output wire                                          out_id_23_reset,
    output wire                                          out_id_24_clk,
    output wire [                                  65:0] out_id_24_if_din,
    input wire  [                                  65:0] out_id_24_if_dout,
    input wire                                           out_id_24_if_empty_n,
    input wire                                           out_id_24_if_full_n,
    output wire                                          out_id_24_if_read,
    output wire                                          out_id_24_if_read_ce,
    output wire                                          out_id_24_if_write,
    output wire                                          out_id_24_if_write_ce,
    output wire                                          out_id_24_reset,
    output wire                                          out_id_25_clk,
    output wire [                                  65:0] out_id_25_if_din,
    input wire  [                                  65:0] out_id_25_if_dout,
    input wire                                           out_id_25_if_empty_n,
    input wire                                           out_id_25_if_full_n,
    output wire                                          out_id_25_if_read,
    output wire                                          out_id_25_if_read_ce,
    output wire                                          out_id_25_if_write,
    output wire                                          out_id_25_if_write_ce,
    output wire                                          out_id_25_reset,
    output wire                                          out_id_26_clk,
    output wire [                                  65:0] out_id_26_if_din,
    input wire  [                                  65:0] out_id_26_if_dout,
    input wire                                           out_id_26_if_empty_n,
    input wire                                           out_id_26_if_full_n,
    output wire                                          out_id_26_if_read,
    output wire                                          out_id_26_if_read_ce,
    output wire                                          out_id_26_if_write,
    output wire                                          out_id_26_if_write_ce,
    output wire                                          out_id_26_reset,
    output wire                                          out_id_27_clk,
    output wire [                                  65:0] out_id_27_if_din,
    input wire  [                                  65:0] out_id_27_if_dout,
    input wire                                           out_id_27_if_empty_n,
    input wire                                           out_id_27_if_full_n,
    output wire                                          out_id_27_if_read,
    output wire                                          out_id_27_if_read_ce,
    output wire                                          out_id_27_if_write,
    output wire                                          out_id_27_if_write_ce,
    output wire                                          out_id_27_reset,
    output wire                                          out_id_28_clk,
    output wire [                                  65:0] out_id_28_if_din,
    input wire  [                                  65:0] out_id_28_if_dout,
    input wire                                           out_id_28_if_empty_n,
    input wire                                           out_id_28_if_full_n,
    output wire                                          out_id_28_if_read,
    output wire                                          out_id_28_if_read_ce,
    output wire                                          out_id_28_if_write,
    output wire                                          out_id_28_if_write_ce,
    output wire                                          out_id_28_reset,
    output wire                                          out_id_29_clk,
    output wire [                                  65:0] out_id_29_if_din,
    input wire  [                                  65:0] out_id_29_if_dout,
    input wire                                           out_id_29_if_empty_n,
    input wire                                           out_id_29_if_full_n,
    output wire                                          out_id_29_if_read,
    output wire                                          out_id_29_if_read_ce,
    output wire                                          out_id_29_if_write,
    output wire                                          out_id_29_if_write_ce,
    output wire                                          out_id_29_reset,
    output wire                                          out_id_2_clk,
    output wire [                                  65:0] out_id_2_if_din,
    input wire  [                                  65:0] out_id_2_if_dout,
    input wire                                           out_id_2_if_empty_n,
    input wire                                           out_id_2_if_full_n,
    output wire                                          out_id_2_if_read,
    output wire                                          out_id_2_if_read_ce,
    output wire                                          out_id_2_if_write,
    output wire                                          out_id_2_if_write_ce,
    output wire                                          out_id_2_reset,
    output wire                                          out_id_30_clk,
    output wire [                                  65:0] out_id_30_if_din,
    input wire  [                                  65:0] out_id_30_if_dout,
    input wire                                           out_id_30_if_empty_n,
    input wire                                           out_id_30_if_full_n,
    output wire                                          out_id_30_if_read,
    output wire                                          out_id_30_if_read_ce,
    output wire                                          out_id_30_if_write,
    output wire                                          out_id_30_if_write_ce,
    output wire                                          out_id_30_reset,
    output wire                                          out_id_31_clk,
    output wire [                                  65:0] out_id_31_if_din,
    input wire  [                                  65:0] out_id_31_if_dout,
    input wire                                           out_id_31_if_empty_n,
    input wire                                           out_id_31_if_full_n,
    output wire                                          out_id_31_if_read,
    output wire                                          out_id_31_if_read_ce,
    output wire                                          out_id_31_if_write,
    output wire                                          out_id_31_if_write_ce,
    output wire                                          out_id_31_reset,
    output wire                                          out_id_32_clk,
    output wire [                                  65:0] out_id_32_if_din,
    input wire  [                                  65:0] out_id_32_if_dout,
    input wire                                           out_id_32_if_empty_n,
    input wire                                           out_id_32_if_full_n,
    output wire                                          out_id_32_if_read,
    output wire                                          out_id_32_if_read_ce,
    output wire                                          out_id_32_if_write,
    output wire                                          out_id_32_if_write_ce,
    output wire                                          out_id_32_reset,
    output wire                                          out_id_33_clk,
    output wire [                                  65:0] out_id_33_if_din,
    input wire  [                                  65:0] out_id_33_if_dout,
    input wire                                           out_id_33_if_empty_n,
    input wire                                           out_id_33_if_full_n,
    output wire                                          out_id_33_if_read,
    output wire                                          out_id_33_if_read_ce,
    output wire                                          out_id_33_if_write,
    output wire                                          out_id_33_if_write_ce,
    output wire                                          out_id_33_reset,
    output wire                                          out_id_34_clk,
    output wire [                                  65:0] out_id_34_if_din,
    input wire  [                                  65:0] out_id_34_if_dout,
    input wire                                           out_id_34_if_empty_n,
    input wire                                           out_id_34_if_full_n,
    output wire                                          out_id_34_if_read,
    output wire                                          out_id_34_if_read_ce,
    output wire                                          out_id_34_if_write,
    output wire                                          out_id_34_if_write_ce,
    output wire                                          out_id_34_reset,
    output wire                                          out_id_35_clk,
    output wire [                                  65:0] out_id_35_if_din,
    input wire  [                                  65:0] out_id_35_if_dout,
    input wire                                           out_id_35_if_empty_n,
    input wire                                           out_id_35_if_full_n,
    output wire                                          out_id_35_if_read,
    output wire                                          out_id_35_if_read_ce,
    output wire                                          out_id_35_if_write,
    output wire                                          out_id_35_if_write_ce,
    output wire                                          out_id_35_reset,
    output wire                                          out_id_36_clk,
    output wire [                                  65:0] out_id_36_if_din,
    input wire  [                                  65:0] out_id_36_if_dout,
    input wire                                           out_id_36_if_empty_n,
    input wire                                           out_id_36_if_full_n,
    output wire                                          out_id_36_if_read,
    output wire                                          out_id_36_if_read_ce,
    output wire                                          out_id_36_if_write,
    output wire                                          out_id_36_if_write_ce,
    output wire                                          out_id_36_reset,
    output wire                                          out_id_37_clk,
    output wire [                                  65:0] out_id_37_if_din,
    input wire  [                                  65:0] out_id_37_if_dout,
    input wire                                           out_id_37_if_empty_n,
    input wire                                           out_id_37_if_full_n,
    output wire                                          out_id_37_if_read,
    output wire                                          out_id_37_if_read_ce,
    output wire                                          out_id_37_if_write,
    output wire                                          out_id_37_if_write_ce,
    output wire                                          out_id_37_reset,
    output wire                                          out_id_38_clk,
    output wire [                                  65:0] out_id_38_if_din,
    input wire  [                                  65:0] out_id_38_if_dout,
    input wire                                           out_id_38_if_empty_n,
    input wire                                           out_id_38_if_full_n,
    output wire                                          out_id_38_if_read,
    output wire                                          out_id_38_if_read_ce,
    output wire                                          out_id_38_if_write,
    output wire                                          out_id_38_if_write_ce,
    output wire                                          out_id_38_reset,
    output wire                                          out_id_39_clk,
    output wire [                                  65:0] out_id_39_if_din,
    input wire  [                                  65:0] out_id_39_if_dout,
    input wire                                           out_id_39_if_empty_n,
    input wire                                           out_id_39_if_full_n,
    output wire                                          out_id_39_if_read,
    output wire                                          out_id_39_if_read_ce,
    output wire                                          out_id_39_if_write,
    output wire                                          out_id_39_if_write_ce,
    output wire                                          out_id_39_reset,
    output wire                                          out_id_3_clk,
    output wire [                                  65:0] out_id_3_if_din,
    input wire  [                                  65:0] out_id_3_if_dout,
    input wire                                           out_id_3_if_empty_n,
    input wire                                           out_id_3_if_full_n,
    output wire                                          out_id_3_if_read,
    output wire                                          out_id_3_if_read_ce,
    output wire                                          out_id_3_if_write,
    output wire                                          out_id_3_if_write_ce,
    output wire                                          out_id_3_reset,
    output wire                                          out_id_40_clk,
    output wire [                                  65:0] out_id_40_if_din,
    input wire  [                                  65:0] out_id_40_if_dout,
    input wire                                           out_id_40_if_empty_n,
    input wire                                           out_id_40_if_full_n,
    output wire                                          out_id_40_if_read,
    output wire                                          out_id_40_if_read_ce,
    output wire                                          out_id_40_if_write,
    output wire                                          out_id_40_if_write_ce,
    output wire                                          out_id_40_reset,
    output wire                                          out_id_41_clk,
    output wire [                                  65:0] out_id_41_if_din,
    input wire  [                                  65:0] out_id_41_if_dout,
    input wire                                           out_id_41_if_empty_n,
    input wire                                           out_id_41_if_full_n,
    output wire                                          out_id_41_if_read,
    output wire                                          out_id_41_if_read_ce,
    output wire                                          out_id_41_if_write,
    output wire                                          out_id_41_if_write_ce,
    output wire                                          out_id_41_reset,
    output wire                                          out_id_42_clk,
    output wire [                                  65:0] out_id_42_if_din,
    input wire  [                                  65:0] out_id_42_if_dout,
    input wire                                           out_id_42_if_empty_n,
    input wire                                           out_id_42_if_full_n,
    output wire                                          out_id_42_if_read,
    output wire                                          out_id_42_if_read_ce,
    output wire                                          out_id_42_if_write,
    output wire                                          out_id_42_if_write_ce,
    output wire                                          out_id_42_reset,
    output wire                                          out_id_43_clk,
    output wire [                                  65:0] out_id_43_if_din,
    input wire  [                                  65:0] out_id_43_if_dout,
    input wire                                           out_id_43_if_empty_n,
    input wire                                           out_id_43_if_full_n,
    output wire                                          out_id_43_if_read,
    output wire                                          out_id_43_if_read_ce,
    output wire                                          out_id_43_if_write,
    output wire                                          out_id_43_if_write_ce,
    output wire                                          out_id_43_reset,
    output wire                                          out_id_44_clk,
    output wire [                                  65:0] out_id_44_if_din,
    input wire  [                                  65:0] out_id_44_if_dout,
    input wire                                           out_id_44_if_empty_n,
    input wire                                           out_id_44_if_full_n,
    output wire                                          out_id_44_if_read,
    output wire                                          out_id_44_if_read_ce,
    output wire                                          out_id_44_if_write,
    output wire                                          out_id_44_if_write_ce,
    output wire                                          out_id_44_reset,
    output wire                                          out_id_45_clk,
    output wire [                                  65:0] out_id_45_if_din,
    input wire  [                                  65:0] out_id_45_if_dout,
    input wire                                           out_id_45_if_empty_n,
    input wire                                           out_id_45_if_full_n,
    output wire                                          out_id_45_if_read,
    output wire                                          out_id_45_if_read_ce,
    output wire                                          out_id_45_if_write,
    output wire                                          out_id_45_if_write_ce,
    output wire                                          out_id_45_reset,
    output wire                                          out_id_46_clk,
    output wire [                                  65:0] out_id_46_if_din,
    input wire  [                                  65:0] out_id_46_if_dout,
    input wire                                           out_id_46_if_empty_n,
    input wire                                           out_id_46_if_full_n,
    output wire                                          out_id_46_if_read,
    output wire                                          out_id_46_if_read_ce,
    output wire                                          out_id_46_if_write,
    output wire                                          out_id_46_if_write_ce,
    output wire                                          out_id_46_reset,
    output wire                                          out_id_47_clk,
    output wire [                                  65:0] out_id_47_if_din,
    input wire  [                                  65:0] out_id_47_if_dout,
    input wire                                           out_id_47_if_empty_n,
    input wire                                           out_id_47_if_full_n,
    output wire                                          out_id_47_if_read,
    output wire                                          out_id_47_if_read_ce,
    output wire                                          out_id_47_if_write,
    output wire                                          out_id_47_if_write_ce,
    output wire                                          out_id_47_reset,
    output wire                                          out_id_48_clk,
    output wire [                                  65:0] out_id_48_if_din,
    input wire  [                                  65:0] out_id_48_if_dout,
    input wire                                           out_id_48_if_empty_n,
    input wire                                           out_id_48_if_full_n,
    output wire                                          out_id_48_if_read,
    output wire                                          out_id_48_if_read_ce,
    output wire                                          out_id_48_if_write,
    output wire                                          out_id_48_if_write_ce,
    output wire                                          out_id_48_reset,
    output wire                                          out_id_49_clk,
    output wire [                                  65:0] out_id_49_if_din,
    input wire  [                                  65:0] out_id_49_if_dout,
    input wire                                           out_id_49_if_empty_n,
    input wire                                           out_id_49_if_full_n,
    output wire                                          out_id_49_if_read,
    output wire                                          out_id_49_if_read_ce,
    output wire                                          out_id_49_if_write,
    output wire                                          out_id_49_if_write_ce,
    output wire                                          out_id_49_reset,
    output wire                                          out_id_4_clk,
    output wire [                                  65:0] out_id_4_if_din,
    input wire  [                                  65:0] out_id_4_if_dout,
    input wire                                           out_id_4_if_empty_n,
    input wire                                           out_id_4_if_full_n,
    output wire                                          out_id_4_if_read,
    output wire                                          out_id_4_if_read_ce,
    output wire                                          out_id_4_if_write,
    output wire                                          out_id_4_if_write_ce,
    output wire                                          out_id_4_reset,
    output wire                                          out_id_50_clk,
    output wire [                                  65:0] out_id_50_if_din,
    input wire  [                                  65:0] out_id_50_if_dout,
    input wire                                           out_id_50_if_empty_n,
    input wire                                           out_id_50_if_full_n,
    output wire                                          out_id_50_if_read,
    output wire                                          out_id_50_if_read_ce,
    output wire                                          out_id_50_if_write,
    output wire                                          out_id_50_if_write_ce,
    output wire                                          out_id_50_reset,
    output wire                                          out_id_51_clk,
    output wire [                                  65:0] out_id_51_if_din,
    input wire  [                                  65:0] out_id_51_if_dout,
    input wire                                           out_id_51_if_empty_n,
    input wire                                           out_id_51_if_full_n,
    output wire                                          out_id_51_if_read,
    output wire                                          out_id_51_if_read_ce,
    output wire                                          out_id_51_if_write,
    output wire                                          out_id_51_if_write_ce,
    output wire                                          out_id_51_reset,
    output wire                                          out_id_52_clk,
    output wire [                                  65:0] out_id_52_if_din,
    input wire  [                                  65:0] out_id_52_if_dout,
    input wire                                           out_id_52_if_empty_n,
    input wire                                           out_id_52_if_full_n,
    output wire                                          out_id_52_if_read,
    output wire                                          out_id_52_if_read_ce,
    output wire                                          out_id_52_if_write,
    output wire                                          out_id_52_if_write_ce,
    output wire                                          out_id_52_reset,
    output wire                                          out_id_53_clk,
    output wire [                                  65:0] out_id_53_if_din,
    input wire  [                                  65:0] out_id_53_if_dout,
    input wire                                           out_id_53_if_empty_n,
    input wire                                           out_id_53_if_full_n,
    output wire                                          out_id_53_if_read,
    output wire                                          out_id_53_if_read_ce,
    output wire                                          out_id_53_if_write,
    output wire                                          out_id_53_if_write_ce,
    output wire                                          out_id_53_reset,
    output wire                                          out_id_5_clk,
    output wire [                                  65:0] out_id_5_if_din,
    input wire  [                                  65:0] out_id_5_if_dout,
    input wire                                           out_id_5_if_empty_n,
    input wire                                           out_id_5_if_full_n,
    output wire                                          out_id_5_if_read,
    output wire                                          out_id_5_if_read_ce,
    output wire                                          out_id_5_if_write,
    output wire                                          out_id_5_if_write_ce,
    output wire                                          out_id_5_reset,
    output wire                                          out_id_6_clk,
    output wire [                                  65:0] out_id_6_if_din,
    input wire  [                                  65:0] out_id_6_if_dout,
    input wire                                           out_id_6_if_empty_n,
    input wire                                           out_id_6_if_full_n,
    output wire                                          out_id_6_if_read,
    output wire                                          out_id_6_if_read_ce,
    output wire                                          out_id_6_if_write,
    output wire                                          out_id_6_if_write_ce,
    output wire                                          out_id_6_reset,
    output wire                                          out_id_7_clk,
    output wire [                                  65:0] out_id_7_if_din,
    input wire  [                                  65:0] out_id_7_if_dout,
    input wire                                           out_id_7_if_empty_n,
    input wire                                           out_id_7_if_full_n,
    output wire                                          out_id_7_if_read,
    output wire                                          out_id_7_if_read_ce,
    output wire                                          out_id_7_if_write,
    output wire                                          out_id_7_if_write_ce,
    output wire                                          out_id_7_reset,
    output wire                                          out_id_8_clk,
    output wire [                                  65:0] out_id_8_if_din,
    input wire  [                                  65:0] out_id_8_if_dout,
    input wire                                           out_id_8_if_empty_n,
    input wire                                           out_id_8_if_full_n,
    output wire                                          out_id_8_if_read,
    output wire                                          out_id_8_if_read_ce,
    output wire                                          out_id_8_if_write,
    output wire                                          out_id_8_if_write_ce,
    output wire                                          out_id_8_reset,
    output wire                                          out_id_9_clk,
    output wire [                                  65:0] out_id_9_if_din,
    input wire  [                                  65:0] out_id_9_if_dout,
    input wire                                           out_id_9_if_empty_n,
    input wire                                           out_id_9_if_full_n,
    output wire                                          out_id_9_if_read,
    output wire                                          out_id_9_if_read_ce,
    output wire                                          out_id_9_if_write,
    output wire                                          out_id_9_if_write_ce,
    output wire                                          out_id_9_reset,
    output wire                                          krnl_globalSort_L1_L2_0_ap_clk,
    input wire                                           krnl_globalSort_L1_L2_0_ap_done,
    input wire                                           krnl_globalSort_L1_L2_0_ap_idle,
    input wire                                           krnl_globalSort_L1_L2_0_ap_ready,
    output wire                                          krnl_globalSort_L1_L2_0_ap_rst_n,
    output wire                                          krnl_globalSort_L1_L2_0_ap_start,
    output wire [                                  65:0] krnl_globalSort_L1_L2_0_in_dist0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_0_in_dist0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_0_in_dist0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_0_in_dist0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_0_in_dist0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_0_in_dist0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_0_in_dist1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_0_in_dist1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_0_in_dist1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_0_in_dist1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_0_in_dist1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_0_in_dist1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_0_in_dist2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_0_in_dist2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_0_in_dist2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_0_in_dist2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_0_in_dist2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_0_in_dist2_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_0_in_id0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_0_in_id0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_0_in_id0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_0_in_id0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_0_in_id0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_0_in_id0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_0_in_id1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_0_in_id1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_0_in_id1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_0_in_id1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_0_in_id1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_0_in_id1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_0_in_id2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_0_in_id2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_0_in_id2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_0_in_id2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_0_in_id2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_0_in_id2_s_read,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_0_out_dist_din,
    output wire                                          krnl_globalSort_L1_L2_0_out_dist_full_n,
    input wire                                           krnl_globalSort_L1_L2_0_out_dist_write,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_0_out_id_din,
    output wire                                          krnl_globalSort_L1_L2_0_out_id_full_n,
    input wire                                           krnl_globalSort_L1_L2_0_out_id_write,
    output wire                                          krnl_globalSort_L1_L2_1_ap_clk,
    input wire                                           krnl_globalSort_L1_L2_1_ap_done,
    input wire                                           krnl_globalSort_L1_L2_1_ap_idle,
    input wire                                           krnl_globalSort_L1_L2_1_ap_ready,
    output wire                                          krnl_globalSort_L1_L2_1_ap_rst_n,
    output wire                                          krnl_globalSort_L1_L2_1_ap_start,
    output wire [                                  65:0] krnl_globalSort_L1_L2_1_in_dist0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_1_in_dist0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_1_in_dist0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_1_in_dist0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_1_in_dist0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_1_in_dist0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_1_in_dist1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_1_in_dist1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_1_in_dist1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_1_in_dist1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_1_in_dist1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_1_in_dist1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_1_in_dist2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_1_in_dist2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_1_in_dist2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_1_in_dist2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_1_in_dist2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_1_in_dist2_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_1_in_id0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_1_in_id0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_1_in_id0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_1_in_id0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_1_in_id0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_1_in_id0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_1_in_id1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_1_in_id1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_1_in_id1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_1_in_id1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_1_in_id1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_1_in_id1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_1_in_id2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_1_in_id2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_1_in_id2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_1_in_id2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_1_in_id2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_1_in_id2_s_read,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_1_out_dist_din,
    output wire                                          krnl_globalSort_L1_L2_1_out_dist_full_n,
    input wire                                           krnl_globalSort_L1_L2_1_out_dist_write,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_1_out_id_din,
    output wire                                          krnl_globalSort_L1_L2_1_out_id_full_n,
    input wire                                           krnl_globalSort_L1_L2_1_out_id_write,
    output wire                                          krnl_globalSort_L1_L2_2_ap_clk,
    input wire                                           krnl_globalSort_L1_L2_2_ap_done,
    input wire                                           krnl_globalSort_L1_L2_2_ap_idle,
    input wire                                           krnl_globalSort_L1_L2_2_ap_ready,
    output wire                                          krnl_globalSort_L1_L2_2_ap_rst_n,
    output wire                                          krnl_globalSort_L1_L2_2_ap_start,
    output wire [                                  65:0] krnl_globalSort_L1_L2_2_in_dist0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_2_in_dist0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_2_in_dist0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_2_in_dist0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_2_in_dist0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_2_in_dist0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_2_in_dist1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_2_in_dist1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_2_in_dist1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_2_in_dist1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_2_in_dist1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_2_in_dist1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_2_in_dist2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_2_in_dist2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_2_in_dist2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_2_in_dist2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_2_in_dist2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_2_in_dist2_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_2_in_id0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_2_in_id0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_2_in_id0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_2_in_id0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_2_in_id0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_2_in_id0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_2_in_id1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_2_in_id1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_2_in_id1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_2_in_id1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_2_in_id1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_2_in_id1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_2_in_id2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_2_in_id2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_2_in_id2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_2_in_id2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_2_in_id2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_2_in_id2_s_read,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_2_out_dist_din,
    output wire                                          krnl_globalSort_L1_L2_2_out_dist_full_n,
    input wire                                           krnl_globalSort_L1_L2_2_out_dist_write,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_2_out_id_din,
    output wire                                          krnl_globalSort_L1_L2_2_out_id_full_n,
    input wire                                           krnl_globalSort_L1_L2_2_out_id_write,
    output wire                                          krnl_globalSort_L1_L2_3_ap_clk,
    input wire                                           krnl_globalSort_L1_L2_3_ap_done,
    input wire                                           krnl_globalSort_L1_L2_3_ap_idle,
    input wire                                           krnl_globalSort_L1_L2_3_ap_ready,
    output wire                                          krnl_globalSort_L1_L2_3_ap_rst_n,
    output wire                                          krnl_globalSort_L1_L2_3_ap_start,
    output wire [                                  65:0] krnl_globalSort_L1_L2_3_in_dist0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_3_in_dist0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_3_in_dist0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_3_in_dist0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_3_in_dist0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_3_in_dist0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_3_in_dist1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_3_in_dist1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_3_in_dist1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_3_in_dist1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_3_in_dist1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_3_in_dist1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_3_in_dist2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_3_in_dist2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_3_in_dist2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_3_in_dist2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_3_in_dist2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_3_in_dist2_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_3_in_id0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_3_in_id0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_3_in_id0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_3_in_id0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_3_in_id0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_3_in_id0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_3_in_id1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_3_in_id1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_3_in_id1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_3_in_id1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_3_in_id1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_3_in_id1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_3_in_id2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_3_in_id2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_3_in_id2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_3_in_id2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_3_in_id2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_3_in_id2_s_read,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_3_out_dist_din,
    output wire                                          krnl_globalSort_L1_L2_3_out_dist_full_n,
    input wire                                           krnl_globalSort_L1_L2_3_out_dist_write,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_3_out_id_din,
    output wire                                          krnl_globalSort_L1_L2_3_out_id_full_n,
    input wire                                           krnl_globalSort_L1_L2_3_out_id_write,
    output wire                                          krnl_globalSort_L1_L2_4_ap_clk,
    input wire                                           krnl_globalSort_L1_L2_4_ap_done,
    input wire                                           krnl_globalSort_L1_L2_4_ap_idle,
    input wire                                           krnl_globalSort_L1_L2_4_ap_ready,
    output wire                                          krnl_globalSort_L1_L2_4_ap_rst_n,
    output wire                                          krnl_globalSort_L1_L2_4_ap_start,
    output wire [                                  65:0] krnl_globalSort_L1_L2_4_in_dist0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_4_in_dist0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_4_in_dist0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_4_in_dist0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_4_in_dist0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_4_in_dist0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_4_in_dist1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_4_in_dist1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_4_in_dist1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_4_in_dist1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_4_in_dist1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_4_in_dist1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_4_in_dist2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_4_in_dist2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_4_in_dist2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_4_in_dist2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_4_in_dist2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_4_in_dist2_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_4_in_id0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_4_in_id0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_4_in_id0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_4_in_id0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_4_in_id0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_4_in_id0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_4_in_id1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_4_in_id1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_4_in_id1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_4_in_id1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_4_in_id1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_4_in_id1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_4_in_id2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_4_in_id2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_4_in_id2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_4_in_id2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_4_in_id2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_4_in_id2_s_read,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_4_out_dist_din,
    output wire                                          krnl_globalSort_L1_L2_4_out_dist_full_n,
    input wire                                           krnl_globalSort_L1_L2_4_out_dist_write,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_4_out_id_din,
    output wire                                          krnl_globalSort_L1_L2_4_out_id_full_n,
    input wire                                           krnl_globalSort_L1_L2_4_out_id_write,
    output wire                                          krnl_globalSort_L1_L2_5_ap_clk,
    input wire                                           krnl_globalSort_L1_L2_5_ap_done,
    input wire                                           krnl_globalSort_L1_L2_5_ap_idle,
    input wire                                           krnl_globalSort_L1_L2_5_ap_ready,
    output wire                                          krnl_globalSort_L1_L2_5_ap_rst_n,
    output wire                                          krnl_globalSort_L1_L2_5_ap_start,
    output wire [                                  65:0] krnl_globalSort_L1_L2_5_in_dist0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_5_in_dist0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_5_in_dist0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_5_in_dist0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_5_in_dist0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_5_in_dist0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_5_in_dist1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_5_in_dist1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_5_in_dist1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_5_in_dist1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_5_in_dist1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_5_in_dist1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_5_in_dist2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_5_in_dist2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_5_in_dist2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_5_in_dist2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_5_in_dist2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_5_in_dist2_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_5_in_id0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_5_in_id0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_5_in_id0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_5_in_id0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_5_in_id0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_5_in_id0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_5_in_id1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_5_in_id1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_5_in_id1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_5_in_id1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_5_in_id1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_5_in_id1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_5_in_id2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_5_in_id2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_5_in_id2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_5_in_id2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_5_in_id2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_5_in_id2_s_read,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_5_out_dist_din,
    output wire                                          krnl_globalSort_L1_L2_5_out_dist_full_n,
    input wire                                           krnl_globalSort_L1_L2_5_out_dist_write,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_5_out_id_din,
    output wire                                          krnl_globalSort_L1_L2_5_out_id_full_n,
    input wire                                           krnl_globalSort_L1_L2_5_out_id_write,
    output wire                                          krnl_globalSort_L1_L2_6_ap_clk,
    input wire                                           krnl_globalSort_L1_L2_6_ap_done,
    input wire                                           krnl_globalSort_L1_L2_6_ap_idle,
    input wire                                           krnl_globalSort_L1_L2_6_ap_ready,
    output wire                                          krnl_globalSort_L1_L2_6_ap_rst_n,
    output wire                                          krnl_globalSort_L1_L2_6_ap_start,
    output wire [                                  65:0] krnl_globalSort_L1_L2_6_in_dist0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_6_in_dist0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_6_in_dist0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_6_in_dist0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_6_in_dist0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_6_in_dist0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_6_in_dist1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_6_in_dist1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_6_in_dist1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_6_in_dist1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_6_in_dist1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_6_in_dist1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_6_in_dist2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_6_in_dist2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_6_in_dist2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_6_in_dist2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_6_in_dist2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_6_in_dist2_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_6_in_id0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_6_in_id0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_6_in_id0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_6_in_id0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_6_in_id0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_6_in_id0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_6_in_id1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_6_in_id1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_6_in_id1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_6_in_id1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_6_in_id1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_6_in_id1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_6_in_id2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_6_in_id2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_6_in_id2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_6_in_id2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_6_in_id2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_6_in_id2_s_read,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_6_out_dist_din,
    output wire                                          krnl_globalSort_L1_L2_6_out_dist_full_n,
    input wire                                           krnl_globalSort_L1_L2_6_out_dist_write,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_6_out_id_din,
    output wire                                          krnl_globalSort_L1_L2_6_out_id_full_n,
    input wire                                           krnl_globalSort_L1_L2_6_out_id_write,
    output wire                                          krnl_globalSort_L1_L2_7_ap_clk,
    input wire                                           krnl_globalSort_L1_L2_7_ap_done,
    input wire                                           krnl_globalSort_L1_L2_7_ap_idle,
    input wire                                           krnl_globalSort_L1_L2_7_ap_ready,
    output wire                                          krnl_globalSort_L1_L2_7_ap_rst_n,
    output wire                                          krnl_globalSort_L1_L2_7_ap_start,
    output wire [                                  65:0] krnl_globalSort_L1_L2_7_in_dist0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_7_in_dist0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_7_in_dist0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_7_in_dist0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_7_in_dist0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_7_in_dist0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_7_in_dist1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_7_in_dist1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_7_in_dist1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_7_in_dist1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_7_in_dist1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_7_in_dist1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_7_in_dist2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_7_in_dist2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_7_in_dist2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_7_in_dist2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_7_in_dist2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_7_in_dist2_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_7_in_id0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_7_in_id0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_7_in_id0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_7_in_id0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_7_in_id0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_7_in_id0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_7_in_id1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_7_in_id1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_7_in_id1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_7_in_id1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_7_in_id1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_7_in_id1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_7_in_id2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_7_in_id2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_7_in_id2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_7_in_id2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_7_in_id2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_7_in_id2_s_read,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_7_out_dist_din,
    output wire                                          krnl_globalSort_L1_L2_7_out_dist_full_n,
    input wire                                           krnl_globalSort_L1_L2_7_out_dist_write,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_7_out_id_din,
    output wire                                          krnl_globalSort_L1_L2_7_out_id_full_n,
    input wire                                           krnl_globalSort_L1_L2_7_out_id_write,
    output wire                                          krnl_globalSort_L1_L2_8_ap_clk,
    input wire                                           krnl_globalSort_L1_L2_8_ap_done,
    input wire                                           krnl_globalSort_L1_L2_8_ap_idle,
    input wire                                           krnl_globalSort_L1_L2_8_ap_ready,
    output wire                                          krnl_globalSort_L1_L2_8_ap_rst_n,
    output wire                                          krnl_globalSort_L1_L2_8_ap_start,
    output wire [                                  65:0] krnl_globalSort_L1_L2_8_in_dist0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_8_in_dist0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_8_in_dist0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_8_in_dist0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_8_in_dist0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_8_in_dist0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_8_in_dist1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_8_in_dist1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_8_in_dist1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_8_in_dist1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_8_in_dist1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_8_in_dist1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_8_in_dist2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_8_in_dist2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_8_in_dist2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_8_in_dist2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_8_in_dist2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_8_in_dist2_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_8_in_id0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_8_in_id0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_8_in_id0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_8_in_id0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_8_in_id0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_8_in_id0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_8_in_id1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_8_in_id1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_8_in_id1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_8_in_id1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_8_in_id1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_8_in_id1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_8_in_id2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_8_in_id2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_8_in_id2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_8_in_id2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_8_in_id2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_8_in_id2_s_read,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_8_out_dist_din,
    output wire                                          krnl_globalSort_L1_L2_8_out_dist_full_n,
    input wire                                           krnl_globalSort_L1_L2_8_out_dist_write,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_8_out_id_din,
    output wire                                          krnl_globalSort_L1_L2_8_out_id_full_n,
    input wire                                           krnl_globalSort_L1_L2_8_out_id_write,
    output wire                                          krnl_globalSort_L1_L2_9_ap_clk,
    input wire                                           krnl_globalSort_L1_L2_9_ap_done,
    input wire                                           krnl_globalSort_L1_L2_9_ap_idle,
    input wire                                           krnl_globalSort_L1_L2_9_ap_ready,
    output wire                                          krnl_globalSort_L1_L2_9_ap_rst_n,
    output wire                                          krnl_globalSort_L1_L2_9_ap_start,
    output wire [                                  65:0] krnl_globalSort_L1_L2_9_in_dist0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_9_in_dist0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_9_in_dist0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_9_in_dist0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_9_in_dist0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_9_in_dist0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_9_in_dist1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_9_in_dist1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_9_in_dist1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_9_in_dist1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_9_in_dist1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_9_in_dist1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_9_in_dist2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_9_in_dist2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_9_in_dist2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_9_in_dist2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_9_in_dist2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_9_in_dist2_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_9_in_id0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_9_in_id0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_9_in_id0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_9_in_id0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_9_in_id0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_9_in_id0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_9_in_id1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_9_in_id1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_9_in_id1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_9_in_id1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_9_in_id1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_9_in_id1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_9_in_id2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_9_in_id2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_9_in_id2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_9_in_id2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_9_in_id2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_9_in_id2_s_read,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_9_out_dist_din,
    output wire                                          krnl_globalSort_L1_L2_9_out_dist_full_n,
    input wire                                           krnl_globalSort_L1_L2_9_out_dist_write,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_9_out_id_din,
    output wire                                          krnl_globalSort_L1_L2_9_out_id_full_n,
    input wire                                           krnl_globalSort_L1_L2_9_out_id_write,
    output wire                                          krnl_globalSort_L1_L2_10_ap_clk,
    input wire                                           krnl_globalSort_L1_L2_10_ap_done,
    input wire                                           krnl_globalSort_L1_L2_10_ap_idle,
    input wire                                           krnl_globalSort_L1_L2_10_ap_ready,
    output wire                                          krnl_globalSort_L1_L2_10_ap_rst_n,
    output wire                                          krnl_globalSort_L1_L2_10_ap_start,
    output wire [                                  65:0] krnl_globalSort_L1_L2_10_in_dist0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_10_in_dist0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_10_in_dist0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_10_in_dist0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_10_in_dist0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_10_in_dist0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_10_in_dist1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_10_in_dist1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_10_in_dist1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_10_in_dist1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_10_in_dist1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_10_in_dist1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_10_in_dist2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_10_in_dist2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_10_in_dist2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_10_in_dist2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_10_in_dist2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_10_in_dist2_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_10_in_id0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_10_in_id0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_10_in_id0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_10_in_id0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_10_in_id0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_10_in_id0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_10_in_id1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_10_in_id1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_10_in_id1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_10_in_id1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_10_in_id1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_10_in_id1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_10_in_id2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_10_in_id2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_10_in_id2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_10_in_id2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_10_in_id2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_10_in_id2_s_read,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_10_out_dist_din,
    output wire                                          krnl_globalSort_L1_L2_10_out_dist_full_n,
    input wire                                           krnl_globalSort_L1_L2_10_out_dist_write,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_10_out_id_din,
    output wire                                          krnl_globalSort_L1_L2_10_out_id_full_n,
    input wire                                           krnl_globalSort_L1_L2_10_out_id_write,
    output wire                                          krnl_globalSort_L1_L2_11_ap_clk,
    input wire                                           krnl_globalSort_L1_L2_11_ap_done,
    input wire                                           krnl_globalSort_L1_L2_11_ap_idle,
    input wire                                           krnl_globalSort_L1_L2_11_ap_ready,
    output wire                                          krnl_globalSort_L1_L2_11_ap_rst_n,
    output wire                                          krnl_globalSort_L1_L2_11_ap_start,
    output wire [                                  65:0] krnl_globalSort_L1_L2_11_in_dist0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_11_in_dist0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_11_in_dist0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_11_in_dist0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_11_in_dist0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_11_in_dist0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_11_in_dist1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_11_in_dist1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_11_in_dist1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_11_in_dist1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_11_in_dist1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_11_in_dist1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_11_in_dist2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_11_in_dist2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_11_in_dist2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_11_in_dist2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_11_in_dist2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_11_in_dist2_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_11_in_id0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_11_in_id0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_11_in_id0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_11_in_id0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_11_in_id0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_11_in_id0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_11_in_id1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_11_in_id1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_11_in_id1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_11_in_id1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_11_in_id1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_11_in_id1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_11_in_id2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_11_in_id2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_11_in_id2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_11_in_id2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_11_in_id2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_11_in_id2_s_read,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_11_out_dist_din,
    output wire                                          krnl_globalSort_L1_L2_11_out_dist_full_n,
    input wire                                           krnl_globalSort_L1_L2_11_out_dist_write,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_11_out_id_din,
    output wire                                          krnl_globalSort_L1_L2_11_out_id_full_n,
    input wire                                           krnl_globalSort_L1_L2_11_out_id_write,
    output wire                                          krnl_globalSort_L1_L2_12_ap_clk,
    input wire                                           krnl_globalSort_L1_L2_12_ap_done,
    input wire                                           krnl_globalSort_L1_L2_12_ap_idle,
    input wire                                           krnl_globalSort_L1_L2_12_ap_ready,
    output wire                                          krnl_globalSort_L1_L2_12_ap_rst_n,
    output wire                                          krnl_globalSort_L1_L2_12_ap_start,
    output wire [                                  65:0] krnl_globalSort_L1_L2_12_in_dist0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_12_in_dist0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_12_in_dist0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_12_in_dist0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_12_in_dist0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_12_in_dist0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_12_in_dist1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_12_in_dist1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_12_in_dist1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_12_in_dist1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_12_in_dist1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_12_in_dist1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_12_in_dist2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_12_in_dist2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_12_in_dist2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_12_in_dist2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_12_in_dist2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_12_in_dist2_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_12_in_id0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_12_in_id0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_12_in_id0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_12_in_id0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_12_in_id0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_12_in_id0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_12_in_id1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_12_in_id1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_12_in_id1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_12_in_id1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_12_in_id1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_12_in_id1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_12_in_id2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_12_in_id2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_12_in_id2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_12_in_id2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_12_in_id2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_12_in_id2_s_read,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_12_out_dist_din,
    output wire                                          krnl_globalSort_L1_L2_12_out_dist_full_n,
    input wire                                           krnl_globalSort_L1_L2_12_out_dist_write,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_12_out_id_din,
    output wire                                          krnl_globalSort_L1_L2_12_out_id_full_n,
    input wire                                           krnl_globalSort_L1_L2_12_out_id_write,
    output wire                                          krnl_globalSort_L1_L2_13_ap_clk,
    input wire                                           krnl_globalSort_L1_L2_13_ap_done,
    input wire                                           krnl_globalSort_L1_L2_13_ap_idle,
    input wire                                           krnl_globalSort_L1_L2_13_ap_ready,
    output wire                                          krnl_globalSort_L1_L2_13_ap_rst_n,
    output wire                                          krnl_globalSort_L1_L2_13_ap_start,
    output wire [                                  65:0] krnl_globalSort_L1_L2_13_in_dist0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_13_in_dist0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_13_in_dist0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_13_in_dist0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_13_in_dist0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_13_in_dist0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_13_in_dist1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_13_in_dist1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_13_in_dist1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_13_in_dist1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_13_in_dist1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_13_in_dist1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_13_in_dist2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_13_in_dist2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_13_in_dist2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_13_in_dist2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_13_in_dist2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_13_in_dist2_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_13_in_id0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_13_in_id0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_13_in_id0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_13_in_id0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_13_in_id0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_13_in_id0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_13_in_id1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_13_in_id1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_13_in_id1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_13_in_id1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_13_in_id1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_13_in_id1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_13_in_id2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_13_in_id2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_13_in_id2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_13_in_id2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_13_in_id2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_13_in_id2_s_read,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_13_out_dist_din,
    output wire                                          krnl_globalSort_L1_L2_13_out_dist_full_n,
    input wire                                           krnl_globalSort_L1_L2_13_out_dist_write,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_13_out_id_din,
    output wire                                          krnl_globalSort_L1_L2_13_out_id_full_n,
    input wire                                           krnl_globalSort_L1_L2_13_out_id_write,
    output wire                                          krnl_globalSort_L1_L2_14_ap_clk,
    input wire                                           krnl_globalSort_L1_L2_14_ap_done,
    input wire                                           krnl_globalSort_L1_L2_14_ap_idle,
    input wire                                           krnl_globalSort_L1_L2_14_ap_ready,
    output wire                                          krnl_globalSort_L1_L2_14_ap_rst_n,
    output wire                                          krnl_globalSort_L1_L2_14_ap_start,
    output wire [                                  65:0] krnl_globalSort_L1_L2_14_in_dist0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_14_in_dist0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_14_in_dist0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_14_in_dist0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_14_in_dist0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_14_in_dist0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_14_in_dist1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_14_in_dist1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_14_in_dist1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_14_in_dist1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_14_in_dist1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_14_in_dist1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_14_in_dist2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_14_in_dist2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_14_in_dist2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_14_in_dist2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_14_in_dist2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_14_in_dist2_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_14_in_id0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_14_in_id0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_14_in_id0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_14_in_id0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_14_in_id0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_14_in_id0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_14_in_id1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_14_in_id1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_14_in_id1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_14_in_id1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_14_in_id1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_14_in_id1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_14_in_id2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_14_in_id2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_14_in_id2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_14_in_id2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_14_in_id2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_14_in_id2_s_read,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_14_out_dist_din,
    output wire                                          krnl_globalSort_L1_L2_14_out_dist_full_n,
    input wire                                           krnl_globalSort_L1_L2_14_out_dist_write,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_14_out_id_din,
    output wire                                          krnl_globalSort_L1_L2_14_out_id_full_n,
    input wire                                           krnl_globalSort_L1_L2_14_out_id_write,
    output wire                                          krnl_globalSort_L1_L2_15_ap_clk,
    input wire                                           krnl_globalSort_L1_L2_15_ap_done,
    input wire                                           krnl_globalSort_L1_L2_15_ap_idle,
    input wire                                           krnl_globalSort_L1_L2_15_ap_ready,
    output wire                                          krnl_globalSort_L1_L2_15_ap_rst_n,
    output wire                                          krnl_globalSort_L1_L2_15_ap_start,
    output wire [                                  65:0] krnl_globalSort_L1_L2_15_in_dist0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_15_in_dist0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_15_in_dist0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_15_in_dist0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_15_in_dist0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_15_in_dist0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_15_in_dist1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_15_in_dist1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_15_in_dist1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_15_in_dist1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_15_in_dist1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_15_in_dist1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_15_in_dist2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_15_in_dist2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_15_in_dist2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_15_in_dist2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_15_in_dist2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_15_in_dist2_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_15_in_id0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_15_in_id0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_15_in_id0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_15_in_id0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_15_in_id0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_15_in_id0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_15_in_id1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_15_in_id1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_15_in_id1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_15_in_id1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_15_in_id1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_15_in_id1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_15_in_id2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_15_in_id2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_15_in_id2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_15_in_id2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_15_in_id2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_15_in_id2_s_read,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_15_out_dist_din,
    output wire                                          krnl_globalSort_L1_L2_15_out_dist_full_n,
    input wire                                           krnl_globalSort_L1_L2_15_out_dist_write,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_15_out_id_din,
    output wire                                          krnl_globalSort_L1_L2_15_out_id_full_n,
    input wire                                           krnl_globalSort_L1_L2_15_out_id_write,
    output wire                                          krnl_globalSort_L1_L2_16_ap_clk,
    input wire                                           krnl_globalSort_L1_L2_16_ap_done,
    input wire                                           krnl_globalSort_L1_L2_16_ap_idle,
    input wire                                           krnl_globalSort_L1_L2_16_ap_ready,
    output wire                                          krnl_globalSort_L1_L2_16_ap_rst_n,
    output wire                                          krnl_globalSort_L1_L2_16_ap_start,
    output wire [                                  65:0] krnl_globalSort_L1_L2_16_in_dist0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_16_in_dist0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_16_in_dist0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_16_in_dist0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_16_in_dist0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_16_in_dist0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_16_in_dist1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_16_in_dist1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_16_in_dist1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_16_in_dist1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_16_in_dist1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_16_in_dist1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_16_in_dist2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_16_in_dist2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_16_in_dist2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_16_in_dist2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_16_in_dist2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_16_in_dist2_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_16_in_id0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_16_in_id0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_16_in_id0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_16_in_id0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_16_in_id0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_16_in_id0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_16_in_id1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_16_in_id1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_16_in_id1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_16_in_id1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_16_in_id1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_16_in_id1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_16_in_id2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_16_in_id2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_16_in_id2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_16_in_id2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_16_in_id2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_16_in_id2_s_read,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_16_out_dist_din,
    output wire                                          krnl_globalSort_L1_L2_16_out_dist_full_n,
    input wire                                           krnl_globalSort_L1_L2_16_out_dist_write,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_16_out_id_din,
    output wire                                          krnl_globalSort_L1_L2_16_out_id_full_n,
    input wire                                           krnl_globalSort_L1_L2_16_out_id_write,
    output wire                                          krnl_globalSort_L1_L2_17_ap_clk,
    input wire                                           krnl_globalSort_L1_L2_17_ap_done,
    input wire                                           krnl_globalSort_L1_L2_17_ap_idle,
    input wire                                           krnl_globalSort_L1_L2_17_ap_ready,
    output wire                                          krnl_globalSort_L1_L2_17_ap_rst_n,
    output wire                                          krnl_globalSort_L1_L2_17_ap_start,
    output wire [                                  65:0] krnl_globalSort_L1_L2_17_in_dist0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_17_in_dist0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_17_in_dist0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_17_in_dist0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_17_in_dist0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_17_in_dist0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_17_in_dist1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_17_in_dist1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_17_in_dist1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_17_in_dist1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_17_in_dist1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_17_in_dist1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_17_in_dist2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_17_in_dist2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_17_in_dist2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_17_in_dist2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_17_in_dist2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_17_in_dist2_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_17_in_id0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_17_in_id0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_17_in_id0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_17_in_id0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_17_in_id0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_17_in_id0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_17_in_id1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_17_in_id1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_17_in_id1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_17_in_id1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_17_in_id1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_17_in_id1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_17_in_id2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_17_in_id2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_17_in_id2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_17_in_id2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_17_in_id2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_17_in_id2_s_read,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_17_out_dist_din,
    output wire                                          krnl_globalSort_L1_L2_17_out_dist_full_n,
    input wire                                           krnl_globalSort_L1_L2_17_out_dist_write,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_17_out_id_din,
    output wire                                          krnl_globalSort_L1_L2_17_out_id_full_n,
    input wire                                           krnl_globalSort_L1_L2_17_out_id_write,
    output wire                                          krnl_globalSort_L1_L2_18_ap_clk,
    input wire                                           krnl_globalSort_L1_L2_18_ap_done,
    input wire                                           krnl_globalSort_L1_L2_18_ap_idle,
    input wire                                           krnl_globalSort_L1_L2_18_ap_ready,
    output wire                                          krnl_globalSort_L1_L2_18_ap_rst_n,
    output wire                                          krnl_globalSort_L1_L2_18_ap_start,
    output wire [                                  65:0] krnl_globalSort_L1_L2_18_in_dist0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_18_in_dist0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_18_in_dist0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_18_in_dist0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_18_in_dist0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_18_in_dist0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_18_in_dist1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_18_in_dist1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_18_in_dist1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_18_in_dist1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_18_in_dist1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_18_in_dist1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_18_in_dist2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_18_in_dist2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_18_in_dist2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_18_in_dist2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_18_in_dist2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_18_in_dist2_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_18_in_id0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_18_in_id0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_18_in_id0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_18_in_id0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_18_in_id0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_18_in_id0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_18_in_id1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_18_in_id1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_18_in_id1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_18_in_id1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_18_in_id1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_18_in_id1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_18_in_id2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_18_in_id2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_18_in_id2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_18_in_id2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_18_in_id2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_18_in_id2_s_read,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_18_out_dist_din,
    output wire                                          krnl_globalSort_L1_L2_18_out_dist_full_n,
    input wire                                           krnl_globalSort_L1_L2_18_out_dist_write,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_18_out_id_din,
    output wire                                          krnl_globalSort_L1_L2_18_out_id_full_n,
    input wire                                           krnl_globalSort_L1_L2_18_out_id_write,
    output wire                                          krnl_globalSort_L1_L2_19_ap_clk,
    input wire                                           krnl_globalSort_L1_L2_19_ap_done,
    input wire                                           krnl_globalSort_L1_L2_19_ap_idle,
    input wire                                           krnl_globalSort_L1_L2_19_ap_ready,
    output wire                                          krnl_globalSort_L1_L2_19_ap_rst_n,
    output wire                                          krnl_globalSort_L1_L2_19_ap_start,
    output wire [                                  65:0] krnl_globalSort_L1_L2_19_in_dist0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_19_in_dist0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_19_in_dist0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_19_in_dist0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_19_in_dist0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_19_in_dist0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_19_in_dist1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_19_in_dist1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_19_in_dist1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_19_in_dist1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_19_in_dist1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_19_in_dist1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_19_in_dist2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_19_in_dist2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_19_in_dist2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_19_in_dist2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_19_in_dist2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_19_in_dist2_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_19_in_id0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_19_in_id0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_19_in_id0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_19_in_id0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_19_in_id0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_19_in_id0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_19_in_id1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_19_in_id1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_19_in_id1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_19_in_id1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_19_in_id1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_19_in_id1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_19_in_id2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_19_in_id2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_19_in_id2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_19_in_id2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_19_in_id2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_19_in_id2_s_read,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_19_out_dist_din,
    output wire                                          krnl_globalSort_L1_L2_19_out_dist_full_n,
    input wire                                           krnl_globalSort_L1_L2_19_out_dist_write,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_19_out_id_din,
    output wire                                          krnl_globalSort_L1_L2_19_out_id_full_n,
    input wire                                           krnl_globalSort_L1_L2_19_out_id_write,
    output wire                                          krnl_globalSort_L1_L2_20_ap_clk,
    input wire                                           krnl_globalSort_L1_L2_20_ap_done,
    input wire                                           krnl_globalSort_L1_L2_20_ap_idle,
    input wire                                           krnl_globalSort_L1_L2_20_ap_ready,
    output wire                                          krnl_globalSort_L1_L2_20_ap_rst_n,
    output wire                                          krnl_globalSort_L1_L2_20_ap_start,
    output wire [                                  65:0] krnl_globalSort_L1_L2_20_in_dist0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_20_in_dist0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_20_in_dist0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_20_in_dist0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_20_in_dist0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_20_in_dist0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_20_in_dist1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_20_in_dist1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_20_in_dist1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_20_in_dist1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_20_in_dist1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_20_in_dist1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_20_in_dist2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_20_in_dist2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_20_in_dist2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_20_in_dist2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_20_in_dist2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_20_in_dist2_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_20_in_id0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_20_in_id0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_20_in_id0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_20_in_id0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_20_in_id0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_20_in_id0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_20_in_id1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_20_in_id1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_20_in_id1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_20_in_id1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_20_in_id1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_20_in_id1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_20_in_id2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_20_in_id2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_20_in_id2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_20_in_id2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_20_in_id2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_20_in_id2_s_read,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_20_out_dist_din,
    output wire                                          krnl_globalSort_L1_L2_20_out_dist_full_n,
    input wire                                           krnl_globalSort_L1_L2_20_out_dist_write,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_20_out_id_din,
    output wire                                          krnl_globalSort_L1_L2_20_out_id_full_n,
    input wire                                           krnl_globalSort_L1_L2_20_out_id_write,
    output wire                                          krnl_globalSort_L1_L2_21_ap_clk,
    input wire                                           krnl_globalSort_L1_L2_21_ap_done,
    input wire                                           krnl_globalSort_L1_L2_21_ap_idle,
    input wire                                           krnl_globalSort_L1_L2_21_ap_ready,
    output wire                                          krnl_globalSort_L1_L2_21_ap_rst_n,
    output wire                                          krnl_globalSort_L1_L2_21_ap_start,
    output wire [                                  65:0] krnl_globalSort_L1_L2_21_in_dist0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_21_in_dist0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_21_in_dist0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_21_in_dist0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_21_in_dist0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_21_in_dist0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_21_in_dist1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_21_in_dist1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_21_in_dist1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_21_in_dist1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_21_in_dist1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_21_in_dist1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_21_in_dist2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_21_in_dist2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_21_in_dist2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_21_in_dist2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_21_in_dist2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_21_in_dist2_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_21_in_id0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_21_in_id0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_21_in_id0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_21_in_id0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_21_in_id0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_21_in_id0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_21_in_id1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_21_in_id1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_21_in_id1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_21_in_id1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_21_in_id1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_21_in_id1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_21_in_id2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_21_in_id2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_21_in_id2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_21_in_id2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_21_in_id2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_21_in_id2_s_read,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_21_out_dist_din,
    output wire                                          krnl_globalSort_L1_L2_21_out_dist_full_n,
    input wire                                           krnl_globalSort_L1_L2_21_out_dist_write,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_21_out_id_din,
    output wire                                          krnl_globalSort_L1_L2_21_out_id_full_n,
    input wire                                           krnl_globalSort_L1_L2_21_out_id_write,
    output wire                                          krnl_globalSort_L1_L2_22_ap_clk,
    input wire                                           krnl_globalSort_L1_L2_22_ap_done,
    input wire                                           krnl_globalSort_L1_L2_22_ap_idle,
    input wire                                           krnl_globalSort_L1_L2_22_ap_ready,
    output wire                                          krnl_globalSort_L1_L2_22_ap_rst_n,
    output wire                                          krnl_globalSort_L1_L2_22_ap_start,
    output wire [                                  65:0] krnl_globalSort_L1_L2_22_in_dist0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_22_in_dist0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_22_in_dist0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_22_in_dist0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_22_in_dist0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_22_in_dist0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_22_in_dist1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_22_in_dist1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_22_in_dist1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_22_in_dist1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_22_in_dist1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_22_in_dist1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_22_in_dist2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_22_in_dist2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_22_in_dist2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_22_in_dist2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_22_in_dist2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_22_in_dist2_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_22_in_id0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_22_in_id0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_22_in_id0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_22_in_id0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_22_in_id0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_22_in_id0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_22_in_id1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_22_in_id1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_22_in_id1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_22_in_id1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_22_in_id1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_22_in_id1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_22_in_id2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_22_in_id2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_22_in_id2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_22_in_id2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_22_in_id2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_22_in_id2_s_read,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_22_out_dist_din,
    output wire                                          krnl_globalSort_L1_L2_22_out_dist_full_n,
    input wire                                           krnl_globalSort_L1_L2_22_out_dist_write,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_22_out_id_din,
    output wire                                          krnl_globalSort_L1_L2_22_out_id_full_n,
    input wire                                           krnl_globalSort_L1_L2_22_out_id_write,
    output wire                                          krnl_globalSort_L1_L2_23_ap_clk,
    input wire                                           krnl_globalSort_L1_L2_23_ap_done,
    input wire                                           krnl_globalSort_L1_L2_23_ap_idle,
    input wire                                           krnl_globalSort_L1_L2_23_ap_ready,
    output wire                                          krnl_globalSort_L1_L2_23_ap_rst_n,
    output wire                                          krnl_globalSort_L1_L2_23_ap_start,
    output wire [                                  65:0] krnl_globalSort_L1_L2_23_in_dist0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_23_in_dist0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_23_in_dist0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_23_in_dist0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_23_in_dist0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_23_in_dist0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_23_in_dist1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_23_in_dist1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_23_in_dist1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_23_in_dist1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_23_in_dist1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_23_in_dist1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_23_in_dist2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_23_in_dist2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_23_in_dist2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_23_in_dist2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_23_in_dist2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_23_in_dist2_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_23_in_id0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_23_in_id0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_23_in_id0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_23_in_id0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_23_in_id0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_23_in_id0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_23_in_id1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_23_in_id1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_23_in_id1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_23_in_id1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_23_in_id1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_23_in_id1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_23_in_id2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_23_in_id2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_23_in_id2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_23_in_id2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_23_in_id2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_23_in_id2_s_read,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_23_out_dist_din,
    output wire                                          krnl_globalSort_L1_L2_23_out_dist_full_n,
    input wire                                           krnl_globalSort_L1_L2_23_out_dist_write,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_23_out_id_din,
    output wire                                          krnl_globalSort_L1_L2_23_out_id_full_n,
    input wire                                           krnl_globalSort_L1_L2_23_out_id_write,
    output wire                                          krnl_globalSort_L1_L2_24_ap_clk,
    input wire                                           krnl_globalSort_L1_L2_24_ap_done,
    input wire                                           krnl_globalSort_L1_L2_24_ap_idle,
    input wire                                           krnl_globalSort_L1_L2_24_ap_ready,
    output wire                                          krnl_globalSort_L1_L2_24_ap_rst_n,
    output wire                                          krnl_globalSort_L1_L2_24_ap_start,
    output wire [                                  65:0] krnl_globalSort_L1_L2_24_in_dist0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_24_in_dist0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_24_in_dist0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_24_in_dist0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_24_in_dist0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_24_in_dist0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_24_in_dist1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_24_in_dist1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_24_in_dist1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_24_in_dist1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_24_in_dist1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_24_in_dist1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_24_in_dist2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_24_in_dist2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_24_in_dist2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_24_in_dist2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_24_in_dist2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_24_in_dist2_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_24_in_id0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_24_in_id0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_24_in_id0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_24_in_id0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_24_in_id0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_24_in_id0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_24_in_id1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_24_in_id1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_24_in_id1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_24_in_id1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_24_in_id1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_24_in_id1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_24_in_id2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_24_in_id2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_24_in_id2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_24_in_id2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_24_in_id2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_24_in_id2_s_read,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_24_out_dist_din,
    output wire                                          krnl_globalSort_L1_L2_24_out_dist_full_n,
    input wire                                           krnl_globalSort_L1_L2_24_out_dist_write,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_24_out_id_din,
    output wire                                          krnl_globalSort_L1_L2_24_out_id_full_n,
    input wire                                           krnl_globalSort_L1_L2_24_out_id_write,
    output wire                                          krnl_globalSort_L1_L2_25_ap_clk,
    input wire                                           krnl_globalSort_L1_L2_25_ap_done,
    input wire                                           krnl_globalSort_L1_L2_25_ap_idle,
    input wire                                           krnl_globalSort_L1_L2_25_ap_ready,
    output wire                                          krnl_globalSort_L1_L2_25_ap_rst_n,
    output wire                                          krnl_globalSort_L1_L2_25_ap_start,
    output wire [                                  65:0] krnl_globalSort_L1_L2_25_in_dist0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_25_in_dist0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_25_in_dist0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_25_in_dist0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_25_in_dist0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_25_in_dist0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_25_in_dist1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_25_in_dist1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_25_in_dist1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_25_in_dist1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_25_in_dist1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_25_in_dist1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_25_in_dist2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_25_in_dist2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_25_in_dist2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_25_in_dist2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_25_in_dist2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_25_in_dist2_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_25_in_id0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_25_in_id0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_25_in_id0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_25_in_id0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_25_in_id0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_25_in_id0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_25_in_id1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_25_in_id1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_25_in_id1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_25_in_id1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_25_in_id1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_25_in_id1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_25_in_id2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_25_in_id2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_25_in_id2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_25_in_id2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_25_in_id2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_25_in_id2_s_read,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_25_out_dist_din,
    output wire                                          krnl_globalSort_L1_L2_25_out_dist_full_n,
    input wire                                           krnl_globalSort_L1_L2_25_out_dist_write,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_25_out_id_din,
    output wire                                          krnl_globalSort_L1_L2_25_out_id_full_n,
    input wire                                           krnl_globalSort_L1_L2_25_out_id_write,
    output wire                                          krnl_globalSort_L3_0_ap_clk,
    input wire                                           krnl_globalSort_L3_0_ap_done,
    input wire                                           krnl_globalSort_L3_0_ap_idle,
    input wire                                           krnl_globalSort_L3_0_ap_ready,
    output wire                                          krnl_globalSort_L3_0_ap_rst_n,
    output wire                                          krnl_globalSort_L3_0_ap_start,
    output wire [                                  65:0] krnl_globalSort_L3_0_in_dist0_peek_dout,
    output wire                                          krnl_globalSort_L3_0_in_dist0_peek_empty_n,
    input wire                                           krnl_globalSort_L3_0_in_dist0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L3_0_in_dist0_s_dout,
    output wire                                          krnl_globalSort_L3_0_in_dist0_s_empty_n,
    input wire                                           krnl_globalSort_L3_0_in_dist0_s_read,
    output wire [                                  65:0] krnl_globalSort_L3_0_in_dist1_peek_dout,
    output wire                                          krnl_globalSort_L3_0_in_dist1_peek_empty_n,
    input wire                                           krnl_globalSort_L3_0_in_dist1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L3_0_in_dist1_s_dout,
    output wire                                          krnl_globalSort_L3_0_in_dist1_s_empty_n,
    input wire                                           krnl_globalSort_L3_0_in_dist1_s_read,
    output wire [                                  65:0] krnl_globalSort_L3_0_in_id0_peek_dout,
    output wire                                          krnl_globalSort_L3_0_in_id0_peek_empty_n,
    input wire                                           krnl_globalSort_L3_0_in_id0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L3_0_in_id0_s_dout,
    output wire                                          krnl_globalSort_L3_0_in_id0_s_empty_n,
    input wire                                           krnl_globalSort_L3_0_in_id0_s_read,
    output wire [                                  65:0] krnl_globalSort_L3_0_in_id1_peek_dout,
    output wire                                          krnl_globalSort_L3_0_in_id1_peek_empty_n,
    input wire                                           krnl_globalSort_L3_0_in_id1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L3_0_in_id1_s_dout,
    output wire                                          krnl_globalSort_L3_0_in_id1_s_empty_n,
    input wire                                           krnl_globalSort_L3_0_in_id1_s_read,
    output wire [                                  63:0] krnl_globalSort_L3_0_output_knnDist_read_addr_offset,
    input wire  [                                  63:0] krnl_globalSort_L3_0_output_knnDist_read_addr_s_din,
    output wire                                          krnl_globalSort_L3_0_output_knnDist_read_addr_s_full_n,
    input wire                                           krnl_globalSort_L3_0_output_knnDist_read_addr_s_write,
    output wire [                                  32:0] krnl_globalSort_L3_0_output_knnDist_read_data_peek_dout,
    output wire                                          krnl_globalSort_L3_0_output_knnDist_read_data_peek_empty_n,
    input wire                                           krnl_globalSort_L3_0_output_knnDist_read_data_peek_read,
    output wire [                                  32:0] krnl_globalSort_L3_0_output_knnDist_read_data_s_dout,
    output wire                                          krnl_globalSort_L3_0_output_knnDist_read_data_s_empty_n,
    input wire                                           krnl_globalSort_L3_0_output_knnDist_read_data_s_read,
    output wire [                                  63:0] krnl_globalSort_L3_0_output_knnDist_write_addr_offset,
    input wire  [                                  63:0] krnl_globalSort_L3_0_output_knnDist_write_addr_s_din,
    output wire                                          krnl_globalSort_L3_0_output_knnDist_write_addr_s_full_n,
    input wire                                           krnl_globalSort_L3_0_output_knnDist_write_addr_s_write,
    input wire  [                                  32:0] krnl_globalSort_L3_0_output_knnDist_write_data_din,
    output wire                                          krnl_globalSort_L3_0_output_knnDist_write_data_full_n,
    input wire                                           krnl_globalSort_L3_0_output_knnDist_write_data_write,
    output wire [                                   8:0] krnl_globalSort_L3_0_output_knnDist_write_resp_peek_dout,
    output wire                                          krnl_globalSort_L3_0_output_knnDist_write_resp_peek_empty_n,
    input wire                                           krnl_globalSort_L3_0_output_knnDist_write_resp_peek_read,
    output wire [                                   8:0] krnl_globalSort_L3_0_output_knnDist_write_resp_s_dout,
    output wire                                          krnl_globalSort_L3_0_output_knnDist_write_resp_s_empty_n,
    input wire                                           krnl_globalSort_L3_0_output_knnDist_write_resp_s_read,
    output wire [                                  63:0] krnl_globalSort_L3_0_output_knnId_read_addr_offset,
    input wire  [                                  63:0] krnl_globalSort_L3_0_output_knnId_read_addr_s_din,
    output wire                                          krnl_globalSort_L3_0_output_knnId_read_addr_s_full_n,
    input wire                                           krnl_globalSort_L3_0_output_knnId_read_addr_s_write,
    output wire [                                  32:0] krnl_globalSort_L3_0_output_knnId_read_data_peek_dout,
    output wire                                          krnl_globalSort_L3_0_output_knnId_read_data_peek_empty_n,
    input wire                                           krnl_globalSort_L3_0_output_knnId_read_data_peek_read,
    output wire [                                  32:0] krnl_globalSort_L3_0_output_knnId_read_data_s_dout,
    output wire                                          krnl_globalSort_L3_0_output_knnId_read_data_s_empty_n,
    input wire                                           krnl_globalSort_L3_0_output_knnId_read_data_s_read,
    output wire [                                  63:0] krnl_globalSort_L3_0_output_knnId_write_addr_offset,
    input wire  [                                  63:0] krnl_globalSort_L3_0_output_knnId_write_addr_s_din,
    output wire                                          krnl_globalSort_L3_0_output_knnId_write_addr_s_full_n,
    input wire                                           krnl_globalSort_L3_0_output_knnId_write_addr_s_write,
    input wire  [                                  32:0] krnl_globalSort_L3_0_output_knnId_write_data_din,
    output wire                                          krnl_globalSort_L3_0_output_knnId_write_data_full_n,
    input wire                                           krnl_globalSort_L3_0_output_knnId_write_data_write,
    output wire [                                   8:0] krnl_globalSort_L3_0_output_knnId_write_resp_peek_dout,
    output wire                                          krnl_globalSort_L3_0_output_knnId_write_resp_peek_empty_n,
    input wire                                           krnl_globalSort_L3_0_output_knnId_write_resp_peek_read,
    output wire [                                   8:0] krnl_globalSort_L3_0_output_knnId_write_resp_s_dout,
    output wire                                          krnl_globalSort_L3_0_output_knnId_write_resp_s_empty_n,
    input wire                                           krnl_globalSort_L3_0_output_knnId_write_resp_s_read,
    output wire                                          krnl_partialKnn_wrapper_0_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_0_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_0_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_0_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_0_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_0_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_0_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_0_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_0_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_0_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_0_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_0_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_0_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_0_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_0_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_0_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_0_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_0_0_searchSpace_0_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_0_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_0_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_0_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_0_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_0_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_0_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_0_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_0_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_0_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_0_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_0_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_0_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_0_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_0_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_0_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_0_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_0_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_0_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_1_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_1_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_1_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_1_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_1_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_1_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_1_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_1_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_1_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_1_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_1_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_1_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_1_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_1_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_1_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_1_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_1_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_1_0_searchSpace_0_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_1_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_1_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_1_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_1_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_1_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_1_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_1_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_1_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_1_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_1_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_1_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_1_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_1_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_1_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_1_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_1_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_1_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_1_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_10_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_10_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_10_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_10_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_10_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_10_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_10_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_10_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_10_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_10_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_10_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_10_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_10_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_10_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_10_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_10_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_10_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_10_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_10_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_10_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_10_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_10_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_10_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_10_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_10_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_10_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_10_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_10_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_10_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_10_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_10_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_10_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_10_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_10_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_10_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_10_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_11_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_11_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_11_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_11_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_11_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_11_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_11_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_11_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_11_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_11_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_11_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_11_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_11_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_11_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_11_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_11_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_11_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_11_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_11_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_11_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_11_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_11_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_11_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_11_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_11_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_11_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_11_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_11_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_11_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_11_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_11_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_11_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_11_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_11_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_11_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_11_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_12_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_12_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_12_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_12_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_12_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_12_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_12_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_12_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_12_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_12_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_12_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_12_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_12_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_12_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_12_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_12_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_12_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_12_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_12_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_12_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_12_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_12_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_12_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_12_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_12_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_12_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_12_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_12_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_12_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_12_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_12_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_12_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_12_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_12_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_12_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_12_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_13_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_13_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_13_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_13_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_13_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_13_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_13_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_13_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_13_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_13_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_13_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_13_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_13_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_13_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_13_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_13_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_13_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_13_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_13_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_13_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_13_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_13_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_13_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_13_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_13_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_13_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_13_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_13_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_13_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_13_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_13_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_13_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_13_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_13_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_13_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_13_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_14_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_14_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_14_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_14_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_14_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_14_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_14_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_14_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_14_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_14_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_14_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_14_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_14_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_14_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_14_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_14_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_14_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_14_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_14_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_14_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_14_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_14_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_14_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_14_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_14_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_14_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_14_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_14_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_14_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_14_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_14_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_14_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_14_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_14_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_14_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_14_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_15_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_15_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_15_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_15_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_15_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_15_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_15_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_15_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_15_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_15_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_15_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_15_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_15_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_15_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_15_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_15_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_15_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_15_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_15_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_15_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_15_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_15_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_15_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_15_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_15_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_15_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_15_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_15_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_15_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_15_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_15_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_15_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_15_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_15_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_15_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_15_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_16_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_16_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_16_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_16_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_16_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_16_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_16_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_16_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_16_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_16_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_16_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_16_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_16_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_16_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_16_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_16_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_16_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_16_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_16_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_16_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_16_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_16_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_16_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_16_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_16_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_16_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_16_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_16_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_16_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_16_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_16_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_16_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_16_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_16_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_16_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_16_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_17_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_17_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_17_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_17_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_17_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_17_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_17_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_17_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_17_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_17_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_17_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_17_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_17_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_17_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_17_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_17_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_17_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_17_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_17_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_17_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_17_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_17_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_17_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_17_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_17_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_17_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_17_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_17_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_17_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_17_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_17_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_17_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_17_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_17_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_17_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_17_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_18_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_18_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_18_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_18_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_18_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_18_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_18_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_18_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_18_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_18_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_18_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_18_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_18_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_18_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_18_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_18_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_18_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_18_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_18_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_18_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_18_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_18_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_18_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_18_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_18_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_18_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_18_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_18_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_18_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_18_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_18_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_18_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_18_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_18_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_18_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_18_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_19_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_19_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_19_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_19_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_19_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_19_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_19_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_19_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_19_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_19_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_19_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_19_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_19_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_19_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_19_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_19_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_19_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_19_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_19_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_19_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_19_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_19_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_19_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_19_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_19_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_19_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_19_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_19_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_19_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_19_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_19_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_19_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_19_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_19_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_19_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_19_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_2_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_2_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_2_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_2_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_2_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_2_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_2_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_2_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_2_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_2_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_2_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_2_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_2_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_2_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_2_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_2_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_2_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_2_0_searchSpace_0_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_2_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_2_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_2_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_2_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_2_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_2_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_2_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_2_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_2_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_2_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_2_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_2_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_2_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_2_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_2_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_2_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_2_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_2_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_20_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_20_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_20_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_20_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_20_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_20_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_20_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_20_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_20_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_20_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_20_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_20_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_20_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_20_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_20_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_20_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_20_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_20_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_20_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_20_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_20_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_20_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_20_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_20_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_20_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_20_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_20_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_20_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_20_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_20_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_20_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_20_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_20_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_20_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_20_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_20_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_21_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_21_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_21_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_21_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_21_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_21_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_21_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_21_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_21_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_21_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_21_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_21_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_21_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_21_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_21_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_21_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_21_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_21_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_21_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_21_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_21_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_21_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_21_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_21_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_21_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_21_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_21_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_21_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_21_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_21_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_21_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_21_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_21_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_21_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_21_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_21_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_22_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_22_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_22_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_22_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_22_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_22_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_22_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_22_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_22_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_22_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_22_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_22_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_22_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_22_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_22_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_22_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_22_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_22_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_22_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_22_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_22_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_22_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_22_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_22_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_22_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_22_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_22_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_22_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_22_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_22_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_22_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_22_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_22_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_22_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_22_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_22_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_23_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_23_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_23_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_23_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_23_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_23_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_23_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_23_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_23_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_23_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_23_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_23_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_23_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_23_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_23_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_23_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_23_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_23_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_23_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_23_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_23_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_23_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_23_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_23_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_23_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_23_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_23_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_23_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_23_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_23_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_23_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_23_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_23_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_23_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_23_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_23_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_24_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_24_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_24_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_24_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_24_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_24_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_24_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_24_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_24_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_24_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_24_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_24_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_24_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_24_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_24_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_24_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_24_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_24_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_24_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_24_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_24_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_24_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_24_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_24_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_24_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_24_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_24_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_24_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_24_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_24_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_24_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_24_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_24_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_24_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_24_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_24_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_25_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_25_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_25_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_25_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_25_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_25_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_25_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_25_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_25_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_25_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_25_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_25_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_25_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_25_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_25_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_25_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_25_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_25_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_25_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_25_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_25_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_25_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_25_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_25_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_25_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_25_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_25_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_25_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_25_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_25_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_25_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_25_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_25_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_25_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_25_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_25_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_26_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_26_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_26_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_26_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_26_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_26_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_26_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_26_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_26_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_26_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_26_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_26_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_26_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_26_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_26_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_26_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_26_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_26_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_26_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_26_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_26_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_26_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_26_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_26_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_26_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_26_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_26_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_26_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_26_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_26_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_26_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_26_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_26_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_26_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_26_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_26_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_27_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_27_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_27_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_27_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_27_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_27_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_27_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_27_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_27_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_27_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_27_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_27_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_27_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_27_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_27_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_27_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_27_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_27_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_27_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_27_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_27_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_27_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_27_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_27_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_27_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_27_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_27_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_27_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_27_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_27_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_27_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_27_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_27_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_27_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_27_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_27_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_28_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_28_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_28_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_28_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_28_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_28_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_28_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_28_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_28_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_28_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_28_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_28_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_28_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_28_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_28_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_28_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_28_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_28_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_28_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_28_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_28_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_28_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_28_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_28_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_28_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_28_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_28_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_28_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_28_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_28_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_28_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_28_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_28_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_28_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_28_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_28_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_29_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_29_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_29_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_29_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_29_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_29_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_29_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_29_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_29_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_29_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_29_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_29_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_29_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_29_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_29_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_29_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_29_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_29_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_29_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_29_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_29_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_29_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_29_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_29_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_29_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_29_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_29_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_29_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_29_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_29_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_29_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_29_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_29_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_29_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_29_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_29_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_3_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_3_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_3_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_3_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_3_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_3_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_3_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_3_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_3_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_3_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_3_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_3_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_3_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_3_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_3_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_3_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_3_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_3_0_searchSpace_0_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_3_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_3_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_3_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_3_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_3_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_3_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_3_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_3_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_3_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_3_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_3_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_3_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_3_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_3_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_3_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_3_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_3_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_3_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_30_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_30_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_30_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_30_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_30_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_30_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_30_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_30_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_30_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_30_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_30_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_30_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_30_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_30_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_30_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_30_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_30_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_30_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_30_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_30_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_30_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_30_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_30_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_30_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_30_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_30_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_30_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_30_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_30_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_30_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_30_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_30_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_30_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_30_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_30_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_30_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_31_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_31_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_31_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_31_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_31_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_31_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_31_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_31_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_31_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_31_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_31_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_31_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_31_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_31_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_31_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_31_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_31_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_31_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_31_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_31_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_31_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_31_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_31_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_31_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_31_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_31_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_31_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_31_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_31_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_31_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_31_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_31_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_31_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_31_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_31_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_31_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_32_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_32_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_32_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_32_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_32_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_32_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_32_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_32_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_32_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_32_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_32_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_32_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_32_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_32_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_32_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_32_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_32_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_32_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_32_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_32_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_32_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_32_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_32_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_32_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_32_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_32_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_32_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_32_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_32_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_32_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_32_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_32_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_32_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_32_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_32_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_32_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_33_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_33_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_33_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_33_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_33_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_33_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_33_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_33_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_33_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_33_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_33_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_33_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_33_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_33_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_33_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_33_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_33_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_33_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_33_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_33_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_33_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_33_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_33_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_33_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_33_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_33_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_33_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_33_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_33_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_33_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_33_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_33_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_33_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_33_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_33_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_33_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_34_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_34_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_34_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_34_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_34_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_34_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_34_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_34_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_34_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_34_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_34_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_34_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_34_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_34_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_34_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_34_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_34_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_34_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_34_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_34_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_34_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_34_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_34_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_34_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_34_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_34_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_34_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_34_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_34_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_34_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_34_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_34_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_34_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_34_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_34_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_34_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_35_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_35_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_35_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_35_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_35_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_35_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_35_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_35_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_35_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_35_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_35_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_35_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_35_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_35_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_35_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_35_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_35_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_35_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_35_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_35_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_35_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_35_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_35_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_35_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_35_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_35_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_35_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_35_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_35_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_35_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_35_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_35_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_35_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_35_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_35_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_35_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_36_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_36_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_36_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_36_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_36_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_36_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_36_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_36_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_36_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_36_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_36_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_36_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_36_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_36_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_36_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_36_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_36_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_36_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_36_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_36_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_36_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_36_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_36_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_36_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_36_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_36_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_36_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_36_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_36_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_36_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_36_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_36_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_36_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_36_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_36_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_36_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_37_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_37_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_37_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_37_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_37_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_37_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_37_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_37_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_37_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_37_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_37_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_37_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_37_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_37_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_37_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_37_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_37_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_37_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_37_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_37_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_37_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_37_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_37_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_37_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_37_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_37_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_37_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_37_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_37_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_37_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_37_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_37_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_37_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_37_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_37_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_37_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_38_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_38_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_38_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_38_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_38_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_38_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_38_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_38_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_38_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_38_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_38_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_38_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_38_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_38_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_38_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_38_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_38_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_38_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_38_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_38_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_38_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_38_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_38_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_38_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_38_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_38_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_38_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_38_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_38_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_38_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_38_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_38_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_38_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_38_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_38_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_38_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_39_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_39_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_39_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_39_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_39_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_39_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_39_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_39_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_39_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_39_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_39_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_39_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_39_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_39_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_39_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_39_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_39_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_39_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_39_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_39_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_39_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_39_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_39_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_39_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_39_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_39_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_39_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_39_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_39_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_39_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_39_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_39_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_39_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_39_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_39_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_39_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_4_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_4_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_4_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_4_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_4_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_4_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_4_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_4_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_4_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_4_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_4_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_4_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_4_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_4_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_4_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_4_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_4_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_4_0_searchSpace_0_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_4_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_4_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_4_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_4_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_4_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_4_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_4_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_4_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_4_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_4_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_4_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_4_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_4_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_4_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_4_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_4_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_4_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_4_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_40_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_40_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_40_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_40_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_40_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_40_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_40_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_40_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_40_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_40_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_40_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_40_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_40_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_40_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_40_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_40_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_40_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_40_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_40_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_40_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_40_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_40_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_40_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_40_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_40_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_40_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_40_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_40_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_40_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_40_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_40_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_40_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_40_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_40_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_40_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_40_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_41_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_41_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_41_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_41_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_41_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_41_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_41_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_41_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_41_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_41_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_41_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_41_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_41_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_41_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_41_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_41_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_41_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_41_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_41_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_41_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_41_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_41_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_41_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_41_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_41_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_41_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_41_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_41_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_41_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_41_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_41_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_41_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_41_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_41_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_41_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_41_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_42_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_42_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_42_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_42_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_42_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_42_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_42_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_42_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_42_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_42_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_42_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_42_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_42_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_42_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_42_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_42_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_42_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_42_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_42_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_42_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_42_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_42_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_42_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_42_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_42_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_42_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_42_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_42_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_42_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_42_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_42_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_42_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_42_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_42_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_42_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_42_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_43_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_43_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_43_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_43_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_43_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_43_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_43_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_43_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_43_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_43_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_43_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_43_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_43_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_43_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_43_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_43_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_43_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_43_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_43_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_43_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_43_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_43_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_43_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_43_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_43_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_43_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_43_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_43_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_43_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_43_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_43_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_43_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_43_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_43_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_43_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_43_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_44_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_44_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_44_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_44_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_44_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_44_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_44_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_44_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_44_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_44_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_44_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_44_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_44_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_44_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_44_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_44_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_44_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_44_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_44_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_44_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_44_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_44_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_44_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_44_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_44_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_44_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_44_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_44_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_44_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_44_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_44_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_44_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_44_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_44_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_44_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_44_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_45_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_45_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_45_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_45_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_45_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_45_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_45_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_45_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_45_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_45_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_45_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_45_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_45_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_45_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_45_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_45_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_45_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_45_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_45_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_45_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_45_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_45_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_45_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_45_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_45_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_45_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_45_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_45_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_45_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_45_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_45_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_45_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_45_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_45_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_45_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_45_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_46_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_46_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_46_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_46_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_46_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_46_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_46_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_46_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_46_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_46_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_46_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_46_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_46_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_46_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_46_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_46_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_46_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_46_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_46_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_46_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_46_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_46_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_46_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_46_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_46_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_46_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_46_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_46_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_46_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_46_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_46_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_46_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_46_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_46_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_46_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_46_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_47_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_47_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_47_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_47_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_47_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_47_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_47_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_47_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_47_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_47_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_47_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_47_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_47_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_47_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_47_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_47_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_47_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_47_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_47_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_47_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_47_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_47_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_47_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_47_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_47_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_47_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_47_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_47_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_47_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_47_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_47_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_47_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_47_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_47_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_47_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_47_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_48_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_48_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_48_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_48_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_48_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_48_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_48_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_48_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_48_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_48_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_48_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_48_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_48_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_48_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_48_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_48_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_48_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_48_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_48_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_48_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_48_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_48_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_48_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_48_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_48_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_48_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_48_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_48_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_48_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_48_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_48_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_48_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_48_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_48_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_48_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_48_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_49_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_49_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_49_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_49_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_49_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_49_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_49_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_49_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_49_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_49_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_49_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_49_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_49_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_49_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_49_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_49_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_49_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_49_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_49_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_49_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_49_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_49_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_49_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_49_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_49_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_49_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_49_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_49_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_49_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_49_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_49_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_49_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_49_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_49_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_49_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_49_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_5_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_5_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_5_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_5_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_5_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_5_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_5_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_5_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_5_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_5_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_5_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_5_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_5_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_5_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_5_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_5_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_5_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_5_0_searchSpace_0_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_5_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_5_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_5_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_5_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_5_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_5_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_5_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_5_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_5_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_5_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_5_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_5_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_5_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_5_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_5_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_5_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_5_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_5_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_50_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_50_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_50_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_50_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_50_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_50_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_50_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_50_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_50_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_50_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_50_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_50_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_50_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_50_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_50_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_50_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_50_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_50_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_50_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_50_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_50_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_50_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_50_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_50_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_50_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_50_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_50_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_50_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_50_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_50_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_50_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_50_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_50_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_50_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_50_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_50_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_51_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_51_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_51_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_51_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_51_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_51_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_51_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_51_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_51_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_51_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_51_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_51_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_51_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_51_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_51_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_51_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_51_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_51_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_51_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_51_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_51_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_51_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_51_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_51_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_51_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_51_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_51_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_51_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_51_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_51_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_51_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_51_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_51_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_51_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_51_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_51_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_52_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_52_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_52_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_52_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_52_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_52_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_52_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_52_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_52_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_52_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_52_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_52_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_52_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_52_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_52_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_52_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_52_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_52_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_52_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_52_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_52_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_52_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_52_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_52_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_52_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_52_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_52_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_52_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_52_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_52_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_52_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_52_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_52_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_52_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_52_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_52_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_53_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_53_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_53_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_53_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_53_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_53_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_53_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_53_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_53_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_53_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_53_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_53_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_53_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_53_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_53_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_53_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_53_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_53_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_53_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_53_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_53_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_53_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_53_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_53_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_53_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_53_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_53_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_53_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_53_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_53_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_53_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_53_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_53_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_53_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_53_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_53_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_6_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_6_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_6_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_6_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_6_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_6_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_6_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_6_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_6_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_6_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_6_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_6_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_6_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_6_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_6_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_6_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_6_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_6_0_searchSpace_0_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_6_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_6_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_6_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_6_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_6_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_6_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_6_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_6_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_6_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_6_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_6_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_6_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_6_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_6_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_6_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_6_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_6_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_6_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_7_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_7_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_7_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_7_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_7_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_7_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_7_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_7_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_7_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_7_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_7_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_7_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_7_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_7_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_7_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_7_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_7_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_7_0_searchSpace_0_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_7_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_7_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_7_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_7_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_7_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_7_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_7_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_7_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_7_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_7_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_7_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_7_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_7_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_7_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_7_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_7_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_7_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_7_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_8_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_8_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_8_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_8_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_8_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_8_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_8_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_8_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_8_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_8_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_8_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_8_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_8_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_8_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_8_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_8_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_8_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_8_0_searchSpace_0_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_8_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_8_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_8_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_8_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_8_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_8_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_8_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_8_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_8_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_8_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_8_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_8_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_8_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_8_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_8_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_8_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_8_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_8_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_9_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_9_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_9_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_9_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_9_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_9_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_9_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_9_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_9_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_9_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_9_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_9_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_9_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_9_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_9_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_9_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_9_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_9_0_searchSpace_0_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_9_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_9_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_9_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_9_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_9_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_9_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_9_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_9_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_9_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_9_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_9_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_9_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_9_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_9_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_9_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_9_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_9_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_9_0_start_id_0,
    output wire                                          L4_out_dist__m_axi_clk,
    input wire  [                                  63:0] L4_out_dist__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] L4_out_dist__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] L4_out_dist__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] L4_out_dist__m_axi_m_axi_ARID,
    input wire  [                                   7:0] L4_out_dist__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] L4_out_dist__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] L4_out_dist__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] L4_out_dist__m_axi_m_axi_ARQOS,
    output wire                                          L4_out_dist__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] L4_out_dist__m_axi_m_axi_ARSIZE,
    input wire                                           L4_out_dist__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] L4_out_dist__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] L4_out_dist__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] L4_out_dist__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] L4_out_dist__m_axi_m_axi_AWID,
    input wire  [                                   7:0] L4_out_dist__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] L4_out_dist__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] L4_out_dist__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] L4_out_dist__m_axi_m_axi_AWQOS,
    output wire                                          L4_out_dist__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] L4_out_dist__m_axi_m_axi_AWSIZE,
    input wire                                           L4_out_dist__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] L4_out_dist__m_axi_m_axi_BID,
    input wire                                           L4_out_dist__m_axi_m_axi_BREADY,
    output wire [                                   1:0] L4_out_dist__m_axi_m_axi_BRESP,
    output wire                                          L4_out_dist__m_axi_m_axi_BVALID,
    output wire [                                  31:0] L4_out_dist__m_axi_m_axi_RDATA,
    output wire [                                   0:0] L4_out_dist__m_axi_m_axi_RID,
    output wire                                          L4_out_dist__m_axi_m_axi_RLAST,
    input wire                                           L4_out_dist__m_axi_m_axi_RREADY,
    output wire [                                   1:0] L4_out_dist__m_axi_m_axi_RRESP,
    output wire                                          L4_out_dist__m_axi_m_axi_RVALID,
    input wire  [                                  31:0] L4_out_dist__m_axi_m_axi_WDATA,
    input wire                                           L4_out_dist__m_axi_m_axi_WLAST,
    output wire                                          L4_out_dist__m_axi_m_axi_WREADY,
    input wire  [                                   3:0] L4_out_dist__m_axi_m_axi_WSTRB,
    input wire                                           L4_out_dist__m_axi_m_axi_WVALID,
    output wire [                                  63:0] L4_out_dist__m_axi_read_addr_din,
    input wire                                           L4_out_dist__m_axi_read_addr_full_n,
    output wire                                          L4_out_dist__m_axi_read_addr_write,
    input wire  [                                  31:0] L4_out_dist__m_axi_read_data_dout,
    input wire                                           L4_out_dist__m_axi_read_data_empty_n,
    output wire                                          L4_out_dist__m_axi_read_data_read,
    output wire                                          L4_out_dist__m_axi_rst,
    output wire [                                  63:0] L4_out_dist__m_axi_write_addr_din,
    input wire                                           L4_out_dist__m_axi_write_addr_full_n,
    output wire                                          L4_out_dist__m_axi_write_addr_write,
    output wire [                                  31:0] L4_out_dist__m_axi_write_data_din,
    input wire                                           L4_out_dist__m_axi_write_data_full_n,
    output wire                                          L4_out_dist__m_axi_write_data_write,
    input wire  [                                   7:0] L4_out_dist__m_axi_write_resp_dout,
    input wire                                           L4_out_dist__m_axi_write_resp_empty_n,
    output wire                                          L4_out_dist__m_axi_write_resp_read,
    output wire                                          L4_out_id__m_axi_clk,
    input wire  [                                  63:0] L4_out_id__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] L4_out_id__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] L4_out_id__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] L4_out_id__m_axi_m_axi_ARID,
    input wire  [                                   7:0] L4_out_id__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] L4_out_id__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] L4_out_id__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] L4_out_id__m_axi_m_axi_ARQOS,
    output wire                                          L4_out_id__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] L4_out_id__m_axi_m_axi_ARSIZE,
    input wire                                           L4_out_id__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] L4_out_id__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] L4_out_id__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] L4_out_id__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] L4_out_id__m_axi_m_axi_AWID,
    input wire  [                                   7:0] L4_out_id__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] L4_out_id__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] L4_out_id__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] L4_out_id__m_axi_m_axi_AWQOS,
    output wire                                          L4_out_id__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] L4_out_id__m_axi_m_axi_AWSIZE,
    input wire                                           L4_out_id__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] L4_out_id__m_axi_m_axi_BID,
    input wire                                           L4_out_id__m_axi_m_axi_BREADY,
    output wire [                                   1:0] L4_out_id__m_axi_m_axi_BRESP,
    output wire                                          L4_out_id__m_axi_m_axi_BVALID,
    output wire [                                  31:0] L4_out_id__m_axi_m_axi_RDATA,
    output wire [                                   0:0] L4_out_id__m_axi_m_axi_RID,
    output wire                                          L4_out_id__m_axi_m_axi_RLAST,
    input wire                                           L4_out_id__m_axi_m_axi_RREADY,
    output wire [                                   1:0] L4_out_id__m_axi_m_axi_RRESP,
    output wire                                          L4_out_id__m_axi_m_axi_RVALID,
    input wire  [                                  31:0] L4_out_id__m_axi_m_axi_WDATA,
    input wire                                           L4_out_id__m_axi_m_axi_WLAST,
    output wire                                          L4_out_id__m_axi_m_axi_WREADY,
    input wire  [                                   3:0] L4_out_id__m_axi_m_axi_WSTRB,
    input wire                                           L4_out_id__m_axi_m_axi_WVALID,
    output wire [                                  63:0] L4_out_id__m_axi_read_addr_din,
    input wire                                           L4_out_id__m_axi_read_addr_full_n,
    output wire                                          L4_out_id__m_axi_read_addr_write,
    input wire  [                                  31:0] L4_out_id__m_axi_read_data_dout,
    input wire                                           L4_out_id__m_axi_read_data_empty_n,
    output wire                                          L4_out_id__m_axi_read_data_read,
    output wire                                          L4_out_id__m_axi_rst,
    output wire [                                  63:0] L4_out_id__m_axi_write_addr_din,
    input wire                                           L4_out_id__m_axi_write_addr_full_n,
    output wire                                          L4_out_id__m_axi_write_addr_write,
    output wire [                                  31:0] L4_out_id__m_axi_write_data_din,
    input wire                                           L4_out_id__m_axi_write_data_full_n,
    output wire                                          L4_out_id__m_axi_write_data_write,
    input wire  [                                   7:0] L4_out_id__m_axi_write_resp_dout,
    input wire                                           L4_out_id__m_axi_write_resp_empty_n,
    output wire                                          L4_out_id__m_axi_write_resp_read,
    output wire                                          in_0__m_axi_clk,
    input wire  [                                  63:0] in_0__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_0__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_0__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_0__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_0__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_0__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_0__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_0__m_axi_m_axi_ARQOS,
    output wire                                          in_0__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_0__m_axi_m_axi_ARSIZE,
    input wire                                           in_0__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_0__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_0__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_0__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_0__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_0__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_0__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_0__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_0__m_axi_m_axi_AWQOS,
    output wire                                          in_0__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_0__m_axi_m_axi_AWSIZE,
    input wire                                           in_0__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_0__m_axi_m_axi_BID,
    input wire                                           in_0__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_0__m_axi_m_axi_BRESP,
    output wire                                          in_0__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_0__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_0__m_axi_m_axi_RID,
    output wire                                          in_0__m_axi_m_axi_RLAST,
    input wire                                           in_0__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_0__m_axi_m_axi_RRESP,
    output wire                                          in_0__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_0__m_axi_m_axi_WDATA,
    input wire                                           in_0__m_axi_m_axi_WLAST,
    output wire                                          in_0__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_0__m_axi_m_axi_WSTRB,
    input wire                                           in_0__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_0__m_axi_read_addr_din,
    input wire                                           in_0__m_axi_read_addr_full_n,
    output wire                                          in_0__m_axi_read_addr_write,
    input wire  [                                 255:0] in_0__m_axi_read_data_dout,
    input wire                                           in_0__m_axi_read_data_empty_n,
    output wire                                          in_0__m_axi_read_data_read,
    output wire                                          in_0__m_axi_rst,
    output wire [                                  63:0] in_0__m_axi_write_addr_din,
    input wire                                           in_0__m_axi_write_addr_full_n,
    output wire                                          in_0__m_axi_write_addr_write,
    output wire [                                 255:0] in_0__m_axi_write_data_din,
    input wire                                           in_0__m_axi_write_data_full_n,
    output wire                                          in_0__m_axi_write_data_write,
    input wire  [                                   7:0] in_0__m_axi_write_resp_dout,
    input wire                                           in_0__m_axi_write_resp_empty_n,
    output wire                                          in_0__m_axi_write_resp_read,
    output wire                                          in_1__m_axi_clk,
    input wire  [                                  63:0] in_1__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_1__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_1__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_1__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_1__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_1__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_1__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_1__m_axi_m_axi_ARQOS,
    output wire                                          in_1__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_1__m_axi_m_axi_ARSIZE,
    input wire                                           in_1__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_1__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_1__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_1__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_1__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_1__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_1__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_1__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_1__m_axi_m_axi_AWQOS,
    output wire                                          in_1__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_1__m_axi_m_axi_AWSIZE,
    input wire                                           in_1__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_1__m_axi_m_axi_BID,
    input wire                                           in_1__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_1__m_axi_m_axi_BRESP,
    output wire                                          in_1__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_1__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_1__m_axi_m_axi_RID,
    output wire                                          in_1__m_axi_m_axi_RLAST,
    input wire                                           in_1__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_1__m_axi_m_axi_RRESP,
    output wire                                          in_1__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_1__m_axi_m_axi_WDATA,
    input wire                                           in_1__m_axi_m_axi_WLAST,
    output wire                                          in_1__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_1__m_axi_m_axi_WSTRB,
    input wire                                           in_1__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_1__m_axi_read_addr_din,
    input wire                                           in_1__m_axi_read_addr_full_n,
    output wire                                          in_1__m_axi_read_addr_write,
    input wire  [                                 255:0] in_1__m_axi_read_data_dout,
    input wire                                           in_1__m_axi_read_data_empty_n,
    output wire                                          in_1__m_axi_read_data_read,
    output wire                                          in_1__m_axi_rst,
    output wire [                                  63:0] in_1__m_axi_write_addr_din,
    input wire                                           in_1__m_axi_write_addr_full_n,
    output wire                                          in_1__m_axi_write_addr_write,
    output wire [                                 255:0] in_1__m_axi_write_data_din,
    input wire                                           in_1__m_axi_write_data_full_n,
    output wire                                          in_1__m_axi_write_data_write,
    input wire  [                                   7:0] in_1__m_axi_write_resp_dout,
    input wire                                           in_1__m_axi_write_resp_empty_n,
    output wire                                          in_1__m_axi_write_resp_read,
    output wire                                          in_10__m_axi_clk,
    input wire  [                                  63:0] in_10__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_10__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_10__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_10__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_10__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_10__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_10__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_10__m_axi_m_axi_ARQOS,
    output wire                                          in_10__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_10__m_axi_m_axi_ARSIZE,
    input wire                                           in_10__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_10__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_10__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_10__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_10__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_10__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_10__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_10__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_10__m_axi_m_axi_AWQOS,
    output wire                                          in_10__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_10__m_axi_m_axi_AWSIZE,
    input wire                                           in_10__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_10__m_axi_m_axi_BID,
    input wire                                           in_10__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_10__m_axi_m_axi_BRESP,
    output wire                                          in_10__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_10__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_10__m_axi_m_axi_RID,
    output wire                                          in_10__m_axi_m_axi_RLAST,
    input wire                                           in_10__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_10__m_axi_m_axi_RRESP,
    output wire                                          in_10__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_10__m_axi_m_axi_WDATA,
    input wire                                           in_10__m_axi_m_axi_WLAST,
    output wire                                          in_10__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_10__m_axi_m_axi_WSTRB,
    input wire                                           in_10__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_10__m_axi_read_addr_din,
    input wire                                           in_10__m_axi_read_addr_full_n,
    output wire                                          in_10__m_axi_read_addr_write,
    input wire  [                                 255:0] in_10__m_axi_read_data_dout,
    input wire                                           in_10__m_axi_read_data_empty_n,
    output wire                                          in_10__m_axi_read_data_read,
    output wire                                          in_10__m_axi_rst,
    output wire [                                  63:0] in_10__m_axi_write_addr_din,
    input wire                                           in_10__m_axi_write_addr_full_n,
    output wire                                          in_10__m_axi_write_addr_write,
    output wire [                                 255:0] in_10__m_axi_write_data_din,
    input wire                                           in_10__m_axi_write_data_full_n,
    output wire                                          in_10__m_axi_write_data_write,
    input wire  [                                   7:0] in_10__m_axi_write_resp_dout,
    input wire                                           in_10__m_axi_write_resp_empty_n,
    output wire                                          in_10__m_axi_write_resp_read,
    output wire                                          in_11__m_axi_clk,
    input wire  [                                  63:0] in_11__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_11__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_11__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_11__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_11__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_11__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_11__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_11__m_axi_m_axi_ARQOS,
    output wire                                          in_11__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_11__m_axi_m_axi_ARSIZE,
    input wire                                           in_11__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_11__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_11__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_11__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_11__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_11__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_11__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_11__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_11__m_axi_m_axi_AWQOS,
    output wire                                          in_11__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_11__m_axi_m_axi_AWSIZE,
    input wire                                           in_11__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_11__m_axi_m_axi_BID,
    input wire                                           in_11__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_11__m_axi_m_axi_BRESP,
    output wire                                          in_11__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_11__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_11__m_axi_m_axi_RID,
    output wire                                          in_11__m_axi_m_axi_RLAST,
    input wire                                           in_11__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_11__m_axi_m_axi_RRESP,
    output wire                                          in_11__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_11__m_axi_m_axi_WDATA,
    input wire                                           in_11__m_axi_m_axi_WLAST,
    output wire                                          in_11__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_11__m_axi_m_axi_WSTRB,
    input wire                                           in_11__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_11__m_axi_read_addr_din,
    input wire                                           in_11__m_axi_read_addr_full_n,
    output wire                                          in_11__m_axi_read_addr_write,
    input wire  [                                 255:0] in_11__m_axi_read_data_dout,
    input wire                                           in_11__m_axi_read_data_empty_n,
    output wire                                          in_11__m_axi_read_data_read,
    output wire                                          in_11__m_axi_rst,
    output wire [                                  63:0] in_11__m_axi_write_addr_din,
    input wire                                           in_11__m_axi_write_addr_full_n,
    output wire                                          in_11__m_axi_write_addr_write,
    output wire [                                 255:0] in_11__m_axi_write_data_din,
    input wire                                           in_11__m_axi_write_data_full_n,
    output wire                                          in_11__m_axi_write_data_write,
    input wire  [                                   7:0] in_11__m_axi_write_resp_dout,
    input wire                                           in_11__m_axi_write_resp_empty_n,
    output wire                                          in_11__m_axi_write_resp_read,
    output wire                                          in_12__m_axi_clk,
    input wire  [                                  63:0] in_12__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_12__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_12__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_12__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_12__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_12__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_12__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_12__m_axi_m_axi_ARQOS,
    output wire                                          in_12__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_12__m_axi_m_axi_ARSIZE,
    input wire                                           in_12__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_12__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_12__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_12__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_12__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_12__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_12__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_12__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_12__m_axi_m_axi_AWQOS,
    output wire                                          in_12__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_12__m_axi_m_axi_AWSIZE,
    input wire                                           in_12__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_12__m_axi_m_axi_BID,
    input wire                                           in_12__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_12__m_axi_m_axi_BRESP,
    output wire                                          in_12__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_12__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_12__m_axi_m_axi_RID,
    output wire                                          in_12__m_axi_m_axi_RLAST,
    input wire                                           in_12__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_12__m_axi_m_axi_RRESP,
    output wire                                          in_12__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_12__m_axi_m_axi_WDATA,
    input wire                                           in_12__m_axi_m_axi_WLAST,
    output wire                                          in_12__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_12__m_axi_m_axi_WSTRB,
    input wire                                           in_12__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_12__m_axi_read_addr_din,
    input wire                                           in_12__m_axi_read_addr_full_n,
    output wire                                          in_12__m_axi_read_addr_write,
    input wire  [                                 255:0] in_12__m_axi_read_data_dout,
    input wire                                           in_12__m_axi_read_data_empty_n,
    output wire                                          in_12__m_axi_read_data_read,
    output wire                                          in_12__m_axi_rst,
    output wire [                                  63:0] in_12__m_axi_write_addr_din,
    input wire                                           in_12__m_axi_write_addr_full_n,
    output wire                                          in_12__m_axi_write_addr_write,
    output wire [                                 255:0] in_12__m_axi_write_data_din,
    input wire                                           in_12__m_axi_write_data_full_n,
    output wire                                          in_12__m_axi_write_data_write,
    input wire  [                                   7:0] in_12__m_axi_write_resp_dout,
    input wire                                           in_12__m_axi_write_resp_empty_n,
    output wire                                          in_12__m_axi_write_resp_read,
    output wire                                          in_13__m_axi_clk,
    input wire  [                                  63:0] in_13__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_13__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_13__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_13__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_13__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_13__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_13__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_13__m_axi_m_axi_ARQOS,
    output wire                                          in_13__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_13__m_axi_m_axi_ARSIZE,
    input wire                                           in_13__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_13__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_13__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_13__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_13__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_13__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_13__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_13__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_13__m_axi_m_axi_AWQOS,
    output wire                                          in_13__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_13__m_axi_m_axi_AWSIZE,
    input wire                                           in_13__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_13__m_axi_m_axi_BID,
    input wire                                           in_13__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_13__m_axi_m_axi_BRESP,
    output wire                                          in_13__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_13__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_13__m_axi_m_axi_RID,
    output wire                                          in_13__m_axi_m_axi_RLAST,
    input wire                                           in_13__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_13__m_axi_m_axi_RRESP,
    output wire                                          in_13__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_13__m_axi_m_axi_WDATA,
    input wire                                           in_13__m_axi_m_axi_WLAST,
    output wire                                          in_13__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_13__m_axi_m_axi_WSTRB,
    input wire                                           in_13__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_13__m_axi_read_addr_din,
    input wire                                           in_13__m_axi_read_addr_full_n,
    output wire                                          in_13__m_axi_read_addr_write,
    input wire  [                                 255:0] in_13__m_axi_read_data_dout,
    input wire                                           in_13__m_axi_read_data_empty_n,
    output wire                                          in_13__m_axi_read_data_read,
    output wire                                          in_13__m_axi_rst,
    output wire [                                  63:0] in_13__m_axi_write_addr_din,
    input wire                                           in_13__m_axi_write_addr_full_n,
    output wire                                          in_13__m_axi_write_addr_write,
    output wire [                                 255:0] in_13__m_axi_write_data_din,
    input wire                                           in_13__m_axi_write_data_full_n,
    output wire                                          in_13__m_axi_write_data_write,
    input wire  [                                   7:0] in_13__m_axi_write_resp_dout,
    input wire                                           in_13__m_axi_write_resp_empty_n,
    output wire                                          in_13__m_axi_write_resp_read,
    output wire                                          in_14__m_axi_clk,
    input wire  [                                  63:0] in_14__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_14__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_14__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_14__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_14__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_14__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_14__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_14__m_axi_m_axi_ARQOS,
    output wire                                          in_14__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_14__m_axi_m_axi_ARSIZE,
    input wire                                           in_14__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_14__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_14__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_14__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_14__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_14__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_14__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_14__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_14__m_axi_m_axi_AWQOS,
    output wire                                          in_14__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_14__m_axi_m_axi_AWSIZE,
    input wire                                           in_14__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_14__m_axi_m_axi_BID,
    input wire                                           in_14__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_14__m_axi_m_axi_BRESP,
    output wire                                          in_14__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_14__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_14__m_axi_m_axi_RID,
    output wire                                          in_14__m_axi_m_axi_RLAST,
    input wire                                           in_14__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_14__m_axi_m_axi_RRESP,
    output wire                                          in_14__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_14__m_axi_m_axi_WDATA,
    input wire                                           in_14__m_axi_m_axi_WLAST,
    output wire                                          in_14__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_14__m_axi_m_axi_WSTRB,
    input wire                                           in_14__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_14__m_axi_read_addr_din,
    input wire                                           in_14__m_axi_read_addr_full_n,
    output wire                                          in_14__m_axi_read_addr_write,
    input wire  [                                 255:0] in_14__m_axi_read_data_dout,
    input wire                                           in_14__m_axi_read_data_empty_n,
    output wire                                          in_14__m_axi_read_data_read,
    output wire                                          in_14__m_axi_rst,
    output wire [                                  63:0] in_14__m_axi_write_addr_din,
    input wire                                           in_14__m_axi_write_addr_full_n,
    output wire                                          in_14__m_axi_write_addr_write,
    output wire [                                 255:0] in_14__m_axi_write_data_din,
    input wire                                           in_14__m_axi_write_data_full_n,
    output wire                                          in_14__m_axi_write_data_write,
    input wire  [                                   7:0] in_14__m_axi_write_resp_dout,
    input wire                                           in_14__m_axi_write_resp_empty_n,
    output wire                                          in_14__m_axi_write_resp_read,
    output wire                                          in_15__m_axi_clk,
    input wire  [                                  63:0] in_15__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_15__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_15__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_15__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_15__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_15__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_15__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_15__m_axi_m_axi_ARQOS,
    output wire                                          in_15__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_15__m_axi_m_axi_ARSIZE,
    input wire                                           in_15__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_15__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_15__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_15__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_15__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_15__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_15__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_15__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_15__m_axi_m_axi_AWQOS,
    output wire                                          in_15__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_15__m_axi_m_axi_AWSIZE,
    input wire                                           in_15__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_15__m_axi_m_axi_BID,
    input wire                                           in_15__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_15__m_axi_m_axi_BRESP,
    output wire                                          in_15__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_15__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_15__m_axi_m_axi_RID,
    output wire                                          in_15__m_axi_m_axi_RLAST,
    input wire                                           in_15__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_15__m_axi_m_axi_RRESP,
    output wire                                          in_15__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_15__m_axi_m_axi_WDATA,
    input wire                                           in_15__m_axi_m_axi_WLAST,
    output wire                                          in_15__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_15__m_axi_m_axi_WSTRB,
    input wire                                           in_15__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_15__m_axi_read_addr_din,
    input wire                                           in_15__m_axi_read_addr_full_n,
    output wire                                          in_15__m_axi_read_addr_write,
    input wire  [                                 255:0] in_15__m_axi_read_data_dout,
    input wire                                           in_15__m_axi_read_data_empty_n,
    output wire                                          in_15__m_axi_read_data_read,
    output wire                                          in_15__m_axi_rst,
    output wire [                                  63:0] in_15__m_axi_write_addr_din,
    input wire                                           in_15__m_axi_write_addr_full_n,
    output wire                                          in_15__m_axi_write_addr_write,
    output wire [                                 255:0] in_15__m_axi_write_data_din,
    input wire                                           in_15__m_axi_write_data_full_n,
    output wire                                          in_15__m_axi_write_data_write,
    input wire  [                                   7:0] in_15__m_axi_write_resp_dout,
    input wire                                           in_15__m_axi_write_resp_empty_n,
    output wire                                          in_15__m_axi_write_resp_read,
    output wire                                          in_16__m_axi_clk,
    input wire  [                                  63:0] in_16__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_16__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_16__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_16__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_16__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_16__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_16__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_16__m_axi_m_axi_ARQOS,
    output wire                                          in_16__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_16__m_axi_m_axi_ARSIZE,
    input wire                                           in_16__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_16__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_16__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_16__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_16__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_16__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_16__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_16__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_16__m_axi_m_axi_AWQOS,
    output wire                                          in_16__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_16__m_axi_m_axi_AWSIZE,
    input wire                                           in_16__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_16__m_axi_m_axi_BID,
    input wire                                           in_16__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_16__m_axi_m_axi_BRESP,
    output wire                                          in_16__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_16__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_16__m_axi_m_axi_RID,
    output wire                                          in_16__m_axi_m_axi_RLAST,
    input wire                                           in_16__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_16__m_axi_m_axi_RRESP,
    output wire                                          in_16__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_16__m_axi_m_axi_WDATA,
    input wire                                           in_16__m_axi_m_axi_WLAST,
    output wire                                          in_16__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_16__m_axi_m_axi_WSTRB,
    input wire                                           in_16__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_16__m_axi_read_addr_din,
    input wire                                           in_16__m_axi_read_addr_full_n,
    output wire                                          in_16__m_axi_read_addr_write,
    input wire  [                                 255:0] in_16__m_axi_read_data_dout,
    input wire                                           in_16__m_axi_read_data_empty_n,
    output wire                                          in_16__m_axi_read_data_read,
    output wire                                          in_16__m_axi_rst,
    output wire [                                  63:0] in_16__m_axi_write_addr_din,
    input wire                                           in_16__m_axi_write_addr_full_n,
    output wire                                          in_16__m_axi_write_addr_write,
    output wire [                                 255:0] in_16__m_axi_write_data_din,
    input wire                                           in_16__m_axi_write_data_full_n,
    output wire                                          in_16__m_axi_write_data_write,
    input wire  [                                   7:0] in_16__m_axi_write_resp_dout,
    input wire                                           in_16__m_axi_write_resp_empty_n,
    output wire                                          in_16__m_axi_write_resp_read,
    output wire                                          in_17__m_axi_clk,
    input wire  [                                  63:0] in_17__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_17__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_17__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_17__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_17__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_17__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_17__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_17__m_axi_m_axi_ARQOS,
    output wire                                          in_17__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_17__m_axi_m_axi_ARSIZE,
    input wire                                           in_17__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_17__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_17__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_17__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_17__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_17__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_17__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_17__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_17__m_axi_m_axi_AWQOS,
    output wire                                          in_17__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_17__m_axi_m_axi_AWSIZE,
    input wire                                           in_17__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_17__m_axi_m_axi_BID,
    input wire                                           in_17__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_17__m_axi_m_axi_BRESP,
    output wire                                          in_17__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_17__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_17__m_axi_m_axi_RID,
    output wire                                          in_17__m_axi_m_axi_RLAST,
    input wire                                           in_17__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_17__m_axi_m_axi_RRESP,
    output wire                                          in_17__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_17__m_axi_m_axi_WDATA,
    input wire                                           in_17__m_axi_m_axi_WLAST,
    output wire                                          in_17__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_17__m_axi_m_axi_WSTRB,
    input wire                                           in_17__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_17__m_axi_read_addr_din,
    input wire                                           in_17__m_axi_read_addr_full_n,
    output wire                                          in_17__m_axi_read_addr_write,
    input wire  [                                 255:0] in_17__m_axi_read_data_dout,
    input wire                                           in_17__m_axi_read_data_empty_n,
    output wire                                          in_17__m_axi_read_data_read,
    output wire                                          in_17__m_axi_rst,
    output wire [                                  63:0] in_17__m_axi_write_addr_din,
    input wire                                           in_17__m_axi_write_addr_full_n,
    output wire                                          in_17__m_axi_write_addr_write,
    output wire [                                 255:0] in_17__m_axi_write_data_din,
    input wire                                           in_17__m_axi_write_data_full_n,
    output wire                                          in_17__m_axi_write_data_write,
    input wire  [                                   7:0] in_17__m_axi_write_resp_dout,
    input wire                                           in_17__m_axi_write_resp_empty_n,
    output wire                                          in_17__m_axi_write_resp_read,
    output wire                                          in_18__m_axi_clk,
    input wire  [                                  63:0] in_18__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_18__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_18__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_18__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_18__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_18__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_18__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_18__m_axi_m_axi_ARQOS,
    output wire                                          in_18__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_18__m_axi_m_axi_ARSIZE,
    input wire                                           in_18__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_18__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_18__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_18__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_18__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_18__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_18__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_18__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_18__m_axi_m_axi_AWQOS,
    output wire                                          in_18__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_18__m_axi_m_axi_AWSIZE,
    input wire                                           in_18__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_18__m_axi_m_axi_BID,
    input wire                                           in_18__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_18__m_axi_m_axi_BRESP,
    output wire                                          in_18__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_18__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_18__m_axi_m_axi_RID,
    output wire                                          in_18__m_axi_m_axi_RLAST,
    input wire                                           in_18__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_18__m_axi_m_axi_RRESP,
    output wire                                          in_18__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_18__m_axi_m_axi_WDATA,
    input wire                                           in_18__m_axi_m_axi_WLAST,
    output wire                                          in_18__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_18__m_axi_m_axi_WSTRB,
    input wire                                           in_18__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_18__m_axi_read_addr_din,
    input wire                                           in_18__m_axi_read_addr_full_n,
    output wire                                          in_18__m_axi_read_addr_write,
    input wire  [                                 255:0] in_18__m_axi_read_data_dout,
    input wire                                           in_18__m_axi_read_data_empty_n,
    output wire                                          in_18__m_axi_read_data_read,
    output wire                                          in_18__m_axi_rst,
    output wire [                                  63:0] in_18__m_axi_write_addr_din,
    input wire                                           in_18__m_axi_write_addr_full_n,
    output wire                                          in_18__m_axi_write_addr_write,
    output wire [                                 255:0] in_18__m_axi_write_data_din,
    input wire                                           in_18__m_axi_write_data_full_n,
    output wire                                          in_18__m_axi_write_data_write,
    input wire  [                                   7:0] in_18__m_axi_write_resp_dout,
    input wire                                           in_18__m_axi_write_resp_empty_n,
    output wire                                          in_18__m_axi_write_resp_read,
    output wire                                          in_19__m_axi_clk,
    input wire  [                                  63:0] in_19__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_19__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_19__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_19__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_19__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_19__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_19__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_19__m_axi_m_axi_ARQOS,
    output wire                                          in_19__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_19__m_axi_m_axi_ARSIZE,
    input wire                                           in_19__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_19__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_19__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_19__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_19__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_19__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_19__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_19__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_19__m_axi_m_axi_AWQOS,
    output wire                                          in_19__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_19__m_axi_m_axi_AWSIZE,
    input wire                                           in_19__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_19__m_axi_m_axi_BID,
    input wire                                           in_19__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_19__m_axi_m_axi_BRESP,
    output wire                                          in_19__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_19__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_19__m_axi_m_axi_RID,
    output wire                                          in_19__m_axi_m_axi_RLAST,
    input wire                                           in_19__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_19__m_axi_m_axi_RRESP,
    output wire                                          in_19__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_19__m_axi_m_axi_WDATA,
    input wire                                           in_19__m_axi_m_axi_WLAST,
    output wire                                          in_19__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_19__m_axi_m_axi_WSTRB,
    input wire                                           in_19__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_19__m_axi_read_addr_din,
    input wire                                           in_19__m_axi_read_addr_full_n,
    output wire                                          in_19__m_axi_read_addr_write,
    input wire  [                                 255:0] in_19__m_axi_read_data_dout,
    input wire                                           in_19__m_axi_read_data_empty_n,
    output wire                                          in_19__m_axi_read_data_read,
    output wire                                          in_19__m_axi_rst,
    output wire [                                  63:0] in_19__m_axi_write_addr_din,
    input wire                                           in_19__m_axi_write_addr_full_n,
    output wire                                          in_19__m_axi_write_addr_write,
    output wire [                                 255:0] in_19__m_axi_write_data_din,
    input wire                                           in_19__m_axi_write_data_full_n,
    output wire                                          in_19__m_axi_write_data_write,
    input wire  [                                   7:0] in_19__m_axi_write_resp_dout,
    input wire                                           in_19__m_axi_write_resp_empty_n,
    output wire                                          in_19__m_axi_write_resp_read,
    output wire                                          in_2__m_axi_clk,
    input wire  [                                  63:0] in_2__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_2__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_2__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_2__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_2__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_2__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_2__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_2__m_axi_m_axi_ARQOS,
    output wire                                          in_2__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_2__m_axi_m_axi_ARSIZE,
    input wire                                           in_2__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_2__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_2__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_2__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_2__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_2__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_2__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_2__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_2__m_axi_m_axi_AWQOS,
    output wire                                          in_2__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_2__m_axi_m_axi_AWSIZE,
    input wire                                           in_2__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_2__m_axi_m_axi_BID,
    input wire                                           in_2__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_2__m_axi_m_axi_BRESP,
    output wire                                          in_2__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_2__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_2__m_axi_m_axi_RID,
    output wire                                          in_2__m_axi_m_axi_RLAST,
    input wire                                           in_2__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_2__m_axi_m_axi_RRESP,
    output wire                                          in_2__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_2__m_axi_m_axi_WDATA,
    input wire                                           in_2__m_axi_m_axi_WLAST,
    output wire                                          in_2__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_2__m_axi_m_axi_WSTRB,
    input wire                                           in_2__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_2__m_axi_read_addr_din,
    input wire                                           in_2__m_axi_read_addr_full_n,
    output wire                                          in_2__m_axi_read_addr_write,
    input wire  [                                 255:0] in_2__m_axi_read_data_dout,
    input wire                                           in_2__m_axi_read_data_empty_n,
    output wire                                          in_2__m_axi_read_data_read,
    output wire                                          in_2__m_axi_rst,
    output wire [                                  63:0] in_2__m_axi_write_addr_din,
    input wire                                           in_2__m_axi_write_addr_full_n,
    output wire                                          in_2__m_axi_write_addr_write,
    output wire [                                 255:0] in_2__m_axi_write_data_din,
    input wire                                           in_2__m_axi_write_data_full_n,
    output wire                                          in_2__m_axi_write_data_write,
    input wire  [                                   7:0] in_2__m_axi_write_resp_dout,
    input wire                                           in_2__m_axi_write_resp_empty_n,
    output wire                                          in_2__m_axi_write_resp_read,
    output wire                                          in_20__m_axi_clk,
    input wire  [                                  63:0] in_20__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_20__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_20__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_20__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_20__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_20__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_20__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_20__m_axi_m_axi_ARQOS,
    output wire                                          in_20__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_20__m_axi_m_axi_ARSIZE,
    input wire                                           in_20__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_20__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_20__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_20__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_20__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_20__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_20__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_20__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_20__m_axi_m_axi_AWQOS,
    output wire                                          in_20__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_20__m_axi_m_axi_AWSIZE,
    input wire                                           in_20__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_20__m_axi_m_axi_BID,
    input wire                                           in_20__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_20__m_axi_m_axi_BRESP,
    output wire                                          in_20__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_20__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_20__m_axi_m_axi_RID,
    output wire                                          in_20__m_axi_m_axi_RLAST,
    input wire                                           in_20__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_20__m_axi_m_axi_RRESP,
    output wire                                          in_20__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_20__m_axi_m_axi_WDATA,
    input wire                                           in_20__m_axi_m_axi_WLAST,
    output wire                                          in_20__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_20__m_axi_m_axi_WSTRB,
    input wire                                           in_20__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_20__m_axi_read_addr_din,
    input wire                                           in_20__m_axi_read_addr_full_n,
    output wire                                          in_20__m_axi_read_addr_write,
    input wire  [                                 255:0] in_20__m_axi_read_data_dout,
    input wire                                           in_20__m_axi_read_data_empty_n,
    output wire                                          in_20__m_axi_read_data_read,
    output wire                                          in_20__m_axi_rst,
    output wire [                                  63:0] in_20__m_axi_write_addr_din,
    input wire                                           in_20__m_axi_write_addr_full_n,
    output wire                                          in_20__m_axi_write_addr_write,
    output wire [                                 255:0] in_20__m_axi_write_data_din,
    input wire                                           in_20__m_axi_write_data_full_n,
    output wire                                          in_20__m_axi_write_data_write,
    input wire  [                                   7:0] in_20__m_axi_write_resp_dout,
    input wire                                           in_20__m_axi_write_resp_empty_n,
    output wire                                          in_20__m_axi_write_resp_read,
    output wire                                          in_21__m_axi_clk,
    input wire  [                                  63:0] in_21__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_21__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_21__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_21__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_21__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_21__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_21__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_21__m_axi_m_axi_ARQOS,
    output wire                                          in_21__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_21__m_axi_m_axi_ARSIZE,
    input wire                                           in_21__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_21__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_21__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_21__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_21__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_21__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_21__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_21__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_21__m_axi_m_axi_AWQOS,
    output wire                                          in_21__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_21__m_axi_m_axi_AWSIZE,
    input wire                                           in_21__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_21__m_axi_m_axi_BID,
    input wire                                           in_21__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_21__m_axi_m_axi_BRESP,
    output wire                                          in_21__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_21__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_21__m_axi_m_axi_RID,
    output wire                                          in_21__m_axi_m_axi_RLAST,
    input wire                                           in_21__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_21__m_axi_m_axi_RRESP,
    output wire                                          in_21__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_21__m_axi_m_axi_WDATA,
    input wire                                           in_21__m_axi_m_axi_WLAST,
    output wire                                          in_21__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_21__m_axi_m_axi_WSTRB,
    input wire                                           in_21__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_21__m_axi_read_addr_din,
    input wire                                           in_21__m_axi_read_addr_full_n,
    output wire                                          in_21__m_axi_read_addr_write,
    input wire  [                                 255:0] in_21__m_axi_read_data_dout,
    input wire                                           in_21__m_axi_read_data_empty_n,
    output wire                                          in_21__m_axi_read_data_read,
    output wire                                          in_21__m_axi_rst,
    output wire [                                  63:0] in_21__m_axi_write_addr_din,
    input wire                                           in_21__m_axi_write_addr_full_n,
    output wire                                          in_21__m_axi_write_addr_write,
    output wire [                                 255:0] in_21__m_axi_write_data_din,
    input wire                                           in_21__m_axi_write_data_full_n,
    output wire                                          in_21__m_axi_write_data_write,
    input wire  [                                   7:0] in_21__m_axi_write_resp_dout,
    input wire                                           in_21__m_axi_write_resp_empty_n,
    output wire                                          in_21__m_axi_write_resp_read,
    output wire                                          in_22__m_axi_clk,
    input wire  [                                  63:0] in_22__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_22__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_22__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_22__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_22__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_22__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_22__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_22__m_axi_m_axi_ARQOS,
    output wire                                          in_22__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_22__m_axi_m_axi_ARSIZE,
    input wire                                           in_22__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_22__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_22__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_22__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_22__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_22__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_22__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_22__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_22__m_axi_m_axi_AWQOS,
    output wire                                          in_22__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_22__m_axi_m_axi_AWSIZE,
    input wire                                           in_22__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_22__m_axi_m_axi_BID,
    input wire                                           in_22__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_22__m_axi_m_axi_BRESP,
    output wire                                          in_22__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_22__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_22__m_axi_m_axi_RID,
    output wire                                          in_22__m_axi_m_axi_RLAST,
    input wire                                           in_22__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_22__m_axi_m_axi_RRESP,
    output wire                                          in_22__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_22__m_axi_m_axi_WDATA,
    input wire                                           in_22__m_axi_m_axi_WLAST,
    output wire                                          in_22__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_22__m_axi_m_axi_WSTRB,
    input wire                                           in_22__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_22__m_axi_read_addr_din,
    input wire                                           in_22__m_axi_read_addr_full_n,
    output wire                                          in_22__m_axi_read_addr_write,
    input wire  [                                 255:0] in_22__m_axi_read_data_dout,
    input wire                                           in_22__m_axi_read_data_empty_n,
    output wire                                          in_22__m_axi_read_data_read,
    output wire                                          in_22__m_axi_rst,
    output wire [                                  63:0] in_22__m_axi_write_addr_din,
    input wire                                           in_22__m_axi_write_addr_full_n,
    output wire                                          in_22__m_axi_write_addr_write,
    output wire [                                 255:0] in_22__m_axi_write_data_din,
    input wire                                           in_22__m_axi_write_data_full_n,
    output wire                                          in_22__m_axi_write_data_write,
    input wire  [                                   7:0] in_22__m_axi_write_resp_dout,
    input wire                                           in_22__m_axi_write_resp_empty_n,
    output wire                                          in_22__m_axi_write_resp_read,
    output wire                                          in_23__m_axi_clk,
    input wire  [                                  63:0] in_23__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_23__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_23__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_23__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_23__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_23__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_23__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_23__m_axi_m_axi_ARQOS,
    output wire                                          in_23__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_23__m_axi_m_axi_ARSIZE,
    input wire                                           in_23__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_23__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_23__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_23__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_23__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_23__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_23__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_23__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_23__m_axi_m_axi_AWQOS,
    output wire                                          in_23__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_23__m_axi_m_axi_AWSIZE,
    input wire                                           in_23__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_23__m_axi_m_axi_BID,
    input wire                                           in_23__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_23__m_axi_m_axi_BRESP,
    output wire                                          in_23__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_23__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_23__m_axi_m_axi_RID,
    output wire                                          in_23__m_axi_m_axi_RLAST,
    input wire                                           in_23__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_23__m_axi_m_axi_RRESP,
    output wire                                          in_23__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_23__m_axi_m_axi_WDATA,
    input wire                                           in_23__m_axi_m_axi_WLAST,
    output wire                                          in_23__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_23__m_axi_m_axi_WSTRB,
    input wire                                           in_23__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_23__m_axi_read_addr_din,
    input wire                                           in_23__m_axi_read_addr_full_n,
    output wire                                          in_23__m_axi_read_addr_write,
    input wire  [                                 255:0] in_23__m_axi_read_data_dout,
    input wire                                           in_23__m_axi_read_data_empty_n,
    output wire                                          in_23__m_axi_read_data_read,
    output wire                                          in_23__m_axi_rst,
    output wire [                                  63:0] in_23__m_axi_write_addr_din,
    input wire                                           in_23__m_axi_write_addr_full_n,
    output wire                                          in_23__m_axi_write_addr_write,
    output wire [                                 255:0] in_23__m_axi_write_data_din,
    input wire                                           in_23__m_axi_write_data_full_n,
    output wire                                          in_23__m_axi_write_data_write,
    input wire  [                                   7:0] in_23__m_axi_write_resp_dout,
    input wire                                           in_23__m_axi_write_resp_empty_n,
    output wire                                          in_23__m_axi_write_resp_read,
    output wire                                          in_24__m_axi_clk,
    input wire  [                                  63:0] in_24__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_24__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_24__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_24__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_24__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_24__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_24__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_24__m_axi_m_axi_ARQOS,
    output wire                                          in_24__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_24__m_axi_m_axi_ARSIZE,
    input wire                                           in_24__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_24__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_24__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_24__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_24__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_24__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_24__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_24__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_24__m_axi_m_axi_AWQOS,
    output wire                                          in_24__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_24__m_axi_m_axi_AWSIZE,
    input wire                                           in_24__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_24__m_axi_m_axi_BID,
    input wire                                           in_24__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_24__m_axi_m_axi_BRESP,
    output wire                                          in_24__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_24__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_24__m_axi_m_axi_RID,
    output wire                                          in_24__m_axi_m_axi_RLAST,
    input wire                                           in_24__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_24__m_axi_m_axi_RRESP,
    output wire                                          in_24__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_24__m_axi_m_axi_WDATA,
    input wire                                           in_24__m_axi_m_axi_WLAST,
    output wire                                          in_24__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_24__m_axi_m_axi_WSTRB,
    input wire                                           in_24__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_24__m_axi_read_addr_din,
    input wire                                           in_24__m_axi_read_addr_full_n,
    output wire                                          in_24__m_axi_read_addr_write,
    input wire  [                                 255:0] in_24__m_axi_read_data_dout,
    input wire                                           in_24__m_axi_read_data_empty_n,
    output wire                                          in_24__m_axi_read_data_read,
    output wire                                          in_24__m_axi_rst,
    output wire [                                  63:0] in_24__m_axi_write_addr_din,
    input wire                                           in_24__m_axi_write_addr_full_n,
    output wire                                          in_24__m_axi_write_addr_write,
    output wire [                                 255:0] in_24__m_axi_write_data_din,
    input wire                                           in_24__m_axi_write_data_full_n,
    output wire                                          in_24__m_axi_write_data_write,
    input wire  [                                   7:0] in_24__m_axi_write_resp_dout,
    input wire                                           in_24__m_axi_write_resp_empty_n,
    output wire                                          in_24__m_axi_write_resp_read,
    output wire                                          in_25__m_axi_clk,
    input wire  [                                  63:0] in_25__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_25__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_25__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_25__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_25__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_25__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_25__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_25__m_axi_m_axi_ARQOS,
    output wire                                          in_25__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_25__m_axi_m_axi_ARSIZE,
    input wire                                           in_25__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_25__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_25__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_25__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_25__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_25__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_25__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_25__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_25__m_axi_m_axi_AWQOS,
    output wire                                          in_25__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_25__m_axi_m_axi_AWSIZE,
    input wire                                           in_25__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_25__m_axi_m_axi_BID,
    input wire                                           in_25__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_25__m_axi_m_axi_BRESP,
    output wire                                          in_25__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_25__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_25__m_axi_m_axi_RID,
    output wire                                          in_25__m_axi_m_axi_RLAST,
    input wire                                           in_25__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_25__m_axi_m_axi_RRESP,
    output wire                                          in_25__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_25__m_axi_m_axi_WDATA,
    input wire                                           in_25__m_axi_m_axi_WLAST,
    output wire                                          in_25__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_25__m_axi_m_axi_WSTRB,
    input wire                                           in_25__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_25__m_axi_read_addr_din,
    input wire                                           in_25__m_axi_read_addr_full_n,
    output wire                                          in_25__m_axi_read_addr_write,
    input wire  [                                 255:0] in_25__m_axi_read_data_dout,
    input wire                                           in_25__m_axi_read_data_empty_n,
    output wire                                          in_25__m_axi_read_data_read,
    output wire                                          in_25__m_axi_rst,
    output wire [                                  63:0] in_25__m_axi_write_addr_din,
    input wire                                           in_25__m_axi_write_addr_full_n,
    output wire                                          in_25__m_axi_write_addr_write,
    output wire [                                 255:0] in_25__m_axi_write_data_din,
    input wire                                           in_25__m_axi_write_data_full_n,
    output wire                                          in_25__m_axi_write_data_write,
    input wire  [                                   7:0] in_25__m_axi_write_resp_dout,
    input wire                                           in_25__m_axi_write_resp_empty_n,
    output wire                                          in_25__m_axi_write_resp_read,
    output wire                                          in_26__m_axi_clk,
    input wire  [                                  63:0] in_26__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_26__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_26__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_26__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_26__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_26__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_26__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_26__m_axi_m_axi_ARQOS,
    output wire                                          in_26__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_26__m_axi_m_axi_ARSIZE,
    input wire                                           in_26__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_26__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_26__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_26__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_26__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_26__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_26__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_26__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_26__m_axi_m_axi_AWQOS,
    output wire                                          in_26__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_26__m_axi_m_axi_AWSIZE,
    input wire                                           in_26__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_26__m_axi_m_axi_BID,
    input wire                                           in_26__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_26__m_axi_m_axi_BRESP,
    output wire                                          in_26__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_26__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_26__m_axi_m_axi_RID,
    output wire                                          in_26__m_axi_m_axi_RLAST,
    input wire                                           in_26__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_26__m_axi_m_axi_RRESP,
    output wire                                          in_26__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_26__m_axi_m_axi_WDATA,
    input wire                                           in_26__m_axi_m_axi_WLAST,
    output wire                                          in_26__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_26__m_axi_m_axi_WSTRB,
    input wire                                           in_26__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_26__m_axi_read_addr_din,
    input wire                                           in_26__m_axi_read_addr_full_n,
    output wire                                          in_26__m_axi_read_addr_write,
    input wire  [                                 255:0] in_26__m_axi_read_data_dout,
    input wire                                           in_26__m_axi_read_data_empty_n,
    output wire                                          in_26__m_axi_read_data_read,
    output wire                                          in_26__m_axi_rst,
    output wire [                                  63:0] in_26__m_axi_write_addr_din,
    input wire                                           in_26__m_axi_write_addr_full_n,
    output wire                                          in_26__m_axi_write_addr_write,
    output wire [                                 255:0] in_26__m_axi_write_data_din,
    input wire                                           in_26__m_axi_write_data_full_n,
    output wire                                          in_26__m_axi_write_data_write,
    input wire  [                                   7:0] in_26__m_axi_write_resp_dout,
    input wire                                           in_26__m_axi_write_resp_empty_n,
    output wire                                          in_26__m_axi_write_resp_read,
    output wire                                          in_27__m_axi_clk,
    input wire  [                                  63:0] in_27__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_27__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_27__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_27__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_27__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_27__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_27__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_27__m_axi_m_axi_ARQOS,
    output wire                                          in_27__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_27__m_axi_m_axi_ARSIZE,
    input wire                                           in_27__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_27__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_27__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_27__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_27__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_27__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_27__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_27__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_27__m_axi_m_axi_AWQOS,
    output wire                                          in_27__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_27__m_axi_m_axi_AWSIZE,
    input wire                                           in_27__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_27__m_axi_m_axi_BID,
    input wire                                           in_27__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_27__m_axi_m_axi_BRESP,
    output wire                                          in_27__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_27__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_27__m_axi_m_axi_RID,
    output wire                                          in_27__m_axi_m_axi_RLAST,
    input wire                                           in_27__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_27__m_axi_m_axi_RRESP,
    output wire                                          in_27__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_27__m_axi_m_axi_WDATA,
    input wire                                           in_27__m_axi_m_axi_WLAST,
    output wire                                          in_27__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_27__m_axi_m_axi_WSTRB,
    input wire                                           in_27__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_27__m_axi_read_addr_din,
    input wire                                           in_27__m_axi_read_addr_full_n,
    output wire                                          in_27__m_axi_read_addr_write,
    input wire  [                                 255:0] in_27__m_axi_read_data_dout,
    input wire                                           in_27__m_axi_read_data_empty_n,
    output wire                                          in_27__m_axi_read_data_read,
    output wire                                          in_27__m_axi_rst,
    output wire [                                  63:0] in_27__m_axi_write_addr_din,
    input wire                                           in_27__m_axi_write_addr_full_n,
    output wire                                          in_27__m_axi_write_addr_write,
    output wire [                                 255:0] in_27__m_axi_write_data_din,
    input wire                                           in_27__m_axi_write_data_full_n,
    output wire                                          in_27__m_axi_write_data_write,
    input wire  [                                   7:0] in_27__m_axi_write_resp_dout,
    input wire                                           in_27__m_axi_write_resp_empty_n,
    output wire                                          in_27__m_axi_write_resp_read,
    output wire                                          in_28__m_axi_clk,
    input wire  [                                  63:0] in_28__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_28__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_28__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_28__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_28__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_28__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_28__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_28__m_axi_m_axi_ARQOS,
    output wire                                          in_28__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_28__m_axi_m_axi_ARSIZE,
    input wire                                           in_28__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_28__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_28__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_28__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_28__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_28__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_28__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_28__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_28__m_axi_m_axi_AWQOS,
    output wire                                          in_28__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_28__m_axi_m_axi_AWSIZE,
    input wire                                           in_28__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_28__m_axi_m_axi_BID,
    input wire                                           in_28__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_28__m_axi_m_axi_BRESP,
    output wire                                          in_28__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_28__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_28__m_axi_m_axi_RID,
    output wire                                          in_28__m_axi_m_axi_RLAST,
    input wire                                           in_28__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_28__m_axi_m_axi_RRESP,
    output wire                                          in_28__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_28__m_axi_m_axi_WDATA,
    input wire                                           in_28__m_axi_m_axi_WLAST,
    output wire                                          in_28__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_28__m_axi_m_axi_WSTRB,
    input wire                                           in_28__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_28__m_axi_read_addr_din,
    input wire                                           in_28__m_axi_read_addr_full_n,
    output wire                                          in_28__m_axi_read_addr_write,
    input wire  [                                 255:0] in_28__m_axi_read_data_dout,
    input wire                                           in_28__m_axi_read_data_empty_n,
    output wire                                          in_28__m_axi_read_data_read,
    output wire                                          in_28__m_axi_rst,
    output wire [                                  63:0] in_28__m_axi_write_addr_din,
    input wire                                           in_28__m_axi_write_addr_full_n,
    output wire                                          in_28__m_axi_write_addr_write,
    output wire [                                 255:0] in_28__m_axi_write_data_din,
    input wire                                           in_28__m_axi_write_data_full_n,
    output wire                                          in_28__m_axi_write_data_write,
    input wire  [                                   7:0] in_28__m_axi_write_resp_dout,
    input wire                                           in_28__m_axi_write_resp_empty_n,
    output wire                                          in_28__m_axi_write_resp_read,
    output wire                                          in_29__m_axi_clk,
    input wire  [                                  63:0] in_29__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_29__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_29__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_29__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_29__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_29__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_29__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_29__m_axi_m_axi_ARQOS,
    output wire                                          in_29__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_29__m_axi_m_axi_ARSIZE,
    input wire                                           in_29__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_29__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_29__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_29__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_29__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_29__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_29__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_29__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_29__m_axi_m_axi_AWQOS,
    output wire                                          in_29__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_29__m_axi_m_axi_AWSIZE,
    input wire                                           in_29__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_29__m_axi_m_axi_BID,
    input wire                                           in_29__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_29__m_axi_m_axi_BRESP,
    output wire                                          in_29__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_29__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_29__m_axi_m_axi_RID,
    output wire                                          in_29__m_axi_m_axi_RLAST,
    input wire                                           in_29__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_29__m_axi_m_axi_RRESP,
    output wire                                          in_29__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_29__m_axi_m_axi_WDATA,
    input wire                                           in_29__m_axi_m_axi_WLAST,
    output wire                                          in_29__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_29__m_axi_m_axi_WSTRB,
    input wire                                           in_29__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_29__m_axi_read_addr_din,
    input wire                                           in_29__m_axi_read_addr_full_n,
    output wire                                          in_29__m_axi_read_addr_write,
    input wire  [                                 255:0] in_29__m_axi_read_data_dout,
    input wire                                           in_29__m_axi_read_data_empty_n,
    output wire                                          in_29__m_axi_read_data_read,
    output wire                                          in_29__m_axi_rst,
    output wire [                                  63:0] in_29__m_axi_write_addr_din,
    input wire                                           in_29__m_axi_write_addr_full_n,
    output wire                                          in_29__m_axi_write_addr_write,
    output wire [                                 255:0] in_29__m_axi_write_data_din,
    input wire                                           in_29__m_axi_write_data_full_n,
    output wire                                          in_29__m_axi_write_data_write,
    input wire  [                                   7:0] in_29__m_axi_write_resp_dout,
    input wire                                           in_29__m_axi_write_resp_empty_n,
    output wire                                          in_29__m_axi_write_resp_read,
    output wire                                          in_3__m_axi_clk,
    input wire  [                                  63:0] in_3__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_3__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_3__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_3__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_3__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_3__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_3__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_3__m_axi_m_axi_ARQOS,
    output wire                                          in_3__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_3__m_axi_m_axi_ARSIZE,
    input wire                                           in_3__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_3__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_3__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_3__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_3__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_3__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_3__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_3__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_3__m_axi_m_axi_AWQOS,
    output wire                                          in_3__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_3__m_axi_m_axi_AWSIZE,
    input wire                                           in_3__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_3__m_axi_m_axi_BID,
    input wire                                           in_3__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_3__m_axi_m_axi_BRESP,
    output wire                                          in_3__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_3__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_3__m_axi_m_axi_RID,
    output wire                                          in_3__m_axi_m_axi_RLAST,
    input wire                                           in_3__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_3__m_axi_m_axi_RRESP,
    output wire                                          in_3__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_3__m_axi_m_axi_WDATA,
    input wire                                           in_3__m_axi_m_axi_WLAST,
    output wire                                          in_3__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_3__m_axi_m_axi_WSTRB,
    input wire                                           in_3__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_3__m_axi_read_addr_din,
    input wire                                           in_3__m_axi_read_addr_full_n,
    output wire                                          in_3__m_axi_read_addr_write,
    input wire  [                                 255:0] in_3__m_axi_read_data_dout,
    input wire                                           in_3__m_axi_read_data_empty_n,
    output wire                                          in_3__m_axi_read_data_read,
    output wire                                          in_3__m_axi_rst,
    output wire [                                  63:0] in_3__m_axi_write_addr_din,
    input wire                                           in_3__m_axi_write_addr_full_n,
    output wire                                          in_3__m_axi_write_addr_write,
    output wire [                                 255:0] in_3__m_axi_write_data_din,
    input wire                                           in_3__m_axi_write_data_full_n,
    output wire                                          in_3__m_axi_write_data_write,
    input wire  [                                   7:0] in_3__m_axi_write_resp_dout,
    input wire                                           in_3__m_axi_write_resp_empty_n,
    output wire                                          in_3__m_axi_write_resp_read,
    output wire                                          in_30__m_axi_clk,
    input wire  [                                  63:0] in_30__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_30__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_30__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_30__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_30__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_30__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_30__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_30__m_axi_m_axi_ARQOS,
    output wire                                          in_30__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_30__m_axi_m_axi_ARSIZE,
    input wire                                           in_30__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_30__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_30__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_30__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_30__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_30__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_30__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_30__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_30__m_axi_m_axi_AWQOS,
    output wire                                          in_30__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_30__m_axi_m_axi_AWSIZE,
    input wire                                           in_30__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_30__m_axi_m_axi_BID,
    input wire                                           in_30__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_30__m_axi_m_axi_BRESP,
    output wire                                          in_30__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_30__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_30__m_axi_m_axi_RID,
    output wire                                          in_30__m_axi_m_axi_RLAST,
    input wire                                           in_30__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_30__m_axi_m_axi_RRESP,
    output wire                                          in_30__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_30__m_axi_m_axi_WDATA,
    input wire                                           in_30__m_axi_m_axi_WLAST,
    output wire                                          in_30__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_30__m_axi_m_axi_WSTRB,
    input wire                                           in_30__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_30__m_axi_read_addr_din,
    input wire                                           in_30__m_axi_read_addr_full_n,
    output wire                                          in_30__m_axi_read_addr_write,
    input wire  [                                 255:0] in_30__m_axi_read_data_dout,
    input wire                                           in_30__m_axi_read_data_empty_n,
    output wire                                          in_30__m_axi_read_data_read,
    output wire                                          in_30__m_axi_rst,
    output wire [                                  63:0] in_30__m_axi_write_addr_din,
    input wire                                           in_30__m_axi_write_addr_full_n,
    output wire                                          in_30__m_axi_write_addr_write,
    output wire [                                 255:0] in_30__m_axi_write_data_din,
    input wire                                           in_30__m_axi_write_data_full_n,
    output wire                                          in_30__m_axi_write_data_write,
    input wire  [                                   7:0] in_30__m_axi_write_resp_dout,
    input wire                                           in_30__m_axi_write_resp_empty_n,
    output wire                                          in_30__m_axi_write_resp_read,
    output wire                                          in_31__m_axi_clk,
    input wire  [                                  63:0] in_31__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_31__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_31__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_31__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_31__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_31__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_31__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_31__m_axi_m_axi_ARQOS,
    output wire                                          in_31__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_31__m_axi_m_axi_ARSIZE,
    input wire                                           in_31__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_31__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_31__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_31__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_31__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_31__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_31__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_31__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_31__m_axi_m_axi_AWQOS,
    output wire                                          in_31__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_31__m_axi_m_axi_AWSIZE,
    input wire                                           in_31__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_31__m_axi_m_axi_BID,
    input wire                                           in_31__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_31__m_axi_m_axi_BRESP,
    output wire                                          in_31__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_31__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_31__m_axi_m_axi_RID,
    output wire                                          in_31__m_axi_m_axi_RLAST,
    input wire                                           in_31__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_31__m_axi_m_axi_RRESP,
    output wire                                          in_31__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_31__m_axi_m_axi_WDATA,
    input wire                                           in_31__m_axi_m_axi_WLAST,
    output wire                                          in_31__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_31__m_axi_m_axi_WSTRB,
    input wire                                           in_31__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_31__m_axi_read_addr_din,
    input wire                                           in_31__m_axi_read_addr_full_n,
    output wire                                          in_31__m_axi_read_addr_write,
    input wire  [                                 255:0] in_31__m_axi_read_data_dout,
    input wire                                           in_31__m_axi_read_data_empty_n,
    output wire                                          in_31__m_axi_read_data_read,
    output wire                                          in_31__m_axi_rst,
    output wire [                                  63:0] in_31__m_axi_write_addr_din,
    input wire                                           in_31__m_axi_write_addr_full_n,
    output wire                                          in_31__m_axi_write_addr_write,
    output wire [                                 255:0] in_31__m_axi_write_data_din,
    input wire                                           in_31__m_axi_write_data_full_n,
    output wire                                          in_31__m_axi_write_data_write,
    input wire  [                                   7:0] in_31__m_axi_write_resp_dout,
    input wire                                           in_31__m_axi_write_resp_empty_n,
    output wire                                          in_31__m_axi_write_resp_read,
    output wire                                          in_32__m_axi_clk,
    input wire  [                                  63:0] in_32__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_32__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_32__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_32__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_32__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_32__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_32__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_32__m_axi_m_axi_ARQOS,
    output wire                                          in_32__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_32__m_axi_m_axi_ARSIZE,
    input wire                                           in_32__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_32__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_32__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_32__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_32__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_32__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_32__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_32__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_32__m_axi_m_axi_AWQOS,
    output wire                                          in_32__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_32__m_axi_m_axi_AWSIZE,
    input wire                                           in_32__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_32__m_axi_m_axi_BID,
    input wire                                           in_32__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_32__m_axi_m_axi_BRESP,
    output wire                                          in_32__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_32__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_32__m_axi_m_axi_RID,
    output wire                                          in_32__m_axi_m_axi_RLAST,
    input wire                                           in_32__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_32__m_axi_m_axi_RRESP,
    output wire                                          in_32__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_32__m_axi_m_axi_WDATA,
    input wire                                           in_32__m_axi_m_axi_WLAST,
    output wire                                          in_32__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_32__m_axi_m_axi_WSTRB,
    input wire                                           in_32__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_32__m_axi_read_addr_din,
    input wire                                           in_32__m_axi_read_addr_full_n,
    output wire                                          in_32__m_axi_read_addr_write,
    input wire  [                                 255:0] in_32__m_axi_read_data_dout,
    input wire                                           in_32__m_axi_read_data_empty_n,
    output wire                                          in_32__m_axi_read_data_read,
    output wire                                          in_32__m_axi_rst,
    output wire [                                  63:0] in_32__m_axi_write_addr_din,
    input wire                                           in_32__m_axi_write_addr_full_n,
    output wire                                          in_32__m_axi_write_addr_write,
    output wire [                                 255:0] in_32__m_axi_write_data_din,
    input wire                                           in_32__m_axi_write_data_full_n,
    output wire                                          in_32__m_axi_write_data_write,
    input wire  [                                   7:0] in_32__m_axi_write_resp_dout,
    input wire                                           in_32__m_axi_write_resp_empty_n,
    output wire                                          in_32__m_axi_write_resp_read,
    output wire                                          in_33__m_axi_clk,
    input wire  [                                  63:0] in_33__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_33__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_33__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_33__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_33__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_33__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_33__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_33__m_axi_m_axi_ARQOS,
    output wire                                          in_33__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_33__m_axi_m_axi_ARSIZE,
    input wire                                           in_33__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_33__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_33__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_33__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_33__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_33__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_33__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_33__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_33__m_axi_m_axi_AWQOS,
    output wire                                          in_33__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_33__m_axi_m_axi_AWSIZE,
    input wire                                           in_33__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_33__m_axi_m_axi_BID,
    input wire                                           in_33__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_33__m_axi_m_axi_BRESP,
    output wire                                          in_33__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_33__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_33__m_axi_m_axi_RID,
    output wire                                          in_33__m_axi_m_axi_RLAST,
    input wire                                           in_33__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_33__m_axi_m_axi_RRESP,
    output wire                                          in_33__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_33__m_axi_m_axi_WDATA,
    input wire                                           in_33__m_axi_m_axi_WLAST,
    output wire                                          in_33__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_33__m_axi_m_axi_WSTRB,
    input wire                                           in_33__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_33__m_axi_read_addr_din,
    input wire                                           in_33__m_axi_read_addr_full_n,
    output wire                                          in_33__m_axi_read_addr_write,
    input wire  [                                 255:0] in_33__m_axi_read_data_dout,
    input wire                                           in_33__m_axi_read_data_empty_n,
    output wire                                          in_33__m_axi_read_data_read,
    output wire                                          in_33__m_axi_rst,
    output wire [                                  63:0] in_33__m_axi_write_addr_din,
    input wire                                           in_33__m_axi_write_addr_full_n,
    output wire                                          in_33__m_axi_write_addr_write,
    output wire [                                 255:0] in_33__m_axi_write_data_din,
    input wire                                           in_33__m_axi_write_data_full_n,
    output wire                                          in_33__m_axi_write_data_write,
    input wire  [                                   7:0] in_33__m_axi_write_resp_dout,
    input wire                                           in_33__m_axi_write_resp_empty_n,
    output wire                                          in_33__m_axi_write_resp_read,
    output wire                                          in_34__m_axi_clk,
    input wire  [                                  63:0] in_34__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_34__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_34__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_34__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_34__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_34__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_34__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_34__m_axi_m_axi_ARQOS,
    output wire                                          in_34__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_34__m_axi_m_axi_ARSIZE,
    input wire                                           in_34__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_34__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_34__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_34__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_34__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_34__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_34__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_34__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_34__m_axi_m_axi_AWQOS,
    output wire                                          in_34__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_34__m_axi_m_axi_AWSIZE,
    input wire                                           in_34__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_34__m_axi_m_axi_BID,
    input wire                                           in_34__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_34__m_axi_m_axi_BRESP,
    output wire                                          in_34__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_34__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_34__m_axi_m_axi_RID,
    output wire                                          in_34__m_axi_m_axi_RLAST,
    input wire                                           in_34__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_34__m_axi_m_axi_RRESP,
    output wire                                          in_34__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_34__m_axi_m_axi_WDATA,
    input wire                                           in_34__m_axi_m_axi_WLAST,
    output wire                                          in_34__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_34__m_axi_m_axi_WSTRB,
    input wire                                           in_34__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_34__m_axi_read_addr_din,
    input wire                                           in_34__m_axi_read_addr_full_n,
    output wire                                          in_34__m_axi_read_addr_write,
    input wire  [                                 255:0] in_34__m_axi_read_data_dout,
    input wire                                           in_34__m_axi_read_data_empty_n,
    output wire                                          in_34__m_axi_read_data_read,
    output wire                                          in_34__m_axi_rst,
    output wire [                                  63:0] in_34__m_axi_write_addr_din,
    input wire                                           in_34__m_axi_write_addr_full_n,
    output wire                                          in_34__m_axi_write_addr_write,
    output wire [                                 255:0] in_34__m_axi_write_data_din,
    input wire                                           in_34__m_axi_write_data_full_n,
    output wire                                          in_34__m_axi_write_data_write,
    input wire  [                                   7:0] in_34__m_axi_write_resp_dout,
    input wire                                           in_34__m_axi_write_resp_empty_n,
    output wire                                          in_34__m_axi_write_resp_read,
    output wire                                          in_35__m_axi_clk,
    input wire  [                                  63:0] in_35__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_35__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_35__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_35__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_35__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_35__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_35__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_35__m_axi_m_axi_ARQOS,
    output wire                                          in_35__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_35__m_axi_m_axi_ARSIZE,
    input wire                                           in_35__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_35__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_35__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_35__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_35__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_35__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_35__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_35__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_35__m_axi_m_axi_AWQOS,
    output wire                                          in_35__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_35__m_axi_m_axi_AWSIZE,
    input wire                                           in_35__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_35__m_axi_m_axi_BID,
    input wire                                           in_35__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_35__m_axi_m_axi_BRESP,
    output wire                                          in_35__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_35__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_35__m_axi_m_axi_RID,
    output wire                                          in_35__m_axi_m_axi_RLAST,
    input wire                                           in_35__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_35__m_axi_m_axi_RRESP,
    output wire                                          in_35__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_35__m_axi_m_axi_WDATA,
    input wire                                           in_35__m_axi_m_axi_WLAST,
    output wire                                          in_35__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_35__m_axi_m_axi_WSTRB,
    input wire                                           in_35__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_35__m_axi_read_addr_din,
    input wire                                           in_35__m_axi_read_addr_full_n,
    output wire                                          in_35__m_axi_read_addr_write,
    input wire  [                                 255:0] in_35__m_axi_read_data_dout,
    input wire                                           in_35__m_axi_read_data_empty_n,
    output wire                                          in_35__m_axi_read_data_read,
    output wire                                          in_35__m_axi_rst,
    output wire [                                  63:0] in_35__m_axi_write_addr_din,
    input wire                                           in_35__m_axi_write_addr_full_n,
    output wire                                          in_35__m_axi_write_addr_write,
    output wire [                                 255:0] in_35__m_axi_write_data_din,
    input wire                                           in_35__m_axi_write_data_full_n,
    output wire                                          in_35__m_axi_write_data_write,
    input wire  [                                   7:0] in_35__m_axi_write_resp_dout,
    input wire                                           in_35__m_axi_write_resp_empty_n,
    output wire                                          in_35__m_axi_write_resp_read,
    output wire                                          in_36__m_axi_clk,
    input wire  [                                  63:0] in_36__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_36__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_36__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_36__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_36__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_36__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_36__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_36__m_axi_m_axi_ARQOS,
    output wire                                          in_36__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_36__m_axi_m_axi_ARSIZE,
    input wire                                           in_36__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_36__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_36__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_36__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_36__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_36__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_36__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_36__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_36__m_axi_m_axi_AWQOS,
    output wire                                          in_36__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_36__m_axi_m_axi_AWSIZE,
    input wire                                           in_36__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_36__m_axi_m_axi_BID,
    input wire                                           in_36__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_36__m_axi_m_axi_BRESP,
    output wire                                          in_36__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_36__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_36__m_axi_m_axi_RID,
    output wire                                          in_36__m_axi_m_axi_RLAST,
    input wire                                           in_36__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_36__m_axi_m_axi_RRESP,
    output wire                                          in_36__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_36__m_axi_m_axi_WDATA,
    input wire                                           in_36__m_axi_m_axi_WLAST,
    output wire                                          in_36__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_36__m_axi_m_axi_WSTRB,
    input wire                                           in_36__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_36__m_axi_read_addr_din,
    input wire                                           in_36__m_axi_read_addr_full_n,
    output wire                                          in_36__m_axi_read_addr_write,
    input wire  [                                 255:0] in_36__m_axi_read_data_dout,
    input wire                                           in_36__m_axi_read_data_empty_n,
    output wire                                          in_36__m_axi_read_data_read,
    output wire                                          in_36__m_axi_rst,
    output wire [                                  63:0] in_36__m_axi_write_addr_din,
    input wire                                           in_36__m_axi_write_addr_full_n,
    output wire                                          in_36__m_axi_write_addr_write,
    output wire [                                 255:0] in_36__m_axi_write_data_din,
    input wire                                           in_36__m_axi_write_data_full_n,
    output wire                                          in_36__m_axi_write_data_write,
    input wire  [                                   7:0] in_36__m_axi_write_resp_dout,
    input wire                                           in_36__m_axi_write_resp_empty_n,
    output wire                                          in_36__m_axi_write_resp_read,
    output wire                                          in_37__m_axi_clk,
    input wire  [                                  63:0] in_37__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_37__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_37__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_37__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_37__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_37__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_37__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_37__m_axi_m_axi_ARQOS,
    output wire                                          in_37__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_37__m_axi_m_axi_ARSIZE,
    input wire                                           in_37__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_37__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_37__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_37__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_37__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_37__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_37__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_37__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_37__m_axi_m_axi_AWQOS,
    output wire                                          in_37__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_37__m_axi_m_axi_AWSIZE,
    input wire                                           in_37__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_37__m_axi_m_axi_BID,
    input wire                                           in_37__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_37__m_axi_m_axi_BRESP,
    output wire                                          in_37__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_37__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_37__m_axi_m_axi_RID,
    output wire                                          in_37__m_axi_m_axi_RLAST,
    input wire                                           in_37__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_37__m_axi_m_axi_RRESP,
    output wire                                          in_37__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_37__m_axi_m_axi_WDATA,
    input wire                                           in_37__m_axi_m_axi_WLAST,
    output wire                                          in_37__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_37__m_axi_m_axi_WSTRB,
    input wire                                           in_37__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_37__m_axi_read_addr_din,
    input wire                                           in_37__m_axi_read_addr_full_n,
    output wire                                          in_37__m_axi_read_addr_write,
    input wire  [                                 255:0] in_37__m_axi_read_data_dout,
    input wire                                           in_37__m_axi_read_data_empty_n,
    output wire                                          in_37__m_axi_read_data_read,
    output wire                                          in_37__m_axi_rst,
    output wire [                                  63:0] in_37__m_axi_write_addr_din,
    input wire                                           in_37__m_axi_write_addr_full_n,
    output wire                                          in_37__m_axi_write_addr_write,
    output wire [                                 255:0] in_37__m_axi_write_data_din,
    input wire                                           in_37__m_axi_write_data_full_n,
    output wire                                          in_37__m_axi_write_data_write,
    input wire  [                                   7:0] in_37__m_axi_write_resp_dout,
    input wire                                           in_37__m_axi_write_resp_empty_n,
    output wire                                          in_37__m_axi_write_resp_read,
    output wire                                          in_38__m_axi_clk,
    input wire  [                                  63:0] in_38__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_38__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_38__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_38__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_38__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_38__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_38__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_38__m_axi_m_axi_ARQOS,
    output wire                                          in_38__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_38__m_axi_m_axi_ARSIZE,
    input wire                                           in_38__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_38__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_38__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_38__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_38__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_38__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_38__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_38__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_38__m_axi_m_axi_AWQOS,
    output wire                                          in_38__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_38__m_axi_m_axi_AWSIZE,
    input wire                                           in_38__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_38__m_axi_m_axi_BID,
    input wire                                           in_38__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_38__m_axi_m_axi_BRESP,
    output wire                                          in_38__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_38__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_38__m_axi_m_axi_RID,
    output wire                                          in_38__m_axi_m_axi_RLAST,
    input wire                                           in_38__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_38__m_axi_m_axi_RRESP,
    output wire                                          in_38__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_38__m_axi_m_axi_WDATA,
    input wire                                           in_38__m_axi_m_axi_WLAST,
    output wire                                          in_38__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_38__m_axi_m_axi_WSTRB,
    input wire                                           in_38__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_38__m_axi_read_addr_din,
    input wire                                           in_38__m_axi_read_addr_full_n,
    output wire                                          in_38__m_axi_read_addr_write,
    input wire  [                                 255:0] in_38__m_axi_read_data_dout,
    input wire                                           in_38__m_axi_read_data_empty_n,
    output wire                                          in_38__m_axi_read_data_read,
    output wire                                          in_38__m_axi_rst,
    output wire [                                  63:0] in_38__m_axi_write_addr_din,
    input wire                                           in_38__m_axi_write_addr_full_n,
    output wire                                          in_38__m_axi_write_addr_write,
    output wire [                                 255:0] in_38__m_axi_write_data_din,
    input wire                                           in_38__m_axi_write_data_full_n,
    output wire                                          in_38__m_axi_write_data_write,
    input wire  [                                   7:0] in_38__m_axi_write_resp_dout,
    input wire                                           in_38__m_axi_write_resp_empty_n,
    output wire                                          in_38__m_axi_write_resp_read,
    output wire                                          in_39__m_axi_clk,
    input wire  [                                  63:0] in_39__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_39__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_39__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_39__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_39__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_39__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_39__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_39__m_axi_m_axi_ARQOS,
    output wire                                          in_39__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_39__m_axi_m_axi_ARSIZE,
    input wire                                           in_39__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_39__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_39__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_39__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_39__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_39__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_39__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_39__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_39__m_axi_m_axi_AWQOS,
    output wire                                          in_39__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_39__m_axi_m_axi_AWSIZE,
    input wire                                           in_39__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_39__m_axi_m_axi_BID,
    input wire                                           in_39__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_39__m_axi_m_axi_BRESP,
    output wire                                          in_39__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_39__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_39__m_axi_m_axi_RID,
    output wire                                          in_39__m_axi_m_axi_RLAST,
    input wire                                           in_39__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_39__m_axi_m_axi_RRESP,
    output wire                                          in_39__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_39__m_axi_m_axi_WDATA,
    input wire                                           in_39__m_axi_m_axi_WLAST,
    output wire                                          in_39__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_39__m_axi_m_axi_WSTRB,
    input wire                                           in_39__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_39__m_axi_read_addr_din,
    input wire                                           in_39__m_axi_read_addr_full_n,
    output wire                                          in_39__m_axi_read_addr_write,
    input wire  [                                 255:0] in_39__m_axi_read_data_dout,
    input wire                                           in_39__m_axi_read_data_empty_n,
    output wire                                          in_39__m_axi_read_data_read,
    output wire                                          in_39__m_axi_rst,
    output wire [                                  63:0] in_39__m_axi_write_addr_din,
    input wire                                           in_39__m_axi_write_addr_full_n,
    output wire                                          in_39__m_axi_write_addr_write,
    output wire [                                 255:0] in_39__m_axi_write_data_din,
    input wire                                           in_39__m_axi_write_data_full_n,
    output wire                                          in_39__m_axi_write_data_write,
    input wire  [                                   7:0] in_39__m_axi_write_resp_dout,
    input wire                                           in_39__m_axi_write_resp_empty_n,
    output wire                                          in_39__m_axi_write_resp_read,
    output wire                                          in_4__m_axi_clk,
    input wire  [                                  63:0] in_4__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_4__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_4__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_4__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_4__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_4__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_4__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_4__m_axi_m_axi_ARQOS,
    output wire                                          in_4__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_4__m_axi_m_axi_ARSIZE,
    input wire                                           in_4__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_4__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_4__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_4__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_4__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_4__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_4__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_4__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_4__m_axi_m_axi_AWQOS,
    output wire                                          in_4__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_4__m_axi_m_axi_AWSIZE,
    input wire                                           in_4__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_4__m_axi_m_axi_BID,
    input wire                                           in_4__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_4__m_axi_m_axi_BRESP,
    output wire                                          in_4__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_4__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_4__m_axi_m_axi_RID,
    output wire                                          in_4__m_axi_m_axi_RLAST,
    input wire                                           in_4__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_4__m_axi_m_axi_RRESP,
    output wire                                          in_4__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_4__m_axi_m_axi_WDATA,
    input wire                                           in_4__m_axi_m_axi_WLAST,
    output wire                                          in_4__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_4__m_axi_m_axi_WSTRB,
    input wire                                           in_4__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_4__m_axi_read_addr_din,
    input wire                                           in_4__m_axi_read_addr_full_n,
    output wire                                          in_4__m_axi_read_addr_write,
    input wire  [                                 255:0] in_4__m_axi_read_data_dout,
    input wire                                           in_4__m_axi_read_data_empty_n,
    output wire                                          in_4__m_axi_read_data_read,
    output wire                                          in_4__m_axi_rst,
    output wire [                                  63:0] in_4__m_axi_write_addr_din,
    input wire                                           in_4__m_axi_write_addr_full_n,
    output wire                                          in_4__m_axi_write_addr_write,
    output wire [                                 255:0] in_4__m_axi_write_data_din,
    input wire                                           in_4__m_axi_write_data_full_n,
    output wire                                          in_4__m_axi_write_data_write,
    input wire  [                                   7:0] in_4__m_axi_write_resp_dout,
    input wire                                           in_4__m_axi_write_resp_empty_n,
    output wire                                          in_4__m_axi_write_resp_read,
    output wire                                          in_40__m_axi_clk,
    input wire  [                                  63:0] in_40__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_40__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_40__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_40__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_40__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_40__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_40__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_40__m_axi_m_axi_ARQOS,
    output wire                                          in_40__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_40__m_axi_m_axi_ARSIZE,
    input wire                                           in_40__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_40__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_40__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_40__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_40__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_40__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_40__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_40__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_40__m_axi_m_axi_AWQOS,
    output wire                                          in_40__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_40__m_axi_m_axi_AWSIZE,
    input wire                                           in_40__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_40__m_axi_m_axi_BID,
    input wire                                           in_40__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_40__m_axi_m_axi_BRESP,
    output wire                                          in_40__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_40__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_40__m_axi_m_axi_RID,
    output wire                                          in_40__m_axi_m_axi_RLAST,
    input wire                                           in_40__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_40__m_axi_m_axi_RRESP,
    output wire                                          in_40__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_40__m_axi_m_axi_WDATA,
    input wire                                           in_40__m_axi_m_axi_WLAST,
    output wire                                          in_40__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_40__m_axi_m_axi_WSTRB,
    input wire                                           in_40__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_40__m_axi_read_addr_din,
    input wire                                           in_40__m_axi_read_addr_full_n,
    output wire                                          in_40__m_axi_read_addr_write,
    input wire  [                                 255:0] in_40__m_axi_read_data_dout,
    input wire                                           in_40__m_axi_read_data_empty_n,
    output wire                                          in_40__m_axi_read_data_read,
    output wire                                          in_40__m_axi_rst,
    output wire [                                  63:0] in_40__m_axi_write_addr_din,
    input wire                                           in_40__m_axi_write_addr_full_n,
    output wire                                          in_40__m_axi_write_addr_write,
    output wire [                                 255:0] in_40__m_axi_write_data_din,
    input wire                                           in_40__m_axi_write_data_full_n,
    output wire                                          in_40__m_axi_write_data_write,
    input wire  [                                   7:0] in_40__m_axi_write_resp_dout,
    input wire                                           in_40__m_axi_write_resp_empty_n,
    output wire                                          in_40__m_axi_write_resp_read,
    output wire                                          in_41__m_axi_clk,
    input wire  [                                  63:0] in_41__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_41__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_41__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_41__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_41__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_41__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_41__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_41__m_axi_m_axi_ARQOS,
    output wire                                          in_41__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_41__m_axi_m_axi_ARSIZE,
    input wire                                           in_41__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_41__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_41__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_41__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_41__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_41__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_41__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_41__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_41__m_axi_m_axi_AWQOS,
    output wire                                          in_41__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_41__m_axi_m_axi_AWSIZE,
    input wire                                           in_41__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_41__m_axi_m_axi_BID,
    input wire                                           in_41__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_41__m_axi_m_axi_BRESP,
    output wire                                          in_41__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_41__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_41__m_axi_m_axi_RID,
    output wire                                          in_41__m_axi_m_axi_RLAST,
    input wire                                           in_41__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_41__m_axi_m_axi_RRESP,
    output wire                                          in_41__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_41__m_axi_m_axi_WDATA,
    input wire                                           in_41__m_axi_m_axi_WLAST,
    output wire                                          in_41__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_41__m_axi_m_axi_WSTRB,
    input wire                                           in_41__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_41__m_axi_read_addr_din,
    input wire                                           in_41__m_axi_read_addr_full_n,
    output wire                                          in_41__m_axi_read_addr_write,
    input wire  [                                 255:0] in_41__m_axi_read_data_dout,
    input wire                                           in_41__m_axi_read_data_empty_n,
    output wire                                          in_41__m_axi_read_data_read,
    output wire                                          in_41__m_axi_rst,
    output wire [                                  63:0] in_41__m_axi_write_addr_din,
    input wire                                           in_41__m_axi_write_addr_full_n,
    output wire                                          in_41__m_axi_write_addr_write,
    output wire [                                 255:0] in_41__m_axi_write_data_din,
    input wire                                           in_41__m_axi_write_data_full_n,
    output wire                                          in_41__m_axi_write_data_write,
    input wire  [                                   7:0] in_41__m_axi_write_resp_dout,
    input wire                                           in_41__m_axi_write_resp_empty_n,
    output wire                                          in_41__m_axi_write_resp_read,
    output wire                                          in_42__m_axi_clk,
    input wire  [                                  63:0] in_42__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_42__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_42__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_42__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_42__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_42__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_42__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_42__m_axi_m_axi_ARQOS,
    output wire                                          in_42__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_42__m_axi_m_axi_ARSIZE,
    input wire                                           in_42__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_42__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_42__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_42__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_42__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_42__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_42__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_42__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_42__m_axi_m_axi_AWQOS,
    output wire                                          in_42__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_42__m_axi_m_axi_AWSIZE,
    input wire                                           in_42__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_42__m_axi_m_axi_BID,
    input wire                                           in_42__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_42__m_axi_m_axi_BRESP,
    output wire                                          in_42__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_42__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_42__m_axi_m_axi_RID,
    output wire                                          in_42__m_axi_m_axi_RLAST,
    input wire                                           in_42__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_42__m_axi_m_axi_RRESP,
    output wire                                          in_42__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_42__m_axi_m_axi_WDATA,
    input wire                                           in_42__m_axi_m_axi_WLAST,
    output wire                                          in_42__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_42__m_axi_m_axi_WSTRB,
    input wire                                           in_42__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_42__m_axi_read_addr_din,
    input wire                                           in_42__m_axi_read_addr_full_n,
    output wire                                          in_42__m_axi_read_addr_write,
    input wire  [                                 255:0] in_42__m_axi_read_data_dout,
    input wire                                           in_42__m_axi_read_data_empty_n,
    output wire                                          in_42__m_axi_read_data_read,
    output wire                                          in_42__m_axi_rst,
    output wire [                                  63:0] in_42__m_axi_write_addr_din,
    input wire                                           in_42__m_axi_write_addr_full_n,
    output wire                                          in_42__m_axi_write_addr_write,
    output wire [                                 255:0] in_42__m_axi_write_data_din,
    input wire                                           in_42__m_axi_write_data_full_n,
    output wire                                          in_42__m_axi_write_data_write,
    input wire  [                                   7:0] in_42__m_axi_write_resp_dout,
    input wire                                           in_42__m_axi_write_resp_empty_n,
    output wire                                          in_42__m_axi_write_resp_read,
    output wire                                          in_43__m_axi_clk,
    input wire  [                                  63:0] in_43__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_43__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_43__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_43__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_43__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_43__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_43__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_43__m_axi_m_axi_ARQOS,
    output wire                                          in_43__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_43__m_axi_m_axi_ARSIZE,
    input wire                                           in_43__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_43__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_43__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_43__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_43__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_43__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_43__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_43__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_43__m_axi_m_axi_AWQOS,
    output wire                                          in_43__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_43__m_axi_m_axi_AWSIZE,
    input wire                                           in_43__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_43__m_axi_m_axi_BID,
    input wire                                           in_43__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_43__m_axi_m_axi_BRESP,
    output wire                                          in_43__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_43__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_43__m_axi_m_axi_RID,
    output wire                                          in_43__m_axi_m_axi_RLAST,
    input wire                                           in_43__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_43__m_axi_m_axi_RRESP,
    output wire                                          in_43__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_43__m_axi_m_axi_WDATA,
    input wire                                           in_43__m_axi_m_axi_WLAST,
    output wire                                          in_43__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_43__m_axi_m_axi_WSTRB,
    input wire                                           in_43__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_43__m_axi_read_addr_din,
    input wire                                           in_43__m_axi_read_addr_full_n,
    output wire                                          in_43__m_axi_read_addr_write,
    input wire  [                                 255:0] in_43__m_axi_read_data_dout,
    input wire                                           in_43__m_axi_read_data_empty_n,
    output wire                                          in_43__m_axi_read_data_read,
    output wire                                          in_43__m_axi_rst,
    output wire [                                  63:0] in_43__m_axi_write_addr_din,
    input wire                                           in_43__m_axi_write_addr_full_n,
    output wire                                          in_43__m_axi_write_addr_write,
    output wire [                                 255:0] in_43__m_axi_write_data_din,
    input wire                                           in_43__m_axi_write_data_full_n,
    output wire                                          in_43__m_axi_write_data_write,
    input wire  [                                   7:0] in_43__m_axi_write_resp_dout,
    input wire                                           in_43__m_axi_write_resp_empty_n,
    output wire                                          in_43__m_axi_write_resp_read,
    output wire                                          in_44__m_axi_clk,
    input wire  [                                  63:0] in_44__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_44__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_44__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_44__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_44__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_44__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_44__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_44__m_axi_m_axi_ARQOS,
    output wire                                          in_44__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_44__m_axi_m_axi_ARSIZE,
    input wire                                           in_44__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_44__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_44__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_44__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_44__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_44__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_44__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_44__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_44__m_axi_m_axi_AWQOS,
    output wire                                          in_44__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_44__m_axi_m_axi_AWSIZE,
    input wire                                           in_44__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_44__m_axi_m_axi_BID,
    input wire                                           in_44__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_44__m_axi_m_axi_BRESP,
    output wire                                          in_44__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_44__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_44__m_axi_m_axi_RID,
    output wire                                          in_44__m_axi_m_axi_RLAST,
    input wire                                           in_44__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_44__m_axi_m_axi_RRESP,
    output wire                                          in_44__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_44__m_axi_m_axi_WDATA,
    input wire                                           in_44__m_axi_m_axi_WLAST,
    output wire                                          in_44__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_44__m_axi_m_axi_WSTRB,
    input wire                                           in_44__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_44__m_axi_read_addr_din,
    input wire                                           in_44__m_axi_read_addr_full_n,
    output wire                                          in_44__m_axi_read_addr_write,
    input wire  [                                 255:0] in_44__m_axi_read_data_dout,
    input wire                                           in_44__m_axi_read_data_empty_n,
    output wire                                          in_44__m_axi_read_data_read,
    output wire                                          in_44__m_axi_rst,
    output wire [                                  63:0] in_44__m_axi_write_addr_din,
    input wire                                           in_44__m_axi_write_addr_full_n,
    output wire                                          in_44__m_axi_write_addr_write,
    output wire [                                 255:0] in_44__m_axi_write_data_din,
    input wire                                           in_44__m_axi_write_data_full_n,
    output wire                                          in_44__m_axi_write_data_write,
    input wire  [                                   7:0] in_44__m_axi_write_resp_dout,
    input wire                                           in_44__m_axi_write_resp_empty_n,
    output wire                                          in_44__m_axi_write_resp_read,
    output wire                                          in_45__m_axi_clk,
    input wire  [                                  63:0] in_45__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_45__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_45__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_45__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_45__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_45__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_45__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_45__m_axi_m_axi_ARQOS,
    output wire                                          in_45__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_45__m_axi_m_axi_ARSIZE,
    input wire                                           in_45__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_45__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_45__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_45__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_45__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_45__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_45__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_45__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_45__m_axi_m_axi_AWQOS,
    output wire                                          in_45__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_45__m_axi_m_axi_AWSIZE,
    input wire                                           in_45__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_45__m_axi_m_axi_BID,
    input wire                                           in_45__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_45__m_axi_m_axi_BRESP,
    output wire                                          in_45__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_45__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_45__m_axi_m_axi_RID,
    output wire                                          in_45__m_axi_m_axi_RLAST,
    input wire                                           in_45__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_45__m_axi_m_axi_RRESP,
    output wire                                          in_45__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_45__m_axi_m_axi_WDATA,
    input wire                                           in_45__m_axi_m_axi_WLAST,
    output wire                                          in_45__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_45__m_axi_m_axi_WSTRB,
    input wire                                           in_45__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_45__m_axi_read_addr_din,
    input wire                                           in_45__m_axi_read_addr_full_n,
    output wire                                          in_45__m_axi_read_addr_write,
    input wire  [                                 255:0] in_45__m_axi_read_data_dout,
    input wire                                           in_45__m_axi_read_data_empty_n,
    output wire                                          in_45__m_axi_read_data_read,
    output wire                                          in_45__m_axi_rst,
    output wire [                                  63:0] in_45__m_axi_write_addr_din,
    input wire                                           in_45__m_axi_write_addr_full_n,
    output wire                                          in_45__m_axi_write_addr_write,
    output wire [                                 255:0] in_45__m_axi_write_data_din,
    input wire                                           in_45__m_axi_write_data_full_n,
    output wire                                          in_45__m_axi_write_data_write,
    input wire  [                                   7:0] in_45__m_axi_write_resp_dout,
    input wire                                           in_45__m_axi_write_resp_empty_n,
    output wire                                          in_45__m_axi_write_resp_read,
    output wire                                          in_46__m_axi_clk,
    input wire  [                                  63:0] in_46__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_46__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_46__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_46__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_46__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_46__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_46__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_46__m_axi_m_axi_ARQOS,
    output wire                                          in_46__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_46__m_axi_m_axi_ARSIZE,
    input wire                                           in_46__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_46__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_46__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_46__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_46__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_46__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_46__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_46__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_46__m_axi_m_axi_AWQOS,
    output wire                                          in_46__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_46__m_axi_m_axi_AWSIZE,
    input wire                                           in_46__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_46__m_axi_m_axi_BID,
    input wire                                           in_46__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_46__m_axi_m_axi_BRESP,
    output wire                                          in_46__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_46__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_46__m_axi_m_axi_RID,
    output wire                                          in_46__m_axi_m_axi_RLAST,
    input wire                                           in_46__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_46__m_axi_m_axi_RRESP,
    output wire                                          in_46__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_46__m_axi_m_axi_WDATA,
    input wire                                           in_46__m_axi_m_axi_WLAST,
    output wire                                          in_46__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_46__m_axi_m_axi_WSTRB,
    input wire                                           in_46__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_46__m_axi_read_addr_din,
    input wire                                           in_46__m_axi_read_addr_full_n,
    output wire                                          in_46__m_axi_read_addr_write,
    input wire  [                                 255:0] in_46__m_axi_read_data_dout,
    input wire                                           in_46__m_axi_read_data_empty_n,
    output wire                                          in_46__m_axi_read_data_read,
    output wire                                          in_46__m_axi_rst,
    output wire [                                  63:0] in_46__m_axi_write_addr_din,
    input wire                                           in_46__m_axi_write_addr_full_n,
    output wire                                          in_46__m_axi_write_addr_write,
    output wire [                                 255:0] in_46__m_axi_write_data_din,
    input wire                                           in_46__m_axi_write_data_full_n,
    output wire                                          in_46__m_axi_write_data_write,
    input wire  [                                   7:0] in_46__m_axi_write_resp_dout,
    input wire                                           in_46__m_axi_write_resp_empty_n,
    output wire                                          in_46__m_axi_write_resp_read,
    output wire                                          in_47__m_axi_clk,
    input wire  [                                  63:0] in_47__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_47__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_47__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_47__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_47__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_47__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_47__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_47__m_axi_m_axi_ARQOS,
    output wire                                          in_47__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_47__m_axi_m_axi_ARSIZE,
    input wire                                           in_47__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_47__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_47__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_47__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_47__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_47__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_47__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_47__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_47__m_axi_m_axi_AWQOS,
    output wire                                          in_47__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_47__m_axi_m_axi_AWSIZE,
    input wire                                           in_47__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_47__m_axi_m_axi_BID,
    input wire                                           in_47__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_47__m_axi_m_axi_BRESP,
    output wire                                          in_47__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_47__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_47__m_axi_m_axi_RID,
    output wire                                          in_47__m_axi_m_axi_RLAST,
    input wire                                           in_47__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_47__m_axi_m_axi_RRESP,
    output wire                                          in_47__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_47__m_axi_m_axi_WDATA,
    input wire                                           in_47__m_axi_m_axi_WLAST,
    output wire                                          in_47__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_47__m_axi_m_axi_WSTRB,
    input wire                                           in_47__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_47__m_axi_read_addr_din,
    input wire                                           in_47__m_axi_read_addr_full_n,
    output wire                                          in_47__m_axi_read_addr_write,
    input wire  [                                 255:0] in_47__m_axi_read_data_dout,
    input wire                                           in_47__m_axi_read_data_empty_n,
    output wire                                          in_47__m_axi_read_data_read,
    output wire                                          in_47__m_axi_rst,
    output wire [                                  63:0] in_47__m_axi_write_addr_din,
    input wire                                           in_47__m_axi_write_addr_full_n,
    output wire                                          in_47__m_axi_write_addr_write,
    output wire [                                 255:0] in_47__m_axi_write_data_din,
    input wire                                           in_47__m_axi_write_data_full_n,
    output wire                                          in_47__m_axi_write_data_write,
    input wire  [                                   7:0] in_47__m_axi_write_resp_dout,
    input wire                                           in_47__m_axi_write_resp_empty_n,
    output wire                                          in_47__m_axi_write_resp_read,
    output wire                                          in_48__m_axi_clk,
    input wire  [                                  63:0] in_48__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_48__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_48__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_48__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_48__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_48__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_48__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_48__m_axi_m_axi_ARQOS,
    output wire                                          in_48__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_48__m_axi_m_axi_ARSIZE,
    input wire                                           in_48__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_48__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_48__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_48__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_48__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_48__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_48__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_48__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_48__m_axi_m_axi_AWQOS,
    output wire                                          in_48__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_48__m_axi_m_axi_AWSIZE,
    input wire                                           in_48__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_48__m_axi_m_axi_BID,
    input wire                                           in_48__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_48__m_axi_m_axi_BRESP,
    output wire                                          in_48__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_48__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_48__m_axi_m_axi_RID,
    output wire                                          in_48__m_axi_m_axi_RLAST,
    input wire                                           in_48__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_48__m_axi_m_axi_RRESP,
    output wire                                          in_48__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_48__m_axi_m_axi_WDATA,
    input wire                                           in_48__m_axi_m_axi_WLAST,
    output wire                                          in_48__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_48__m_axi_m_axi_WSTRB,
    input wire                                           in_48__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_48__m_axi_read_addr_din,
    input wire                                           in_48__m_axi_read_addr_full_n,
    output wire                                          in_48__m_axi_read_addr_write,
    input wire  [                                 255:0] in_48__m_axi_read_data_dout,
    input wire                                           in_48__m_axi_read_data_empty_n,
    output wire                                          in_48__m_axi_read_data_read,
    output wire                                          in_48__m_axi_rst,
    output wire [                                  63:0] in_48__m_axi_write_addr_din,
    input wire                                           in_48__m_axi_write_addr_full_n,
    output wire                                          in_48__m_axi_write_addr_write,
    output wire [                                 255:0] in_48__m_axi_write_data_din,
    input wire                                           in_48__m_axi_write_data_full_n,
    output wire                                          in_48__m_axi_write_data_write,
    input wire  [                                   7:0] in_48__m_axi_write_resp_dout,
    input wire                                           in_48__m_axi_write_resp_empty_n,
    output wire                                          in_48__m_axi_write_resp_read,
    output wire                                          in_49__m_axi_clk,
    input wire  [                                  63:0] in_49__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_49__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_49__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_49__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_49__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_49__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_49__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_49__m_axi_m_axi_ARQOS,
    output wire                                          in_49__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_49__m_axi_m_axi_ARSIZE,
    input wire                                           in_49__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_49__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_49__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_49__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_49__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_49__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_49__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_49__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_49__m_axi_m_axi_AWQOS,
    output wire                                          in_49__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_49__m_axi_m_axi_AWSIZE,
    input wire                                           in_49__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_49__m_axi_m_axi_BID,
    input wire                                           in_49__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_49__m_axi_m_axi_BRESP,
    output wire                                          in_49__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_49__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_49__m_axi_m_axi_RID,
    output wire                                          in_49__m_axi_m_axi_RLAST,
    input wire                                           in_49__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_49__m_axi_m_axi_RRESP,
    output wire                                          in_49__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_49__m_axi_m_axi_WDATA,
    input wire                                           in_49__m_axi_m_axi_WLAST,
    output wire                                          in_49__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_49__m_axi_m_axi_WSTRB,
    input wire                                           in_49__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_49__m_axi_read_addr_din,
    input wire                                           in_49__m_axi_read_addr_full_n,
    output wire                                          in_49__m_axi_read_addr_write,
    input wire  [                                 255:0] in_49__m_axi_read_data_dout,
    input wire                                           in_49__m_axi_read_data_empty_n,
    output wire                                          in_49__m_axi_read_data_read,
    output wire                                          in_49__m_axi_rst,
    output wire [                                  63:0] in_49__m_axi_write_addr_din,
    input wire                                           in_49__m_axi_write_addr_full_n,
    output wire                                          in_49__m_axi_write_addr_write,
    output wire [                                 255:0] in_49__m_axi_write_data_din,
    input wire                                           in_49__m_axi_write_data_full_n,
    output wire                                          in_49__m_axi_write_data_write,
    input wire  [                                   7:0] in_49__m_axi_write_resp_dout,
    input wire                                           in_49__m_axi_write_resp_empty_n,
    output wire                                          in_49__m_axi_write_resp_read,
    output wire                                          in_5__m_axi_clk,
    input wire  [                                  63:0] in_5__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_5__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_5__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_5__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_5__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_5__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_5__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_5__m_axi_m_axi_ARQOS,
    output wire                                          in_5__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_5__m_axi_m_axi_ARSIZE,
    input wire                                           in_5__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_5__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_5__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_5__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_5__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_5__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_5__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_5__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_5__m_axi_m_axi_AWQOS,
    output wire                                          in_5__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_5__m_axi_m_axi_AWSIZE,
    input wire                                           in_5__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_5__m_axi_m_axi_BID,
    input wire                                           in_5__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_5__m_axi_m_axi_BRESP,
    output wire                                          in_5__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_5__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_5__m_axi_m_axi_RID,
    output wire                                          in_5__m_axi_m_axi_RLAST,
    input wire                                           in_5__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_5__m_axi_m_axi_RRESP,
    output wire                                          in_5__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_5__m_axi_m_axi_WDATA,
    input wire                                           in_5__m_axi_m_axi_WLAST,
    output wire                                          in_5__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_5__m_axi_m_axi_WSTRB,
    input wire                                           in_5__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_5__m_axi_read_addr_din,
    input wire                                           in_5__m_axi_read_addr_full_n,
    output wire                                          in_5__m_axi_read_addr_write,
    input wire  [                                 255:0] in_5__m_axi_read_data_dout,
    input wire                                           in_5__m_axi_read_data_empty_n,
    output wire                                          in_5__m_axi_read_data_read,
    output wire                                          in_5__m_axi_rst,
    output wire [                                  63:0] in_5__m_axi_write_addr_din,
    input wire                                           in_5__m_axi_write_addr_full_n,
    output wire                                          in_5__m_axi_write_addr_write,
    output wire [                                 255:0] in_5__m_axi_write_data_din,
    input wire                                           in_5__m_axi_write_data_full_n,
    output wire                                          in_5__m_axi_write_data_write,
    input wire  [                                   7:0] in_5__m_axi_write_resp_dout,
    input wire                                           in_5__m_axi_write_resp_empty_n,
    output wire                                          in_5__m_axi_write_resp_read,
    output wire                                          in_50__m_axi_clk,
    input wire  [                                  63:0] in_50__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_50__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_50__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_50__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_50__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_50__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_50__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_50__m_axi_m_axi_ARQOS,
    output wire                                          in_50__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_50__m_axi_m_axi_ARSIZE,
    input wire                                           in_50__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_50__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_50__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_50__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_50__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_50__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_50__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_50__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_50__m_axi_m_axi_AWQOS,
    output wire                                          in_50__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_50__m_axi_m_axi_AWSIZE,
    input wire                                           in_50__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_50__m_axi_m_axi_BID,
    input wire                                           in_50__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_50__m_axi_m_axi_BRESP,
    output wire                                          in_50__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_50__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_50__m_axi_m_axi_RID,
    output wire                                          in_50__m_axi_m_axi_RLAST,
    input wire                                           in_50__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_50__m_axi_m_axi_RRESP,
    output wire                                          in_50__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_50__m_axi_m_axi_WDATA,
    input wire                                           in_50__m_axi_m_axi_WLAST,
    output wire                                          in_50__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_50__m_axi_m_axi_WSTRB,
    input wire                                           in_50__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_50__m_axi_read_addr_din,
    input wire                                           in_50__m_axi_read_addr_full_n,
    output wire                                          in_50__m_axi_read_addr_write,
    input wire  [                                 255:0] in_50__m_axi_read_data_dout,
    input wire                                           in_50__m_axi_read_data_empty_n,
    output wire                                          in_50__m_axi_read_data_read,
    output wire                                          in_50__m_axi_rst,
    output wire [                                  63:0] in_50__m_axi_write_addr_din,
    input wire                                           in_50__m_axi_write_addr_full_n,
    output wire                                          in_50__m_axi_write_addr_write,
    output wire [                                 255:0] in_50__m_axi_write_data_din,
    input wire                                           in_50__m_axi_write_data_full_n,
    output wire                                          in_50__m_axi_write_data_write,
    input wire  [                                   7:0] in_50__m_axi_write_resp_dout,
    input wire                                           in_50__m_axi_write_resp_empty_n,
    output wire                                          in_50__m_axi_write_resp_read,
    output wire                                          in_51__m_axi_clk,
    input wire  [                                  63:0] in_51__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_51__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_51__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_51__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_51__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_51__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_51__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_51__m_axi_m_axi_ARQOS,
    output wire                                          in_51__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_51__m_axi_m_axi_ARSIZE,
    input wire                                           in_51__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_51__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_51__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_51__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_51__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_51__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_51__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_51__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_51__m_axi_m_axi_AWQOS,
    output wire                                          in_51__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_51__m_axi_m_axi_AWSIZE,
    input wire                                           in_51__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_51__m_axi_m_axi_BID,
    input wire                                           in_51__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_51__m_axi_m_axi_BRESP,
    output wire                                          in_51__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_51__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_51__m_axi_m_axi_RID,
    output wire                                          in_51__m_axi_m_axi_RLAST,
    input wire                                           in_51__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_51__m_axi_m_axi_RRESP,
    output wire                                          in_51__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_51__m_axi_m_axi_WDATA,
    input wire                                           in_51__m_axi_m_axi_WLAST,
    output wire                                          in_51__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_51__m_axi_m_axi_WSTRB,
    input wire                                           in_51__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_51__m_axi_read_addr_din,
    input wire                                           in_51__m_axi_read_addr_full_n,
    output wire                                          in_51__m_axi_read_addr_write,
    input wire  [                                 255:0] in_51__m_axi_read_data_dout,
    input wire                                           in_51__m_axi_read_data_empty_n,
    output wire                                          in_51__m_axi_read_data_read,
    output wire                                          in_51__m_axi_rst,
    output wire [                                  63:0] in_51__m_axi_write_addr_din,
    input wire                                           in_51__m_axi_write_addr_full_n,
    output wire                                          in_51__m_axi_write_addr_write,
    output wire [                                 255:0] in_51__m_axi_write_data_din,
    input wire                                           in_51__m_axi_write_data_full_n,
    output wire                                          in_51__m_axi_write_data_write,
    input wire  [                                   7:0] in_51__m_axi_write_resp_dout,
    input wire                                           in_51__m_axi_write_resp_empty_n,
    output wire                                          in_51__m_axi_write_resp_read,
    output wire                                          in_52__m_axi_clk,
    input wire  [                                  63:0] in_52__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_52__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_52__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_52__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_52__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_52__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_52__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_52__m_axi_m_axi_ARQOS,
    output wire                                          in_52__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_52__m_axi_m_axi_ARSIZE,
    input wire                                           in_52__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_52__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_52__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_52__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_52__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_52__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_52__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_52__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_52__m_axi_m_axi_AWQOS,
    output wire                                          in_52__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_52__m_axi_m_axi_AWSIZE,
    input wire                                           in_52__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_52__m_axi_m_axi_BID,
    input wire                                           in_52__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_52__m_axi_m_axi_BRESP,
    output wire                                          in_52__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_52__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_52__m_axi_m_axi_RID,
    output wire                                          in_52__m_axi_m_axi_RLAST,
    input wire                                           in_52__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_52__m_axi_m_axi_RRESP,
    output wire                                          in_52__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_52__m_axi_m_axi_WDATA,
    input wire                                           in_52__m_axi_m_axi_WLAST,
    output wire                                          in_52__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_52__m_axi_m_axi_WSTRB,
    input wire                                           in_52__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_52__m_axi_read_addr_din,
    input wire                                           in_52__m_axi_read_addr_full_n,
    output wire                                          in_52__m_axi_read_addr_write,
    input wire  [                                 255:0] in_52__m_axi_read_data_dout,
    input wire                                           in_52__m_axi_read_data_empty_n,
    output wire                                          in_52__m_axi_read_data_read,
    output wire                                          in_52__m_axi_rst,
    output wire [                                  63:0] in_52__m_axi_write_addr_din,
    input wire                                           in_52__m_axi_write_addr_full_n,
    output wire                                          in_52__m_axi_write_addr_write,
    output wire [                                 255:0] in_52__m_axi_write_data_din,
    input wire                                           in_52__m_axi_write_data_full_n,
    output wire                                          in_52__m_axi_write_data_write,
    input wire  [                                   7:0] in_52__m_axi_write_resp_dout,
    input wire                                           in_52__m_axi_write_resp_empty_n,
    output wire                                          in_52__m_axi_write_resp_read,
    output wire                                          in_53__m_axi_clk,
    input wire  [                                  63:0] in_53__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_53__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_53__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_53__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_53__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_53__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_53__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_53__m_axi_m_axi_ARQOS,
    output wire                                          in_53__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_53__m_axi_m_axi_ARSIZE,
    input wire                                           in_53__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_53__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_53__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_53__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_53__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_53__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_53__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_53__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_53__m_axi_m_axi_AWQOS,
    output wire                                          in_53__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_53__m_axi_m_axi_AWSIZE,
    input wire                                           in_53__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_53__m_axi_m_axi_BID,
    input wire                                           in_53__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_53__m_axi_m_axi_BRESP,
    output wire                                          in_53__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_53__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_53__m_axi_m_axi_RID,
    output wire                                          in_53__m_axi_m_axi_RLAST,
    input wire                                           in_53__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_53__m_axi_m_axi_RRESP,
    output wire                                          in_53__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_53__m_axi_m_axi_WDATA,
    input wire                                           in_53__m_axi_m_axi_WLAST,
    output wire                                          in_53__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_53__m_axi_m_axi_WSTRB,
    input wire                                           in_53__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_53__m_axi_read_addr_din,
    input wire                                           in_53__m_axi_read_addr_full_n,
    output wire                                          in_53__m_axi_read_addr_write,
    input wire  [                                 255:0] in_53__m_axi_read_data_dout,
    input wire                                           in_53__m_axi_read_data_empty_n,
    output wire                                          in_53__m_axi_read_data_read,
    output wire                                          in_53__m_axi_rst,
    output wire [                                  63:0] in_53__m_axi_write_addr_din,
    input wire                                           in_53__m_axi_write_addr_full_n,
    output wire                                          in_53__m_axi_write_addr_write,
    output wire [                                 255:0] in_53__m_axi_write_data_din,
    input wire                                           in_53__m_axi_write_data_full_n,
    output wire                                          in_53__m_axi_write_data_write,
    input wire  [                                   7:0] in_53__m_axi_write_resp_dout,
    input wire                                           in_53__m_axi_write_resp_empty_n,
    output wire                                          in_53__m_axi_write_resp_read,
    output wire                                          in_6__m_axi_clk,
    input wire  [                                  63:0] in_6__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_6__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_6__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_6__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_6__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_6__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_6__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_6__m_axi_m_axi_ARQOS,
    output wire                                          in_6__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_6__m_axi_m_axi_ARSIZE,
    input wire                                           in_6__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_6__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_6__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_6__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_6__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_6__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_6__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_6__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_6__m_axi_m_axi_AWQOS,
    output wire                                          in_6__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_6__m_axi_m_axi_AWSIZE,
    input wire                                           in_6__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_6__m_axi_m_axi_BID,
    input wire                                           in_6__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_6__m_axi_m_axi_BRESP,
    output wire                                          in_6__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_6__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_6__m_axi_m_axi_RID,
    output wire                                          in_6__m_axi_m_axi_RLAST,
    input wire                                           in_6__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_6__m_axi_m_axi_RRESP,
    output wire                                          in_6__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_6__m_axi_m_axi_WDATA,
    input wire                                           in_6__m_axi_m_axi_WLAST,
    output wire                                          in_6__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_6__m_axi_m_axi_WSTRB,
    input wire                                           in_6__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_6__m_axi_read_addr_din,
    input wire                                           in_6__m_axi_read_addr_full_n,
    output wire                                          in_6__m_axi_read_addr_write,
    input wire  [                                 255:0] in_6__m_axi_read_data_dout,
    input wire                                           in_6__m_axi_read_data_empty_n,
    output wire                                          in_6__m_axi_read_data_read,
    output wire                                          in_6__m_axi_rst,
    output wire [                                  63:0] in_6__m_axi_write_addr_din,
    input wire                                           in_6__m_axi_write_addr_full_n,
    output wire                                          in_6__m_axi_write_addr_write,
    output wire [                                 255:0] in_6__m_axi_write_data_din,
    input wire                                           in_6__m_axi_write_data_full_n,
    output wire                                          in_6__m_axi_write_data_write,
    input wire  [                                   7:0] in_6__m_axi_write_resp_dout,
    input wire                                           in_6__m_axi_write_resp_empty_n,
    output wire                                          in_6__m_axi_write_resp_read,
    output wire                                          in_7__m_axi_clk,
    input wire  [                                  63:0] in_7__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_7__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_7__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_7__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_7__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_7__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_7__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_7__m_axi_m_axi_ARQOS,
    output wire                                          in_7__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_7__m_axi_m_axi_ARSIZE,
    input wire                                           in_7__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_7__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_7__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_7__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_7__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_7__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_7__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_7__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_7__m_axi_m_axi_AWQOS,
    output wire                                          in_7__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_7__m_axi_m_axi_AWSIZE,
    input wire                                           in_7__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_7__m_axi_m_axi_BID,
    input wire                                           in_7__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_7__m_axi_m_axi_BRESP,
    output wire                                          in_7__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_7__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_7__m_axi_m_axi_RID,
    output wire                                          in_7__m_axi_m_axi_RLAST,
    input wire                                           in_7__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_7__m_axi_m_axi_RRESP,
    output wire                                          in_7__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_7__m_axi_m_axi_WDATA,
    input wire                                           in_7__m_axi_m_axi_WLAST,
    output wire                                          in_7__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_7__m_axi_m_axi_WSTRB,
    input wire                                           in_7__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_7__m_axi_read_addr_din,
    input wire                                           in_7__m_axi_read_addr_full_n,
    output wire                                          in_7__m_axi_read_addr_write,
    input wire  [                                 255:0] in_7__m_axi_read_data_dout,
    input wire                                           in_7__m_axi_read_data_empty_n,
    output wire                                          in_7__m_axi_read_data_read,
    output wire                                          in_7__m_axi_rst,
    output wire [                                  63:0] in_7__m_axi_write_addr_din,
    input wire                                           in_7__m_axi_write_addr_full_n,
    output wire                                          in_7__m_axi_write_addr_write,
    output wire [                                 255:0] in_7__m_axi_write_data_din,
    input wire                                           in_7__m_axi_write_data_full_n,
    output wire                                          in_7__m_axi_write_data_write,
    input wire  [                                   7:0] in_7__m_axi_write_resp_dout,
    input wire                                           in_7__m_axi_write_resp_empty_n,
    output wire                                          in_7__m_axi_write_resp_read,
    output wire                                          in_8__m_axi_clk,
    input wire  [                                  63:0] in_8__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_8__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_8__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_8__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_8__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_8__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_8__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_8__m_axi_m_axi_ARQOS,
    output wire                                          in_8__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_8__m_axi_m_axi_ARSIZE,
    input wire                                           in_8__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_8__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_8__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_8__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_8__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_8__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_8__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_8__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_8__m_axi_m_axi_AWQOS,
    output wire                                          in_8__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_8__m_axi_m_axi_AWSIZE,
    input wire                                           in_8__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_8__m_axi_m_axi_BID,
    input wire                                           in_8__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_8__m_axi_m_axi_BRESP,
    output wire                                          in_8__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_8__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_8__m_axi_m_axi_RID,
    output wire                                          in_8__m_axi_m_axi_RLAST,
    input wire                                           in_8__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_8__m_axi_m_axi_RRESP,
    output wire                                          in_8__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_8__m_axi_m_axi_WDATA,
    input wire                                           in_8__m_axi_m_axi_WLAST,
    output wire                                          in_8__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_8__m_axi_m_axi_WSTRB,
    input wire                                           in_8__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_8__m_axi_read_addr_din,
    input wire                                           in_8__m_axi_read_addr_full_n,
    output wire                                          in_8__m_axi_read_addr_write,
    input wire  [                                 255:0] in_8__m_axi_read_data_dout,
    input wire                                           in_8__m_axi_read_data_empty_n,
    output wire                                          in_8__m_axi_read_data_read,
    output wire                                          in_8__m_axi_rst,
    output wire [                                  63:0] in_8__m_axi_write_addr_din,
    input wire                                           in_8__m_axi_write_addr_full_n,
    output wire                                          in_8__m_axi_write_addr_write,
    output wire [                                 255:0] in_8__m_axi_write_data_din,
    input wire                                           in_8__m_axi_write_data_full_n,
    output wire                                          in_8__m_axi_write_data_write,
    input wire  [                                   7:0] in_8__m_axi_write_resp_dout,
    input wire                                           in_8__m_axi_write_resp_empty_n,
    output wire                                          in_8__m_axi_write_resp_read,
    output wire                                          in_9__m_axi_clk,
    input wire  [                                  63:0] in_9__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_9__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_9__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_9__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_9__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_9__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_9__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_9__m_axi_m_axi_ARQOS,
    output wire                                          in_9__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_9__m_axi_m_axi_ARSIZE,
    input wire                                           in_9__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_9__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_9__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_9__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_9__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_9__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_9__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_9__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_9__m_axi_m_axi_AWQOS,
    output wire                                          in_9__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_9__m_axi_m_axi_AWSIZE,
    input wire                                           in_9__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_9__m_axi_m_axi_BID,
    input wire                                           in_9__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_9__m_axi_m_axi_BRESP,
    output wire                                          in_9__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_9__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_9__m_axi_m_axi_RID,
    output wire                                          in_9__m_axi_m_axi_RLAST,
    input wire                                           in_9__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_9__m_axi_m_axi_RRESP,
    output wire                                          in_9__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_9__m_axi_m_axi_WDATA,
    input wire                                           in_9__m_axi_m_axi_WLAST,
    output wire                                          in_9__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_9__m_axi_m_axi_WSTRB,
    input wire                                           in_9__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_9__m_axi_read_addr_din,
    input wire                                           in_9__m_axi_read_addr_full_n,
    output wire                                          in_9__m_axi_read_addr_write,
    input wire  [                                 255:0] in_9__m_axi_read_data_dout,
    input wire                                           in_9__m_axi_read_data_empty_n,
    output wire                                          in_9__m_axi_read_data_read,
    output wire                                          in_9__m_axi_rst,
    output wire [                                  63:0] in_9__m_axi_write_addr_din,
    input wire                                           in_9__m_axi_write_addr_full_n,
    output wire                                          in_9__m_axi_write_addr_write,
    output wire [                                 255:0] in_9__m_axi_write_data_din,
    input wire                                           in_9__m_axi_write_data_full_n,
    output wire                                          in_9__m_axi_write_data_write,
    input wire  [                                   7:0] in_9__m_axi_write_resp_dout,
    input wire                                           in_9__m_axi_write_resp_empty_n,
    output wire                                          in_9__m_axi_write_resp_read,
    output wire [                                  63:0] __tapa_fsm_unit_L4_out_dist,
    output wire [                                  63:0] __tapa_fsm_unit_L4_out_id,
    output wire                                          __tapa_fsm_unit_ap_clk,
    input wire                                           __tapa_fsm_unit_ap_done,
    input wire                                           __tapa_fsm_unit_ap_idle,
    input wire                                           __tapa_fsm_unit_ap_ready,
    output wire                                          __tapa_fsm_unit_ap_rst_n,
    output wire                                          __tapa_fsm_unit_ap_start,
    output wire [                                  63:0] __tapa_fsm_unit_in_0,
    output wire [                                  63:0] __tapa_fsm_unit_in_1,
    output wire [                                  63:0] __tapa_fsm_unit_in_10,
    output wire [                                  63:0] __tapa_fsm_unit_in_11,
    output wire [                                  63:0] __tapa_fsm_unit_in_12,
    output wire [                                  63:0] __tapa_fsm_unit_in_13,
    output wire [                                  63:0] __tapa_fsm_unit_in_14,
    output wire [                                  63:0] __tapa_fsm_unit_in_15,
    output wire [                                  63:0] __tapa_fsm_unit_in_16,
    output wire [                                  63:0] __tapa_fsm_unit_in_17,
    output wire [                                  63:0] __tapa_fsm_unit_in_18,
    output wire [                                  63:0] __tapa_fsm_unit_in_19,
    output wire [                                  63:0] __tapa_fsm_unit_in_2,
    output wire [                                  63:0] __tapa_fsm_unit_in_20,
    output wire [                                  63:0] __tapa_fsm_unit_in_21,
    output wire [                                  63:0] __tapa_fsm_unit_in_22,
    output wire [                                  63:0] __tapa_fsm_unit_in_23,
    output wire [                                  63:0] __tapa_fsm_unit_in_24,
    output wire [                                  63:0] __tapa_fsm_unit_in_25,
    output wire [                                  63:0] __tapa_fsm_unit_in_26,
    output wire [                                  63:0] __tapa_fsm_unit_in_27,
    output wire [                                  63:0] __tapa_fsm_unit_in_28,
    output wire [                                  63:0] __tapa_fsm_unit_in_29,
    output wire [                                  63:0] __tapa_fsm_unit_in_3,
    output wire [                                  63:0] __tapa_fsm_unit_in_30,
    output wire [                                  63:0] __tapa_fsm_unit_in_31,
    output wire [                                  63:0] __tapa_fsm_unit_in_32,
    output wire [                                  63:0] __tapa_fsm_unit_in_33,
    output wire [                                  63:0] __tapa_fsm_unit_in_34,
    output wire [                                  63:0] __tapa_fsm_unit_in_35,
    output wire [                                  63:0] __tapa_fsm_unit_in_36,
    output wire [                                  63:0] __tapa_fsm_unit_in_37,
    output wire [                                  63:0] __tapa_fsm_unit_in_38,
    output wire [                                  63:0] __tapa_fsm_unit_in_39,
    output wire [                                  63:0] __tapa_fsm_unit_in_4,
    output wire [                                  63:0] __tapa_fsm_unit_in_40,
    output wire [                                  63:0] __tapa_fsm_unit_in_41,
    output wire [                                  63:0] __tapa_fsm_unit_in_42,
    output wire [                                  63:0] __tapa_fsm_unit_in_43,
    output wire [                                  63:0] __tapa_fsm_unit_in_44,
    output wire [                                  63:0] __tapa_fsm_unit_in_45,
    output wire [                                  63:0] __tapa_fsm_unit_in_46,
    output wire [                                  63:0] __tapa_fsm_unit_in_47,
    output wire [                                  63:0] __tapa_fsm_unit_in_48,
    output wire [                                  63:0] __tapa_fsm_unit_in_49,
    output wire [                                  63:0] __tapa_fsm_unit_in_5,
    output wire [                                  63:0] __tapa_fsm_unit_in_50,
    output wire [                                  63:0] __tapa_fsm_unit_in_51,
    output wire [                                  63:0] __tapa_fsm_unit_in_52,
    output wire [                                  63:0] __tapa_fsm_unit_in_53,
    output wire [                                  63:0] __tapa_fsm_unit_in_6,
    output wire [                                  63:0] __tapa_fsm_unit_in_7,
    output wire [                                  63:0] __tapa_fsm_unit_in_8,
    output wire [                                  63:0] __tapa_fsm_unit_in_9,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_globalSort_L1_L2_0__ap_start,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_10__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_10__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_10__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_globalSort_L1_L2_10__ap_start,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_11__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_11__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_11__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_globalSort_L1_L2_11__ap_start,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_12__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_12__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_12__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_globalSort_L1_L2_12__ap_start,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_13__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_13__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_13__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_globalSort_L1_L2_13__ap_start,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_14__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_14__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_14__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_globalSort_L1_L2_14__ap_start,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_15__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_15__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_15__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_globalSort_L1_L2_15__ap_start,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_16__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_16__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_16__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_globalSort_L1_L2_16__ap_start,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_17__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_17__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_17__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_globalSort_L1_L2_17__ap_start,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_18__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_18__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_18__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_globalSort_L1_L2_18__ap_start,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_19__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_19__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_19__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_globalSort_L1_L2_19__ap_start,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_1__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_1__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_1__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_globalSort_L1_L2_1__ap_start,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_20__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_20__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_20__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_globalSort_L1_L2_20__ap_start,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_21__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_21__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_21__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_globalSort_L1_L2_21__ap_start,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_22__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_22__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_22__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_globalSort_L1_L2_22__ap_start,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_23__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_23__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_23__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_globalSort_L1_L2_23__ap_start,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_24__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_24__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_24__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_globalSort_L1_L2_24__ap_start,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_25__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_25__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_25__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_globalSort_L1_L2_25__ap_start,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_2__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_2__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_2__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_globalSort_L1_L2_2__ap_start,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_3__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_3__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_3__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_globalSort_L1_L2_3__ap_start,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_4__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_4__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_4__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_globalSort_L1_L2_4__ap_start,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_5__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_5__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_5__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_globalSort_L1_L2_5__ap_start,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_6__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_6__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_6__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_globalSort_L1_L2_6__ap_start,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_7__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_7__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_7__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_globalSort_L1_L2_7__ap_start,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_8__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_8__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_8__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_globalSort_L1_L2_8__ap_start,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_9__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_9__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_9__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_globalSort_L1_L2_9__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_globalSort_L3_0___L4_out_dist__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_globalSort_L3_0___L4_out_id__q0,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L3_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L3_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L3_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_globalSort_L3_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_0_0___in_0__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_0_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_0_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_0_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_0_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_10_0___in_10__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_10_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_10_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_10_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_10_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_11_0___in_11__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_11_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_11_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_11_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_11_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_12_0___in_12__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_12_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_12_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_12_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_12_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_13_0___in_13__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_13_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_13_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_13_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_13_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_14_0___in_14__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_14_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_14_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_14_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_14_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_15_0___in_15__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_15_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_15_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_15_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_15_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_16_0___in_16__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_16_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_16_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_16_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_16_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_17_0___in_17__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_17_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_17_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_17_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_17_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_18_0___in_18__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_18_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_18_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_18_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_18_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_19_0___in_19__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_19_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_19_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_19_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_19_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_1_0___in_1__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_1_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_1_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_1_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_1_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_20_0___in_20__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_20_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_20_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_20_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_20_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_21_0___in_21__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_21_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_21_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_21_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_21_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_22_0___in_22__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_22_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_22_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_22_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_22_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_23_0___in_23__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_23_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_23_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_23_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_23_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_24_0___in_24__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_24_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_24_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_24_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_24_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_25_0___in_25__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_25_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_25_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_25_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_25_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_26_0___in_26__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_26_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_26_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_26_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_26_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_27_0___in_27__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_27_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_27_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_27_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_27_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_28_0___in_28__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_28_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_28_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_28_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_28_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_29_0___in_29__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_29_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_29_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_29_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_29_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_2_0___in_2__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_2_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_2_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_2_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_2_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_30_0___in_30__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_30_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_30_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_30_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_30_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_31_0___in_31__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_31_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_31_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_31_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_31_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_32_0___in_32__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_32_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_32_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_32_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_32_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_33_0___in_33__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_33_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_33_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_33_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_33_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_34_0___in_34__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_34_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_34_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_34_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_34_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_35_0___in_35__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_35_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_35_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_35_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_35_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_36_0___in_36__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_36_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_36_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_36_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_36_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_37_0___in_37__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_37_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_37_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_37_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_37_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_38_0___in_38__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_38_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_38_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_38_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_38_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_39_0___in_39__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_39_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_39_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_39_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_39_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_3_0___in_3__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_3_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_3_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_3_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_3_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_40_0___in_40__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_40_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_40_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_40_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_40_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_41_0___in_41__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_41_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_41_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_41_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_41_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_42_0___in_42__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_42_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_42_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_42_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_42_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_43_0___in_43__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_43_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_43_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_43_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_43_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_44_0___in_44__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_44_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_44_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_44_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_44_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_45_0___in_45__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_45_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_45_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_45_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_45_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_46_0___in_46__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_46_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_46_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_46_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_46_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_47_0___in_47__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_47_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_47_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_47_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_47_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_48_0___in_48__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_48_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_48_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_48_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_48_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_49_0___in_49__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_49_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_49_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_49_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_49_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_4_0___in_4__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_4_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_4_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_4_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_4_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_50_0___in_50__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_50_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_50_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_50_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_50_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_51_0___in_51__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_51_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_51_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_51_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_51_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_52_0___in_52__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_52_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_52_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_52_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_52_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_53_0___in_53__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_53_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_53_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_53_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_53_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_5_0___in_5__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_5_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_5_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_5_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_5_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_6_0___in_6__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_6_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_6_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_6_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_6_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_7_0___in_7__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_7_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_7_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_7_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_7_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_8_0___in_8__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_8_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_8_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_8_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_8_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_9_0___in_9__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_9_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_9_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_9_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_9_0__ap_start
);
  wire ap_start;
  wire [63:0] in_0;
  wire [63:0] in_1;
  wire [63:0] in_2;
  wire [63:0] in_3;
  wire [63:0] in_4;
  wire [63:0] in_5;
  wire [63:0] in_6;
  wire [63:0] in_7;
  wire [63:0] in_8;
  wire [63:0] in_9;
  wire [63:0] in_10;
  wire [63:0] in_11;
  wire [63:0] in_12;
  wire [63:0] in_13;
  wire [63:0] in_14;
  wire [63:0] in_15;
  wire [63:0] in_16;
  wire [63:0] in_17;
  wire [63:0] in_18;
  wire [63:0] in_19;
  wire [63:0] in_20;
  wire [63:0] in_21;
  wire [63:0] in_22;
  wire [63:0] in_23;
  wire [63:0] in_24;
  wire [63:0] in_25;
  wire [63:0] in_26;
  wire [63:0] in_27;
  wire [63:0] in_28;
  wire [63:0] in_29;
  wire [63:0] in_30;
  wire [63:0] in_31;
  wire [63:0] in_32;
  wire [63:0] in_33;
  wire [63:0] in_34;
  wire [63:0] in_35;
  wire [63:0] in_36;
  wire [63:0] in_37;
  wire [63:0] in_38;
  wire [63:0] in_39;
  wire [63:0] in_40;
  wire [63:0] in_41;
  wire [63:0] in_42;
  wire [63:0] in_43;
  wire [63:0] in_44;
  wire [63:0] in_45;
  wire [63:0] in_46;
  wire [63:0] in_47;
  wire [63:0] in_48;
  wire [63:0] in_49;
  wire [63:0] in_50;
  wire [63:0] in_51;
  wire [63:0] in_52;
  wire [63:0] in_53;
  wire [63:0] L4_out_dist;
  wire [63:0] L4_out_id;
  wire [65:0] L1_out_dist_0__dout;
  wire L1_out_dist_0__empty_n;
  wire L1_out_dist_0__read;
  wire [65:0] L1_out_dist_0__din;
  wire L1_out_dist_0__full_n;
  wire L1_out_dist_0__write;
  wire [65:0] L1_out_dist_10__dout;
  wire L1_out_dist_10__empty_n;
  wire L1_out_dist_10__read;
  wire [65:0] L1_out_dist_10__din;
  wire L1_out_dist_10__full_n;
  wire L1_out_dist_10__write;
  wire [65:0] L1_out_dist_11__dout;
  wire L1_out_dist_11__empty_n;
  wire L1_out_dist_11__read;
  wire [65:0] L1_out_dist_11__din;
  wire L1_out_dist_11__full_n;
  wire L1_out_dist_11__write;
  wire [65:0] L1_out_dist_12__dout;
  wire L1_out_dist_12__empty_n;
  wire L1_out_dist_12__read;
  wire [65:0] L1_out_dist_12__din;
  wire L1_out_dist_12__full_n;
  wire L1_out_dist_12__write;
  wire [65:0] L1_out_dist_13__dout;
  wire L1_out_dist_13__empty_n;
  wire L1_out_dist_13__read;
  wire [65:0] L1_out_dist_13__din;
  wire L1_out_dist_13__full_n;
  wire L1_out_dist_13__write;
  wire [65:0] L1_out_dist_14__dout;
  wire L1_out_dist_14__empty_n;
  wire L1_out_dist_14__read;
  wire [65:0] L1_out_dist_14__din;
  wire L1_out_dist_14__full_n;
  wire L1_out_dist_14__write;
  wire [65:0] L1_out_dist_15__dout;
  wire L1_out_dist_15__empty_n;
  wire L1_out_dist_15__read;
  wire [65:0] L1_out_dist_15__din;
  wire L1_out_dist_15__full_n;
  wire L1_out_dist_15__write;
  wire [65:0] L1_out_dist_16__dout;
  wire L1_out_dist_16__empty_n;
  wire L1_out_dist_16__read;
  wire [65:0] L1_out_dist_16__din;
  wire L1_out_dist_16__full_n;
  wire L1_out_dist_16__write;
  wire [65:0] L1_out_dist_17__dout;
  wire L1_out_dist_17__empty_n;
  wire L1_out_dist_17__read;
  wire [65:0] L1_out_dist_17__din;
  wire L1_out_dist_17__full_n;
  wire L1_out_dist_17__write;
  wire [65:0] L1_out_dist_1__dout;
  wire L1_out_dist_1__empty_n;
  wire L1_out_dist_1__read;
  wire [65:0] L1_out_dist_1__din;
  wire L1_out_dist_1__full_n;
  wire L1_out_dist_1__write;
  wire [65:0] L1_out_dist_2__dout;
  wire L1_out_dist_2__empty_n;
  wire L1_out_dist_2__read;
  wire [65:0] L1_out_dist_2__din;
  wire L1_out_dist_2__full_n;
  wire L1_out_dist_2__write;
  wire [65:0] L1_out_dist_3__dout;
  wire L1_out_dist_3__empty_n;
  wire L1_out_dist_3__read;
  wire [65:0] L1_out_dist_3__din;
  wire L1_out_dist_3__full_n;
  wire L1_out_dist_3__write;
  wire [65:0] L1_out_dist_4__dout;
  wire L1_out_dist_4__empty_n;
  wire L1_out_dist_4__read;
  wire [65:0] L1_out_dist_4__din;
  wire L1_out_dist_4__full_n;
  wire L1_out_dist_4__write;
  wire [65:0] L1_out_dist_5__dout;
  wire L1_out_dist_5__empty_n;
  wire L1_out_dist_5__read;
  wire [65:0] L1_out_dist_5__din;
  wire L1_out_dist_5__full_n;
  wire L1_out_dist_5__write;
  wire [65:0] L1_out_dist_6__dout;
  wire L1_out_dist_6__empty_n;
  wire L1_out_dist_6__read;
  wire [65:0] L1_out_dist_6__din;
  wire L1_out_dist_6__full_n;
  wire L1_out_dist_6__write;
  wire [65:0] L1_out_dist_7__dout;
  wire L1_out_dist_7__empty_n;
  wire L1_out_dist_7__read;
  wire [65:0] L1_out_dist_7__din;
  wire L1_out_dist_7__full_n;
  wire L1_out_dist_7__write;
  wire [65:0] L1_out_dist_8__dout;
  wire L1_out_dist_8__empty_n;
  wire L1_out_dist_8__read;
  wire [65:0] L1_out_dist_8__din;
  wire L1_out_dist_8__full_n;
  wire L1_out_dist_8__write;
  wire [65:0] L1_out_dist_9__dout;
  wire L1_out_dist_9__empty_n;
  wire L1_out_dist_9__read;
  wire [65:0] L1_out_dist_9__din;
  wire L1_out_dist_9__full_n;
  wire L1_out_dist_9__write;
  wire [65:0] L1_out_id_0__dout;
  wire L1_out_id_0__empty_n;
  wire L1_out_id_0__read;
  wire [65:0] L1_out_id_0__din;
  wire L1_out_id_0__full_n;
  wire L1_out_id_0__write;
  wire [65:0] L1_out_id_10__dout;
  wire L1_out_id_10__empty_n;
  wire L1_out_id_10__read;
  wire [65:0] L1_out_id_10__din;
  wire L1_out_id_10__full_n;
  wire L1_out_id_10__write;
  wire [65:0] L1_out_id_11__dout;
  wire L1_out_id_11__empty_n;
  wire L1_out_id_11__read;
  wire [65:0] L1_out_id_11__din;
  wire L1_out_id_11__full_n;
  wire L1_out_id_11__write;
  wire [65:0] L1_out_id_12__dout;
  wire L1_out_id_12__empty_n;
  wire L1_out_id_12__read;
  wire [65:0] L1_out_id_12__din;
  wire L1_out_id_12__full_n;
  wire L1_out_id_12__write;
  wire [65:0] L1_out_id_13__dout;
  wire L1_out_id_13__empty_n;
  wire L1_out_id_13__read;
  wire [65:0] L1_out_id_13__din;
  wire L1_out_id_13__full_n;
  wire L1_out_id_13__write;
  wire [65:0] L1_out_id_14__dout;
  wire L1_out_id_14__empty_n;
  wire L1_out_id_14__read;
  wire [65:0] L1_out_id_14__din;
  wire L1_out_id_14__full_n;
  wire L1_out_id_14__write;
  wire [65:0] L1_out_id_15__dout;
  wire L1_out_id_15__empty_n;
  wire L1_out_id_15__read;
  wire [65:0] L1_out_id_15__din;
  wire L1_out_id_15__full_n;
  wire L1_out_id_15__write;
  wire [65:0] L1_out_id_16__dout;
  wire L1_out_id_16__empty_n;
  wire L1_out_id_16__read;
  wire [65:0] L1_out_id_16__din;
  wire L1_out_id_16__full_n;
  wire L1_out_id_16__write;
  wire [65:0] L1_out_id_17__dout;
  wire L1_out_id_17__empty_n;
  wire L1_out_id_17__read;
  wire [65:0] L1_out_id_17__din;
  wire L1_out_id_17__full_n;
  wire L1_out_id_17__write;
  wire [65:0] L1_out_id_1__dout;
  wire L1_out_id_1__empty_n;
  wire L1_out_id_1__read;
  wire [65:0] L1_out_id_1__din;
  wire L1_out_id_1__full_n;
  wire L1_out_id_1__write;
  wire [65:0] L1_out_id_2__dout;
  wire L1_out_id_2__empty_n;
  wire L1_out_id_2__read;
  wire [65:0] L1_out_id_2__din;
  wire L1_out_id_2__full_n;
  wire L1_out_id_2__write;
  wire [65:0] L1_out_id_3__dout;
  wire L1_out_id_3__empty_n;
  wire L1_out_id_3__read;
  wire [65:0] L1_out_id_3__din;
  wire L1_out_id_3__full_n;
  wire L1_out_id_3__write;
  wire [65:0] L1_out_id_4__dout;
  wire L1_out_id_4__empty_n;
  wire L1_out_id_4__read;
  wire [65:0] L1_out_id_4__din;
  wire L1_out_id_4__full_n;
  wire L1_out_id_4__write;
  wire [65:0] L1_out_id_5__dout;
  wire L1_out_id_5__empty_n;
  wire L1_out_id_5__read;
  wire [65:0] L1_out_id_5__din;
  wire L1_out_id_5__full_n;
  wire L1_out_id_5__write;
  wire [65:0] L1_out_id_6__dout;
  wire L1_out_id_6__empty_n;
  wire L1_out_id_6__read;
  wire [65:0] L1_out_id_6__din;
  wire L1_out_id_6__full_n;
  wire L1_out_id_6__write;
  wire [65:0] L1_out_id_7__dout;
  wire L1_out_id_7__empty_n;
  wire L1_out_id_7__read;
  wire [65:0] L1_out_id_7__din;
  wire L1_out_id_7__full_n;
  wire L1_out_id_7__write;
  wire [65:0] L1_out_id_8__dout;
  wire L1_out_id_8__empty_n;
  wire L1_out_id_8__read;
  wire [65:0] L1_out_id_8__din;
  wire L1_out_id_8__full_n;
  wire L1_out_id_8__write;
  wire [65:0] L1_out_id_9__dout;
  wire L1_out_id_9__empty_n;
  wire L1_out_id_9__read;
  wire [65:0] L1_out_id_9__din;
  wire L1_out_id_9__full_n;
  wire L1_out_id_9__write;
  wire [65:0] L2_out_dist0__dout;
  wire L2_out_dist0__empty_n;
  wire L2_out_dist0__read;
  wire [65:0] L2_out_dist0__din;
  wire L2_out_dist0__full_n;
  wire L2_out_dist0__write;
  wire [65:0] L2_out_dist1__dout;
  wire L2_out_dist1__empty_n;
  wire L2_out_dist1__read;
  wire [65:0] L2_out_dist1__din;
  wire L2_out_dist1__full_n;
  wire L2_out_dist1__write;
  wire [65:0] L2_out_dist2__dout;
  wire L2_out_dist2__empty_n;
  wire L2_out_dist2__read;
  wire [65:0] L2_out_dist2__din;
  wire L2_out_dist2__full_n;
  wire L2_out_dist2__write;
  wire [65:0] L2_out_dist3__dout;
  wire L2_out_dist3__empty_n;
  wire L2_out_dist3__read;
  wire [65:0] L2_out_dist3__din;
  wire L2_out_dist3__full_n;
  wire L2_out_dist3__write;
  wire [65:0] L2_out_dist4__dout;
  wire L2_out_dist4__empty_n;
  wire L2_out_dist4__read;
  wire [65:0] L2_out_dist4__din;
  wire L2_out_dist4__full_n;
  wire L2_out_dist4__write;
  wire [65:0] L2_out_dist5__dout;
  wire L2_out_dist5__empty_n;
  wire L2_out_dist5__read;
  wire [65:0] L2_out_dist5__din;
  wire L2_out_dist5__full_n;
  wire L2_out_dist5__write;
  wire [65:0] L2_out_id0__dout;
  wire L2_out_id0__empty_n;
  wire L2_out_id0__read;
  wire [65:0] L2_out_id0__din;
  wire L2_out_id0__full_n;
  wire L2_out_id0__write;
  wire [65:0] L2_out_id1__dout;
  wire L2_out_id1__empty_n;
  wire L2_out_id1__read;
  wire [65:0] L2_out_id1__din;
  wire L2_out_id1__full_n;
  wire L2_out_id1__write;
  wire [65:0] L2_out_id2__dout;
  wire L2_out_id2__empty_n;
  wire L2_out_id2__read;
  wire [65:0] L2_out_id2__din;
  wire L2_out_id2__full_n;
  wire L2_out_id2__write;
  wire [65:0] L2_out_id3__dout;
  wire L2_out_id3__empty_n;
  wire L2_out_id3__read;
  wire [65:0] L2_out_id3__din;
  wire L2_out_id3__full_n;
  wire L2_out_id3__write;
  wire [65:0] L2_out_id4__dout;
  wire L2_out_id4__empty_n;
  wire L2_out_id4__read;
  wire [65:0] L2_out_id4__din;
  wire L2_out_id4__full_n;
  wire L2_out_id4__write;
  wire [65:0] L2_out_id5__dout;
  wire L2_out_id5__empty_n;
  wire L2_out_id5__read;
  wire [65:0] L2_out_id5__din;
  wire L2_out_id5__full_n;
  wire L2_out_id5__write;
  wire [65:0] L3_out_dist0__dout;
  wire L3_out_dist0__empty_n;
  wire L3_out_dist0__read;
  wire [65:0] L3_out_dist0__din;
  wire L3_out_dist0__full_n;
  wire L3_out_dist0__write;
  wire [65:0] L3_out_dist1__dout;
  wire L3_out_dist1__empty_n;
  wire L3_out_dist1__read;
  wire [65:0] L3_out_dist1__din;
  wire L3_out_dist1__full_n;
  wire L3_out_dist1__write;
  wire [65:0] L3_out_id0__dout;
  wire L3_out_id0__empty_n;
  wire L3_out_id0__read;
  wire [65:0] L3_out_id0__din;
  wire L3_out_id0__full_n;
  wire L3_out_id0__write;
  wire [65:0] L3_out_id1__dout;
  wire L3_out_id1__empty_n;
  wire L3_out_id1__read;
  wire [65:0] L3_out_id1__din;
  wire L3_out_id1__full_n;
  wire L3_out_id1__write;
  wire [65:0] out_dist_0__dout;
  wire out_dist_0__empty_n;
  wire out_dist_0__read;
  wire [65:0] out_dist_0__din;
  wire out_dist_0__full_n;
  wire out_dist_0__write;
  wire [65:0] out_dist_10__dout;
  wire out_dist_10__empty_n;
  wire out_dist_10__read;
  wire [65:0] out_dist_10__din;
  wire out_dist_10__full_n;
  wire out_dist_10__write;
  wire [65:0] out_dist_11__dout;
  wire out_dist_11__empty_n;
  wire out_dist_11__read;
  wire [65:0] out_dist_11__din;
  wire out_dist_11__full_n;
  wire out_dist_11__write;
  wire [65:0] out_dist_12__dout;
  wire out_dist_12__empty_n;
  wire out_dist_12__read;
  wire [65:0] out_dist_12__din;
  wire out_dist_12__full_n;
  wire out_dist_12__write;
  wire [65:0] out_dist_13__dout;
  wire out_dist_13__empty_n;
  wire out_dist_13__read;
  wire [65:0] out_dist_13__din;
  wire out_dist_13__full_n;
  wire out_dist_13__write;
  wire [65:0] out_dist_14__dout;
  wire out_dist_14__empty_n;
  wire out_dist_14__read;
  wire [65:0] out_dist_14__din;
  wire out_dist_14__full_n;
  wire out_dist_14__write;
  wire [65:0] out_dist_15__dout;
  wire out_dist_15__empty_n;
  wire out_dist_15__read;
  wire [65:0] out_dist_15__din;
  wire out_dist_15__full_n;
  wire out_dist_15__write;
  wire [65:0] out_dist_16__dout;
  wire out_dist_16__empty_n;
  wire out_dist_16__read;
  wire [65:0] out_dist_16__din;
  wire out_dist_16__full_n;
  wire out_dist_16__write;
  wire [65:0] out_dist_17__dout;
  wire out_dist_17__empty_n;
  wire out_dist_17__read;
  wire [65:0] out_dist_17__din;
  wire out_dist_17__full_n;
  wire out_dist_17__write;
  wire [65:0] out_dist_18__dout;
  wire out_dist_18__empty_n;
  wire out_dist_18__read;
  wire [65:0] out_dist_18__din;
  wire out_dist_18__full_n;
  wire out_dist_18__write;
  wire [65:0] out_dist_19__dout;
  wire out_dist_19__empty_n;
  wire out_dist_19__read;
  wire [65:0] out_dist_19__din;
  wire out_dist_19__full_n;
  wire out_dist_19__write;
  wire [65:0] out_dist_1__dout;
  wire out_dist_1__empty_n;
  wire out_dist_1__read;
  wire [65:0] out_dist_1__din;
  wire out_dist_1__full_n;
  wire out_dist_1__write;
  wire [65:0] out_dist_20__dout;
  wire out_dist_20__empty_n;
  wire out_dist_20__read;
  wire [65:0] out_dist_20__din;
  wire out_dist_20__full_n;
  wire out_dist_20__write;
  wire [65:0] out_dist_21__dout;
  wire out_dist_21__empty_n;
  wire out_dist_21__read;
  wire [65:0] out_dist_21__din;
  wire out_dist_21__full_n;
  wire out_dist_21__write;
  wire [65:0] out_dist_22__dout;
  wire out_dist_22__empty_n;
  wire out_dist_22__read;
  wire [65:0] out_dist_22__din;
  wire out_dist_22__full_n;
  wire out_dist_22__write;
  wire [65:0] out_dist_23__dout;
  wire out_dist_23__empty_n;
  wire out_dist_23__read;
  wire [65:0] out_dist_23__din;
  wire out_dist_23__full_n;
  wire out_dist_23__write;
  wire [65:0] out_dist_24__dout;
  wire out_dist_24__empty_n;
  wire out_dist_24__read;
  wire [65:0] out_dist_24__din;
  wire out_dist_24__full_n;
  wire out_dist_24__write;
  wire [65:0] out_dist_25__dout;
  wire out_dist_25__empty_n;
  wire out_dist_25__read;
  wire [65:0] out_dist_25__din;
  wire out_dist_25__full_n;
  wire out_dist_25__write;
  wire [65:0] out_dist_26__dout;
  wire out_dist_26__empty_n;
  wire out_dist_26__read;
  wire [65:0] out_dist_26__din;
  wire out_dist_26__full_n;
  wire out_dist_26__write;
  wire [65:0] out_dist_27__dout;
  wire out_dist_27__empty_n;
  wire out_dist_27__read;
  wire [65:0] out_dist_27__din;
  wire out_dist_27__full_n;
  wire out_dist_27__write;
  wire [65:0] out_dist_28__dout;
  wire out_dist_28__empty_n;
  wire out_dist_28__read;
  wire [65:0] out_dist_28__din;
  wire out_dist_28__full_n;
  wire out_dist_28__write;
  wire [65:0] out_dist_29__dout;
  wire out_dist_29__empty_n;
  wire out_dist_29__read;
  wire [65:0] out_dist_29__din;
  wire out_dist_29__full_n;
  wire out_dist_29__write;
  wire [65:0] out_dist_2__dout;
  wire out_dist_2__empty_n;
  wire out_dist_2__read;
  wire [65:0] out_dist_2__din;
  wire out_dist_2__full_n;
  wire out_dist_2__write;
  wire [65:0] out_dist_30__dout;
  wire out_dist_30__empty_n;
  wire out_dist_30__read;
  wire [65:0] out_dist_30__din;
  wire out_dist_30__full_n;
  wire out_dist_30__write;
  wire [65:0] out_dist_31__dout;
  wire out_dist_31__empty_n;
  wire out_dist_31__read;
  wire [65:0] out_dist_31__din;
  wire out_dist_31__full_n;
  wire out_dist_31__write;
  wire [65:0] out_dist_32__dout;
  wire out_dist_32__empty_n;
  wire out_dist_32__read;
  wire [65:0] out_dist_32__din;
  wire out_dist_32__full_n;
  wire out_dist_32__write;
  wire [65:0] out_dist_33__dout;
  wire out_dist_33__empty_n;
  wire out_dist_33__read;
  wire [65:0] out_dist_33__din;
  wire out_dist_33__full_n;
  wire out_dist_33__write;
  wire [65:0] out_dist_34__dout;
  wire out_dist_34__empty_n;
  wire out_dist_34__read;
  wire [65:0] out_dist_34__din;
  wire out_dist_34__full_n;
  wire out_dist_34__write;
  wire [65:0] out_dist_35__dout;
  wire out_dist_35__empty_n;
  wire out_dist_35__read;
  wire [65:0] out_dist_35__din;
  wire out_dist_35__full_n;
  wire out_dist_35__write;
  wire [65:0] out_dist_36__dout;
  wire out_dist_36__empty_n;
  wire out_dist_36__read;
  wire [65:0] out_dist_36__din;
  wire out_dist_36__full_n;
  wire out_dist_36__write;
  wire [65:0] out_dist_37__dout;
  wire out_dist_37__empty_n;
  wire out_dist_37__read;
  wire [65:0] out_dist_37__din;
  wire out_dist_37__full_n;
  wire out_dist_37__write;
  wire [65:0] out_dist_38__dout;
  wire out_dist_38__empty_n;
  wire out_dist_38__read;
  wire [65:0] out_dist_38__din;
  wire out_dist_38__full_n;
  wire out_dist_38__write;
  wire [65:0] out_dist_39__dout;
  wire out_dist_39__empty_n;
  wire out_dist_39__read;
  wire [65:0] out_dist_39__din;
  wire out_dist_39__full_n;
  wire out_dist_39__write;
  wire [65:0] out_dist_3__dout;
  wire out_dist_3__empty_n;
  wire out_dist_3__read;
  wire [65:0] out_dist_3__din;
  wire out_dist_3__full_n;
  wire out_dist_3__write;
  wire [65:0] out_dist_40__dout;
  wire out_dist_40__empty_n;
  wire out_dist_40__read;
  wire [65:0] out_dist_40__din;
  wire out_dist_40__full_n;
  wire out_dist_40__write;
  wire [65:0] out_dist_41__dout;
  wire out_dist_41__empty_n;
  wire out_dist_41__read;
  wire [65:0] out_dist_41__din;
  wire out_dist_41__full_n;
  wire out_dist_41__write;
  wire [65:0] out_dist_42__dout;
  wire out_dist_42__empty_n;
  wire out_dist_42__read;
  wire [65:0] out_dist_42__din;
  wire out_dist_42__full_n;
  wire out_dist_42__write;
  wire [65:0] out_dist_43__dout;
  wire out_dist_43__empty_n;
  wire out_dist_43__read;
  wire [65:0] out_dist_43__din;
  wire out_dist_43__full_n;
  wire out_dist_43__write;
  wire [65:0] out_dist_44__dout;
  wire out_dist_44__empty_n;
  wire out_dist_44__read;
  wire [65:0] out_dist_44__din;
  wire out_dist_44__full_n;
  wire out_dist_44__write;
  wire [65:0] out_dist_45__dout;
  wire out_dist_45__empty_n;
  wire out_dist_45__read;
  wire [65:0] out_dist_45__din;
  wire out_dist_45__full_n;
  wire out_dist_45__write;
  wire [65:0] out_dist_46__dout;
  wire out_dist_46__empty_n;
  wire out_dist_46__read;
  wire [65:0] out_dist_46__din;
  wire out_dist_46__full_n;
  wire out_dist_46__write;
  wire [65:0] out_dist_47__dout;
  wire out_dist_47__empty_n;
  wire out_dist_47__read;
  wire [65:0] out_dist_47__din;
  wire out_dist_47__full_n;
  wire out_dist_47__write;
  wire [65:0] out_dist_48__dout;
  wire out_dist_48__empty_n;
  wire out_dist_48__read;
  wire [65:0] out_dist_48__din;
  wire out_dist_48__full_n;
  wire out_dist_48__write;
  wire [65:0] out_dist_49__dout;
  wire out_dist_49__empty_n;
  wire out_dist_49__read;
  wire [65:0] out_dist_49__din;
  wire out_dist_49__full_n;
  wire out_dist_49__write;
  wire [65:0] out_dist_4__dout;
  wire out_dist_4__empty_n;
  wire out_dist_4__read;
  wire [65:0] out_dist_4__din;
  wire out_dist_4__full_n;
  wire out_dist_4__write;
  wire [65:0] out_dist_50__dout;
  wire out_dist_50__empty_n;
  wire out_dist_50__read;
  wire [65:0] out_dist_50__din;
  wire out_dist_50__full_n;
  wire out_dist_50__write;
  wire [65:0] out_dist_51__dout;
  wire out_dist_51__empty_n;
  wire out_dist_51__read;
  wire [65:0] out_dist_51__din;
  wire out_dist_51__full_n;
  wire out_dist_51__write;
  wire [65:0] out_dist_52__dout;
  wire out_dist_52__empty_n;
  wire out_dist_52__read;
  wire [65:0] out_dist_52__din;
  wire out_dist_52__full_n;
  wire out_dist_52__write;
  wire [65:0] out_dist_53__dout;
  wire out_dist_53__empty_n;
  wire out_dist_53__read;
  wire [65:0] out_dist_53__din;
  wire out_dist_53__full_n;
  wire out_dist_53__write;
  wire [65:0] out_dist_5__dout;
  wire out_dist_5__empty_n;
  wire out_dist_5__read;
  wire [65:0] out_dist_5__din;
  wire out_dist_5__full_n;
  wire out_dist_5__write;
  wire [65:0] out_dist_6__dout;
  wire out_dist_6__empty_n;
  wire out_dist_6__read;
  wire [65:0] out_dist_6__din;
  wire out_dist_6__full_n;
  wire out_dist_6__write;
  wire [65:0] out_dist_7__dout;
  wire out_dist_7__empty_n;
  wire out_dist_7__read;
  wire [65:0] out_dist_7__din;
  wire out_dist_7__full_n;
  wire out_dist_7__write;
  wire [65:0] out_dist_8__dout;
  wire out_dist_8__empty_n;
  wire out_dist_8__read;
  wire [65:0] out_dist_8__din;
  wire out_dist_8__full_n;
  wire out_dist_8__write;
  wire [65:0] out_dist_9__dout;
  wire out_dist_9__empty_n;
  wire out_dist_9__read;
  wire [65:0] out_dist_9__din;
  wire out_dist_9__full_n;
  wire out_dist_9__write;
  wire [65:0] out_id_0__dout;
  wire out_id_0__empty_n;
  wire out_id_0__read;
  wire [65:0] out_id_0__din;
  wire out_id_0__full_n;
  wire out_id_0__write;
  wire [65:0] out_id_10__dout;
  wire out_id_10__empty_n;
  wire out_id_10__read;
  wire [65:0] out_id_10__din;
  wire out_id_10__full_n;
  wire out_id_10__write;
  wire [65:0] out_id_11__dout;
  wire out_id_11__empty_n;
  wire out_id_11__read;
  wire [65:0] out_id_11__din;
  wire out_id_11__full_n;
  wire out_id_11__write;
  wire [65:0] out_id_12__dout;
  wire out_id_12__empty_n;
  wire out_id_12__read;
  wire [65:0] out_id_12__din;
  wire out_id_12__full_n;
  wire out_id_12__write;
  wire [65:0] out_id_13__dout;
  wire out_id_13__empty_n;
  wire out_id_13__read;
  wire [65:0] out_id_13__din;
  wire out_id_13__full_n;
  wire out_id_13__write;
  wire [65:0] out_id_14__dout;
  wire out_id_14__empty_n;
  wire out_id_14__read;
  wire [65:0] out_id_14__din;
  wire out_id_14__full_n;
  wire out_id_14__write;
  wire [65:0] out_id_15__dout;
  wire out_id_15__empty_n;
  wire out_id_15__read;
  wire [65:0] out_id_15__din;
  wire out_id_15__full_n;
  wire out_id_15__write;
  wire [65:0] out_id_16__dout;
  wire out_id_16__empty_n;
  wire out_id_16__read;
  wire [65:0] out_id_16__din;
  wire out_id_16__full_n;
  wire out_id_16__write;
  wire [65:0] out_id_17__dout;
  wire out_id_17__empty_n;
  wire out_id_17__read;
  wire [65:0] out_id_17__din;
  wire out_id_17__full_n;
  wire out_id_17__write;
  wire [65:0] out_id_18__dout;
  wire out_id_18__empty_n;
  wire out_id_18__read;
  wire [65:0] out_id_18__din;
  wire out_id_18__full_n;
  wire out_id_18__write;
  wire [65:0] out_id_19__dout;
  wire out_id_19__empty_n;
  wire out_id_19__read;
  wire [65:0] out_id_19__din;
  wire out_id_19__full_n;
  wire out_id_19__write;
  wire [65:0] out_id_1__dout;
  wire out_id_1__empty_n;
  wire out_id_1__read;
  wire [65:0] out_id_1__din;
  wire out_id_1__full_n;
  wire out_id_1__write;
  wire [65:0] out_id_20__dout;
  wire out_id_20__empty_n;
  wire out_id_20__read;
  wire [65:0] out_id_20__din;
  wire out_id_20__full_n;
  wire out_id_20__write;
  wire [65:0] out_id_21__dout;
  wire out_id_21__empty_n;
  wire out_id_21__read;
  wire [65:0] out_id_21__din;
  wire out_id_21__full_n;
  wire out_id_21__write;
  wire [65:0] out_id_22__dout;
  wire out_id_22__empty_n;
  wire out_id_22__read;
  wire [65:0] out_id_22__din;
  wire out_id_22__full_n;
  wire out_id_22__write;
  wire [65:0] out_id_23__dout;
  wire out_id_23__empty_n;
  wire out_id_23__read;
  wire [65:0] out_id_23__din;
  wire out_id_23__full_n;
  wire out_id_23__write;
  wire [65:0] out_id_24__dout;
  wire out_id_24__empty_n;
  wire out_id_24__read;
  wire [65:0] out_id_24__din;
  wire out_id_24__full_n;
  wire out_id_24__write;
  wire [65:0] out_id_25__dout;
  wire out_id_25__empty_n;
  wire out_id_25__read;
  wire [65:0] out_id_25__din;
  wire out_id_25__full_n;
  wire out_id_25__write;
  wire [65:0] out_id_26__dout;
  wire out_id_26__empty_n;
  wire out_id_26__read;
  wire [65:0] out_id_26__din;
  wire out_id_26__full_n;
  wire out_id_26__write;
  wire [65:0] out_id_27__dout;
  wire out_id_27__empty_n;
  wire out_id_27__read;
  wire [65:0] out_id_27__din;
  wire out_id_27__full_n;
  wire out_id_27__write;
  wire [65:0] out_id_28__dout;
  wire out_id_28__empty_n;
  wire out_id_28__read;
  wire [65:0] out_id_28__din;
  wire out_id_28__full_n;
  wire out_id_28__write;
  wire [65:0] out_id_29__dout;
  wire out_id_29__empty_n;
  wire out_id_29__read;
  wire [65:0] out_id_29__din;
  wire out_id_29__full_n;
  wire out_id_29__write;
  wire [65:0] out_id_2__dout;
  wire out_id_2__empty_n;
  wire out_id_2__read;
  wire [65:0] out_id_2__din;
  wire out_id_2__full_n;
  wire out_id_2__write;
  wire [65:0] out_id_30__dout;
  wire out_id_30__empty_n;
  wire out_id_30__read;
  wire [65:0] out_id_30__din;
  wire out_id_30__full_n;
  wire out_id_30__write;
  wire [65:0] out_id_31__dout;
  wire out_id_31__empty_n;
  wire out_id_31__read;
  wire [65:0] out_id_31__din;
  wire out_id_31__full_n;
  wire out_id_31__write;
  wire [65:0] out_id_32__dout;
  wire out_id_32__empty_n;
  wire out_id_32__read;
  wire [65:0] out_id_32__din;
  wire out_id_32__full_n;
  wire out_id_32__write;
  wire [65:0] out_id_33__dout;
  wire out_id_33__empty_n;
  wire out_id_33__read;
  wire [65:0] out_id_33__din;
  wire out_id_33__full_n;
  wire out_id_33__write;
  wire [65:0] out_id_34__dout;
  wire out_id_34__empty_n;
  wire out_id_34__read;
  wire [65:0] out_id_34__din;
  wire out_id_34__full_n;
  wire out_id_34__write;
  wire [65:0] out_id_35__dout;
  wire out_id_35__empty_n;
  wire out_id_35__read;
  wire [65:0] out_id_35__din;
  wire out_id_35__full_n;
  wire out_id_35__write;
  wire [65:0] out_id_36__dout;
  wire out_id_36__empty_n;
  wire out_id_36__read;
  wire [65:0] out_id_36__din;
  wire out_id_36__full_n;
  wire out_id_36__write;
  wire [65:0] out_id_37__dout;
  wire out_id_37__empty_n;
  wire out_id_37__read;
  wire [65:0] out_id_37__din;
  wire out_id_37__full_n;
  wire out_id_37__write;
  wire [65:0] out_id_38__dout;
  wire out_id_38__empty_n;
  wire out_id_38__read;
  wire [65:0] out_id_38__din;
  wire out_id_38__full_n;
  wire out_id_38__write;
  wire [65:0] out_id_39__dout;
  wire out_id_39__empty_n;
  wire out_id_39__read;
  wire [65:0] out_id_39__din;
  wire out_id_39__full_n;
  wire out_id_39__write;
  wire [65:0] out_id_3__dout;
  wire out_id_3__empty_n;
  wire out_id_3__read;
  wire [65:0] out_id_3__din;
  wire out_id_3__full_n;
  wire out_id_3__write;
  wire [65:0] out_id_40__dout;
  wire out_id_40__empty_n;
  wire out_id_40__read;
  wire [65:0] out_id_40__din;
  wire out_id_40__full_n;
  wire out_id_40__write;
  wire [65:0] out_id_41__dout;
  wire out_id_41__empty_n;
  wire out_id_41__read;
  wire [65:0] out_id_41__din;
  wire out_id_41__full_n;
  wire out_id_41__write;
  wire [65:0] out_id_42__dout;
  wire out_id_42__empty_n;
  wire out_id_42__read;
  wire [65:0] out_id_42__din;
  wire out_id_42__full_n;
  wire out_id_42__write;
  wire [65:0] out_id_43__dout;
  wire out_id_43__empty_n;
  wire out_id_43__read;
  wire [65:0] out_id_43__din;
  wire out_id_43__full_n;
  wire out_id_43__write;
  wire [65:0] out_id_44__dout;
  wire out_id_44__empty_n;
  wire out_id_44__read;
  wire [65:0] out_id_44__din;
  wire out_id_44__full_n;
  wire out_id_44__write;
  wire [65:0] out_id_45__dout;
  wire out_id_45__empty_n;
  wire out_id_45__read;
  wire [65:0] out_id_45__din;
  wire out_id_45__full_n;
  wire out_id_45__write;
  wire [65:0] out_id_46__dout;
  wire out_id_46__empty_n;
  wire out_id_46__read;
  wire [65:0] out_id_46__din;
  wire out_id_46__full_n;
  wire out_id_46__write;
  wire [65:0] out_id_47__dout;
  wire out_id_47__empty_n;
  wire out_id_47__read;
  wire [65:0] out_id_47__din;
  wire out_id_47__full_n;
  wire out_id_47__write;
  wire [65:0] out_id_48__dout;
  wire out_id_48__empty_n;
  wire out_id_48__read;
  wire [65:0] out_id_48__din;
  wire out_id_48__full_n;
  wire out_id_48__write;
  wire [65:0] out_id_49__dout;
  wire out_id_49__empty_n;
  wire out_id_49__read;
  wire [65:0] out_id_49__din;
  wire out_id_49__full_n;
  wire out_id_49__write;
  wire [65:0] out_id_4__dout;
  wire out_id_4__empty_n;
  wire out_id_4__read;
  wire [65:0] out_id_4__din;
  wire out_id_4__full_n;
  wire out_id_4__write;
  wire [65:0] out_id_50__dout;
  wire out_id_50__empty_n;
  wire out_id_50__read;
  wire [65:0] out_id_50__din;
  wire out_id_50__full_n;
  wire out_id_50__write;
  wire [65:0] out_id_51__dout;
  wire out_id_51__empty_n;
  wire out_id_51__read;
  wire [65:0] out_id_51__din;
  wire out_id_51__full_n;
  wire out_id_51__write;
  wire [65:0] out_id_52__dout;
  wire out_id_52__empty_n;
  wire out_id_52__read;
  wire [65:0] out_id_52__din;
  wire out_id_52__full_n;
  wire out_id_52__write;
  wire [65:0] out_id_53__dout;
  wire out_id_53__empty_n;
  wire out_id_53__read;
  wire [65:0] out_id_53__din;
  wire out_id_53__full_n;
  wire out_id_53__write;
  wire [65:0] out_id_5__dout;
  wire out_id_5__empty_n;
  wire out_id_5__read;
  wire [65:0] out_id_5__din;
  wire out_id_5__full_n;
  wire out_id_5__write;
  wire [65:0] out_id_6__dout;
  wire out_id_6__empty_n;
  wire out_id_6__read;
  wire [65:0] out_id_6__din;
  wire out_id_6__full_n;
  wire out_id_6__write;
  wire [65:0] out_id_7__dout;
  wire out_id_7__empty_n;
  wire out_id_7__read;
  wire [65:0] out_id_7__din;
  wire out_id_7__full_n;
  wire out_id_7__write;
  wire [65:0] out_id_8__dout;
  wire out_id_8__empty_n;
  wire out_id_8__read;
  wire [65:0] out_id_8__din;
  wire out_id_8__full_n;
  wire out_id_8__write;
  wire [65:0] out_id_9__dout;
  wire out_id_9__empty_n;
  wire out_id_9__read;
  wire [65:0] out_id_9__din;
  wire out_id_9__full_n;
  wire out_id_9__write;
  wire krnl_globalSort_L1_L2_0__ap_start;
  wire krnl_globalSort_L1_L2_0__ap_ready;
  wire krnl_globalSort_L1_L2_0__ap_done;
  wire krnl_globalSort_L1_L2_0__ap_idle;
  wire krnl_globalSort_L1_L2_1__ap_start;
  wire krnl_globalSort_L1_L2_1__ap_ready;
  wire krnl_globalSort_L1_L2_1__ap_done;
  wire krnl_globalSort_L1_L2_1__ap_idle;
  wire krnl_globalSort_L1_L2_2__ap_start;
  wire krnl_globalSort_L1_L2_2__ap_ready;
  wire krnl_globalSort_L1_L2_2__ap_done;
  wire krnl_globalSort_L1_L2_2__ap_idle;
  wire krnl_globalSort_L1_L2_3__ap_start;
  wire krnl_globalSort_L1_L2_3__ap_ready;
  wire krnl_globalSort_L1_L2_3__ap_done;
  wire krnl_globalSort_L1_L2_3__ap_idle;
  wire krnl_globalSort_L1_L2_4__ap_start;
  wire krnl_globalSort_L1_L2_4__ap_ready;
  wire krnl_globalSort_L1_L2_4__ap_done;
  wire krnl_globalSort_L1_L2_4__ap_idle;
  wire krnl_globalSort_L1_L2_5__ap_start;
  wire krnl_globalSort_L1_L2_5__ap_ready;
  wire krnl_globalSort_L1_L2_5__ap_done;
  wire krnl_globalSort_L1_L2_5__ap_idle;
  wire krnl_globalSort_L1_L2_6__ap_start;
  wire krnl_globalSort_L1_L2_6__ap_ready;
  wire krnl_globalSort_L1_L2_6__ap_done;
  wire krnl_globalSort_L1_L2_6__ap_idle;
  wire krnl_globalSort_L1_L2_7__ap_start;
  wire krnl_globalSort_L1_L2_7__ap_ready;
  wire krnl_globalSort_L1_L2_7__ap_done;
  wire krnl_globalSort_L1_L2_7__ap_idle;
  wire krnl_globalSort_L1_L2_8__ap_start;
  wire krnl_globalSort_L1_L2_8__ap_ready;
  wire krnl_globalSort_L1_L2_8__ap_done;
  wire krnl_globalSort_L1_L2_8__ap_idle;
  wire krnl_globalSort_L1_L2_9__ap_start;
  wire krnl_globalSort_L1_L2_9__ap_ready;
  wire krnl_globalSort_L1_L2_9__ap_done;
  wire krnl_globalSort_L1_L2_9__ap_idle;
  wire krnl_globalSort_L1_L2_10__ap_start;
  wire krnl_globalSort_L1_L2_10__ap_ready;
  wire krnl_globalSort_L1_L2_10__ap_done;
  wire krnl_globalSort_L1_L2_10__ap_idle;
  wire krnl_globalSort_L1_L2_11__ap_start;
  wire krnl_globalSort_L1_L2_11__ap_ready;
  wire krnl_globalSort_L1_L2_11__ap_done;
  wire krnl_globalSort_L1_L2_11__ap_idle;
  wire krnl_globalSort_L1_L2_12__ap_start;
  wire krnl_globalSort_L1_L2_12__ap_ready;
  wire krnl_globalSort_L1_L2_12__ap_done;
  wire krnl_globalSort_L1_L2_12__ap_idle;
  wire krnl_globalSort_L1_L2_13__ap_start;
  wire krnl_globalSort_L1_L2_13__ap_ready;
  wire krnl_globalSort_L1_L2_13__ap_done;
  wire krnl_globalSort_L1_L2_13__ap_idle;
  wire krnl_globalSort_L1_L2_14__ap_start;
  wire krnl_globalSort_L1_L2_14__ap_ready;
  wire krnl_globalSort_L1_L2_14__ap_done;
  wire krnl_globalSort_L1_L2_14__ap_idle;
  wire krnl_globalSort_L1_L2_15__ap_start;
  wire krnl_globalSort_L1_L2_15__ap_ready;
  wire krnl_globalSort_L1_L2_15__ap_done;
  wire krnl_globalSort_L1_L2_15__ap_idle;
  wire krnl_globalSort_L1_L2_16__ap_start;
  wire krnl_globalSort_L1_L2_16__ap_ready;
  wire krnl_globalSort_L1_L2_16__ap_done;
  wire krnl_globalSort_L1_L2_16__ap_idle;
  wire krnl_globalSort_L1_L2_17__ap_start;
  wire krnl_globalSort_L1_L2_17__ap_ready;
  wire krnl_globalSort_L1_L2_17__ap_done;
  wire krnl_globalSort_L1_L2_17__ap_idle;
  wire krnl_globalSort_L1_L2_18__ap_start;
  wire krnl_globalSort_L1_L2_18__ap_ready;
  wire krnl_globalSort_L1_L2_18__ap_done;
  wire krnl_globalSort_L1_L2_18__ap_idle;
  wire krnl_globalSort_L1_L2_19__ap_start;
  wire krnl_globalSort_L1_L2_19__ap_ready;
  wire krnl_globalSort_L1_L2_19__ap_done;
  wire krnl_globalSort_L1_L2_19__ap_idle;
  wire krnl_globalSort_L1_L2_20__ap_start;
  wire krnl_globalSort_L1_L2_20__ap_ready;
  wire krnl_globalSort_L1_L2_20__ap_done;
  wire krnl_globalSort_L1_L2_20__ap_idle;
  wire krnl_globalSort_L1_L2_21__ap_start;
  wire krnl_globalSort_L1_L2_21__ap_ready;
  wire krnl_globalSort_L1_L2_21__ap_done;
  wire krnl_globalSort_L1_L2_21__ap_idle;
  wire krnl_globalSort_L1_L2_22__ap_start;
  wire krnl_globalSort_L1_L2_22__ap_ready;
  wire krnl_globalSort_L1_L2_22__ap_done;
  wire krnl_globalSort_L1_L2_22__ap_idle;
  wire krnl_globalSort_L1_L2_23__ap_start;
  wire krnl_globalSort_L1_L2_23__ap_ready;
  wire krnl_globalSort_L1_L2_23__ap_done;
  wire krnl_globalSort_L1_L2_23__ap_idle;
  wire krnl_globalSort_L1_L2_24__ap_start;
  wire krnl_globalSort_L1_L2_24__ap_ready;
  wire krnl_globalSort_L1_L2_24__ap_done;
  wire krnl_globalSort_L1_L2_24__ap_idle;
  wire krnl_globalSort_L1_L2_25__ap_start;
  wire krnl_globalSort_L1_L2_25__ap_ready;
  wire krnl_globalSort_L1_L2_25__ap_done;
  wire krnl_globalSort_L1_L2_25__ap_idle;
  wire [63:0] krnl_globalSort_L3_0___L4_out_dist__q0;
  wire [63:0] L4_out_dist_read_addr__din;
  wire L4_out_dist_read_addr__full_n;
  wire L4_out_dist_read_addr__write;
  wire [31:0] L4_out_dist_read_data__dout;
  wire L4_out_dist_read_data__empty_n;
  wire L4_out_dist_read_data__read;
  wire [63:0] L4_out_dist_write_addr__din;
  wire L4_out_dist_write_addr__full_n;
  wire L4_out_dist_write_addr__write;
  wire [31:0] L4_out_dist_write_data__din;
  wire L4_out_dist_write_data__full_n;
  wire L4_out_dist_write_data__write;
  wire [7:0] L4_out_dist_write_resp__dout;
  wire L4_out_dist_write_resp__empty_n;
  wire L4_out_dist_write_resp__read;
  wire [63:0] krnl_globalSort_L3_0___L4_out_id__q0;
  wire [63:0] L4_out_id_read_addr__din;
  wire L4_out_id_read_addr__full_n;
  wire L4_out_id_read_addr__write;
  wire [31:0] L4_out_id_read_data__dout;
  wire L4_out_id_read_data__empty_n;
  wire L4_out_id_read_data__read;
  wire [63:0] L4_out_id_write_addr__din;
  wire L4_out_id_write_addr__full_n;
  wire L4_out_id_write_addr__write;
  wire [31:0] L4_out_id_write_data__din;
  wire L4_out_id_write_data__full_n;
  wire L4_out_id_write_data__write;
  wire [7:0] L4_out_id_write_resp__dout;
  wire L4_out_id_write_resp__empty_n;
  wire L4_out_id_write_resp__read;
  wire krnl_globalSort_L3_0__ap_start;
  wire krnl_globalSort_L3_0__ap_ready;
  wire krnl_globalSort_L3_0__ap_done;
  wire krnl_globalSort_L3_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_0_0___in_0__q0;
  wire [63:0] in_0_read_addr__din;
  wire in_0_read_addr__full_n;
  wire in_0_read_addr__write;
  wire [255:0] in_0_read_data__dout;
  wire in_0_read_data__empty_n;
  wire in_0_read_data__read;
  wire [63:0] in_0_write_addr__din;
  wire in_0_write_addr__full_n;
  wire in_0_write_addr__write;
  wire [255:0] in_0_write_data__din;
  wire in_0_write_data__full_n;
  wire in_0_write_data__write;
  wire [7:0] in_0_write_resp__dout;
  wire in_0_write_resp__empty_n;
  wire in_0_write_resp__read;
  wire krnl_partialKnn_wrapper_0_0__ap_start;
  wire krnl_partialKnn_wrapper_0_0__ap_ready;
  wire krnl_partialKnn_wrapper_0_0__ap_done;
  wire krnl_partialKnn_wrapper_0_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_1_0___in_1__q0;
  wire [63:0] in_1_read_addr__din;
  wire in_1_read_addr__full_n;
  wire in_1_read_addr__write;
  wire [255:0] in_1_read_data__dout;
  wire in_1_read_data__empty_n;
  wire in_1_read_data__read;
  wire [63:0] in_1_write_addr__din;
  wire in_1_write_addr__full_n;
  wire in_1_write_addr__write;
  wire [255:0] in_1_write_data__din;
  wire in_1_write_data__full_n;
  wire in_1_write_data__write;
  wire [7:0] in_1_write_resp__dout;
  wire in_1_write_resp__empty_n;
  wire in_1_write_resp__read;
  wire krnl_partialKnn_wrapper_1_0__ap_start;
  wire krnl_partialKnn_wrapper_1_0__ap_ready;
  wire krnl_partialKnn_wrapper_1_0__ap_done;
  wire krnl_partialKnn_wrapper_1_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_10_0___in_10__q0;
  wire [63:0] in_10_read_addr__din;
  wire in_10_read_addr__full_n;
  wire in_10_read_addr__write;
  wire [255:0] in_10_read_data__dout;
  wire in_10_read_data__empty_n;
  wire in_10_read_data__read;
  wire [63:0] in_10_write_addr__din;
  wire in_10_write_addr__full_n;
  wire in_10_write_addr__write;
  wire [255:0] in_10_write_data__din;
  wire in_10_write_data__full_n;
  wire in_10_write_data__write;
  wire [7:0] in_10_write_resp__dout;
  wire in_10_write_resp__empty_n;
  wire in_10_write_resp__read;
  wire krnl_partialKnn_wrapper_10_0__ap_start;
  wire krnl_partialKnn_wrapper_10_0__ap_ready;
  wire krnl_partialKnn_wrapper_10_0__ap_done;
  wire krnl_partialKnn_wrapper_10_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_11_0___in_11__q0;
  wire [63:0] in_11_read_addr__din;
  wire in_11_read_addr__full_n;
  wire in_11_read_addr__write;
  wire [255:0] in_11_read_data__dout;
  wire in_11_read_data__empty_n;
  wire in_11_read_data__read;
  wire [63:0] in_11_write_addr__din;
  wire in_11_write_addr__full_n;
  wire in_11_write_addr__write;
  wire [255:0] in_11_write_data__din;
  wire in_11_write_data__full_n;
  wire in_11_write_data__write;
  wire [7:0] in_11_write_resp__dout;
  wire in_11_write_resp__empty_n;
  wire in_11_write_resp__read;
  wire krnl_partialKnn_wrapper_11_0__ap_start;
  wire krnl_partialKnn_wrapper_11_0__ap_ready;
  wire krnl_partialKnn_wrapper_11_0__ap_done;
  wire krnl_partialKnn_wrapper_11_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_12_0___in_12__q0;
  wire [63:0] in_12_read_addr__din;
  wire in_12_read_addr__full_n;
  wire in_12_read_addr__write;
  wire [255:0] in_12_read_data__dout;
  wire in_12_read_data__empty_n;
  wire in_12_read_data__read;
  wire [63:0] in_12_write_addr__din;
  wire in_12_write_addr__full_n;
  wire in_12_write_addr__write;
  wire [255:0] in_12_write_data__din;
  wire in_12_write_data__full_n;
  wire in_12_write_data__write;
  wire [7:0] in_12_write_resp__dout;
  wire in_12_write_resp__empty_n;
  wire in_12_write_resp__read;
  wire krnl_partialKnn_wrapper_12_0__ap_start;
  wire krnl_partialKnn_wrapper_12_0__ap_ready;
  wire krnl_partialKnn_wrapper_12_0__ap_done;
  wire krnl_partialKnn_wrapper_12_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_13_0___in_13__q0;
  wire [63:0] in_13_read_addr__din;
  wire in_13_read_addr__full_n;
  wire in_13_read_addr__write;
  wire [255:0] in_13_read_data__dout;
  wire in_13_read_data__empty_n;
  wire in_13_read_data__read;
  wire [63:0] in_13_write_addr__din;
  wire in_13_write_addr__full_n;
  wire in_13_write_addr__write;
  wire [255:0] in_13_write_data__din;
  wire in_13_write_data__full_n;
  wire in_13_write_data__write;
  wire [7:0] in_13_write_resp__dout;
  wire in_13_write_resp__empty_n;
  wire in_13_write_resp__read;
  wire krnl_partialKnn_wrapper_13_0__ap_start;
  wire krnl_partialKnn_wrapper_13_0__ap_ready;
  wire krnl_partialKnn_wrapper_13_0__ap_done;
  wire krnl_partialKnn_wrapper_13_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_14_0___in_14__q0;
  wire [63:0] in_14_read_addr__din;
  wire in_14_read_addr__full_n;
  wire in_14_read_addr__write;
  wire [255:0] in_14_read_data__dout;
  wire in_14_read_data__empty_n;
  wire in_14_read_data__read;
  wire [63:0] in_14_write_addr__din;
  wire in_14_write_addr__full_n;
  wire in_14_write_addr__write;
  wire [255:0] in_14_write_data__din;
  wire in_14_write_data__full_n;
  wire in_14_write_data__write;
  wire [7:0] in_14_write_resp__dout;
  wire in_14_write_resp__empty_n;
  wire in_14_write_resp__read;
  wire krnl_partialKnn_wrapper_14_0__ap_start;
  wire krnl_partialKnn_wrapper_14_0__ap_ready;
  wire krnl_partialKnn_wrapper_14_0__ap_done;
  wire krnl_partialKnn_wrapper_14_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_15_0___in_15__q0;
  wire [63:0] in_15_read_addr__din;
  wire in_15_read_addr__full_n;
  wire in_15_read_addr__write;
  wire [255:0] in_15_read_data__dout;
  wire in_15_read_data__empty_n;
  wire in_15_read_data__read;
  wire [63:0] in_15_write_addr__din;
  wire in_15_write_addr__full_n;
  wire in_15_write_addr__write;
  wire [255:0] in_15_write_data__din;
  wire in_15_write_data__full_n;
  wire in_15_write_data__write;
  wire [7:0] in_15_write_resp__dout;
  wire in_15_write_resp__empty_n;
  wire in_15_write_resp__read;
  wire krnl_partialKnn_wrapper_15_0__ap_start;
  wire krnl_partialKnn_wrapper_15_0__ap_ready;
  wire krnl_partialKnn_wrapper_15_0__ap_done;
  wire krnl_partialKnn_wrapper_15_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_16_0___in_16__q0;
  wire [63:0] in_16_read_addr__din;
  wire in_16_read_addr__full_n;
  wire in_16_read_addr__write;
  wire [255:0] in_16_read_data__dout;
  wire in_16_read_data__empty_n;
  wire in_16_read_data__read;
  wire [63:0] in_16_write_addr__din;
  wire in_16_write_addr__full_n;
  wire in_16_write_addr__write;
  wire [255:0] in_16_write_data__din;
  wire in_16_write_data__full_n;
  wire in_16_write_data__write;
  wire [7:0] in_16_write_resp__dout;
  wire in_16_write_resp__empty_n;
  wire in_16_write_resp__read;
  wire krnl_partialKnn_wrapper_16_0__ap_start;
  wire krnl_partialKnn_wrapper_16_0__ap_ready;
  wire krnl_partialKnn_wrapper_16_0__ap_done;
  wire krnl_partialKnn_wrapper_16_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_17_0___in_17__q0;
  wire [63:0] in_17_read_addr__din;
  wire in_17_read_addr__full_n;
  wire in_17_read_addr__write;
  wire [255:0] in_17_read_data__dout;
  wire in_17_read_data__empty_n;
  wire in_17_read_data__read;
  wire [63:0] in_17_write_addr__din;
  wire in_17_write_addr__full_n;
  wire in_17_write_addr__write;
  wire [255:0] in_17_write_data__din;
  wire in_17_write_data__full_n;
  wire in_17_write_data__write;
  wire [7:0] in_17_write_resp__dout;
  wire in_17_write_resp__empty_n;
  wire in_17_write_resp__read;
  wire krnl_partialKnn_wrapper_17_0__ap_start;
  wire krnl_partialKnn_wrapper_17_0__ap_ready;
  wire krnl_partialKnn_wrapper_17_0__ap_done;
  wire krnl_partialKnn_wrapper_17_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_18_0___in_18__q0;
  wire [63:0] in_18_read_addr__din;
  wire in_18_read_addr__full_n;
  wire in_18_read_addr__write;
  wire [255:0] in_18_read_data__dout;
  wire in_18_read_data__empty_n;
  wire in_18_read_data__read;
  wire [63:0] in_18_write_addr__din;
  wire in_18_write_addr__full_n;
  wire in_18_write_addr__write;
  wire [255:0] in_18_write_data__din;
  wire in_18_write_data__full_n;
  wire in_18_write_data__write;
  wire [7:0] in_18_write_resp__dout;
  wire in_18_write_resp__empty_n;
  wire in_18_write_resp__read;
  wire krnl_partialKnn_wrapper_18_0__ap_start;
  wire krnl_partialKnn_wrapper_18_0__ap_ready;
  wire krnl_partialKnn_wrapper_18_0__ap_done;
  wire krnl_partialKnn_wrapper_18_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_19_0___in_19__q0;
  wire [63:0] in_19_read_addr__din;
  wire in_19_read_addr__full_n;
  wire in_19_read_addr__write;
  wire [255:0] in_19_read_data__dout;
  wire in_19_read_data__empty_n;
  wire in_19_read_data__read;
  wire [63:0] in_19_write_addr__din;
  wire in_19_write_addr__full_n;
  wire in_19_write_addr__write;
  wire [255:0] in_19_write_data__din;
  wire in_19_write_data__full_n;
  wire in_19_write_data__write;
  wire [7:0] in_19_write_resp__dout;
  wire in_19_write_resp__empty_n;
  wire in_19_write_resp__read;
  wire krnl_partialKnn_wrapper_19_0__ap_start;
  wire krnl_partialKnn_wrapper_19_0__ap_ready;
  wire krnl_partialKnn_wrapper_19_0__ap_done;
  wire krnl_partialKnn_wrapper_19_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_2_0___in_2__q0;
  wire [63:0] in_2_read_addr__din;
  wire in_2_read_addr__full_n;
  wire in_2_read_addr__write;
  wire [255:0] in_2_read_data__dout;
  wire in_2_read_data__empty_n;
  wire in_2_read_data__read;
  wire [63:0] in_2_write_addr__din;
  wire in_2_write_addr__full_n;
  wire in_2_write_addr__write;
  wire [255:0] in_2_write_data__din;
  wire in_2_write_data__full_n;
  wire in_2_write_data__write;
  wire [7:0] in_2_write_resp__dout;
  wire in_2_write_resp__empty_n;
  wire in_2_write_resp__read;
  wire krnl_partialKnn_wrapper_2_0__ap_start;
  wire krnl_partialKnn_wrapper_2_0__ap_ready;
  wire krnl_partialKnn_wrapper_2_0__ap_done;
  wire krnl_partialKnn_wrapper_2_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_20_0___in_20__q0;
  wire [63:0] in_20_read_addr__din;
  wire in_20_read_addr__full_n;
  wire in_20_read_addr__write;
  wire [255:0] in_20_read_data__dout;
  wire in_20_read_data__empty_n;
  wire in_20_read_data__read;
  wire [63:0] in_20_write_addr__din;
  wire in_20_write_addr__full_n;
  wire in_20_write_addr__write;
  wire [255:0] in_20_write_data__din;
  wire in_20_write_data__full_n;
  wire in_20_write_data__write;
  wire [7:0] in_20_write_resp__dout;
  wire in_20_write_resp__empty_n;
  wire in_20_write_resp__read;
  wire krnl_partialKnn_wrapper_20_0__ap_start;
  wire krnl_partialKnn_wrapper_20_0__ap_ready;
  wire krnl_partialKnn_wrapper_20_0__ap_done;
  wire krnl_partialKnn_wrapper_20_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_21_0___in_21__q0;
  wire [63:0] in_21_read_addr__din;
  wire in_21_read_addr__full_n;
  wire in_21_read_addr__write;
  wire [255:0] in_21_read_data__dout;
  wire in_21_read_data__empty_n;
  wire in_21_read_data__read;
  wire [63:0] in_21_write_addr__din;
  wire in_21_write_addr__full_n;
  wire in_21_write_addr__write;
  wire [255:0] in_21_write_data__din;
  wire in_21_write_data__full_n;
  wire in_21_write_data__write;
  wire [7:0] in_21_write_resp__dout;
  wire in_21_write_resp__empty_n;
  wire in_21_write_resp__read;
  wire krnl_partialKnn_wrapper_21_0__ap_start;
  wire krnl_partialKnn_wrapper_21_0__ap_ready;
  wire krnl_partialKnn_wrapper_21_0__ap_done;
  wire krnl_partialKnn_wrapper_21_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_22_0___in_22__q0;
  wire [63:0] in_22_read_addr__din;
  wire in_22_read_addr__full_n;
  wire in_22_read_addr__write;
  wire [255:0] in_22_read_data__dout;
  wire in_22_read_data__empty_n;
  wire in_22_read_data__read;
  wire [63:0] in_22_write_addr__din;
  wire in_22_write_addr__full_n;
  wire in_22_write_addr__write;
  wire [255:0] in_22_write_data__din;
  wire in_22_write_data__full_n;
  wire in_22_write_data__write;
  wire [7:0] in_22_write_resp__dout;
  wire in_22_write_resp__empty_n;
  wire in_22_write_resp__read;
  wire krnl_partialKnn_wrapper_22_0__ap_start;
  wire krnl_partialKnn_wrapper_22_0__ap_ready;
  wire krnl_partialKnn_wrapper_22_0__ap_done;
  wire krnl_partialKnn_wrapper_22_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_23_0___in_23__q0;
  wire [63:0] in_23_read_addr__din;
  wire in_23_read_addr__full_n;
  wire in_23_read_addr__write;
  wire [255:0] in_23_read_data__dout;
  wire in_23_read_data__empty_n;
  wire in_23_read_data__read;
  wire [63:0] in_23_write_addr__din;
  wire in_23_write_addr__full_n;
  wire in_23_write_addr__write;
  wire [255:0] in_23_write_data__din;
  wire in_23_write_data__full_n;
  wire in_23_write_data__write;
  wire [7:0] in_23_write_resp__dout;
  wire in_23_write_resp__empty_n;
  wire in_23_write_resp__read;
  wire krnl_partialKnn_wrapper_23_0__ap_start;
  wire krnl_partialKnn_wrapper_23_0__ap_ready;
  wire krnl_partialKnn_wrapper_23_0__ap_done;
  wire krnl_partialKnn_wrapper_23_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_24_0___in_24__q0;
  wire [63:0] in_24_read_addr__din;
  wire in_24_read_addr__full_n;
  wire in_24_read_addr__write;
  wire [255:0] in_24_read_data__dout;
  wire in_24_read_data__empty_n;
  wire in_24_read_data__read;
  wire [63:0] in_24_write_addr__din;
  wire in_24_write_addr__full_n;
  wire in_24_write_addr__write;
  wire [255:0] in_24_write_data__din;
  wire in_24_write_data__full_n;
  wire in_24_write_data__write;
  wire [7:0] in_24_write_resp__dout;
  wire in_24_write_resp__empty_n;
  wire in_24_write_resp__read;
  wire krnl_partialKnn_wrapper_24_0__ap_start;
  wire krnl_partialKnn_wrapper_24_0__ap_ready;
  wire krnl_partialKnn_wrapper_24_0__ap_done;
  wire krnl_partialKnn_wrapper_24_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_25_0___in_25__q0;
  wire [63:0] in_25_read_addr__din;
  wire in_25_read_addr__full_n;
  wire in_25_read_addr__write;
  wire [255:0] in_25_read_data__dout;
  wire in_25_read_data__empty_n;
  wire in_25_read_data__read;
  wire [63:0] in_25_write_addr__din;
  wire in_25_write_addr__full_n;
  wire in_25_write_addr__write;
  wire [255:0] in_25_write_data__din;
  wire in_25_write_data__full_n;
  wire in_25_write_data__write;
  wire [7:0] in_25_write_resp__dout;
  wire in_25_write_resp__empty_n;
  wire in_25_write_resp__read;
  wire krnl_partialKnn_wrapper_25_0__ap_start;
  wire krnl_partialKnn_wrapper_25_0__ap_ready;
  wire krnl_partialKnn_wrapper_25_0__ap_done;
  wire krnl_partialKnn_wrapper_25_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_26_0___in_26__q0;
  wire [63:0] in_26_read_addr__din;
  wire in_26_read_addr__full_n;
  wire in_26_read_addr__write;
  wire [255:0] in_26_read_data__dout;
  wire in_26_read_data__empty_n;
  wire in_26_read_data__read;
  wire [63:0] in_26_write_addr__din;
  wire in_26_write_addr__full_n;
  wire in_26_write_addr__write;
  wire [255:0] in_26_write_data__din;
  wire in_26_write_data__full_n;
  wire in_26_write_data__write;
  wire [7:0] in_26_write_resp__dout;
  wire in_26_write_resp__empty_n;
  wire in_26_write_resp__read;
  wire krnl_partialKnn_wrapper_26_0__ap_start;
  wire krnl_partialKnn_wrapper_26_0__ap_ready;
  wire krnl_partialKnn_wrapper_26_0__ap_done;
  wire krnl_partialKnn_wrapper_26_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_27_0___in_27__q0;
  wire [63:0] in_27_read_addr__din;
  wire in_27_read_addr__full_n;
  wire in_27_read_addr__write;
  wire [255:0] in_27_read_data__dout;
  wire in_27_read_data__empty_n;
  wire in_27_read_data__read;
  wire [63:0] in_27_write_addr__din;
  wire in_27_write_addr__full_n;
  wire in_27_write_addr__write;
  wire [255:0] in_27_write_data__din;
  wire in_27_write_data__full_n;
  wire in_27_write_data__write;
  wire [7:0] in_27_write_resp__dout;
  wire in_27_write_resp__empty_n;
  wire in_27_write_resp__read;
  wire krnl_partialKnn_wrapper_27_0__ap_start;
  wire krnl_partialKnn_wrapper_27_0__ap_ready;
  wire krnl_partialKnn_wrapper_27_0__ap_done;
  wire krnl_partialKnn_wrapper_27_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_28_0___in_28__q0;
  wire [63:0] in_28_read_addr__din;
  wire in_28_read_addr__full_n;
  wire in_28_read_addr__write;
  wire [255:0] in_28_read_data__dout;
  wire in_28_read_data__empty_n;
  wire in_28_read_data__read;
  wire [63:0] in_28_write_addr__din;
  wire in_28_write_addr__full_n;
  wire in_28_write_addr__write;
  wire [255:0] in_28_write_data__din;
  wire in_28_write_data__full_n;
  wire in_28_write_data__write;
  wire [7:0] in_28_write_resp__dout;
  wire in_28_write_resp__empty_n;
  wire in_28_write_resp__read;
  wire krnl_partialKnn_wrapper_28_0__ap_start;
  wire krnl_partialKnn_wrapper_28_0__ap_ready;
  wire krnl_partialKnn_wrapper_28_0__ap_done;
  wire krnl_partialKnn_wrapper_28_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_29_0___in_29__q0;
  wire [63:0] in_29_read_addr__din;
  wire in_29_read_addr__full_n;
  wire in_29_read_addr__write;
  wire [255:0] in_29_read_data__dout;
  wire in_29_read_data__empty_n;
  wire in_29_read_data__read;
  wire [63:0] in_29_write_addr__din;
  wire in_29_write_addr__full_n;
  wire in_29_write_addr__write;
  wire [255:0] in_29_write_data__din;
  wire in_29_write_data__full_n;
  wire in_29_write_data__write;
  wire [7:0] in_29_write_resp__dout;
  wire in_29_write_resp__empty_n;
  wire in_29_write_resp__read;
  wire krnl_partialKnn_wrapper_29_0__ap_start;
  wire krnl_partialKnn_wrapper_29_0__ap_ready;
  wire krnl_partialKnn_wrapper_29_0__ap_done;
  wire krnl_partialKnn_wrapper_29_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_3_0___in_3__q0;
  wire [63:0] in_3_read_addr__din;
  wire in_3_read_addr__full_n;
  wire in_3_read_addr__write;
  wire [255:0] in_3_read_data__dout;
  wire in_3_read_data__empty_n;
  wire in_3_read_data__read;
  wire [63:0] in_3_write_addr__din;
  wire in_3_write_addr__full_n;
  wire in_3_write_addr__write;
  wire [255:0] in_3_write_data__din;
  wire in_3_write_data__full_n;
  wire in_3_write_data__write;
  wire [7:0] in_3_write_resp__dout;
  wire in_3_write_resp__empty_n;
  wire in_3_write_resp__read;
  wire krnl_partialKnn_wrapper_3_0__ap_start;
  wire krnl_partialKnn_wrapper_3_0__ap_ready;
  wire krnl_partialKnn_wrapper_3_0__ap_done;
  wire krnl_partialKnn_wrapper_3_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_30_0___in_30__q0;
  wire [63:0] in_30_read_addr__din;
  wire in_30_read_addr__full_n;
  wire in_30_read_addr__write;
  wire [255:0] in_30_read_data__dout;
  wire in_30_read_data__empty_n;
  wire in_30_read_data__read;
  wire [63:0] in_30_write_addr__din;
  wire in_30_write_addr__full_n;
  wire in_30_write_addr__write;
  wire [255:0] in_30_write_data__din;
  wire in_30_write_data__full_n;
  wire in_30_write_data__write;
  wire [7:0] in_30_write_resp__dout;
  wire in_30_write_resp__empty_n;
  wire in_30_write_resp__read;
  wire krnl_partialKnn_wrapper_30_0__ap_start;
  wire krnl_partialKnn_wrapper_30_0__ap_ready;
  wire krnl_partialKnn_wrapper_30_0__ap_done;
  wire krnl_partialKnn_wrapper_30_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_31_0___in_31__q0;
  wire [63:0] in_31_read_addr__din;
  wire in_31_read_addr__full_n;
  wire in_31_read_addr__write;
  wire [255:0] in_31_read_data__dout;
  wire in_31_read_data__empty_n;
  wire in_31_read_data__read;
  wire [63:0] in_31_write_addr__din;
  wire in_31_write_addr__full_n;
  wire in_31_write_addr__write;
  wire [255:0] in_31_write_data__din;
  wire in_31_write_data__full_n;
  wire in_31_write_data__write;
  wire [7:0] in_31_write_resp__dout;
  wire in_31_write_resp__empty_n;
  wire in_31_write_resp__read;
  wire krnl_partialKnn_wrapper_31_0__ap_start;
  wire krnl_partialKnn_wrapper_31_0__ap_ready;
  wire krnl_partialKnn_wrapper_31_0__ap_done;
  wire krnl_partialKnn_wrapper_31_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_32_0___in_32__q0;
  wire [63:0] in_32_read_addr__din;
  wire in_32_read_addr__full_n;
  wire in_32_read_addr__write;
  wire [255:0] in_32_read_data__dout;
  wire in_32_read_data__empty_n;
  wire in_32_read_data__read;
  wire [63:0] in_32_write_addr__din;
  wire in_32_write_addr__full_n;
  wire in_32_write_addr__write;
  wire [255:0] in_32_write_data__din;
  wire in_32_write_data__full_n;
  wire in_32_write_data__write;
  wire [7:0] in_32_write_resp__dout;
  wire in_32_write_resp__empty_n;
  wire in_32_write_resp__read;
  wire krnl_partialKnn_wrapper_32_0__ap_start;
  wire krnl_partialKnn_wrapper_32_0__ap_ready;
  wire krnl_partialKnn_wrapper_32_0__ap_done;
  wire krnl_partialKnn_wrapper_32_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_33_0___in_33__q0;
  wire [63:0] in_33_read_addr__din;
  wire in_33_read_addr__full_n;
  wire in_33_read_addr__write;
  wire [255:0] in_33_read_data__dout;
  wire in_33_read_data__empty_n;
  wire in_33_read_data__read;
  wire [63:0] in_33_write_addr__din;
  wire in_33_write_addr__full_n;
  wire in_33_write_addr__write;
  wire [255:0] in_33_write_data__din;
  wire in_33_write_data__full_n;
  wire in_33_write_data__write;
  wire [7:0] in_33_write_resp__dout;
  wire in_33_write_resp__empty_n;
  wire in_33_write_resp__read;
  wire krnl_partialKnn_wrapper_33_0__ap_start;
  wire krnl_partialKnn_wrapper_33_0__ap_ready;
  wire krnl_partialKnn_wrapper_33_0__ap_done;
  wire krnl_partialKnn_wrapper_33_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_34_0___in_34__q0;
  wire [63:0] in_34_read_addr__din;
  wire in_34_read_addr__full_n;
  wire in_34_read_addr__write;
  wire [255:0] in_34_read_data__dout;
  wire in_34_read_data__empty_n;
  wire in_34_read_data__read;
  wire [63:0] in_34_write_addr__din;
  wire in_34_write_addr__full_n;
  wire in_34_write_addr__write;
  wire [255:0] in_34_write_data__din;
  wire in_34_write_data__full_n;
  wire in_34_write_data__write;
  wire [7:0] in_34_write_resp__dout;
  wire in_34_write_resp__empty_n;
  wire in_34_write_resp__read;
  wire krnl_partialKnn_wrapper_34_0__ap_start;
  wire krnl_partialKnn_wrapper_34_0__ap_ready;
  wire krnl_partialKnn_wrapper_34_0__ap_done;
  wire krnl_partialKnn_wrapper_34_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_35_0___in_35__q0;
  wire [63:0] in_35_read_addr__din;
  wire in_35_read_addr__full_n;
  wire in_35_read_addr__write;
  wire [255:0] in_35_read_data__dout;
  wire in_35_read_data__empty_n;
  wire in_35_read_data__read;
  wire [63:0] in_35_write_addr__din;
  wire in_35_write_addr__full_n;
  wire in_35_write_addr__write;
  wire [255:0] in_35_write_data__din;
  wire in_35_write_data__full_n;
  wire in_35_write_data__write;
  wire [7:0] in_35_write_resp__dout;
  wire in_35_write_resp__empty_n;
  wire in_35_write_resp__read;
  wire krnl_partialKnn_wrapper_35_0__ap_start;
  wire krnl_partialKnn_wrapper_35_0__ap_ready;
  wire krnl_partialKnn_wrapper_35_0__ap_done;
  wire krnl_partialKnn_wrapper_35_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_36_0___in_36__q0;
  wire [63:0] in_36_read_addr__din;
  wire in_36_read_addr__full_n;
  wire in_36_read_addr__write;
  wire [255:0] in_36_read_data__dout;
  wire in_36_read_data__empty_n;
  wire in_36_read_data__read;
  wire [63:0] in_36_write_addr__din;
  wire in_36_write_addr__full_n;
  wire in_36_write_addr__write;
  wire [255:0] in_36_write_data__din;
  wire in_36_write_data__full_n;
  wire in_36_write_data__write;
  wire [7:0] in_36_write_resp__dout;
  wire in_36_write_resp__empty_n;
  wire in_36_write_resp__read;
  wire krnl_partialKnn_wrapper_36_0__ap_start;
  wire krnl_partialKnn_wrapper_36_0__ap_ready;
  wire krnl_partialKnn_wrapper_36_0__ap_done;
  wire krnl_partialKnn_wrapper_36_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_37_0___in_37__q0;
  wire [63:0] in_37_read_addr__din;
  wire in_37_read_addr__full_n;
  wire in_37_read_addr__write;
  wire [255:0] in_37_read_data__dout;
  wire in_37_read_data__empty_n;
  wire in_37_read_data__read;
  wire [63:0] in_37_write_addr__din;
  wire in_37_write_addr__full_n;
  wire in_37_write_addr__write;
  wire [255:0] in_37_write_data__din;
  wire in_37_write_data__full_n;
  wire in_37_write_data__write;
  wire [7:0] in_37_write_resp__dout;
  wire in_37_write_resp__empty_n;
  wire in_37_write_resp__read;
  wire krnl_partialKnn_wrapper_37_0__ap_start;
  wire krnl_partialKnn_wrapper_37_0__ap_ready;
  wire krnl_partialKnn_wrapper_37_0__ap_done;
  wire krnl_partialKnn_wrapper_37_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_38_0___in_38__q0;
  wire [63:0] in_38_read_addr__din;
  wire in_38_read_addr__full_n;
  wire in_38_read_addr__write;
  wire [255:0] in_38_read_data__dout;
  wire in_38_read_data__empty_n;
  wire in_38_read_data__read;
  wire [63:0] in_38_write_addr__din;
  wire in_38_write_addr__full_n;
  wire in_38_write_addr__write;
  wire [255:0] in_38_write_data__din;
  wire in_38_write_data__full_n;
  wire in_38_write_data__write;
  wire [7:0] in_38_write_resp__dout;
  wire in_38_write_resp__empty_n;
  wire in_38_write_resp__read;
  wire krnl_partialKnn_wrapper_38_0__ap_start;
  wire krnl_partialKnn_wrapper_38_0__ap_ready;
  wire krnl_partialKnn_wrapper_38_0__ap_done;
  wire krnl_partialKnn_wrapper_38_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_39_0___in_39__q0;
  wire [63:0] in_39_read_addr__din;
  wire in_39_read_addr__full_n;
  wire in_39_read_addr__write;
  wire [255:0] in_39_read_data__dout;
  wire in_39_read_data__empty_n;
  wire in_39_read_data__read;
  wire [63:0] in_39_write_addr__din;
  wire in_39_write_addr__full_n;
  wire in_39_write_addr__write;
  wire [255:0] in_39_write_data__din;
  wire in_39_write_data__full_n;
  wire in_39_write_data__write;
  wire [7:0] in_39_write_resp__dout;
  wire in_39_write_resp__empty_n;
  wire in_39_write_resp__read;
  wire krnl_partialKnn_wrapper_39_0__ap_start;
  wire krnl_partialKnn_wrapper_39_0__ap_ready;
  wire krnl_partialKnn_wrapper_39_0__ap_done;
  wire krnl_partialKnn_wrapper_39_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_4_0___in_4__q0;
  wire [63:0] in_4_read_addr__din;
  wire in_4_read_addr__full_n;
  wire in_4_read_addr__write;
  wire [255:0] in_4_read_data__dout;
  wire in_4_read_data__empty_n;
  wire in_4_read_data__read;
  wire [63:0] in_4_write_addr__din;
  wire in_4_write_addr__full_n;
  wire in_4_write_addr__write;
  wire [255:0] in_4_write_data__din;
  wire in_4_write_data__full_n;
  wire in_4_write_data__write;
  wire [7:0] in_4_write_resp__dout;
  wire in_4_write_resp__empty_n;
  wire in_4_write_resp__read;
  wire krnl_partialKnn_wrapper_4_0__ap_start;
  wire krnl_partialKnn_wrapper_4_0__ap_ready;
  wire krnl_partialKnn_wrapper_4_0__ap_done;
  wire krnl_partialKnn_wrapper_4_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_40_0___in_40__q0;
  wire [63:0] in_40_read_addr__din;
  wire in_40_read_addr__full_n;
  wire in_40_read_addr__write;
  wire [255:0] in_40_read_data__dout;
  wire in_40_read_data__empty_n;
  wire in_40_read_data__read;
  wire [63:0] in_40_write_addr__din;
  wire in_40_write_addr__full_n;
  wire in_40_write_addr__write;
  wire [255:0] in_40_write_data__din;
  wire in_40_write_data__full_n;
  wire in_40_write_data__write;
  wire [7:0] in_40_write_resp__dout;
  wire in_40_write_resp__empty_n;
  wire in_40_write_resp__read;
  wire krnl_partialKnn_wrapper_40_0__ap_start;
  wire krnl_partialKnn_wrapper_40_0__ap_ready;
  wire krnl_partialKnn_wrapper_40_0__ap_done;
  wire krnl_partialKnn_wrapper_40_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_41_0___in_41__q0;
  wire [63:0] in_41_read_addr__din;
  wire in_41_read_addr__full_n;
  wire in_41_read_addr__write;
  wire [255:0] in_41_read_data__dout;
  wire in_41_read_data__empty_n;
  wire in_41_read_data__read;
  wire [63:0] in_41_write_addr__din;
  wire in_41_write_addr__full_n;
  wire in_41_write_addr__write;
  wire [255:0] in_41_write_data__din;
  wire in_41_write_data__full_n;
  wire in_41_write_data__write;
  wire [7:0] in_41_write_resp__dout;
  wire in_41_write_resp__empty_n;
  wire in_41_write_resp__read;
  wire krnl_partialKnn_wrapper_41_0__ap_start;
  wire krnl_partialKnn_wrapper_41_0__ap_ready;
  wire krnl_partialKnn_wrapper_41_0__ap_done;
  wire krnl_partialKnn_wrapper_41_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_42_0___in_42__q0;
  wire [63:0] in_42_read_addr__din;
  wire in_42_read_addr__full_n;
  wire in_42_read_addr__write;
  wire [255:0] in_42_read_data__dout;
  wire in_42_read_data__empty_n;
  wire in_42_read_data__read;
  wire [63:0] in_42_write_addr__din;
  wire in_42_write_addr__full_n;
  wire in_42_write_addr__write;
  wire [255:0] in_42_write_data__din;
  wire in_42_write_data__full_n;
  wire in_42_write_data__write;
  wire [7:0] in_42_write_resp__dout;
  wire in_42_write_resp__empty_n;
  wire in_42_write_resp__read;
  wire krnl_partialKnn_wrapper_42_0__ap_start;
  wire krnl_partialKnn_wrapper_42_0__ap_ready;
  wire krnl_partialKnn_wrapper_42_0__ap_done;
  wire krnl_partialKnn_wrapper_42_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_43_0___in_43__q0;
  wire [63:0] in_43_read_addr__din;
  wire in_43_read_addr__full_n;
  wire in_43_read_addr__write;
  wire [255:0] in_43_read_data__dout;
  wire in_43_read_data__empty_n;
  wire in_43_read_data__read;
  wire [63:0] in_43_write_addr__din;
  wire in_43_write_addr__full_n;
  wire in_43_write_addr__write;
  wire [255:0] in_43_write_data__din;
  wire in_43_write_data__full_n;
  wire in_43_write_data__write;
  wire [7:0] in_43_write_resp__dout;
  wire in_43_write_resp__empty_n;
  wire in_43_write_resp__read;
  wire krnl_partialKnn_wrapper_43_0__ap_start;
  wire krnl_partialKnn_wrapper_43_0__ap_ready;
  wire krnl_partialKnn_wrapper_43_0__ap_done;
  wire krnl_partialKnn_wrapper_43_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_44_0___in_44__q0;
  wire [63:0] in_44_read_addr__din;
  wire in_44_read_addr__full_n;
  wire in_44_read_addr__write;
  wire [255:0] in_44_read_data__dout;
  wire in_44_read_data__empty_n;
  wire in_44_read_data__read;
  wire [63:0] in_44_write_addr__din;
  wire in_44_write_addr__full_n;
  wire in_44_write_addr__write;
  wire [255:0] in_44_write_data__din;
  wire in_44_write_data__full_n;
  wire in_44_write_data__write;
  wire [7:0] in_44_write_resp__dout;
  wire in_44_write_resp__empty_n;
  wire in_44_write_resp__read;
  wire krnl_partialKnn_wrapper_44_0__ap_start;
  wire krnl_partialKnn_wrapper_44_0__ap_ready;
  wire krnl_partialKnn_wrapper_44_0__ap_done;
  wire krnl_partialKnn_wrapper_44_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_45_0___in_45__q0;
  wire [63:0] in_45_read_addr__din;
  wire in_45_read_addr__full_n;
  wire in_45_read_addr__write;
  wire [255:0] in_45_read_data__dout;
  wire in_45_read_data__empty_n;
  wire in_45_read_data__read;
  wire [63:0] in_45_write_addr__din;
  wire in_45_write_addr__full_n;
  wire in_45_write_addr__write;
  wire [255:0] in_45_write_data__din;
  wire in_45_write_data__full_n;
  wire in_45_write_data__write;
  wire [7:0] in_45_write_resp__dout;
  wire in_45_write_resp__empty_n;
  wire in_45_write_resp__read;
  wire krnl_partialKnn_wrapper_45_0__ap_start;
  wire krnl_partialKnn_wrapper_45_0__ap_ready;
  wire krnl_partialKnn_wrapper_45_0__ap_done;
  wire krnl_partialKnn_wrapper_45_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_46_0___in_46__q0;
  wire [63:0] in_46_read_addr__din;
  wire in_46_read_addr__full_n;
  wire in_46_read_addr__write;
  wire [255:0] in_46_read_data__dout;
  wire in_46_read_data__empty_n;
  wire in_46_read_data__read;
  wire [63:0] in_46_write_addr__din;
  wire in_46_write_addr__full_n;
  wire in_46_write_addr__write;
  wire [255:0] in_46_write_data__din;
  wire in_46_write_data__full_n;
  wire in_46_write_data__write;
  wire [7:0] in_46_write_resp__dout;
  wire in_46_write_resp__empty_n;
  wire in_46_write_resp__read;
  wire krnl_partialKnn_wrapper_46_0__ap_start;
  wire krnl_partialKnn_wrapper_46_0__ap_ready;
  wire krnl_partialKnn_wrapper_46_0__ap_done;
  wire krnl_partialKnn_wrapper_46_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_47_0___in_47__q0;
  wire [63:0] in_47_read_addr__din;
  wire in_47_read_addr__full_n;
  wire in_47_read_addr__write;
  wire [255:0] in_47_read_data__dout;
  wire in_47_read_data__empty_n;
  wire in_47_read_data__read;
  wire [63:0] in_47_write_addr__din;
  wire in_47_write_addr__full_n;
  wire in_47_write_addr__write;
  wire [255:0] in_47_write_data__din;
  wire in_47_write_data__full_n;
  wire in_47_write_data__write;
  wire [7:0] in_47_write_resp__dout;
  wire in_47_write_resp__empty_n;
  wire in_47_write_resp__read;
  wire krnl_partialKnn_wrapper_47_0__ap_start;
  wire krnl_partialKnn_wrapper_47_0__ap_ready;
  wire krnl_partialKnn_wrapper_47_0__ap_done;
  wire krnl_partialKnn_wrapper_47_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_48_0___in_48__q0;
  wire [63:0] in_48_read_addr__din;
  wire in_48_read_addr__full_n;
  wire in_48_read_addr__write;
  wire [255:0] in_48_read_data__dout;
  wire in_48_read_data__empty_n;
  wire in_48_read_data__read;
  wire [63:0] in_48_write_addr__din;
  wire in_48_write_addr__full_n;
  wire in_48_write_addr__write;
  wire [255:0] in_48_write_data__din;
  wire in_48_write_data__full_n;
  wire in_48_write_data__write;
  wire [7:0] in_48_write_resp__dout;
  wire in_48_write_resp__empty_n;
  wire in_48_write_resp__read;
  wire krnl_partialKnn_wrapper_48_0__ap_start;
  wire krnl_partialKnn_wrapper_48_0__ap_ready;
  wire krnl_partialKnn_wrapper_48_0__ap_done;
  wire krnl_partialKnn_wrapper_48_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_49_0___in_49__q0;
  wire [63:0] in_49_read_addr__din;
  wire in_49_read_addr__full_n;
  wire in_49_read_addr__write;
  wire [255:0] in_49_read_data__dout;
  wire in_49_read_data__empty_n;
  wire in_49_read_data__read;
  wire [63:0] in_49_write_addr__din;
  wire in_49_write_addr__full_n;
  wire in_49_write_addr__write;
  wire [255:0] in_49_write_data__din;
  wire in_49_write_data__full_n;
  wire in_49_write_data__write;
  wire [7:0] in_49_write_resp__dout;
  wire in_49_write_resp__empty_n;
  wire in_49_write_resp__read;
  wire krnl_partialKnn_wrapper_49_0__ap_start;
  wire krnl_partialKnn_wrapper_49_0__ap_ready;
  wire krnl_partialKnn_wrapper_49_0__ap_done;
  wire krnl_partialKnn_wrapper_49_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_5_0___in_5__q0;
  wire [63:0] in_5_read_addr__din;
  wire in_5_read_addr__full_n;
  wire in_5_read_addr__write;
  wire [255:0] in_5_read_data__dout;
  wire in_5_read_data__empty_n;
  wire in_5_read_data__read;
  wire [63:0] in_5_write_addr__din;
  wire in_5_write_addr__full_n;
  wire in_5_write_addr__write;
  wire [255:0] in_5_write_data__din;
  wire in_5_write_data__full_n;
  wire in_5_write_data__write;
  wire [7:0] in_5_write_resp__dout;
  wire in_5_write_resp__empty_n;
  wire in_5_write_resp__read;
  wire krnl_partialKnn_wrapper_5_0__ap_start;
  wire krnl_partialKnn_wrapper_5_0__ap_ready;
  wire krnl_partialKnn_wrapper_5_0__ap_done;
  wire krnl_partialKnn_wrapper_5_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_50_0___in_50__q0;
  wire [63:0] in_50_read_addr__din;
  wire in_50_read_addr__full_n;
  wire in_50_read_addr__write;
  wire [255:0] in_50_read_data__dout;
  wire in_50_read_data__empty_n;
  wire in_50_read_data__read;
  wire [63:0] in_50_write_addr__din;
  wire in_50_write_addr__full_n;
  wire in_50_write_addr__write;
  wire [255:0] in_50_write_data__din;
  wire in_50_write_data__full_n;
  wire in_50_write_data__write;
  wire [7:0] in_50_write_resp__dout;
  wire in_50_write_resp__empty_n;
  wire in_50_write_resp__read;
  wire krnl_partialKnn_wrapper_50_0__ap_start;
  wire krnl_partialKnn_wrapper_50_0__ap_ready;
  wire krnl_partialKnn_wrapper_50_0__ap_done;
  wire krnl_partialKnn_wrapper_50_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_51_0___in_51__q0;
  wire [63:0] in_51_read_addr__din;
  wire in_51_read_addr__full_n;
  wire in_51_read_addr__write;
  wire [255:0] in_51_read_data__dout;
  wire in_51_read_data__empty_n;
  wire in_51_read_data__read;
  wire [63:0] in_51_write_addr__din;
  wire in_51_write_addr__full_n;
  wire in_51_write_addr__write;
  wire [255:0] in_51_write_data__din;
  wire in_51_write_data__full_n;
  wire in_51_write_data__write;
  wire [7:0] in_51_write_resp__dout;
  wire in_51_write_resp__empty_n;
  wire in_51_write_resp__read;
  wire krnl_partialKnn_wrapper_51_0__ap_start;
  wire krnl_partialKnn_wrapper_51_0__ap_ready;
  wire krnl_partialKnn_wrapper_51_0__ap_done;
  wire krnl_partialKnn_wrapper_51_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_52_0___in_52__q0;
  wire [63:0] in_52_read_addr__din;
  wire in_52_read_addr__full_n;
  wire in_52_read_addr__write;
  wire [255:0] in_52_read_data__dout;
  wire in_52_read_data__empty_n;
  wire in_52_read_data__read;
  wire [63:0] in_52_write_addr__din;
  wire in_52_write_addr__full_n;
  wire in_52_write_addr__write;
  wire [255:0] in_52_write_data__din;
  wire in_52_write_data__full_n;
  wire in_52_write_data__write;
  wire [7:0] in_52_write_resp__dout;
  wire in_52_write_resp__empty_n;
  wire in_52_write_resp__read;
  wire krnl_partialKnn_wrapper_52_0__ap_start;
  wire krnl_partialKnn_wrapper_52_0__ap_ready;
  wire krnl_partialKnn_wrapper_52_0__ap_done;
  wire krnl_partialKnn_wrapper_52_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_53_0___in_53__q0;
  wire [63:0] in_53_read_addr__din;
  wire in_53_read_addr__full_n;
  wire in_53_read_addr__write;
  wire [255:0] in_53_read_data__dout;
  wire in_53_read_data__empty_n;
  wire in_53_read_data__read;
  wire [63:0] in_53_write_addr__din;
  wire in_53_write_addr__full_n;
  wire in_53_write_addr__write;
  wire [255:0] in_53_write_data__din;
  wire in_53_write_data__full_n;
  wire in_53_write_data__write;
  wire [7:0] in_53_write_resp__dout;
  wire in_53_write_resp__empty_n;
  wire in_53_write_resp__read;
  wire krnl_partialKnn_wrapper_53_0__ap_start;
  wire krnl_partialKnn_wrapper_53_0__ap_ready;
  wire krnl_partialKnn_wrapper_53_0__ap_done;
  wire krnl_partialKnn_wrapper_53_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_6_0___in_6__q0;
  wire [63:0] in_6_read_addr__din;
  wire in_6_read_addr__full_n;
  wire in_6_read_addr__write;
  wire [255:0] in_6_read_data__dout;
  wire in_6_read_data__empty_n;
  wire in_6_read_data__read;
  wire [63:0] in_6_write_addr__din;
  wire in_6_write_addr__full_n;
  wire in_6_write_addr__write;
  wire [255:0] in_6_write_data__din;
  wire in_6_write_data__full_n;
  wire in_6_write_data__write;
  wire [7:0] in_6_write_resp__dout;
  wire in_6_write_resp__empty_n;
  wire in_6_write_resp__read;
  wire krnl_partialKnn_wrapper_6_0__ap_start;
  wire krnl_partialKnn_wrapper_6_0__ap_ready;
  wire krnl_partialKnn_wrapper_6_0__ap_done;
  wire krnl_partialKnn_wrapper_6_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_7_0___in_7__q0;
  wire [63:0] in_7_read_addr__din;
  wire in_7_read_addr__full_n;
  wire in_7_read_addr__write;
  wire [255:0] in_7_read_data__dout;
  wire in_7_read_data__empty_n;
  wire in_7_read_data__read;
  wire [63:0] in_7_write_addr__din;
  wire in_7_write_addr__full_n;
  wire in_7_write_addr__write;
  wire [255:0] in_7_write_data__din;
  wire in_7_write_data__full_n;
  wire in_7_write_data__write;
  wire [7:0] in_7_write_resp__dout;
  wire in_7_write_resp__empty_n;
  wire in_7_write_resp__read;
  wire krnl_partialKnn_wrapper_7_0__ap_start;
  wire krnl_partialKnn_wrapper_7_0__ap_ready;
  wire krnl_partialKnn_wrapper_7_0__ap_done;
  wire krnl_partialKnn_wrapper_7_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_8_0___in_8__q0;
  wire [63:0] in_8_read_addr__din;
  wire in_8_read_addr__full_n;
  wire in_8_read_addr__write;
  wire [255:0] in_8_read_data__dout;
  wire in_8_read_data__empty_n;
  wire in_8_read_data__read;
  wire [63:0] in_8_write_addr__din;
  wire in_8_write_addr__full_n;
  wire in_8_write_addr__write;
  wire [255:0] in_8_write_data__din;
  wire in_8_write_data__full_n;
  wire in_8_write_data__write;
  wire [7:0] in_8_write_resp__dout;
  wire in_8_write_resp__empty_n;
  wire in_8_write_resp__read;
  wire krnl_partialKnn_wrapper_8_0__ap_start;
  wire krnl_partialKnn_wrapper_8_0__ap_ready;
  wire krnl_partialKnn_wrapper_8_0__ap_done;
  wire krnl_partialKnn_wrapper_8_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_9_0___in_9__q0;
  wire [63:0] in_9_read_addr__din;
  wire in_9_read_addr__full_n;
  wire in_9_read_addr__write;
  wire [255:0] in_9_read_data__dout;
  wire in_9_read_data__empty_n;
  wire in_9_read_data__read;
  wire [63:0] in_9_write_addr__din;
  wire in_9_write_addr__full_n;
  wire in_9_write_addr__write;
  wire [255:0] in_9_write_data__din;
  wire in_9_write_data__full_n;
  wire in_9_write_data__write;
  wire [7:0] in_9_write_resp__dout;
  wire in_9_write_resp__empty_n;
  wire in_9_write_resp__read;
  wire krnl_partialKnn_wrapper_9_0__ap_start;
  wire krnl_partialKnn_wrapper_9_0__ap_ready;
  wire krnl_partialKnn_wrapper_9_0__ap_done;
  wire krnl_partialKnn_wrapper_9_0__ap_idle;
  wire ap_rst_n_inv;
  wire ap_done;
  wire ap_idle;
  wire ap_ready;
  assign ap_rst_n_inv = (~ap_rst_n);
  assign control_s_axi_U_ACLK = ap_clk;
  assign control_s_axi_U_ACLK_EN = 1'b1;
  assign control_s_axi_U_ARADDR = s_axi_control_ARADDR;
  assign control_s_axi_U_ARESET = ap_rst_n_inv;
  assign s_axi_control_ARREADY = control_s_axi_U_ARREADY;
  assign control_s_axi_U_ARVALID = s_axi_control_ARVALID;
  assign control_s_axi_U_AWADDR = s_axi_control_AWADDR;
  assign s_axi_control_AWREADY = control_s_axi_U_AWREADY;
  assign control_s_axi_U_AWVALID = s_axi_control_AWVALID;
  assign control_s_axi_U_BREADY = s_axi_control_BREADY;
  assign s_axi_control_BRESP = control_s_axi_U_BRESP;
  assign s_axi_control_BVALID = control_s_axi_U_BVALID;
  assign L4_out_dist = control_s_axi_U_L4_out_dist;
  assign L4_out_id = control_s_axi_U_L4_out_id;
  assign s_axi_control_RDATA = control_s_axi_U_RDATA;
  assign control_s_axi_U_RREADY = s_axi_control_RREADY;
  assign s_axi_control_RRESP = control_s_axi_U_RRESP;
  assign s_axi_control_RVALID = control_s_axi_U_RVALID;
  assign control_s_axi_U_WDATA = s_axi_control_WDATA;
  assign s_axi_control_WREADY = control_s_axi_U_WREADY;
  assign control_s_axi_U_WSTRB = s_axi_control_WSTRB;
  assign control_s_axi_U_WVALID = s_axi_control_WVALID;
  assign control_s_axi_U_ap_done = ap_done;
  assign control_s_axi_U_ap_idle = ap_idle;
  assign control_s_axi_U_ap_ready = ap_ready;
  assign ap_start = control_s_axi_U_ap_start;
  assign in_0 = control_s_axi_U_in_0;
  assign in_1 = control_s_axi_U_in_1;
  assign in_10 = control_s_axi_U_in_10;
  assign in_11 = control_s_axi_U_in_11;
  assign in_12 = control_s_axi_U_in_12;
  assign in_13 = control_s_axi_U_in_13;
  assign in_14 = control_s_axi_U_in_14;
  assign in_15 = control_s_axi_U_in_15;
  assign in_16 = control_s_axi_U_in_16;
  assign in_17 = control_s_axi_U_in_17;
  assign in_18 = control_s_axi_U_in_18;
  assign in_19 = control_s_axi_U_in_19;
  assign in_2 = control_s_axi_U_in_2;
  assign in_20 = control_s_axi_U_in_20;
  assign in_21 = control_s_axi_U_in_21;
  assign in_22 = control_s_axi_U_in_22;
  assign in_23 = control_s_axi_U_in_23;
  assign in_24 = control_s_axi_U_in_24;
  assign in_25 = control_s_axi_U_in_25;
  assign in_26 = control_s_axi_U_in_26;
  assign in_27 = control_s_axi_U_in_27;
  assign in_28 = control_s_axi_U_in_28;
  assign in_29 = control_s_axi_U_in_29;
  assign in_3 = control_s_axi_U_in_3;
  assign in_30 = control_s_axi_U_in_30;
  assign in_31 = control_s_axi_U_in_31;
  assign in_32 = control_s_axi_U_in_32;
  assign in_33 = control_s_axi_U_in_33;
  assign in_34 = control_s_axi_U_in_34;
  assign in_35 = control_s_axi_U_in_35;
  assign in_36 = control_s_axi_U_in_36;
  assign in_37 = control_s_axi_U_in_37;
  assign in_38 = control_s_axi_U_in_38;
  assign in_39 = control_s_axi_U_in_39;
  assign in_4 = control_s_axi_U_in_4;
  assign in_40 = control_s_axi_U_in_40;
  assign in_41 = control_s_axi_U_in_41;
  assign in_42 = control_s_axi_U_in_42;
  assign in_43 = control_s_axi_U_in_43;
  assign in_44 = control_s_axi_U_in_44;
  assign in_45 = control_s_axi_U_in_45;
  assign in_46 = control_s_axi_U_in_46;
  assign in_47 = control_s_axi_U_in_47;
  assign in_48 = control_s_axi_U_in_48;
  assign in_49 = control_s_axi_U_in_49;
  assign in_5 = control_s_axi_U_in_5;
  assign in_50 = control_s_axi_U_in_50;
  assign in_51 = control_s_axi_U_in_51;
  assign in_52 = control_s_axi_U_in_52;
  assign in_53 = control_s_axi_U_in_53;
  assign in_6 = control_s_axi_U_in_6;
  assign in_7 = control_s_axi_U_in_7;
  assign in_8 = control_s_axi_U_in_8;
  assign in_9 = control_s_axi_U_in_9;
  assign interrupt = control_s_axi_U_interrupt;
  assign L1_out_dist_0_clk = ap_clk;
  assign L1_out_dist_0_if_din = L1_out_dist_0__din;
  assign L1_out_dist_0__dout = L1_out_dist_0_if_dout;
  assign L1_out_dist_0__empty_n = L1_out_dist_0_if_empty_n;
  assign L1_out_dist_0__full_n = L1_out_dist_0_if_full_n;
  assign L1_out_dist_0_if_read = L1_out_dist_0__read;
  assign L1_out_dist_0_if_read_ce = 1'b1;
  assign L1_out_dist_0_if_write = L1_out_dist_0__write;
  assign L1_out_dist_0_if_write_ce = 1'b1;
  assign L1_out_dist_0_reset = ~ ap_rst_n;
  assign L1_out_dist_10_clk = ap_clk;
  assign L1_out_dist_10_if_din = L1_out_dist_10__din;
  assign L1_out_dist_10__dout = L1_out_dist_10_if_dout;
  assign L1_out_dist_10__empty_n = L1_out_dist_10_if_empty_n;
  assign L1_out_dist_10__full_n = L1_out_dist_10_if_full_n;
  assign L1_out_dist_10_if_read = L1_out_dist_10__read;
  assign L1_out_dist_10_if_read_ce = 1'b1;
  assign L1_out_dist_10_if_write = L1_out_dist_10__write;
  assign L1_out_dist_10_if_write_ce = 1'b1;
  assign L1_out_dist_10_reset = ~ ap_rst_n;
  assign L1_out_dist_11_clk = ap_clk;
  assign L1_out_dist_11_if_din = L1_out_dist_11__din;
  assign L1_out_dist_11__dout = L1_out_dist_11_if_dout;
  assign L1_out_dist_11__empty_n = L1_out_dist_11_if_empty_n;
  assign L1_out_dist_11__full_n = L1_out_dist_11_if_full_n;
  assign L1_out_dist_11_if_read = L1_out_dist_11__read;
  assign L1_out_dist_11_if_read_ce = 1'b1;
  assign L1_out_dist_11_if_write = L1_out_dist_11__write;
  assign L1_out_dist_11_if_write_ce = 1'b1;
  assign L1_out_dist_11_reset = ~ ap_rst_n;
  assign L1_out_dist_12_clk = ap_clk;
  assign L1_out_dist_12_if_din = L1_out_dist_12__din;
  assign L1_out_dist_12__dout = L1_out_dist_12_if_dout;
  assign L1_out_dist_12__empty_n = L1_out_dist_12_if_empty_n;
  assign L1_out_dist_12__full_n = L1_out_dist_12_if_full_n;
  assign L1_out_dist_12_if_read = L1_out_dist_12__read;
  assign L1_out_dist_12_if_read_ce = 1'b1;
  assign L1_out_dist_12_if_write = L1_out_dist_12__write;
  assign L1_out_dist_12_if_write_ce = 1'b1;
  assign L1_out_dist_12_reset = ~ ap_rst_n;
  assign L1_out_dist_13_clk = ap_clk;
  assign L1_out_dist_13_if_din = L1_out_dist_13__din;
  assign L1_out_dist_13__dout = L1_out_dist_13_if_dout;
  assign L1_out_dist_13__empty_n = L1_out_dist_13_if_empty_n;
  assign L1_out_dist_13__full_n = L1_out_dist_13_if_full_n;
  assign L1_out_dist_13_if_read = L1_out_dist_13__read;
  assign L1_out_dist_13_if_read_ce = 1'b1;
  assign L1_out_dist_13_if_write = L1_out_dist_13__write;
  assign L1_out_dist_13_if_write_ce = 1'b1;
  assign L1_out_dist_13_reset = ~ ap_rst_n;
  assign L1_out_dist_14_clk = ap_clk;
  assign L1_out_dist_14_if_din = L1_out_dist_14__din;
  assign L1_out_dist_14__dout = L1_out_dist_14_if_dout;
  assign L1_out_dist_14__empty_n = L1_out_dist_14_if_empty_n;
  assign L1_out_dist_14__full_n = L1_out_dist_14_if_full_n;
  assign L1_out_dist_14_if_read = L1_out_dist_14__read;
  assign L1_out_dist_14_if_read_ce = 1'b1;
  assign L1_out_dist_14_if_write = L1_out_dist_14__write;
  assign L1_out_dist_14_if_write_ce = 1'b1;
  assign L1_out_dist_14_reset = ~ ap_rst_n;
  assign L1_out_dist_15_clk = ap_clk;
  assign L1_out_dist_15_if_din = L1_out_dist_15__din;
  assign L1_out_dist_15__dout = L1_out_dist_15_if_dout;
  assign L1_out_dist_15__empty_n = L1_out_dist_15_if_empty_n;
  assign L1_out_dist_15__full_n = L1_out_dist_15_if_full_n;
  assign L1_out_dist_15_if_read = L1_out_dist_15__read;
  assign L1_out_dist_15_if_read_ce = 1'b1;
  assign L1_out_dist_15_if_write = L1_out_dist_15__write;
  assign L1_out_dist_15_if_write_ce = 1'b1;
  assign L1_out_dist_15_reset = ~ ap_rst_n;
  assign L1_out_dist_16_clk = ap_clk;
  assign L1_out_dist_16_if_din = L1_out_dist_16__din;
  assign L1_out_dist_16__dout = L1_out_dist_16_if_dout;
  assign L1_out_dist_16__empty_n = L1_out_dist_16_if_empty_n;
  assign L1_out_dist_16__full_n = L1_out_dist_16_if_full_n;
  assign L1_out_dist_16_if_read = L1_out_dist_16__read;
  assign L1_out_dist_16_if_read_ce = 1'b1;
  assign L1_out_dist_16_if_write = L1_out_dist_16__write;
  assign L1_out_dist_16_if_write_ce = 1'b1;
  assign L1_out_dist_16_reset = ~ ap_rst_n;
  assign L1_out_dist_17_clk = ap_clk;
  assign L1_out_dist_17_if_din = L1_out_dist_17__din;
  assign L1_out_dist_17__dout = L1_out_dist_17_if_dout;
  assign L1_out_dist_17__empty_n = L1_out_dist_17_if_empty_n;
  assign L1_out_dist_17__full_n = L1_out_dist_17_if_full_n;
  assign L1_out_dist_17_if_read = L1_out_dist_17__read;
  assign L1_out_dist_17_if_read_ce = 1'b1;
  assign L1_out_dist_17_if_write = L1_out_dist_17__write;
  assign L1_out_dist_17_if_write_ce = 1'b1;
  assign L1_out_dist_17_reset = ~ ap_rst_n;
  assign L1_out_dist_1_clk = ap_clk;
  assign L1_out_dist_1_if_din = L1_out_dist_1__din;
  assign L1_out_dist_1__dout = L1_out_dist_1_if_dout;
  assign L1_out_dist_1__empty_n = L1_out_dist_1_if_empty_n;
  assign L1_out_dist_1__full_n = L1_out_dist_1_if_full_n;
  assign L1_out_dist_1_if_read = L1_out_dist_1__read;
  assign L1_out_dist_1_if_read_ce = 1'b1;
  assign L1_out_dist_1_if_write = L1_out_dist_1__write;
  assign L1_out_dist_1_if_write_ce = 1'b1;
  assign L1_out_dist_1_reset = ~ ap_rst_n;
  assign L1_out_dist_2_clk = ap_clk;
  assign L1_out_dist_2_if_din = L1_out_dist_2__din;
  assign L1_out_dist_2__dout = L1_out_dist_2_if_dout;
  assign L1_out_dist_2__empty_n = L1_out_dist_2_if_empty_n;
  assign L1_out_dist_2__full_n = L1_out_dist_2_if_full_n;
  assign L1_out_dist_2_if_read = L1_out_dist_2__read;
  assign L1_out_dist_2_if_read_ce = 1'b1;
  assign L1_out_dist_2_if_write = L1_out_dist_2__write;
  assign L1_out_dist_2_if_write_ce = 1'b1;
  assign L1_out_dist_2_reset = ~ ap_rst_n;
  assign L1_out_dist_3_clk = ap_clk;
  assign L1_out_dist_3_if_din = L1_out_dist_3__din;
  assign L1_out_dist_3__dout = L1_out_dist_3_if_dout;
  assign L1_out_dist_3__empty_n = L1_out_dist_3_if_empty_n;
  assign L1_out_dist_3__full_n = L1_out_dist_3_if_full_n;
  assign L1_out_dist_3_if_read = L1_out_dist_3__read;
  assign L1_out_dist_3_if_read_ce = 1'b1;
  assign L1_out_dist_3_if_write = L1_out_dist_3__write;
  assign L1_out_dist_3_if_write_ce = 1'b1;
  assign L1_out_dist_3_reset = ~ ap_rst_n;
  assign L1_out_dist_4_clk = ap_clk;
  assign L1_out_dist_4_if_din = L1_out_dist_4__din;
  assign L1_out_dist_4__dout = L1_out_dist_4_if_dout;
  assign L1_out_dist_4__empty_n = L1_out_dist_4_if_empty_n;
  assign L1_out_dist_4__full_n = L1_out_dist_4_if_full_n;
  assign L1_out_dist_4_if_read = L1_out_dist_4__read;
  assign L1_out_dist_4_if_read_ce = 1'b1;
  assign L1_out_dist_4_if_write = L1_out_dist_4__write;
  assign L1_out_dist_4_if_write_ce = 1'b1;
  assign L1_out_dist_4_reset = ~ ap_rst_n;
  assign L1_out_dist_5_clk = ap_clk;
  assign L1_out_dist_5_if_din = L1_out_dist_5__din;
  assign L1_out_dist_5__dout = L1_out_dist_5_if_dout;
  assign L1_out_dist_5__empty_n = L1_out_dist_5_if_empty_n;
  assign L1_out_dist_5__full_n = L1_out_dist_5_if_full_n;
  assign L1_out_dist_5_if_read = L1_out_dist_5__read;
  assign L1_out_dist_5_if_read_ce = 1'b1;
  assign L1_out_dist_5_if_write = L1_out_dist_5__write;
  assign L1_out_dist_5_if_write_ce = 1'b1;
  assign L1_out_dist_5_reset = ~ ap_rst_n;
  assign L1_out_dist_6_clk = ap_clk;
  assign L1_out_dist_6_if_din = L1_out_dist_6__din;
  assign L1_out_dist_6__dout = L1_out_dist_6_if_dout;
  assign L1_out_dist_6__empty_n = L1_out_dist_6_if_empty_n;
  assign L1_out_dist_6__full_n = L1_out_dist_6_if_full_n;
  assign L1_out_dist_6_if_read = L1_out_dist_6__read;
  assign L1_out_dist_6_if_read_ce = 1'b1;
  assign L1_out_dist_6_if_write = L1_out_dist_6__write;
  assign L1_out_dist_6_if_write_ce = 1'b1;
  assign L1_out_dist_6_reset = ~ ap_rst_n;
  assign L1_out_dist_7_clk = ap_clk;
  assign L1_out_dist_7_if_din = L1_out_dist_7__din;
  assign L1_out_dist_7__dout = L1_out_dist_7_if_dout;
  assign L1_out_dist_7__empty_n = L1_out_dist_7_if_empty_n;
  assign L1_out_dist_7__full_n = L1_out_dist_7_if_full_n;
  assign L1_out_dist_7_if_read = L1_out_dist_7__read;
  assign L1_out_dist_7_if_read_ce = 1'b1;
  assign L1_out_dist_7_if_write = L1_out_dist_7__write;
  assign L1_out_dist_7_if_write_ce = 1'b1;
  assign L1_out_dist_7_reset = ~ ap_rst_n;
  assign L1_out_dist_8_clk = ap_clk;
  assign L1_out_dist_8_if_din = L1_out_dist_8__din;
  assign L1_out_dist_8__dout = L1_out_dist_8_if_dout;
  assign L1_out_dist_8__empty_n = L1_out_dist_8_if_empty_n;
  assign L1_out_dist_8__full_n = L1_out_dist_8_if_full_n;
  assign L1_out_dist_8_if_read = L1_out_dist_8__read;
  assign L1_out_dist_8_if_read_ce = 1'b1;
  assign L1_out_dist_8_if_write = L1_out_dist_8__write;
  assign L1_out_dist_8_if_write_ce = 1'b1;
  assign L1_out_dist_8_reset = ~ ap_rst_n;
  assign L1_out_dist_9_clk = ap_clk;
  assign L1_out_dist_9_if_din = L1_out_dist_9__din;
  assign L1_out_dist_9__dout = L1_out_dist_9_if_dout;
  assign L1_out_dist_9__empty_n = L1_out_dist_9_if_empty_n;
  assign L1_out_dist_9__full_n = L1_out_dist_9_if_full_n;
  assign L1_out_dist_9_if_read = L1_out_dist_9__read;
  assign L1_out_dist_9_if_read_ce = 1'b1;
  assign L1_out_dist_9_if_write = L1_out_dist_9__write;
  assign L1_out_dist_9_if_write_ce = 1'b1;
  assign L1_out_dist_9_reset = ~ ap_rst_n;
  assign L1_out_id_0_clk = ap_clk;
  assign L1_out_id_0_if_din = L1_out_id_0__din;
  assign L1_out_id_0__dout = L1_out_id_0_if_dout;
  assign L1_out_id_0__empty_n = L1_out_id_0_if_empty_n;
  assign L1_out_id_0__full_n = L1_out_id_0_if_full_n;
  assign L1_out_id_0_if_read = L1_out_id_0__read;
  assign L1_out_id_0_if_read_ce = 1'b1;
  assign L1_out_id_0_if_write = L1_out_id_0__write;
  assign L1_out_id_0_if_write_ce = 1'b1;
  assign L1_out_id_0_reset = ~ ap_rst_n;
  assign L1_out_id_10_clk = ap_clk;
  assign L1_out_id_10_if_din = L1_out_id_10__din;
  assign L1_out_id_10__dout = L1_out_id_10_if_dout;
  assign L1_out_id_10__empty_n = L1_out_id_10_if_empty_n;
  assign L1_out_id_10__full_n = L1_out_id_10_if_full_n;
  assign L1_out_id_10_if_read = L1_out_id_10__read;
  assign L1_out_id_10_if_read_ce = 1'b1;
  assign L1_out_id_10_if_write = L1_out_id_10__write;
  assign L1_out_id_10_if_write_ce = 1'b1;
  assign L1_out_id_10_reset = ~ ap_rst_n;
  assign L1_out_id_11_clk = ap_clk;
  assign L1_out_id_11_if_din = L1_out_id_11__din;
  assign L1_out_id_11__dout = L1_out_id_11_if_dout;
  assign L1_out_id_11__empty_n = L1_out_id_11_if_empty_n;
  assign L1_out_id_11__full_n = L1_out_id_11_if_full_n;
  assign L1_out_id_11_if_read = L1_out_id_11__read;
  assign L1_out_id_11_if_read_ce = 1'b1;
  assign L1_out_id_11_if_write = L1_out_id_11__write;
  assign L1_out_id_11_if_write_ce = 1'b1;
  assign L1_out_id_11_reset = ~ ap_rst_n;
  assign L1_out_id_12_clk = ap_clk;
  assign L1_out_id_12_if_din = L1_out_id_12__din;
  assign L1_out_id_12__dout = L1_out_id_12_if_dout;
  assign L1_out_id_12__empty_n = L1_out_id_12_if_empty_n;
  assign L1_out_id_12__full_n = L1_out_id_12_if_full_n;
  assign L1_out_id_12_if_read = L1_out_id_12__read;
  assign L1_out_id_12_if_read_ce = 1'b1;
  assign L1_out_id_12_if_write = L1_out_id_12__write;
  assign L1_out_id_12_if_write_ce = 1'b1;
  assign L1_out_id_12_reset = ~ ap_rst_n;
  assign L1_out_id_13_clk = ap_clk;
  assign L1_out_id_13_if_din = L1_out_id_13__din;
  assign L1_out_id_13__dout = L1_out_id_13_if_dout;
  assign L1_out_id_13__empty_n = L1_out_id_13_if_empty_n;
  assign L1_out_id_13__full_n = L1_out_id_13_if_full_n;
  assign L1_out_id_13_if_read = L1_out_id_13__read;
  assign L1_out_id_13_if_read_ce = 1'b1;
  assign L1_out_id_13_if_write = L1_out_id_13__write;
  assign L1_out_id_13_if_write_ce = 1'b1;
  assign L1_out_id_13_reset = ~ ap_rst_n;
  assign L1_out_id_14_clk = ap_clk;
  assign L1_out_id_14_if_din = L1_out_id_14__din;
  assign L1_out_id_14__dout = L1_out_id_14_if_dout;
  assign L1_out_id_14__empty_n = L1_out_id_14_if_empty_n;
  assign L1_out_id_14__full_n = L1_out_id_14_if_full_n;
  assign L1_out_id_14_if_read = L1_out_id_14__read;
  assign L1_out_id_14_if_read_ce = 1'b1;
  assign L1_out_id_14_if_write = L1_out_id_14__write;
  assign L1_out_id_14_if_write_ce = 1'b1;
  assign L1_out_id_14_reset = ~ ap_rst_n;
  assign L1_out_id_15_clk = ap_clk;
  assign L1_out_id_15_if_din = L1_out_id_15__din;
  assign L1_out_id_15__dout = L1_out_id_15_if_dout;
  assign L1_out_id_15__empty_n = L1_out_id_15_if_empty_n;
  assign L1_out_id_15__full_n = L1_out_id_15_if_full_n;
  assign L1_out_id_15_if_read = L1_out_id_15__read;
  assign L1_out_id_15_if_read_ce = 1'b1;
  assign L1_out_id_15_if_write = L1_out_id_15__write;
  assign L1_out_id_15_if_write_ce = 1'b1;
  assign L1_out_id_15_reset = ~ ap_rst_n;
  assign L1_out_id_16_clk = ap_clk;
  assign L1_out_id_16_if_din = L1_out_id_16__din;
  assign L1_out_id_16__dout = L1_out_id_16_if_dout;
  assign L1_out_id_16__empty_n = L1_out_id_16_if_empty_n;
  assign L1_out_id_16__full_n = L1_out_id_16_if_full_n;
  assign L1_out_id_16_if_read = L1_out_id_16__read;
  assign L1_out_id_16_if_read_ce = 1'b1;
  assign L1_out_id_16_if_write = L1_out_id_16__write;
  assign L1_out_id_16_if_write_ce = 1'b1;
  assign L1_out_id_16_reset = ~ ap_rst_n;
  assign L1_out_id_17_clk = ap_clk;
  assign L1_out_id_17_if_din = L1_out_id_17__din;
  assign L1_out_id_17__dout = L1_out_id_17_if_dout;
  assign L1_out_id_17__empty_n = L1_out_id_17_if_empty_n;
  assign L1_out_id_17__full_n = L1_out_id_17_if_full_n;
  assign L1_out_id_17_if_read = L1_out_id_17__read;
  assign L1_out_id_17_if_read_ce = 1'b1;
  assign L1_out_id_17_if_write = L1_out_id_17__write;
  assign L1_out_id_17_if_write_ce = 1'b1;
  assign L1_out_id_17_reset = ~ ap_rst_n;
  assign L1_out_id_1_clk = ap_clk;
  assign L1_out_id_1_if_din = L1_out_id_1__din;
  assign L1_out_id_1__dout = L1_out_id_1_if_dout;
  assign L1_out_id_1__empty_n = L1_out_id_1_if_empty_n;
  assign L1_out_id_1__full_n = L1_out_id_1_if_full_n;
  assign L1_out_id_1_if_read = L1_out_id_1__read;
  assign L1_out_id_1_if_read_ce = 1'b1;
  assign L1_out_id_1_if_write = L1_out_id_1__write;
  assign L1_out_id_1_if_write_ce = 1'b1;
  assign L1_out_id_1_reset = ~ ap_rst_n;
  assign L1_out_id_2_clk = ap_clk;
  assign L1_out_id_2_if_din = L1_out_id_2__din;
  assign L1_out_id_2__dout = L1_out_id_2_if_dout;
  assign L1_out_id_2__empty_n = L1_out_id_2_if_empty_n;
  assign L1_out_id_2__full_n = L1_out_id_2_if_full_n;
  assign L1_out_id_2_if_read = L1_out_id_2__read;
  assign L1_out_id_2_if_read_ce = 1'b1;
  assign L1_out_id_2_if_write = L1_out_id_2__write;
  assign L1_out_id_2_if_write_ce = 1'b1;
  assign L1_out_id_2_reset = ~ ap_rst_n;
  assign L1_out_id_3_clk = ap_clk;
  assign L1_out_id_3_if_din = L1_out_id_3__din;
  assign L1_out_id_3__dout = L1_out_id_3_if_dout;
  assign L1_out_id_3__empty_n = L1_out_id_3_if_empty_n;
  assign L1_out_id_3__full_n = L1_out_id_3_if_full_n;
  assign L1_out_id_3_if_read = L1_out_id_3__read;
  assign L1_out_id_3_if_read_ce = 1'b1;
  assign L1_out_id_3_if_write = L1_out_id_3__write;
  assign L1_out_id_3_if_write_ce = 1'b1;
  assign L1_out_id_3_reset = ~ ap_rst_n;
  assign L1_out_id_4_clk = ap_clk;
  assign L1_out_id_4_if_din = L1_out_id_4__din;
  assign L1_out_id_4__dout = L1_out_id_4_if_dout;
  assign L1_out_id_4__empty_n = L1_out_id_4_if_empty_n;
  assign L1_out_id_4__full_n = L1_out_id_4_if_full_n;
  assign L1_out_id_4_if_read = L1_out_id_4__read;
  assign L1_out_id_4_if_read_ce = 1'b1;
  assign L1_out_id_4_if_write = L1_out_id_4__write;
  assign L1_out_id_4_if_write_ce = 1'b1;
  assign L1_out_id_4_reset = ~ ap_rst_n;
  assign L1_out_id_5_clk = ap_clk;
  assign L1_out_id_5_if_din = L1_out_id_5__din;
  assign L1_out_id_5__dout = L1_out_id_5_if_dout;
  assign L1_out_id_5__empty_n = L1_out_id_5_if_empty_n;
  assign L1_out_id_5__full_n = L1_out_id_5_if_full_n;
  assign L1_out_id_5_if_read = L1_out_id_5__read;
  assign L1_out_id_5_if_read_ce = 1'b1;
  assign L1_out_id_5_if_write = L1_out_id_5__write;
  assign L1_out_id_5_if_write_ce = 1'b1;
  assign L1_out_id_5_reset = ~ ap_rst_n;
  assign L1_out_id_6_clk = ap_clk;
  assign L1_out_id_6_if_din = L1_out_id_6__din;
  assign L1_out_id_6__dout = L1_out_id_6_if_dout;
  assign L1_out_id_6__empty_n = L1_out_id_6_if_empty_n;
  assign L1_out_id_6__full_n = L1_out_id_6_if_full_n;
  assign L1_out_id_6_if_read = L1_out_id_6__read;
  assign L1_out_id_6_if_read_ce = 1'b1;
  assign L1_out_id_6_if_write = L1_out_id_6__write;
  assign L1_out_id_6_if_write_ce = 1'b1;
  assign L1_out_id_6_reset = ~ ap_rst_n;
  assign L1_out_id_7_clk = ap_clk;
  assign L1_out_id_7_if_din = L1_out_id_7__din;
  assign L1_out_id_7__dout = L1_out_id_7_if_dout;
  assign L1_out_id_7__empty_n = L1_out_id_7_if_empty_n;
  assign L1_out_id_7__full_n = L1_out_id_7_if_full_n;
  assign L1_out_id_7_if_read = L1_out_id_7__read;
  assign L1_out_id_7_if_read_ce = 1'b1;
  assign L1_out_id_7_if_write = L1_out_id_7__write;
  assign L1_out_id_7_if_write_ce = 1'b1;
  assign L1_out_id_7_reset = ~ ap_rst_n;
  assign L1_out_id_8_clk = ap_clk;
  assign L1_out_id_8_if_din = L1_out_id_8__din;
  assign L1_out_id_8__dout = L1_out_id_8_if_dout;
  assign L1_out_id_8__empty_n = L1_out_id_8_if_empty_n;
  assign L1_out_id_8__full_n = L1_out_id_8_if_full_n;
  assign L1_out_id_8_if_read = L1_out_id_8__read;
  assign L1_out_id_8_if_read_ce = 1'b1;
  assign L1_out_id_8_if_write = L1_out_id_8__write;
  assign L1_out_id_8_if_write_ce = 1'b1;
  assign L1_out_id_8_reset = ~ ap_rst_n;
  assign L1_out_id_9_clk = ap_clk;
  assign L1_out_id_9_if_din = L1_out_id_9__din;
  assign L1_out_id_9__dout = L1_out_id_9_if_dout;
  assign L1_out_id_9__empty_n = L1_out_id_9_if_empty_n;
  assign L1_out_id_9__full_n = L1_out_id_9_if_full_n;
  assign L1_out_id_9_if_read = L1_out_id_9__read;
  assign L1_out_id_9_if_read_ce = 1'b1;
  assign L1_out_id_9_if_write = L1_out_id_9__write;
  assign L1_out_id_9_if_write_ce = 1'b1;
  assign L1_out_id_9_reset = ~ ap_rst_n;
  assign L2_out_dist0_clk = ap_clk;
  assign L2_out_dist0_if_din = L2_out_dist0__din;
  assign L2_out_dist0__dout = L2_out_dist0_if_dout;
  assign L2_out_dist0__empty_n = L2_out_dist0_if_empty_n;
  assign L2_out_dist0__full_n = L2_out_dist0_if_full_n;
  assign L2_out_dist0_if_read = L2_out_dist0__read;
  assign L2_out_dist0_if_read_ce = 1'b1;
  assign L2_out_dist0_if_write = L2_out_dist0__write;
  assign L2_out_dist0_if_write_ce = 1'b1;
  assign L2_out_dist0_reset = ~ ap_rst_n;
  assign L2_out_dist1_clk = ap_clk;
  assign L2_out_dist1_if_din = L2_out_dist1__din;
  assign L2_out_dist1__dout = L2_out_dist1_if_dout;
  assign L2_out_dist1__empty_n = L2_out_dist1_if_empty_n;
  assign L2_out_dist1__full_n = L2_out_dist1_if_full_n;
  assign L2_out_dist1_if_read = L2_out_dist1__read;
  assign L2_out_dist1_if_read_ce = 1'b1;
  assign L2_out_dist1_if_write = L2_out_dist1__write;
  assign L2_out_dist1_if_write_ce = 1'b1;
  assign L2_out_dist1_reset = ~ ap_rst_n;
  assign L2_out_dist2_clk = ap_clk;
  assign L2_out_dist2_if_din = L2_out_dist2__din;
  assign L2_out_dist2__dout = L2_out_dist2_if_dout;
  assign L2_out_dist2__empty_n = L2_out_dist2_if_empty_n;
  assign L2_out_dist2__full_n = L2_out_dist2_if_full_n;
  assign L2_out_dist2_if_read = L2_out_dist2__read;
  assign L2_out_dist2_if_read_ce = 1'b1;
  assign L2_out_dist2_if_write = L2_out_dist2__write;
  assign L2_out_dist2_if_write_ce = 1'b1;
  assign L2_out_dist2_reset = ~ ap_rst_n;
  assign L2_out_dist3_clk = ap_clk;
  assign L2_out_dist3_if_din = L2_out_dist3__din;
  assign L2_out_dist3__dout = L2_out_dist3_if_dout;
  assign L2_out_dist3__empty_n = L2_out_dist3_if_empty_n;
  assign L2_out_dist3__full_n = L2_out_dist3_if_full_n;
  assign L2_out_dist3_if_read = L2_out_dist3__read;
  assign L2_out_dist3_if_read_ce = 1'b1;
  assign L2_out_dist3_if_write = L2_out_dist3__write;
  assign L2_out_dist3_if_write_ce = 1'b1;
  assign L2_out_dist3_reset = ~ ap_rst_n;
  assign L2_out_dist4_clk = ap_clk;
  assign L2_out_dist4_if_din = L2_out_dist4__din;
  assign L2_out_dist4__dout = L2_out_dist4_if_dout;
  assign L2_out_dist4__empty_n = L2_out_dist4_if_empty_n;
  assign L2_out_dist4__full_n = L2_out_dist4_if_full_n;
  assign L2_out_dist4_if_read = L2_out_dist4__read;
  assign L2_out_dist4_if_read_ce = 1'b1;
  assign L2_out_dist4_if_write = L2_out_dist4__write;
  assign L2_out_dist4_if_write_ce = 1'b1;
  assign L2_out_dist4_reset = ~ ap_rst_n;
  assign L2_out_dist5_clk = ap_clk;
  assign L2_out_dist5_if_din = L2_out_dist5__din;
  assign L2_out_dist5__dout = L2_out_dist5_if_dout;
  assign L2_out_dist5__empty_n = L2_out_dist5_if_empty_n;
  assign L2_out_dist5__full_n = L2_out_dist5_if_full_n;
  assign L2_out_dist5_if_read = L2_out_dist5__read;
  assign L2_out_dist5_if_read_ce = 1'b1;
  assign L2_out_dist5_if_write = L2_out_dist5__write;
  assign L2_out_dist5_if_write_ce = 1'b1;
  assign L2_out_dist5_reset = ~ ap_rst_n;
  assign L2_out_id0_clk = ap_clk;
  assign L2_out_id0_if_din = L2_out_id0__din;
  assign L2_out_id0__dout = L2_out_id0_if_dout;
  assign L2_out_id0__empty_n = L2_out_id0_if_empty_n;
  assign L2_out_id0__full_n = L2_out_id0_if_full_n;
  assign L2_out_id0_if_read = L2_out_id0__read;
  assign L2_out_id0_if_read_ce = 1'b1;
  assign L2_out_id0_if_write = L2_out_id0__write;
  assign L2_out_id0_if_write_ce = 1'b1;
  assign L2_out_id0_reset = ~ ap_rst_n;
  assign L2_out_id1_clk = ap_clk;
  assign L2_out_id1_if_din = L2_out_id1__din;
  assign L2_out_id1__dout = L2_out_id1_if_dout;
  assign L2_out_id1__empty_n = L2_out_id1_if_empty_n;
  assign L2_out_id1__full_n = L2_out_id1_if_full_n;
  assign L2_out_id1_if_read = L2_out_id1__read;
  assign L2_out_id1_if_read_ce = 1'b1;
  assign L2_out_id1_if_write = L2_out_id1__write;
  assign L2_out_id1_if_write_ce = 1'b1;
  assign L2_out_id1_reset = ~ ap_rst_n;
  assign L2_out_id2_clk = ap_clk;
  assign L2_out_id2_if_din = L2_out_id2__din;
  assign L2_out_id2__dout = L2_out_id2_if_dout;
  assign L2_out_id2__empty_n = L2_out_id2_if_empty_n;
  assign L2_out_id2__full_n = L2_out_id2_if_full_n;
  assign L2_out_id2_if_read = L2_out_id2__read;
  assign L2_out_id2_if_read_ce = 1'b1;
  assign L2_out_id2_if_write = L2_out_id2__write;
  assign L2_out_id2_if_write_ce = 1'b1;
  assign L2_out_id2_reset = ~ ap_rst_n;
  assign L2_out_id3_clk = ap_clk;
  assign L2_out_id3_if_din = L2_out_id3__din;
  assign L2_out_id3__dout = L2_out_id3_if_dout;
  assign L2_out_id3__empty_n = L2_out_id3_if_empty_n;
  assign L2_out_id3__full_n = L2_out_id3_if_full_n;
  assign L2_out_id3_if_read = L2_out_id3__read;
  assign L2_out_id3_if_read_ce = 1'b1;
  assign L2_out_id3_if_write = L2_out_id3__write;
  assign L2_out_id3_if_write_ce = 1'b1;
  assign L2_out_id3_reset = ~ ap_rst_n;
  assign L2_out_id4_clk = ap_clk;
  assign L2_out_id4_if_din = L2_out_id4__din;
  assign L2_out_id4__dout = L2_out_id4_if_dout;
  assign L2_out_id4__empty_n = L2_out_id4_if_empty_n;
  assign L2_out_id4__full_n = L2_out_id4_if_full_n;
  assign L2_out_id4_if_read = L2_out_id4__read;
  assign L2_out_id4_if_read_ce = 1'b1;
  assign L2_out_id4_if_write = L2_out_id4__write;
  assign L2_out_id4_if_write_ce = 1'b1;
  assign L2_out_id4_reset = ~ ap_rst_n;
  assign L2_out_id5_clk = ap_clk;
  assign L2_out_id5_if_din = L2_out_id5__din;
  assign L2_out_id5__dout = L2_out_id5_if_dout;
  assign L2_out_id5__empty_n = L2_out_id5_if_empty_n;
  assign L2_out_id5__full_n = L2_out_id5_if_full_n;
  assign L2_out_id5_if_read = L2_out_id5__read;
  assign L2_out_id5_if_read_ce = 1'b1;
  assign L2_out_id5_if_write = L2_out_id5__write;
  assign L2_out_id5_if_write_ce = 1'b1;
  assign L2_out_id5_reset = ~ ap_rst_n;
  assign L3_out_dist0_clk = ap_clk;
  assign L3_out_dist0_if_din = L3_out_dist0__din;
  assign L3_out_dist0__dout = L3_out_dist0_if_dout;
  assign L3_out_dist0__empty_n = L3_out_dist0_if_empty_n;
  assign L3_out_dist0__full_n = L3_out_dist0_if_full_n;
  assign L3_out_dist0_if_read = L3_out_dist0__read;
  assign L3_out_dist0_if_read_ce = 1'b1;
  assign L3_out_dist0_if_write = L3_out_dist0__write;
  assign L3_out_dist0_if_write_ce = 1'b1;
  assign L3_out_dist0_reset = ~ ap_rst_n;
  assign L3_out_dist1_clk = ap_clk;
  assign L3_out_dist1_if_din = L3_out_dist1__din;
  assign L3_out_dist1__dout = L3_out_dist1_if_dout;
  assign L3_out_dist1__empty_n = L3_out_dist1_if_empty_n;
  assign L3_out_dist1__full_n = L3_out_dist1_if_full_n;
  assign L3_out_dist1_if_read = L3_out_dist1__read;
  assign L3_out_dist1_if_read_ce = 1'b1;
  assign L3_out_dist1_if_write = L3_out_dist1__write;
  assign L3_out_dist1_if_write_ce = 1'b1;
  assign L3_out_dist1_reset = ~ ap_rst_n;
  assign L3_out_id0_clk = ap_clk;
  assign L3_out_id0_if_din = L3_out_id0__din;
  assign L3_out_id0__dout = L3_out_id0_if_dout;
  assign L3_out_id0__empty_n = L3_out_id0_if_empty_n;
  assign L3_out_id0__full_n = L3_out_id0_if_full_n;
  assign L3_out_id0_if_read = L3_out_id0__read;
  assign L3_out_id0_if_read_ce = 1'b1;
  assign L3_out_id0_if_write = L3_out_id0__write;
  assign L3_out_id0_if_write_ce = 1'b1;
  assign L3_out_id0_reset = ~ ap_rst_n;
  assign L3_out_id1_clk = ap_clk;
  assign L3_out_id1_if_din = L3_out_id1__din;
  assign L3_out_id1__dout = L3_out_id1_if_dout;
  assign L3_out_id1__empty_n = L3_out_id1_if_empty_n;
  assign L3_out_id1__full_n = L3_out_id1_if_full_n;
  assign L3_out_id1_if_read = L3_out_id1__read;
  assign L3_out_id1_if_read_ce = 1'b1;
  assign L3_out_id1_if_write = L3_out_id1__write;
  assign L3_out_id1_if_write_ce = 1'b1;
  assign L3_out_id1_reset = ~ ap_rst_n;
  assign out_dist_0_clk = ap_clk;
  assign out_dist_0_if_din = out_dist_0__din;
  assign out_dist_0__dout = out_dist_0_if_dout;
  assign out_dist_0__empty_n = out_dist_0_if_empty_n;
  assign out_dist_0__full_n = out_dist_0_if_full_n;
  assign out_dist_0_if_read = out_dist_0__read;
  assign out_dist_0_if_read_ce = 1'b1;
  assign out_dist_0_if_write = out_dist_0__write;
  assign out_dist_0_if_write_ce = 1'b1;
  assign out_dist_0_reset = ~ ap_rst_n;
  assign out_dist_10_clk = ap_clk;
  assign out_dist_10_if_din = out_dist_10__din;
  assign out_dist_10__dout = out_dist_10_if_dout;
  assign out_dist_10__empty_n = out_dist_10_if_empty_n;
  assign out_dist_10__full_n = out_dist_10_if_full_n;
  assign out_dist_10_if_read = out_dist_10__read;
  assign out_dist_10_if_read_ce = 1'b1;
  assign out_dist_10_if_write = out_dist_10__write;
  assign out_dist_10_if_write_ce = 1'b1;
  assign out_dist_10_reset = ~ ap_rst_n;
  assign out_dist_11_clk = ap_clk;
  assign out_dist_11_if_din = out_dist_11__din;
  assign out_dist_11__dout = out_dist_11_if_dout;
  assign out_dist_11__empty_n = out_dist_11_if_empty_n;
  assign out_dist_11__full_n = out_dist_11_if_full_n;
  assign out_dist_11_if_read = out_dist_11__read;
  assign out_dist_11_if_read_ce = 1'b1;
  assign out_dist_11_if_write = out_dist_11__write;
  assign out_dist_11_if_write_ce = 1'b1;
  assign out_dist_11_reset = ~ ap_rst_n;
  assign out_dist_12_clk = ap_clk;
  assign out_dist_12_if_din = out_dist_12__din;
  assign out_dist_12__dout = out_dist_12_if_dout;
  assign out_dist_12__empty_n = out_dist_12_if_empty_n;
  assign out_dist_12__full_n = out_dist_12_if_full_n;
  assign out_dist_12_if_read = out_dist_12__read;
  assign out_dist_12_if_read_ce = 1'b1;
  assign out_dist_12_if_write = out_dist_12__write;
  assign out_dist_12_if_write_ce = 1'b1;
  assign out_dist_12_reset = ~ ap_rst_n;
  assign out_dist_13_clk = ap_clk;
  assign out_dist_13_if_din = out_dist_13__din;
  assign out_dist_13__dout = out_dist_13_if_dout;
  assign out_dist_13__empty_n = out_dist_13_if_empty_n;
  assign out_dist_13__full_n = out_dist_13_if_full_n;
  assign out_dist_13_if_read = out_dist_13__read;
  assign out_dist_13_if_read_ce = 1'b1;
  assign out_dist_13_if_write = out_dist_13__write;
  assign out_dist_13_if_write_ce = 1'b1;
  assign out_dist_13_reset = ~ ap_rst_n;
  assign out_dist_14_clk = ap_clk;
  assign out_dist_14_if_din = out_dist_14__din;
  assign out_dist_14__dout = out_dist_14_if_dout;
  assign out_dist_14__empty_n = out_dist_14_if_empty_n;
  assign out_dist_14__full_n = out_dist_14_if_full_n;
  assign out_dist_14_if_read = out_dist_14__read;
  assign out_dist_14_if_read_ce = 1'b1;
  assign out_dist_14_if_write = out_dist_14__write;
  assign out_dist_14_if_write_ce = 1'b1;
  assign out_dist_14_reset = ~ ap_rst_n;
  assign out_dist_15_clk = ap_clk;
  assign out_dist_15_if_din = out_dist_15__din;
  assign out_dist_15__dout = out_dist_15_if_dout;
  assign out_dist_15__empty_n = out_dist_15_if_empty_n;
  assign out_dist_15__full_n = out_dist_15_if_full_n;
  assign out_dist_15_if_read = out_dist_15__read;
  assign out_dist_15_if_read_ce = 1'b1;
  assign out_dist_15_if_write = out_dist_15__write;
  assign out_dist_15_if_write_ce = 1'b1;
  assign out_dist_15_reset = ~ ap_rst_n;
  assign out_dist_16_clk = ap_clk;
  assign out_dist_16_if_din = out_dist_16__din;
  assign out_dist_16__dout = out_dist_16_if_dout;
  assign out_dist_16__empty_n = out_dist_16_if_empty_n;
  assign out_dist_16__full_n = out_dist_16_if_full_n;
  assign out_dist_16_if_read = out_dist_16__read;
  assign out_dist_16_if_read_ce = 1'b1;
  assign out_dist_16_if_write = out_dist_16__write;
  assign out_dist_16_if_write_ce = 1'b1;
  assign out_dist_16_reset = ~ ap_rst_n;
  assign out_dist_17_clk = ap_clk;
  assign out_dist_17_if_din = out_dist_17__din;
  assign out_dist_17__dout = out_dist_17_if_dout;
  assign out_dist_17__empty_n = out_dist_17_if_empty_n;
  assign out_dist_17__full_n = out_dist_17_if_full_n;
  assign out_dist_17_if_read = out_dist_17__read;
  assign out_dist_17_if_read_ce = 1'b1;
  assign out_dist_17_if_write = out_dist_17__write;
  assign out_dist_17_if_write_ce = 1'b1;
  assign out_dist_17_reset = ~ ap_rst_n;
  assign out_dist_18_clk = ap_clk;
  assign out_dist_18_if_din = out_dist_18__din;
  assign out_dist_18__dout = out_dist_18_if_dout;
  assign out_dist_18__empty_n = out_dist_18_if_empty_n;
  assign out_dist_18__full_n = out_dist_18_if_full_n;
  assign out_dist_18_if_read = out_dist_18__read;
  assign out_dist_18_if_read_ce = 1'b1;
  assign out_dist_18_if_write = out_dist_18__write;
  assign out_dist_18_if_write_ce = 1'b1;
  assign out_dist_18_reset = ~ ap_rst_n;
  assign out_dist_19_clk = ap_clk;
  assign out_dist_19_if_din = out_dist_19__din;
  assign out_dist_19__dout = out_dist_19_if_dout;
  assign out_dist_19__empty_n = out_dist_19_if_empty_n;
  assign out_dist_19__full_n = out_dist_19_if_full_n;
  assign out_dist_19_if_read = out_dist_19__read;
  assign out_dist_19_if_read_ce = 1'b1;
  assign out_dist_19_if_write = out_dist_19__write;
  assign out_dist_19_if_write_ce = 1'b1;
  assign out_dist_19_reset = ~ ap_rst_n;
  assign out_dist_1_clk = ap_clk;
  assign out_dist_1_if_din = out_dist_1__din;
  assign out_dist_1__dout = out_dist_1_if_dout;
  assign out_dist_1__empty_n = out_dist_1_if_empty_n;
  assign out_dist_1__full_n = out_dist_1_if_full_n;
  assign out_dist_1_if_read = out_dist_1__read;
  assign out_dist_1_if_read_ce = 1'b1;
  assign out_dist_1_if_write = out_dist_1__write;
  assign out_dist_1_if_write_ce = 1'b1;
  assign out_dist_1_reset = ~ ap_rst_n;
  assign out_dist_20_clk = ap_clk;
  assign out_dist_20_if_din = out_dist_20__din;
  assign out_dist_20__dout = out_dist_20_if_dout;
  assign out_dist_20__empty_n = out_dist_20_if_empty_n;
  assign out_dist_20__full_n = out_dist_20_if_full_n;
  assign out_dist_20_if_read = out_dist_20__read;
  assign out_dist_20_if_read_ce = 1'b1;
  assign out_dist_20_if_write = out_dist_20__write;
  assign out_dist_20_if_write_ce = 1'b1;
  assign out_dist_20_reset = ~ ap_rst_n;
  assign out_dist_21_clk = ap_clk;
  assign out_dist_21_if_din = out_dist_21__din;
  assign out_dist_21__dout = out_dist_21_if_dout;
  assign out_dist_21__empty_n = out_dist_21_if_empty_n;
  assign out_dist_21__full_n = out_dist_21_if_full_n;
  assign out_dist_21_if_read = out_dist_21__read;
  assign out_dist_21_if_read_ce = 1'b1;
  assign out_dist_21_if_write = out_dist_21__write;
  assign out_dist_21_if_write_ce = 1'b1;
  assign out_dist_21_reset = ~ ap_rst_n;
  assign out_dist_22_clk = ap_clk;
  assign out_dist_22_if_din = out_dist_22__din;
  assign out_dist_22__dout = out_dist_22_if_dout;
  assign out_dist_22__empty_n = out_dist_22_if_empty_n;
  assign out_dist_22__full_n = out_dist_22_if_full_n;
  assign out_dist_22_if_read = out_dist_22__read;
  assign out_dist_22_if_read_ce = 1'b1;
  assign out_dist_22_if_write = out_dist_22__write;
  assign out_dist_22_if_write_ce = 1'b1;
  assign out_dist_22_reset = ~ ap_rst_n;
  assign out_dist_23_clk = ap_clk;
  assign out_dist_23_if_din = out_dist_23__din;
  assign out_dist_23__dout = out_dist_23_if_dout;
  assign out_dist_23__empty_n = out_dist_23_if_empty_n;
  assign out_dist_23__full_n = out_dist_23_if_full_n;
  assign out_dist_23_if_read = out_dist_23__read;
  assign out_dist_23_if_read_ce = 1'b1;
  assign out_dist_23_if_write = out_dist_23__write;
  assign out_dist_23_if_write_ce = 1'b1;
  assign out_dist_23_reset = ~ ap_rst_n;
  assign out_dist_24_clk = ap_clk;
  assign out_dist_24_if_din = out_dist_24__din;
  assign out_dist_24__dout = out_dist_24_if_dout;
  assign out_dist_24__empty_n = out_dist_24_if_empty_n;
  assign out_dist_24__full_n = out_dist_24_if_full_n;
  assign out_dist_24_if_read = out_dist_24__read;
  assign out_dist_24_if_read_ce = 1'b1;
  assign out_dist_24_if_write = out_dist_24__write;
  assign out_dist_24_if_write_ce = 1'b1;
  assign out_dist_24_reset = ~ ap_rst_n;
  assign out_dist_25_clk = ap_clk;
  assign out_dist_25_if_din = out_dist_25__din;
  assign out_dist_25__dout = out_dist_25_if_dout;
  assign out_dist_25__empty_n = out_dist_25_if_empty_n;
  assign out_dist_25__full_n = out_dist_25_if_full_n;
  assign out_dist_25_if_read = out_dist_25__read;
  assign out_dist_25_if_read_ce = 1'b1;
  assign out_dist_25_if_write = out_dist_25__write;
  assign out_dist_25_if_write_ce = 1'b1;
  assign out_dist_25_reset = ~ ap_rst_n;
  assign out_dist_26_clk = ap_clk;
  assign out_dist_26_if_din = out_dist_26__din;
  assign out_dist_26__dout = out_dist_26_if_dout;
  assign out_dist_26__empty_n = out_dist_26_if_empty_n;
  assign out_dist_26__full_n = out_dist_26_if_full_n;
  assign out_dist_26_if_read = out_dist_26__read;
  assign out_dist_26_if_read_ce = 1'b1;
  assign out_dist_26_if_write = out_dist_26__write;
  assign out_dist_26_if_write_ce = 1'b1;
  assign out_dist_26_reset = ~ ap_rst_n;
  assign out_dist_27_clk = ap_clk;
  assign out_dist_27_if_din = out_dist_27__din;
  assign out_dist_27__dout = out_dist_27_if_dout;
  assign out_dist_27__empty_n = out_dist_27_if_empty_n;
  assign out_dist_27__full_n = out_dist_27_if_full_n;
  assign out_dist_27_if_read = out_dist_27__read;
  assign out_dist_27_if_read_ce = 1'b1;
  assign out_dist_27_if_write = out_dist_27__write;
  assign out_dist_27_if_write_ce = 1'b1;
  assign out_dist_27_reset = ~ ap_rst_n;
  assign out_dist_28_clk = ap_clk;
  assign out_dist_28_if_din = out_dist_28__din;
  assign out_dist_28__dout = out_dist_28_if_dout;
  assign out_dist_28__empty_n = out_dist_28_if_empty_n;
  assign out_dist_28__full_n = out_dist_28_if_full_n;
  assign out_dist_28_if_read = out_dist_28__read;
  assign out_dist_28_if_read_ce = 1'b1;
  assign out_dist_28_if_write = out_dist_28__write;
  assign out_dist_28_if_write_ce = 1'b1;
  assign out_dist_28_reset = ~ ap_rst_n;
  assign out_dist_29_clk = ap_clk;
  assign out_dist_29_if_din = out_dist_29__din;
  assign out_dist_29__dout = out_dist_29_if_dout;
  assign out_dist_29__empty_n = out_dist_29_if_empty_n;
  assign out_dist_29__full_n = out_dist_29_if_full_n;
  assign out_dist_29_if_read = out_dist_29__read;
  assign out_dist_29_if_read_ce = 1'b1;
  assign out_dist_29_if_write = out_dist_29__write;
  assign out_dist_29_if_write_ce = 1'b1;
  assign out_dist_29_reset = ~ ap_rst_n;
  assign out_dist_2_clk = ap_clk;
  assign out_dist_2_if_din = out_dist_2__din;
  assign out_dist_2__dout = out_dist_2_if_dout;
  assign out_dist_2__empty_n = out_dist_2_if_empty_n;
  assign out_dist_2__full_n = out_dist_2_if_full_n;
  assign out_dist_2_if_read = out_dist_2__read;
  assign out_dist_2_if_read_ce = 1'b1;
  assign out_dist_2_if_write = out_dist_2__write;
  assign out_dist_2_if_write_ce = 1'b1;
  assign out_dist_2_reset = ~ ap_rst_n;
  assign out_dist_30_clk = ap_clk;
  assign out_dist_30_if_din = out_dist_30__din;
  assign out_dist_30__dout = out_dist_30_if_dout;
  assign out_dist_30__empty_n = out_dist_30_if_empty_n;
  assign out_dist_30__full_n = out_dist_30_if_full_n;
  assign out_dist_30_if_read = out_dist_30__read;
  assign out_dist_30_if_read_ce = 1'b1;
  assign out_dist_30_if_write = out_dist_30__write;
  assign out_dist_30_if_write_ce = 1'b1;
  assign out_dist_30_reset = ~ ap_rst_n;
  assign out_dist_31_clk = ap_clk;
  assign out_dist_31_if_din = out_dist_31__din;
  assign out_dist_31__dout = out_dist_31_if_dout;
  assign out_dist_31__empty_n = out_dist_31_if_empty_n;
  assign out_dist_31__full_n = out_dist_31_if_full_n;
  assign out_dist_31_if_read = out_dist_31__read;
  assign out_dist_31_if_read_ce = 1'b1;
  assign out_dist_31_if_write = out_dist_31__write;
  assign out_dist_31_if_write_ce = 1'b1;
  assign out_dist_31_reset = ~ ap_rst_n;
  assign out_dist_32_clk = ap_clk;
  assign out_dist_32_if_din = out_dist_32__din;
  assign out_dist_32__dout = out_dist_32_if_dout;
  assign out_dist_32__empty_n = out_dist_32_if_empty_n;
  assign out_dist_32__full_n = out_dist_32_if_full_n;
  assign out_dist_32_if_read = out_dist_32__read;
  assign out_dist_32_if_read_ce = 1'b1;
  assign out_dist_32_if_write = out_dist_32__write;
  assign out_dist_32_if_write_ce = 1'b1;
  assign out_dist_32_reset = ~ ap_rst_n;
  assign out_dist_33_clk = ap_clk;
  assign out_dist_33_if_din = out_dist_33__din;
  assign out_dist_33__dout = out_dist_33_if_dout;
  assign out_dist_33__empty_n = out_dist_33_if_empty_n;
  assign out_dist_33__full_n = out_dist_33_if_full_n;
  assign out_dist_33_if_read = out_dist_33__read;
  assign out_dist_33_if_read_ce = 1'b1;
  assign out_dist_33_if_write = out_dist_33__write;
  assign out_dist_33_if_write_ce = 1'b1;
  assign out_dist_33_reset = ~ ap_rst_n;
  assign out_dist_34_clk = ap_clk;
  assign out_dist_34_if_din = out_dist_34__din;
  assign out_dist_34__dout = out_dist_34_if_dout;
  assign out_dist_34__empty_n = out_dist_34_if_empty_n;
  assign out_dist_34__full_n = out_dist_34_if_full_n;
  assign out_dist_34_if_read = out_dist_34__read;
  assign out_dist_34_if_read_ce = 1'b1;
  assign out_dist_34_if_write = out_dist_34__write;
  assign out_dist_34_if_write_ce = 1'b1;
  assign out_dist_34_reset = ~ ap_rst_n;
  assign out_dist_35_clk = ap_clk;
  assign out_dist_35_if_din = out_dist_35__din;
  assign out_dist_35__dout = out_dist_35_if_dout;
  assign out_dist_35__empty_n = out_dist_35_if_empty_n;
  assign out_dist_35__full_n = out_dist_35_if_full_n;
  assign out_dist_35_if_read = out_dist_35__read;
  assign out_dist_35_if_read_ce = 1'b1;
  assign out_dist_35_if_write = out_dist_35__write;
  assign out_dist_35_if_write_ce = 1'b1;
  assign out_dist_35_reset = ~ ap_rst_n;
  assign out_dist_36_clk = ap_clk;
  assign out_dist_36_if_din = out_dist_36__din;
  assign out_dist_36__dout = out_dist_36_if_dout;
  assign out_dist_36__empty_n = out_dist_36_if_empty_n;
  assign out_dist_36__full_n = out_dist_36_if_full_n;
  assign out_dist_36_if_read = out_dist_36__read;
  assign out_dist_36_if_read_ce = 1'b1;
  assign out_dist_36_if_write = out_dist_36__write;
  assign out_dist_36_if_write_ce = 1'b1;
  assign out_dist_36_reset = ~ ap_rst_n;
  assign out_dist_37_clk = ap_clk;
  assign out_dist_37_if_din = out_dist_37__din;
  assign out_dist_37__dout = out_dist_37_if_dout;
  assign out_dist_37__empty_n = out_dist_37_if_empty_n;
  assign out_dist_37__full_n = out_dist_37_if_full_n;
  assign out_dist_37_if_read = out_dist_37__read;
  assign out_dist_37_if_read_ce = 1'b1;
  assign out_dist_37_if_write = out_dist_37__write;
  assign out_dist_37_if_write_ce = 1'b1;
  assign out_dist_37_reset = ~ ap_rst_n;
  assign out_dist_38_clk = ap_clk;
  assign out_dist_38_if_din = out_dist_38__din;
  assign out_dist_38__dout = out_dist_38_if_dout;
  assign out_dist_38__empty_n = out_dist_38_if_empty_n;
  assign out_dist_38__full_n = out_dist_38_if_full_n;
  assign out_dist_38_if_read = out_dist_38__read;
  assign out_dist_38_if_read_ce = 1'b1;
  assign out_dist_38_if_write = out_dist_38__write;
  assign out_dist_38_if_write_ce = 1'b1;
  assign out_dist_38_reset = ~ ap_rst_n;
  assign out_dist_39_clk = ap_clk;
  assign out_dist_39_if_din = out_dist_39__din;
  assign out_dist_39__dout = out_dist_39_if_dout;
  assign out_dist_39__empty_n = out_dist_39_if_empty_n;
  assign out_dist_39__full_n = out_dist_39_if_full_n;
  assign out_dist_39_if_read = out_dist_39__read;
  assign out_dist_39_if_read_ce = 1'b1;
  assign out_dist_39_if_write = out_dist_39__write;
  assign out_dist_39_if_write_ce = 1'b1;
  assign out_dist_39_reset = ~ ap_rst_n;
  assign out_dist_3_clk = ap_clk;
  assign out_dist_3_if_din = out_dist_3__din;
  assign out_dist_3__dout = out_dist_3_if_dout;
  assign out_dist_3__empty_n = out_dist_3_if_empty_n;
  assign out_dist_3__full_n = out_dist_3_if_full_n;
  assign out_dist_3_if_read = out_dist_3__read;
  assign out_dist_3_if_read_ce = 1'b1;
  assign out_dist_3_if_write = out_dist_3__write;
  assign out_dist_3_if_write_ce = 1'b1;
  assign out_dist_3_reset = ~ ap_rst_n;
  assign out_dist_40_clk = ap_clk;
  assign out_dist_40_if_din = out_dist_40__din;
  assign out_dist_40__dout = out_dist_40_if_dout;
  assign out_dist_40__empty_n = out_dist_40_if_empty_n;
  assign out_dist_40__full_n = out_dist_40_if_full_n;
  assign out_dist_40_if_read = out_dist_40__read;
  assign out_dist_40_if_read_ce = 1'b1;
  assign out_dist_40_if_write = out_dist_40__write;
  assign out_dist_40_if_write_ce = 1'b1;
  assign out_dist_40_reset = ~ ap_rst_n;
  assign out_dist_41_clk = ap_clk;
  assign out_dist_41_if_din = out_dist_41__din;
  assign out_dist_41__dout = out_dist_41_if_dout;
  assign out_dist_41__empty_n = out_dist_41_if_empty_n;
  assign out_dist_41__full_n = out_dist_41_if_full_n;
  assign out_dist_41_if_read = out_dist_41__read;
  assign out_dist_41_if_read_ce = 1'b1;
  assign out_dist_41_if_write = out_dist_41__write;
  assign out_dist_41_if_write_ce = 1'b1;
  assign out_dist_41_reset = ~ ap_rst_n;
  assign out_dist_42_clk = ap_clk;
  assign out_dist_42_if_din = out_dist_42__din;
  assign out_dist_42__dout = out_dist_42_if_dout;
  assign out_dist_42__empty_n = out_dist_42_if_empty_n;
  assign out_dist_42__full_n = out_dist_42_if_full_n;
  assign out_dist_42_if_read = out_dist_42__read;
  assign out_dist_42_if_read_ce = 1'b1;
  assign out_dist_42_if_write = out_dist_42__write;
  assign out_dist_42_if_write_ce = 1'b1;
  assign out_dist_42_reset = ~ ap_rst_n;
  assign out_dist_43_clk = ap_clk;
  assign out_dist_43_if_din = out_dist_43__din;
  assign out_dist_43__dout = out_dist_43_if_dout;
  assign out_dist_43__empty_n = out_dist_43_if_empty_n;
  assign out_dist_43__full_n = out_dist_43_if_full_n;
  assign out_dist_43_if_read = out_dist_43__read;
  assign out_dist_43_if_read_ce = 1'b1;
  assign out_dist_43_if_write = out_dist_43__write;
  assign out_dist_43_if_write_ce = 1'b1;
  assign out_dist_43_reset = ~ ap_rst_n;
  assign out_dist_44_clk = ap_clk;
  assign out_dist_44_if_din = out_dist_44__din;
  assign out_dist_44__dout = out_dist_44_if_dout;
  assign out_dist_44__empty_n = out_dist_44_if_empty_n;
  assign out_dist_44__full_n = out_dist_44_if_full_n;
  assign out_dist_44_if_read = out_dist_44__read;
  assign out_dist_44_if_read_ce = 1'b1;
  assign out_dist_44_if_write = out_dist_44__write;
  assign out_dist_44_if_write_ce = 1'b1;
  assign out_dist_44_reset = ~ ap_rst_n;
  assign out_dist_45_clk = ap_clk;
  assign out_dist_45_if_din = out_dist_45__din;
  assign out_dist_45__dout = out_dist_45_if_dout;
  assign out_dist_45__empty_n = out_dist_45_if_empty_n;
  assign out_dist_45__full_n = out_dist_45_if_full_n;
  assign out_dist_45_if_read = out_dist_45__read;
  assign out_dist_45_if_read_ce = 1'b1;
  assign out_dist_45_if_write = out_dist_45__write;
  assign out_dist_45_if_write_ce = 1'b1;
  assign out_dist_45_reset = ~ ap_rst_n;
  assign out_dist_46_clk = ap_clk;
  assign out_dist_46_if_din = out_dist_46__din;
  assign out_dist_46__dout = out_dist_46_if_dout;
  assign out_dist_46__empty_n = out_dist_46_if_empty_n;
  assign out_dist_46__full_n = out_dist_46_if_full_n;
  assign out_dist_46_if_read = out_dist_46__read;
  assign out_dist_46_if_read_ce = 1'b1;
  assign out_dist_46_if_write = out_dist_46__write;
  assign out_dist_46_if_write_ce = 1'b1;
  assign out_dist_46_reset = ~ ap_rst_n;
  assign out_dist_47_clk = ap_clk;
  assign out_dist_47_if_din = out_dist_47__din;
  assign out_dist_47__dout = out_dist_47_if_dout;
  assign out_dist_47__empty_n = out_dist_47_if_empty_n;
  assign out_dist_47__full_n = out_dist_47_if_full_n;
  assign out_dist_47_if_read = out_dist_47__read;
  assign out_dist_47_if_read_ce = 1'b1;
  assign out_dist_47_if_write = out_dist_47__write;
  assign out_dist_47_if_write_ce = 1'b1;
  assign out_dist_47_reset = ~ ap_rst_n;
  assign out_dist_48_clk = ap_clk;
  assign out_dist_48_if_din = out_dist_48__din;
  assign out_dist_48__dout = out_dist_48_if_dout;
  assign out_dist_48__empty_n = out_dist_48_if_empty_n;
  assign out_dist_48__full_n = out_dist_48_if_full_n;
  assign out_dist_48_if_read = out_dist_48__read;
  assign out_dist_48_if_read_ce = 1'b1;
  assign out_dist_48_if_write = out_dist_48__write;
  assign out_dist_48_if_write_ce = 1'b1;
  assign out_dist_48_reset = ~ ap_rst_n;
  assign out_dist_49_clk = ap_clk;
  assign out_dist_49_if_din = out_dist_49__din;
  assign out_dist_49__dout = out_dist_49_if_dout;
  assign out_dist_49__empty_n = out_dist_49_if_empty_n;
  assign out_dist_49__full_n = out_dist_49_if_full_n;
  assign out_dist_49_if_read = out_dist_49__read;
  assign out_dist_49_if_read_ce = 1'b1;
  assign out_dist_49_if_write = out_dist_49__write;
  assign out_dist_49_if_write_ce = 1'b1;
  assign out_dist_49_reset = ~ ap_rst_n;
  assign out_dist_4_clk = ap_clk;
  assign out_dist_4_if_din = out_dist_4__din;
  assign out_dist_4__dout = out_dist_4_if_dout;
  assign out_dist_4__empty_n = out_dist_4_if_empty_n;
  assign out_dist_4__full_n = out_dist_4_if_full_n;
  assign out_dist_4_if_read = out_dist_4__read;
  assign out_dist_4_if_read_ce = 1'b1;
  assign out_dist_4_if_write = out_dist_4__write;
  assign out_dist_4_if_write_ce = 1'b1;
  assign out_dist_4_reset = ~ ap_rst_n;
  assign out_dist_50_clk = ap_clk;
  assign out_dist_50_if_din = out_dist_50__din;
  assign out_dist_50__dout = out_dist_50_if_dout;
  assign out_dist_50__empty_n = out_dist_50_if_empty_n;
  assign out_dist_50__full_n = out_dist_50_if_full_n;
  assign out_dist_50_if_read = out_dist_50__read;
  assign out_dist_50_if_read_ce = 1'b1;
  assign out_dist_50_if_write = out_dist_50__write;
  assign out_dist_50_if_write_ce = 1'b1;
  assign out_dist_50_reset = ~ ap_rst_n;
  assign out_dist_51_clk = ap_clk;
  assign out_dist_51_if_din = out_dist_51__din;
  assign out_dist_51__dout = out_dist_51_if_dout;
  assign out_dist_51__empty_n = out_dist_51_if_empty_n;
  assign out_dist_51__full_n = out_dist_51_if_full_n;
  assign out_dist_51_if_read = out_dist_51__read;
  assign out_dist_51_if_read_ce = 1'b1;
  assign out_dist_51_if_write = out_dist_51__write;
  assign out_dist_51_if_write_ce = 1'b1;
  assign out_dist_51_reset = ~ ap_rst_n;
  assign out_dist_52_clk = ap_clk;
  assign out_dist_52_if_din = out_dist_52__din;
  assign out_dist_52__dout = out_dist_52_if_dout;
  assign out_dist_52__empty_n = out_dist_52_if_empty_n;
  assign out_dist_52__full_n = out_dist_52_if_full_n;
  assign out_dist_52_if_read = out_dist_52__read;
  assign out_dist_52_if_read_ce = 1'b1;
  assign out_dist_52_if_write = out_dist_52__write;
  assign out_dist_52_if_write_ce = 1'b1;
  assign out_dist_52_reset = ~ ap_rst_n;
  assign out_dist_53_clk = ap_clk;
  assign out_dist_53_if_din = out_dist_53__din;
  assign out_dist_53__dout = out_dist_53_if_dout;
  assign out_dist_53__empty_n = out_dist_53_if_empty_n;
  assign out_dist_53__full_n = out_dist_53_if_full_n;
  assign out_dist_53_if_read = out_dist_53__read;
  assign out_dist_53_if_read_ce = 1'b1;
  assign out_dist_53_if_write = out_dist_53__write;
  assign out_dist_53_if_write_ce = 1'b1;
  assign out_dist_53_reset = ~ ap_rst_n;
  assign out_dist_5_clk = ap_clk;
  assign out_dist_5_if_din = out_dist_5__din;
  assign out_dist_5__dout = out_dist_5_if_dout;
  assign out_dist_5__empty_n = out_dist_5_if_empty_n;
  assign out_dist_5__full_n = out_dist_5_if_full_n;
  assign out_dist_5_if_read = out_dist_5__read;
  assign out_dist_5_if_read_ce = 1'b1;
  assign out_dist_5_if_write = out_dist_5__write;
  assign out_dist_5_if_write_ce = 1'b1;
  assign out_dist_5_reset = ~ ap_rst_n;
  assign out_dist_6_clk = ap_clk;
  assign out_dist_6_if_din = out_dist_6__din;
  assign out_dist_6__dout = out_dist_6_if_dout;
  assign out_dist_6__empty_n = out_dist_6_if_empty_n;
  assign out_dist_6__full_n = out_dist_6_if_full_n;
  assign out_dist_6_if_read = out_dist_6__read;
  assign out_dist_6_if_read_ce = 1'b1;
  assign out_dist_6_if_write = out_dist_6__write;
  assign out_dist_6_if_write_ce = 1'b1;
  assign out_dist_6_reset = ~ ap_rst_n;
  assign out_dist_7_clk = ap_clk;
  assign out_dist_7_if_din = out_dist_7__din;
  assign out_dist_7__dout = out_dist_7_if_dout;
  assign out_dist_7__empty_n = out_dist_7_if_empty_n;
  assign out_dist_7__full_n = out_dist_7_if_full_n;
  assign out_dist_7_if_read = out_dist_7__read;
  assign out_dist_7_if_read_ce = 1'b1;
  assign out_dist_7_if_write = out_dist_7__write;
  assign out_dist_7_if_write_ce = 1'b1;
  assign out_dist_7_reset = ~ ap_rst_n;
  assign out_dist_8_clk = ap_clk;
  assign out_dist_8_if_din = out_dist_8__din;
  assign out_dist_8__dout = out_dist_8_if_dout;
  assign out_dist_8__empty_n = out_dist_8_if_empty_n;
  assign out_dist_8__full_n = out_dist_8_if_full_n;
  assign out_dist_8_if_read = out_dist_8__read;
  assign out_dist_8_if_read_ce = 1'b1;
  assign out_dist_8_if_write = out_dist_8__write;
  assign out_dist_8_if_write_ce = 1'b1;
  assign out_dist_8_reset = ~ ap_rst_n;
  assign out_dist_9_clk = ap_clk;
  assign out_dist_9_if_din = out_dist_9__din;
  assign out_dist_9__dout = out_dist_9_if_dout;
  assign out_dist_9__empty_n = out_dist_9_if_empty_n;
  assign out_dist_9__full_n = out_dist_9_if_full_n;
  assign out_dist_9_if_read = out_dist_9__read;
  assign out_dist_9_if_read_ce = 1'b1;
  assign out_dist_9_if_write = out_dist_9__write;
  assign out_dist_9_if_write_ce = 1'b1;
  assign out_dist_9_reset = ~ ap_rst_n;
  assign out_id_0_clk = ap_clk;
  assign out_id_0_if_din = out_id_0__din;
  assign out_id_0__dout = out_id_0_if_dout;
  assign out_id_0__empty_n = out_id_0_if_empty_n;
  assign out_id_0__full_n = out_id_0_if_full_n;
  assign out_id_0_if_read = out_id_0__read;
  assign out_id_0_if_read_ce = 1'b1;
  assign out_id_0_if_write = out_id_0__write;
  assign out_id_0_if_write_ce = 1'b1;
  assign out_id_0_reset = ~ ap_rst_n;
  assign out_id_10_clk = ap_clk;
  assign out_id_10_if_din = out_id_10__din;
  assign out_id_10__dout = out_id_10_if_dout;
  assign out_id_10__empty_n = out_id_10_if_empty_n;
  assign out_id_10__full_n = out_id_10_if_full_n;
  assign out_id_10_if_read = out_id_10__read;
  assign out_id_10_if_read_ce = 1'b1;
  assign out_id_10_if_write = out_id_10__write;
  assign out_id_10_if_write_ce = 1'b1;
  assign out_id_10_reset = ~ ap_rst_n;
  assign out_id_11_clk = ap_clk;
  assign out_id_11_if_din = out_id_11__din;
  assign out_id_11__dout = out_id_11_if_dout;
  assign out_id_11__empty_n = out_id_11_if_empty_n;
  assign out_id_11__full_n = out_id_11_if_full_n;
  assign out_id_11_if_read = out_id_11__read;
  assign out_id_11_if_read_ce = 1'b1;
  assign out_id_11_if_write = out_id_11__write;
  assign out_id_11_if_write_ce = 1'b1;
  assign out_id_11_reset = ~ ap_rst_n;
  assign out_id_12_clk = ap_clk;
  assign out_id_12_if_din = out_id_12__din;
  assign out_id_12__dout = out_id_12_if_dout;
  assign out_id_12__empty_n = out_id_12_if_empty_n;
  assign out_id_12__full_n = out_id_12_if_full_n;
  assign out_id_12_if_read = out_id_12__read;
  assign out_id_12_if_read_ce = 1'b1;
  assign out_id_12_if_write = out_id_12__write;
  assign out_id_12_if_write_ce = 1'b1;
  assign out_id_12_reset = ~ ap_rst_n;
  assign out_id_13_clk = ap_clk;
  assign out_id_13_if_din = out_id_13__din;
  assign out_id_13__dout = out_id_13_if_dout;
  assign out_id_13__empty_n = out_id_13_if_empty_n;
  assign out_id_13__full_n = out_id_13_if_full_n;
  assign out_id_13_if_read = out_id_13__read;
  assign out_id_13_if_read_ce = 1'b1;
  assign out_id_13_if_write = out_id_13__write;
  assign out_id_13_if_write_ce = 1'b1;
  assign out_id_13_reset = ~ ap_rst_n;
  assign out_id_14_clk = ap_clk;
  assign out_id_14_if_din = out_id_14__din;
  assign out_id_14__dout = out_id_14_if_dout;
  assign out_id_14__empty_n = out_id_14_if_empty_n;
  assign out_id_14__full_n = out_id_14_if_full_n;
  assign out_id_14_if_read = out_id_14__read;
  assign out_id_14_if_read_ce = 1'b1;
  assign out_id_14_if_write = out_id_14__write;
  assign out_id_14_if_write_ce = 1'b1;
  assign out_id_14_reset = ~ ap_rst_n;
  assign out_id_15_clk = ap_clk;
  assign out_id_15_if_din = out_id_15__din;
  assign out_id_15__dout = out_id_15_if_dout;
  assign out_id_15__empty_n = out_id_15_if_empty_n;
  assign out_id_15__full_n = out_id_15_if_full_n;
  assign out_id_15_if_read = out_id_15__read;
  assign out_id_15_if_read_ce = 1'b1;
  assign out_id_15_if_write = out_id_15__write;
  assign out_id_15_if_write_ce = 1'b1;
  assign out_id_15_reset = ~ ap_rst_n;
  assign out_id_16_clk = ap_clk;
  assign out_id_16_if_din = out_id_16__din;
  assign out_id_16__dout = out_id_16_if_dout;
  assign out_id_16__empty_n = out_id_16_if_empty_n;
  assign out_id_16__full_n = out_id_16_if_full_n;
  assign out_id_16_if_read = out_id_16__read;
  assign out_id_16_if_read_ce = 1'b1;
  assign out_id_16_if_write = out_id_16__write;
  assign out_id_16_if_write_ce = 1'b1;
  assign out_id_16_reset = ~ ap_rst_n;
  assign out_id_17_clk = ap_clk;
  assign out_id_17_if_din = out_id_17__din;
  assign out_id_17__dout = out_id_17_if_dout;
  assign out_id_17__empty_n = out_id_17_if_empty_n;
  assign out_id_17__full_n = out_id_17_if_full_n;
  assign out_id_17_if_read = out_id_17__read;
  assign out_id_17_if_read_ce = 1'b1;
  assign out_id_17_if_write = out_id_17__write;
  assign out_id_17_if_write_ce = 1'b1;
  assign out_id_17_reset = ~ ap_rst_n;
  assign out_id_18_clk = ap_clk;
  assign out_id_18_if_din = out_id_18__din;
  assign out_id_18__dout = out_id_18_if_dout;
  assign out_id_18__empty_n = out_id_18_if_empty_n;
  assign out_id_18__full_n = out_id_18_if_full_n;
  assign out_id_18_if_read = out_id_18__read;
  assign out_id_18_if_read_ce = 1'b1;
  assign out_id_18_if_write = out_id_18__write;
  assign out_id_18_if_write_ce = 1'b1;
  assign out_id_18_reset = ~ ap_rst_n;
  assign out_id_19_clk = ap_clk;
  assign out_id_19_if_din = out_id_19__din;
  assign out_id_19__dout = out_id_19_if_dout;
  assign out_id_19__empty_n = out_id_19_if_empty_n;
  assign out_id_19__full_n = out_id_19_if_full_n;
  assign out_id_19_if_read = out_id_19__read;
  assign out_id_19_if_read_ce = 1'b1;
  assign out_id_19_if_write = out_id_19__write;
  assign out_id_19_if_write_ce = 1'b1;
  assign out_id_19_reset = ~ ap_rst_n;
  assign out_id_1_clk = ap_clk;
  assign out_id_1_if_din = out_id_1__din;
  assign out_id_1__dout = out_id_1_if_dout;
  assign out_id_1__empty_n = out_id_1_if_empty_n;
  assign out_id_1__full_n = out_id_1_if_full_n;
  assign out_id_1_if_read = out_id_1__read;
  assign out_id_1_if_read_ce = 1'b1;
  assign out_id_1_if_write = out_id_1__write;
  assign out_id_1_if_write_ce = 1'b1;
  assign out_id_1_reset = ~ ap_rst_n;
  assign out_id_20_clk = ap_clk;
  assign out_id_20_if_din = out_id_20__din;
  assign out_id_20__dout = out_id_20_if_dout;
  assign out_id_20__empty_n = out_id_20_if_empty_n;
  assign out_id_20__full_n = out_id_20_if_full_n;
  assign out_id_20_if_read = out_id_20__read;
  assign out_id_20_if_read_ce = 1'b1;
  assign out_id_20_if_write = out_id_20__write;
  assign out_id_20_if_write_ce = 1'b1;
  assign out_id_20_reset = ~ ap_rst_n;
  assign out_id_21_clk = ap_clk;
  assign out_id_21_if_din = out_id_21__din;
  assign out_id_21__dout = out_id_21_if_dout;
  assign out_id_21__empty_n = out_id_21_if_empty_n;
  assign out_id_21__full_n = out_id_21_if_full_n;
  assign out_id_21_if_read = out_id_21__read;
  assign out_id_21_if_read_ce = 1'b1;
  assign out_id_21_if_write = out_id_21__write;
  assign out_id_21_if_write_ce = 1'b1;
  assign out_id_21_reset = ~ ap_rst_n;
  assign out_id_22_clk = ap_clk;
  assign out_id_22_if_din = out_id_22__din;
  assign out_id_22__dout = out_id_22_if_dout;
  assign out_id_22__empty_n = out_id_22_if_empty_n;
  assign out_id_22__full_n = out_id_22_if_full_n;
  assign out_id_22_if_read = out_id_22__read;
  assign out_id_22_if_read_ce = 1'b1;
  assign out_id_22_if_write = out_id_22__write;
  assign out_id_22_if_write_ce = 1'b1;
  assign out_id_22_reset = ~ ap_rst_n;
  assign out_id_23_clk = ap_clk;
  assign out_id_23_if_din = out_id_23__din;
  assign out_id_23__dout = out_id_23_if_dout;
  assign out_id_23__empty_n = out_id_23_if_empty_n;
  assign out_id_23__full_n = out_id_23_if_full_n;
  assign out_id_23_if_read = out_id_23__read;
  assign out_id_23_if_read_ce = 1'b1;
  assign out_id_23_if_write = out_id_23__write;
  assign out_id_23_if_write_ce = 1'b1;
  assign out_id_23_reset = ~ ap_rst_n;
  assign out_id_24_clk = ap_clk;
  assign out_id_24_if_din = out_id_24__din;
  assign out_id_24__dout = out_id_24_if_dout;
  assign out_id_24__empty_n = out_id_24_if_empty_n;
  assign out_id_24__full_n = out_id_24_if_full_n;
  assign out_id_24_if_read = out_id_24__read;
  assign out_id_24_if_read_ce = 1'b1;
  assign out_id_24_if_write = out_id_24__write;
  assign out_id_24_if_write_ce = 1'b1;
  assign out_id_24_reset = ~ ap_rst_n;
  assign out_id_25_clk = ap_clk;
  assign out_id_25_if_din = out_id_25__din;
  assign out_id_25__dout = out_id_25_if_dout;
  assign out_id_25__empty_n = out_id_25_if_empty_n;
  assign out_id_25__full_n = out_id_25_if_full_n;
  assign out_id_25_if_read = out_id_25__read;
  assign out_id_25_if_read_ce = 1'b1;
  assign out_id_25_if_write = out_id_25__write;
  assign out_id_25_if_write_ce = 1'b1;
  assign out_id_25_reset = ~ ap_rst_n;
  assign out_id_26_clk = ap_clk;
  assign out_id_26_if_din = out_id_26__din;
  assign out_id_26__dout = out_id_26_if_dout;
  assign out_id_26__empty_n = out_id_26_if_empty_n;
  assign out_id_26__full_n = out_id_26_if_full_n;
  assign out_id_26_if_read = out_id_26__read;
  assign out_id_26_if_read_ce = 1'b1;
  assign out_id_26_if_write = out_id_26__write;
  assign out_id_26_if_write_ce = 1'b1;
  assign out_id_26_reset = ~ ap_rst_n;
  assign out_id_27_clk = ap_clk;
  assign out_id_27_if_din = out_id_27__din;
  assign out_id_27__dout = out_id_27_if_dout;
  assign out_id_27__empty_n = out_id_27_if_empty_n;
  assign out_id_27__full_n = out_id_27_if_full_n;
  assign out_id_27_if_read = out_id_27__read;
  assign out_id_27_if_read_ce = 1'b1;
  assign out_id_27_if_write = out_id_27__write;
  assign out_id_27_if_write_ce = 1'b1;
  assign out_id_27_reset = ~ ap_rst_n;
  assign out_id_28_clk = ap_clk;
  assign out_id_28_if_din = out_id_28__din;
  assign out_id_28__dout = out_id_28_if_dout;
  assign out_id_28__empty_n = out_id_28_if_empty_n;
  assign out_id_28__full_n = out_id_28_if_full_n;
  assign out_id_28_if_read = out_id_28__read;
  assign out_id_28_if_read_ce = 1'b1;
  assign out_id_28_if_write = out_id_28__write;
  assign out_id_28_if_write_ce = 1'b1;
  assign out_id_28_reset = ~ ap_rst_n;
  assign out_id_29_clk = ap_clk;
  assign out_id_29_if_din = out_id_29__din;
  assign out_id_29__dout = out_id_29_if_dout;
  assign out_id_29__empty_n = out_id_29_if_empty_n;
  assign out_id_29__full_n = out_id_29_if_full_n;
  assign out_id_29_if_read = out_id_29__read;
  assign out_id_29_if_read_ce = 1'b1;
  assign out_id_29_if_write = out_id_29__write;
  assign out_id_29_if_write_ce = 1'b1;
  assign out_id_29_reset = ~ ap_rst_n;
  assign out_id_2_clk = ap_clk;
  assign out_id_2_if_din = out_id_2__din;
  assign out_id_2__dout = out_id_2_if_dout;
  assign out_id_2__empty_n = out_id_2_if_empty_n;
  assign out_id_2__full_n = out_id_2_if_full_n;
  assign out_id_2_if_read = out_id_2__read;
  assign out_id_2_if_read_ce = 1'b1;
  assign out_id_2_if_write = out_id_2__write;
  assign out_id_2_if_write_ce = 1'b1;
  assign out_id_2_reset = ~ ap_rst_n;
  assign out_id_30_clk = ap_clk;
  assign out_id_30_if_din = out_id_30__din;
  assign out_id_30__dout = out_id_30_if_dout;
  assign out_id_30__empty_n = out_id_30_if_empty_n;
  assign out_id_30__full_n = out_id_30_if_full_n;
  assign out_id_30_if_read = out_id_30__read;
  assign out_id_30_if_read_ce = 1'b1;
  assign out_id_30_if_write = out_id_30__write;
  assign out_id_30_if_write_ce = 1'b1;
  assign out_id_30_reset = ~ ap_rst_n;
  assign out_id_31_clk = ap_clk;
  assign out_id_31_if_din = out_id_31__din;
  assign out_id_31__dout = out_id_31_if_dout;
  assign out_id_31__empty_n = out_id_31_if_empty_n;
  assign out_id_31__full_n = out_id_31_if_full_n;
  assign out_id_31_if_read = out_id_31__read;
  assign out_id_31_if_read_ce = 1'b1;
  assign out_id_31_if_write = out_id_31__write;
  assign out_id_31_if_write_ce = 1'b1;
  assign out_id_31_reset = ~ ap_rst_n;
  assign out_id_32_clk = ap_clk;
  assign out_id_32_if_din = out_id_32__din;
  assign out_id_32__dout = out_id_32_if_dout;
  assign out_id_32__empty_n = out_id_32_if_empty_n;
  assign out_id_32__full_n = out_id_32_if_full_n;
  assign out_id_32_if_read = out_id_32__read;
  assign out_id_32_if_read_ce = 1'b1;
  assign out_id_32_if_write = out_id_32__write;
  assign out_id_32_if_write_ce = 1'b1;
  assign out_id_32_reset = ~ ap_rst_n;
  assign out_id_33_clk = ap_clk;
  assign out_id_33_if_din = out_id_33__din;
  assign out_id_33__dout = out_id_33_if_dout;
  assign out_id_33__empty_n = out_id_33_if_empty_n;
  assign out_id_33__full_n = out_id_33_if_full_n;
  assign out_id_33_if_read = out_id_33__read;
  assign out_id_33_if_read_ce = 1'b1;
  assign out_id_33_if_write = out_id_33__write;
  assign out_id_33_if_write_ce = 1'b1;
  assign out_id_33_reset = ~ ap_rst_n;
  assign out_id_34_clk = ap_clk;
  assign out_id_34_if_din = out_id_34__din;
  assign out_id_34__dout = out_id_34_if_dout;
  assign out_id_34__empty_n = out_id_34_if_empty_n;
  assign out_id_34__full_n = out_id_34_if_full_n;
  assign out_id_34_if_read = out_id_34__read;
  assign out_id_34_if_read_ce = 1'b1;
  assign out_id_34_if_write = out_id_34__write;
  assign out_id_34_if_write_ce = 1'b1;
  assign out_id_34_reset = ~ ap_rst_n;
  assign out_id_35_clk = ap_clk;
  assign out_id_35_if_din = out_id_35__din;
  assign out_id_35__dout = out_id_35_if_dout;
  assign out_id_35__empty_n = out_id_35_if_empty_n;
  assign out_id_35__full_n = out_id_35_if_full_n;
  assign out_id_35_if_read = out_id_35__read;
  assign out_id_35_if_read_ce = 1'b1;
  assign out_id_35_if_write = out_id_35__write;
  assign out_id_35_if_write_ce = 1'b1;
  assign out_id_35_reset = ~ ap_rst_n;
  assign out_id_36_clk = ap_clk;
  assign out_id_36_if_din = out_id_36__din;
  assign out_id_36__dout = out_id_36_if_dout;
  assign out_id_36__empty_n = out_id_36_if_empty_n;
  assign out_id_36__full_n = out_id_36_if_full_n;
  assign out_id_36_if_read = out_id_36__read;
  assign out_id_36_if_read_ce = 1'b1;
  assign out_id_36_if_write = out_id_36__write;
  assign out_id_36_if_write_ce = 1'b1;
  assign out_id_36_reset = ~ ap_rst_n;
  assign out_id_37_clk = ap_clk;
  assign out_id_37_if_din = out_id_37__din;
  assign out_id_37__dout = out_id_37_if_dout;
  assign out_id_37__empty_n = out_id_37_if_empty_n;
  assign out_id_37__full_n = out_id_37_if_full_n;
  assign out_id_37_if_read = out_id_37__read;
  assign out_id_37_if_read_ce = 1'b1;
  assign out_id_37_if_write = out_id_37__write;
  assign out_id_37_if_write_ce = 1'b1;
  assign out_id_37_reset = ~ ap_rst_n;
  assign out_id_38_clk = ap_clk;
  assign out_id_38_if_din = out_id_38__din;
  assign out_id_38__dout = out_id_38_if_dout;
  assign out_id_38__empty_n = out_id_38_if_empty_n;
  assign out_id_38__full_n = out_id_38_if_full_n;
  assign out_id_38_if_read = out_id_38__read;
  assign out_id_38_if_read_ce = 1'b1;
  assign out_id_38_if_write = out_id_38__write;
  assign out_id_38_if_write_ce = 1'b1;
  assign out_id_38_reset = ~ ap_rst_n;
  assign out_id_39_clk = ap_clk;
  assign out_id_39_if_din = out_id_39__din;
  assign out_id_39__dout = out_id_39_if_dout;
  assign out_id_39__empty_n = out_id_39_if_empty_n;
  assign out_id_39__full_n = out_id_39_if_full_n;
  assign out_id_39_if_read = out_id_39__read;
  assign out_id_39_if_read_ce = 1'b1;
  assign out_id_39_if_write = out_id_39__write;
  assign out_id_39_if_write_ce = 1'b1;
  assign out_id_39_reset = ~ ap_rst_n;
  assign out_id_3_clk = ap_clk;
  assign out_id_3_if_din = out_id_3__din;
  assign out_id_3__dout = out_id_3_if_dout;
  assign out_id_3__empty_n = out_id_3_if_empty_n;
  assign out_id_3__full_n = out_id_3_if_full_n;
  assign out_id_3_if_read = out_id_3__read;
  assign out_id_3_if_read_ce = 1'b1;
  assign out_id_3_if_write = out_id_3__write;
  assign out_id_3_if_write_ce = 1'b1;
  assign out_id_3_reset = ~ ap_rst_n;
  assign out_id_40_clk = ap_clk;
  assign out_id_40_if_din = out_id_40__din;
  assign out_id_40__dout = out_id_40_if_dout;
  assign out_id_40__empty_n = out_id_40_if_empty_n;
  assign out_id_40__full_n = out_id_40_if_full_n;
  assign out_id_40_if_read = out_id_40__read;
  assign out_id_40_if_read_ce = 1'b1;
  assign out_id_40_if_write = out_id_40__write;
  assign out_id_40_if_write_ce = 1'b1;
  assign out_id_40_reset = ~ ap_rst_n;
  assign out_id_41_clk = ap_clk;
  assign out_id_41_if_din = out_id_41__din;
  assign out_id_41__dout = out_id_41_if_dout;
  assign out_id_41__empty_n = out_id_41_if_empty_n;
  assign out_id_41__full_n = out_id_41_if_full_n;
  assign out_id_41_if_read = out_id_41__read;
  assign out_id_41_if_read_ce = 1'b1;
  assign out_id_41_if_write = out_id_41__write;
  assign out_id_41_if_write_ce = 1'b1;
  assign out_id_41_reset = ~ ap_rst_n;
  assign out_id_42_clk = ap_clk;
  assign out_id_42_if_din = out_id_42__din;
  assign out_id_42__dout = out_id_42_if_dout;
  assign out_id_42__empty_n = out_id_42_if_empty_n;
  assign out_id_42__full_n = out_id_42_if_full_n;
  assign out_id_42_if_read = out_id_42__read;
  assign out_id_42_if_read_ce = 1'b1;
  assign out_id_42_if_write = out_id_42__write;
  assign out_id_42_if_write_ce = 1'b1;
  assign out_id_42_reset = ~ ap_rst_n;
  assign out_id_43_clk = ap_clk;
  assign out_id_43_if_din = out_id_43__din;
  assign out_id_43__dout = out_id_43_if_dout;
  assign out_id_43__empty_n = out_id_43_if_empty_n;
  assign out_id_43__full_n = out_id_43_if_full_n;
  assign out_id_43_if_read = out_id_43__read;
  assign out_id_43_if_read_ce = 1'b1;
  assign out_id_43_if_write = out_id_43__write;
  assign out_id_43_if_write_ce = 1'b1;
  assign out_id_43_reset = ~ ap_rst_n;
  assign out_id_44_clk = ap_clk;
  assign out_id_44_if_din = out_id_44__din;
  assign out_id_44__dout = out_id_44_if_dout;
  assign out_id_44__empty_n = out_id_44_if_empty_n;
  assign out_id_44__full_n = out_id_44_if_full_n;
  assign out_id_44_if_read = out_id_44__read;
  assign out_id_44_if_read_ce = 1'b1;
  assign out_id_44_if_write = out_id_44__write;
  assign out_id_44_if_write_ce = 1'b1;
  assign out_id_44_reset = ~ ap_rst_n;
  assign out_id_45_clk = ap_clk;
  assign out_id_45_if_din = out_id_45__din;
  assign out_id_45__dout = out_id_45_if_dout;
  assign out_id_45__empty_n = out_id_45_if_empty_n;
  assign out_id_45__full_n = out_id_45_if_full_n;
  assign out_id_45_if_read = out_id_45__read;
  assign out_id_45_if_read_ce = 1'b1;
  assign out_id_45_if_write = out_id_45__write;
  assign out_id_45_if_write_ce = 1'b1;
  assign out_id_45_reset = ~ ap_rst_n;
  assign out_id_46_clk = ap_clk;
  assign out_id_46_if_din = out_id_46__din;
  assign out_id_46__dout = out_id_46_if_dout;
  assign out_id_46__empty_n = out_id_46_if_empty_n;
  assign out_id_46__full_n = out_id_46_if_full_n;
  assign out_id_46_if_read = out_id_46__read;
  assign out_id_46_if_read_ce = 1'b1;
  assign out_id_46_if_write = out_id_46__write;
  assign out_id_46_if_write_ce = 1'b1;
  assign out_id_46_reset = ~ ap_rst_n;
  assign out_id_47_clk = ap_clk;
  assign out_id_47_if_din = out_id_47__din;
  assign out_id_47__dout = out_id_47_if_dout;
  assign out_id_47__empty_n = out_id_47_if_empty_n;
  assign out_id_47__full_n = out_id_47_if_full_n;
  assign out_id_47_if_read = out_id_47__read;
  assign out_id_47_if_read_ce = 1'b1;
  assign out_id_47_if_write = out_id_47__write;
  assign out_id_47_if_write_ce = 1'b1;
  assign out_id_47_reset = ~ ap_rst_n;
  assign out_id_48_clk = ap_clk;
  assign out_id_48_if_din = out_id_48__din;
  assign out_id_48__dout = out_id_48_if_dout;
  assign out_id_48__empty_n = out_id_48_if_empty_n;
  assign out_id_48__full_n = out_id_48_if_full_n;
  assign out_id_48_if_read = out_id_48__read;
  assign out_id_48_if_read_ce = 1'b1;
  assign out_id_48_if_write = out_id_48__write;
  assign out_id_48_if_write_ce = 1'b1;
  assign out_id_48_reset = ~ ap_rst_n;
  assign out_id_49_clk = ap_clk;
  assign out_id_49_if_din = out_id_49__din;
  assign out_id_49__dout = out_id_49_if_dout;
  assign out_id_49__empty_n = out_id_49_if_empty_n;
  assign out_id_49__full_n = out_id_49_if_full_n;
  assign out_id_49_if_read = out_id_49__read;
  assign out_id_49_if_read_ce = 1'b1;
  assign out_id_49_if_write = out_id_49__write;
  assign out_id_49_if_write_ce = 1'b1;
  assign out_id_49_reset = ~ ap_rst_n;
  assign out_id_4_clk = ap_clk;
  assign out_id_4_if_din = out_id_4__din;
  assign out_id_4__dout = out_id_4_if_dout;
  assign out_id_4__empty_n = out_id_4_if_empty_n;
  assign out_id_4__full_n = out_id_4_if_full_n;
  assign out_id_4_if_read = out_id_4__read;
  assign out_id_4_if_read_ce = 1'b1;
  assign out_id_4_if_write = out_id_4__write;
  assign out_id_4_if_write_ce = 1'b1;
  assign out_id_4_reset = ~ ap_rst_n;
  assign out_id_50_clk = ap_clk;
  assign out_id_50_if_din = out_id_50__din;
  assign out_id_50__dout = out_id_50_if_dout;
  assign out_id_50__empty_n = out_id_50_if_empty_n;
  assign out_id_50__full_n = out_id_50_if_full_n;
  assign out_id_50_if_read = out_id_50__read;
  assign out_id_50_if_read_ce = 1'b1;
  assign out_id_50_if_write = out_id_50__write;
  assign out_id_50_if_write_ce = 1'b1;
  assign out_id_50_reset = ~ ap_rst_n;
  assign out_id_51_clk = ap_clk;
  assign out_id_51_if_din = out_id_51__din;
  assign out_id_51__dout = out_id_51_if_dout;
  assign out_id_51__empty_n = out_id_51_if_empty_n;
  assign out_id_51__full_n = out_id_51_if_full_n;
  assign out_id_51_if_read = out_id_51__read;
  assign out_id_51_if_read_ce = 1'b1;
  assign out_id_51_if_write = out_id_51__write;
  assign out_id_51_if_write_ce = 1'b1;
  assign out_id_51_reset = ~ ap_rst_n;
  assign out_id_52_clk = ap_clk;
  assign out_id_52_if_din = out_id_52__din;
  assign out_id_52__dout = out_id_52_if_dout;
  assign out_id_52__empty_n = out_id_52_if_empty_n;
  assign out_id_52__full_n = out_id_52_if_full_n;
  assign out_id_52_if_read = out_id_52__read;
  assign out_id_52_if_read_ce = 1'b1;
  assign out_id_52_if_write = out_id_52__write;
  assign out_id_52_if_write_ce = 1'b1;
  assign out_id_52_reset = ~ ap_rst_n;
  assign out_id_53_clk = ap_clk;
  assign out_id_53_if_din = out_id_53__din;
  assign out_id_53__dout = out_id_53_if_dout;
  assign out_id_53__empty_n = out_id_53_if_empty_n;
  assign out_id_53__full_n = out_id_53_if_full_n;
  assign out_id_53_if_read = out_id_53__read;
  assign out_id_53_if_read_ce = 1'b1;
  assign out_id_53_if_write = out_id_53__write;
  assign out_id_53_if_write_ce = 1'b1;
  assign out_id_53_reset = ~ ap_rst_n;
  assign out_id_5_clk = ap_clk;
  assign out_id_5_if_din = out_id_5__din;
  assign out_id_5__dout = out_id_5_if_dout;
  assign out_id_5__empty_n = out_id_5_if_empty_n;
  assign out_id_5__full_n = out_id_5_if_full_n;
  assign out_id_5_if_read = out_id_5__read;
  assign out_id_5_if_read_ce = 1'b1;
  assign out_id_5_if_write = out_id_5__write;
  assign out_id_5_if_write_ce = 1'b1;
  assign out_id_5_reset = ~ ap_rst_n;
  assign out_id_6_clk = ap_clk;
  assign out_id_6_if_din = out_id_6__din;
  assign out_id_6__dout = out_id_6_if_dout;
  assign out_id_6__empty_n = out_id_6_if_empty_n;
  assign out_id_6__full_n = out_id_6_if_full_n;
  assign out_id_6_if_read = out_id_6__read;
  assign out_id_6_if_read_ce = 1'b1;
  assign out_id_6_if_write = out_id_6__write;
  assign out_id_6_if_write_ce = 1'b1;
  assign out_id_6_reset = ~ ap_rst_n;
  assign out_id_7_clk = ap_clk;
  assign out_id_7_if_din = out_id_7__din;
  assign out_id_7__dout = out_id_7_if_dout;
  assign out_id_7__empty_n = out_id_7_if_empty_n;
  assign out_id_7__full_n = out_id_7_if_full_n;
  assign out_id_7_if_read = out_id_7__read;
  assign out_id_7_if_read_ce = 1'b1;
  assign out_id_7_if_write = out_id_7__write;
  assign out_id_7_if_write_ce = 1'b1;
  assign out_id_7_reset = ~ ap_rst_n;
  assign out_id_8_clk = ap_clk;
  assign out_id_8_if_din = out_id_8__din;
  assign out_id_8__dout = out_id_8_if_dout;
  assign out_id_8__empty_n = out_id_8_if_empty_n;
  assign out_id_8__full_n = out_id_8_if_full_n;
  assign out_id_8_if_read = out_id_8__read;
  assign out_id_8_if_read_ce = 1'b1;
  assign out_id_8_if_write = out_id_8__write;
  assign out_id_8_if_write_ce = 1'b1;
  assign out_id_8_reset = ~ ap_rst_n;
  assign out_id_9_clk = ap_clk;
  assign out_id_9_if_din = out_id_9__din;
  assign out_id_9__dout = out_id_9_if_dout;
  assign out_id_9__empty_n = out_id_9_if_empty_n;
  assign out_id_9__full_n = out_id_9_if_full_n;
  assign out_id_9_if_read = out_id_9__read;
  assign out_id_9_if_read_ce = 1'b1;
  assign out_id_9_if_write = out_id_9__write;
  assign out_id_9_if_write_ce = 1'b1;
  assign out_id_9_reset = ~ ap_rst_n;
  assign krnl_globalSort_L1_L2_0_ap_clk = ap_clk;
  assign krnl_globalSort_L1_L2_0__ap_done = krnl_globalSort_L1_L2_0_ap_done;
  assign krnl_globalSort_L1_L2_0__ap_idle = krnl_globalSort_L1_L2_0_ap_idle;
  assign krnl_globalSort_L1_L2_0__ap_ready = krnl_globalSort_L1_L2_0_ap_ready;
  assign krnl_globalSort_L1_L2_0_ap_rst_n = ap_rst_n;
  assign krnl_globalSort_L1_L2_0_ap_start = krnl_globalSort_L1_L2_0__ap_start;
  assign krnl_globalSort_L1_L2_0_in_dist0_peek_dout = out_dist_0__dout;
  assign krnl_globalSort_L1_L2_0_in_dist0_peek_empty_n = out_dist_0__empty_n;
  assign krnl_globalSort_L1_L2_0_in_dist0_s_dout = out_dist_0__dout;
  assign krnl_globalSort_L1_L2_0_in_dist0_s_empty_n = out_dist_0__empty_n;
  assign out_dist_0__read = krnl_globalSort_L1_L2_0_in_dist0_s_read;
  assign krnl_globalSort_L1_L2_0_in_dist1_peek_dout = out_dist_1__dout;
  assign krnl_globalSort_L1_L2_0_in_dist1_peek_empty_n = out_dist_1__empty_n;
  assign krnl_globalSort_L1_L2_0_in_dist1_s_dout = out_dist_1__dout;
  assign krnl_globalSort_L1_L2_0_in_dist1_s_empty_n = out_dist_1__empty_n;
  assign out_dist_1__read = krnl_globalSort_L1_L2_0_in_dist1_s_read;
  assign krnl_globalSort_L1_L2_0_in_dist2_peek_dout = out_dist_2__dout;
  assign krnl_globalSort_L1_L2_0_in_dist2_peek_empty_n = out_dist_2__empty_n;
  assign krnl_globalSort_L1_L2_0_in_dist2_s_dout = out_dist_2__dout;
  assign krnl_globalSort_L1_L2_0_in_dist2_s_empty_n = out_dist_2__empty_n;
  assign out_dist_2__read = krnl_globalSort_L1_L2_0_in_dist2_s_read;
  assign krnl_globalSort_L1_L2_0_in_id0_peek_dout = out_id_0__dout;
  assign krnl_globalSort_L1_L2_0_in_id0_peek_empty_n = out_id_0__empty_n;
  assign krnl_globalSort_L1_L2_0_in_id0_s_dout = out_id_0__dout;
  assign krnl_globalSort_L1_L2_0_in_id0_s_empty_n = out_id_0__empty_n;
  assign out_id_0__read = krnl_globalSort_L1_L2_0_in_id0_s_read;
  assign krnl_globalSort_L1_L2_0_in_id1_peek_dout = out_id_1__dout;
  assign krnl_globalSort_L1_L2_0_in_id1_peek_empty_n = out_id_1__empty_n;
  assign krnl_globalSort_L1_L2_0_in_id1_s_dout = out_id_1__dout;
  assign krnl_globalSort_L1_L2_0_in_id1_s_empty_n = out_id_1__empty_n;
  assign out_id_1__read = krnl_globalSort_L1_L2_0_in_id1_s_read;
  assign krnl_globalSort_L1_L2_0_in_id2_peek_dout = out_id_2__dout;
  assign krnl_globalSort_L1_L2_0_in_id2_peek_empty_n = out_id_2__empty_n;
  assign krnl_globalSort_L1_L2_0_in_id2_s_dout = out_id_2__dout;
  assign krnl_globalSort_L1_L2_0_in_id2_s_empty_n = out_id_2__empty_n;
  assign out_id_2__read = krnl_globalSort_L1_L2_0_in_id2_s_read;
  assign L1_out_dist_0__din = krnl_globalSort_L1_L2_0_out_dist_din;
  assign krnl_globalSort_L1_L2_0_out_dist_full_n = L1_out_dist_0__full_n;
  assign L1_out_dist_0__write = krnl_globalSort_L1_L2_0_out_dist_write;
  assign L1_out_id_0__din = krnl_globalSort_L1_L2_0_out_id_din;
  assign krnl_globalSort_L1_L2_0_out_id_full_n = L1_out_id_0__full_n;
  assign L1_out_id_0__write = krnl_globalSort_L1_L2_0_out_id_write;
  assign krnl_globalSort_L1_L2_1_ap_clk = ap_clk;
  assign krnl_globalSort_L1_L2_1__ap_done = krnl_globalSort_L1_L2_1_ap_done;
  assign krnl_globalSort_L1_L2_1__ap_idle = krnl_globalSort_L1_L2_1_ap_idle;
  assign krnl_globalSort_L1_L2_1__ap_ready = krnl_globalSort_L1_L2_1_ap_ready;
  assign krnl_globalSort_L1_L2_1_ap_rst_n = ap_rst_n;
  assign krnl_globalSort_L1_L2_1_ap_start = krnl_globalSort_L1_L2_1__ap_start;
  assign krnl_globalSort_L1_L2_1_in_dist0_peek_dout = out_dist_3__dout;
  assign krnl_globalSort_L1_L2_1_in_dist0_peek_empty_n = out_dist_3__empty_n;
  assign krnl_globalSort_L1_L2_1_in_dist0_s_dout = out_dist_3__dout;
  assign krnl_globalSort_L1_L2_1_in_dist0_s_empty_n = out_dist_3__empty_n;
  assign out_dist_3__read = krnl_globalSort_L1_L2_1_in_dist0_s_read;
  assign krnl_globalSort_L1_L2_1_in_dist1_peek_dout = out_dist_4__dout;
  assign krnl_globalSort_L1_L2_1_in_dist1_peek_empty_n = out_dist_4__empty_n;
  assign krnl_globalSort_L1_L2_1_in_dist1_s_dout = out_dist_4__dout;
  assign krnl_globalSort_L1_L2_1_in_dist1_s_empty_n = out_dist_4__empty_n;
  assign out_dist_4__read = krnl_globalSort_L1_L2_1_in_dist1_s_read;
  assign krnl_globalSort_L1_L2_1_in_dist2_peek_dout = out_dist_5__dout;
  assign krnl_globalSort_L1_L2_1_in_dist2_peek_empty_n = out_dist_5__empty_n;
  assign krnl_globalSort_L1_L2_1_in_dist2_s_dout = out_dist_5__dout;
  assign krnl_globalSort_L1_L2_1_in_dist2_s_empty_n = out_dist_5__empty_n;
  assign out_dist_5__read = krnl_globalSort_L1_L2_1_in_dist2_s_read;
  assign krnl_globalSort_L1_L2_1_in_id0_peek_dout = out_id_3__dout;
  assign krnl_globalSort_L1_L2_1_in_id0_peek_empty_n = out_id_3__empty_n;
  assign krnl_globalSort_L1_L2_1_in_id0_s_dout = out_id_3__dout;
  assign krnl_globalSort_L1_L2_1_in_id0_s_empty_n = out_id_3__empty_n;
  assign out_id_3__read = krnl_globalSort_L1_L2_1_in_id0_s_read;
  assign krnl_globalSort_L1_L2_1_in_id1_peek_dout = out_id_4__dout;
  assign krnl_globalSort_L1_L2_1_in_id1_peek_empty_n = out_id_4__empty_n;
  assign krnl_globalSort_L1_L2_1_in_id1_s_dout = out_id_4__dout;
  assign krnl_globalSort_L1_L2_1_in_id1_s_empty_n = out_id_4__empty_n;
  assign out_id_4__read = krnl_globalSort_L1_L2_1_in_id1_s_read;
  assign krnl_globalSort_L1_L2_1_in_id2_peek_dout = out_id_5__dout;
  assign krnl_globalSort_L1_L2_1_in_id2_peek_empty_n = out_id_5__empty_n;
  assign krnl_globalSort_L1_L2_1_in_id2_s_dout = out_id_5__dout;
  assign krnl_globalSort_L1_L2_1_in_id2_s_empty_n = out_id_5__empty_n;
  assign out_id_5__read = krnl_globalSort_L1_L2_1_in_id2_s_read;
  assign L1_out_dist_1__din = krnl_globalSort_L1_L2_1_out_dist_din;
  assign krnl_globalSort_L1_L2_1_out_dist_full_n = L1_out_dist_1__full_n;
  assign L1_out_dist_1__write = krnl_globalSort_L1_L2_1_out_dist_write;
  assign L1_out_id_1__din = krnl_globalSort_L1_L2_1_out_id_din;
  assign krnl_globalSort_L1_L2_1_out_id_full_n = L1_out_id_1__full_n;
  assign L1_out_id_1__write = krnl_globalSort_L1_L2_1_out_id_write;
  assign krnl_globalSort_L1_L2_2_ap_clk = ap_clk;
  assign krnl_globalSort_L1_L2_2__ap_done = krnl_globalSort_L1_L2_2_ap_done;
  assign krnl_globalSort_L1_L2_2__ap_idle = krnl_globalSort_L1_L2_2_ap_idle;
  assign krnl_globalSort_L1_L2_2__ap_ready = krnl_globalSort_L1_L2_2_ap_ready;
  assign krnl_globalSort_L1_L2_2_ap_rst_n = ap_rst_n;
  assign krnl_globalSort_L1_L2_2_ap_start = krnl_globalSort_L1_L2_2__ap_start;
  assign krnl_globalSort_L1_L2_2_in_dist0_peek_dout = out_dist_6__dout;
  assign krnl_globalSort_L1_L2_2_in_dist0_peek_empty_n = out_dist_6__empty_n;
  assign krnl_globalSort_L1_L2_2_in_dist0_s_dout = out_dist_6__dout;
  assign krnl_globalSort_L1_L2_2_in_dist0_s_empty_n = out_dist_6__empty_n;
  assign out_dist_6__read = krnl_globalSort_L1_L2_2_in_dist0_s_read;
  assign krnl_globalSort_L1_L2_2_in_dist1_peek_dout = out_dist_7__dout;
  assign krnl_globalSort_L1_L2_2_in_dist1_peek_empty_n = out_dist_7__empty_n;
  assign krnl_globalSort_L1_L2_2_in_dist1_s_dout = out_dist_7__dout;
  assign krnl_globalSort_L1_L2_2_in_dist1_s_empty_n = out_dist_7__empty_n;
  assign out_dist_7__read = krnl_globalSort_L1_L2_2_in_dist1_s_read;
  assign krnl_globalSort_L1_L2_2_in_dist2_peek_dout = out_dist_8__dout;
  assign krnl_globalSort_L1_L2_2_in_dist2_peek_empty_n = out_dist_8__empty_n;
  assign krnl_globalSort_L1_L2_2_in_dist2_s_dout = out_dist_8__dout;
  assign krnl_globalSort_L1_L2_2_in_dist2_s_empty_n = out_dist_8__empty_n;
  assign out_dist_8__read = krnl_globalSort_L1_L2_2_in_dist2_s_read;
  assign krnl_globalSort_L1_L2_2_in_id0_peek_dout = out_id_6__dout;
  assign krnl_globalSort_L1_L2_2_in_id0_peek_empty_n = out_id_6__empty_n;
  assign krnl_globalSort_L1_L2_2_in_id0_s_dout = out_id_6__dout;
  assign krnl_globalSort_L1_L2_2_in_id0_s_empty_n = out_id_6__empty_n;
  assign out_id_6__read = krnl_globalSort_L1_L2_2_in_id0_s_read;
  assign krnl_globalSort_L1_L2_2_in_id1_peek_dout = out_id_7__dout;
  assign krnl_globalSort_L1_L2_2_in_id1_peek_empty_n = out_id_7__empty_n;
  assign krnl_globalSort_L1_L2_2_in_id1_s_dout = out_id_7__dout;
  assign krnl_globalSort_L1_L2_2_in_id1_s_empty_n = out_id_7__empty_n;
  assign out_id_7__read = krnl_globalSort_L1_L2_2_in_id1_s_read;
  assign krnl_globalSort_L1_L2_2_in_id2_peek_dout = out_id_8__dout;
  assign krnl_globalSort_L1_L2_2_in_id2_peek_empty_n = out_id_8__empty_n;
  assign krnl_globalSort_L1_L2_2_in_id2_s_dout = out_id_8__dout;
  assign krnl_globalSort_L1_L2_2_in_id2_s_empty_n = out_id_8__empty_n;
  assign out_id_8__read = krnl_globalSort_L1_L2_2_in_id2_s_read;
  assign L1_out_dist_2__din = krnl_globalSort_L1_L2_2_out_dist_din;
  assign krnl_globalSort_L1_L2_2_out_dist_full_n = L1_out_dist_2__full_n;
  assign L1_out_dist_2__write = krnl_globalSort_L1_L2_2_out_dist_write;
  assign L1_out_id_2__din = krnl_globalSort_L1_L2_2_out_id_din;
  assign krnl_globalSort_L1_L2_2_out_id_full_n = L1_out_id_2__full_n;
  assign L1_out_id_2__write = krnl_globalSort_L1_L2_2_out_id_write;
  assign krnl_globalSort_L1_L2_3_ap_clk = ap_clk;
  assign krnl_globalSort_L1_L2_3__ap_done = krnl_globalSort_L1_L2_3_ap_done;
  assign krnl_globalSort_L1_L2_3__ap_idle = krnl_globalSort_L1_L2_3_ap_idle;
  assign krnl_globalSort_L1_L2_3__ap_ready = krnl_globalSort_L1_L2_3_ap_ready;
  assign krnl_globalSort_L1_L2_3_ap_rst_n = ap_rst_n;
  assign krnl_globalSort_L1_L2_3_ap_start = krnl_globalSort_L1_L2_3__ap_start;
  assign krnl_globalSort_L1_L2_3_in_dist0_peek_dout = out_dist_9__dout;
  assign krnl_globalSort_L1_L2_3_in_dist0_peek_empty_n = out_dist_9__empty_n;
  assign krnl_globalSort_L1_L2_3_in_dist0_s_dout = out_dist_9__dout;
  assign krnl_globalSort_L1_L2_3_in_dist0_s_empty_n = out_dist_9__empty_n;
  assign out_dist_9__read = krnl_globalSort_L1_L2_3_in_dist0_s_read;
  assign krnl_globalSort_L1_L2_3_in_dist1_peek_dout = out_dist_10__dout;
  assign krnl_globalSort_L1_L2_3_in_dist1_peek_empty_n = out_dist_10__empty_n;
  assign krnl_globalSort_L1_L2_3_in_dist1_s_dout = out_dist_10__dout;
  assign krnl_globalSort_L1_L2_3_in_dist1_s_empty_n = out_dist_10__empty_n;
  assign out_dist_10__read = krnl_globalSort_L1_L2_3_in_dist1_s_read;
  assign krnl_globalSort_L1_L2_3_in_dist2_peek_dout = out_dist_11__dout;
  assign krnl_globalSort_L1_L2_3_in_dist2_peek_empty_n = out_dist_11__empty_n;
  assign krnl_globalSort_L1_L2_3_in_dist2_s_dout = out_dist_11__dout;
  assign krnl_globalSort_L1_L2_3_in_dist2_s_empty_n = out_dist_11__empty_n;
  assign out_dist_11__read = krnl_globalSort_L1_L2_3_in_dist2_s_read;
  assign krnl_globalSort_L1_L2_3_in_id0_peek_dout = out_id_9__dout;
  assign krnl_globalSort_L1_L2_3_in_id0_peek_empty_n = out_id_9__empty_n;
  assign krnl_globalSort_L1_L2_3_in_id0_s_dout = out_id_9__dout;
  assign krnl_globalSort_L1_L2_3_in_id0_s_empty_n = out_id_9__empty_n;
  assign out_id_9__read = krnl_globalSort_L1_L2_3_in_id0_s_read;
  assign krnl_globalSort_L1_L2_3_in_id1_peek_dout = out_id_10__dout;
  assign krnl_globalSort_L1_L2_3_in_id1_peek_empty_n = out_id_10__empty_n;
  assign krnl_globalSort_L1_L2_3_in_id1_s_dout = out_id_10__dout;
  assign krnl_globalSort_L1_L2_3_in_id1_s_empty_n = out_id_10__empty_n;
  assign out_id_10__read = krnl_globalSort_L1_L2_3_in_id1_s_read;
  assign krnl_globalSort_L1_L2_3_in_id2_peek_dout = out_id_11__dout;
  assign krnl_globalSort_L1_L2_3_in_id2_peek_empty_n = out_id_11__empty_n;
  assign krnl_globalSort_L1_L2_3_in_id2_s_dout = out_id_11__dout;
  assign krnl_globalSort_L1_L2_3_in_id2_s_empty_n = out_id_11__empty_n;
  assign out_id_11__read = krnl_globalSort_L1_L2_3_in_id2_s_read;
  assign L1_out_dist_3__din = krnl_globalSort_L1_L2_3_out_dist_din;
  assign krnl_globalSort_L1_L2_3_out_dist_full_n = L1_out_dist_3__full_n;
  assign L1_out_dist_3__write = krnl_globalSort_L1_L2_3_out_dist_write;
  assign L1_out_id_3__din = krnl_globalSort_L1_L2_3_out_id_din;
  assign krnl_globalSort_L1_L2_3_out_id_full_n = L1_out_id_3__full_n;
  assign L1_out_id_3__write = krnl_globalSort_L1_L2_3_out_id_write;
  assign krnl_globalSort_L1_L2_4_ap_clk = ap_clk;
  assign krnl_globalSort_L1_L2_4__ap_done = krnl_globalSort_L1_L2_4_ap_done;
  assign krnl_globalSort_L1_L2_4__ap_idle = krnl_globalSort_L1_L2_4_ap_idle;
  assign krnl_globalSort_L1_L2_4__ap_ready = krnl_globalSort_L1_L2_4_ap_ready;
  assign krnl_globalSort_L1_L2_4_ap_rst_n = ap_rst_n;
  assign krnl_globalSort_L1_L2_4_ap_start = krnl_globalSort_L1_L2_4__ap_start;
  assign krnl_globalSort_L1_L2_4_in_dist0_peek_dout = out_dist_12__dout;
  assign krnl_globalSort_L1_L2_4_in_dist0_peek_empty_n = out_dist_12__empty_n;
  assign krnl_globalSort_L1_L2_4_in_dist0_s_dout = out_dist_12__dout;
  assign krnl_globalSort_L1_L2_4_in_dist0_s_empty_n = out_dist_12__empty_n;
  assign out_dist_12__read = krnl_globalSort_L1_L2_4_in_dist0_s_read;
  assign krnl_globalSort_L1_L2_4_in_dist1_peek_dout = out_dist_13__dout;
  assign krnl_globalSort_L1_L2_4_in_dist1_peek_empty_n = out_dist_13__empty_n;
  assign krnl_globalSort_L1_L2_4_in_dist1_s_dout = out_dist_13__dout;
  assign krnl_globalSort_L1_L2_4_in_dist1_s_empty_n = out_dist_13__empty_n;
  assign out_dist_13__read = krnl_globalSort_L1_L2_4_in_dist1_s_read;
  assign krnl_globalSort_L1_L2_4_in_dist2_peek_dout = out_dist_14__dout;
  assign krnl_globalSort_L1_L2_4_in_dist2_peek_empty_n = out_dist_14__empty_n;
  assign krnl_globalSort_L1_L2_4_in_dist2_s_dout = out_dist_14__dout;
  assign krnl_globalSort_L1_L2_4_in_dist2_s_empty_n = out_dist_14__empty_n;
  assign out_dist_14__read = krnl_globalSort_L1_L2_4_in_dist2_s_read;
  assign krnl_globalSort_L1_L2_4_in_id0_peek_dout = out_id_12__dout;
  assign krnl_globalSort_L1_L2_4_in_id0_peek_empty_n = out_id_12__empty_n;
  assign krnl_globalSort_L1_L2_4_in_id0_s_dout = out_id_12__dout;
  assign krnl_globalSort_L1_L2_4_in_id0_s_empty_n = out_id_12__empty_n;
  assign out_id_12__read = krnl_globalSort_L1_L2_4_in_id0_s_read;
  assign krnl_globalSort_L1_L2_4_in_id1_peek_dout = out_id_13__dout;
  assign krnl_globalSort_L1_L2_4_in_id1_peek_empty_n = out_id_13__empty_n;
  assign krnl_globalSort_L1_L2_4_in_id1_s_dout = out_id_13__dout;
  assign krnl_globalSort_L1_L2_4_in_id1_s_empty_n = out_id_13__empty_n;
  assign out_id_13__read = krnl_globalSort_L1_L2_4_in_id1_s_read;
  assign krnl_globalSort_L1_L2_4_in_id2_peek_dout = out_id_14__dout;
  assign krnl_globalSort_L1_L2_4_in_id2_peek_empty_n = out_id_14__empty_n;
  assign krnl_globalSort_L1_L2_4_in_id2_s_dout = out_id_14__dout;
  assign krnl_globalSort_L1_L2_4_in_id2_s_empty_n = out_id_14__empty_n;
  assign out_id_14__read = krnl_globalSort_L1_L2_4_in_id2_s_read;
  assign L1_out_dist_4__din = krnl_globalSort_L1_L2_4_out_dist_din;
  assign krnl_globalSort_L1_L2_4_out_dist_full_n = L1_out_dist_4__full_n;
  assign L1_out_dist_4__write = krnl_globalSort_L1_L2_4_out_dist_write;
  assign L1_out_id_4__din = krnl_globalSort_L1_L2_4_out_id_din;
  assign krnl_globalSort_L1_L2_4_out_id_full_n = L1_out_id_4__full_n;
  assign L1_out_id_4__write = krnl_globalSort_L1_L2_4_out_id_write;
  assign krnl_globalSort_L1_L2_5_ap_clk = ap_clk;
  assign krnl_globalSort_L1_L2_5__ap_done = krnl_globalSort_L1_L2_5_ap_done;
  assign krnl_globalSort_L1_L2_5__ap_idle = krnl_globalSort_L1_L2_5_ap_idle;
  assign krnl_globalSort_L1_L2_5__ap_ready = krnl_globalSort_L1_L2_5_ap_ready;
  assign krnl_globalSort_L1_L2_5_ap_rst_n = ap_rst_n;
  assign krnl_globalSort_L1_L2_5_ap_start = krnl_globalSort_L1_L2_5__ap_start;
  assign krnl_globalSort_L1_L2_5_in_dist0_peek_dout = out_dist_15__dout;
  assign krnl_globalSort_L1_L2_5_in_dist0_peek_empty_n = out_dist_15__empty_n;
  assign krnl_globalSort_L1_L2_5_in_dist0_s_dout = out_dist_15__dout;
  assign krnl_globalSort_L1_L2_5_in_dist0_s_empty_n = out_dist_15__empty_n;
  assign out_dist_15__read = krnl_globalSort_L1_L2_5_in_dist0_s_read;
  assign krnl_globalSort_L1_L2_5_in_dist1_peek_dout = out_dist_16__dout;
  assign krnl_globalSort_L1_L2_5_in_dist1_peek_empty_n = out_dist_16__empty_n;
  assign krnl_globalSort_L1_L2_5_in_dist1_s_dout = out_dist_16__dout;
  assign krnl_globalSort_L1_L2_5_in_dist1_s_empty_n = out_dist_16__empty_n;
  assign out_dist_16__read = krnl_globalSort_L1_L2_5_in_dist1_s_read;
  assign krnl_globalSort_L1_L2_5_in_dist2_peek_dout = out_dist_17__dout;
  assign krnl_globalSort_L1_L2_5_in_dist2_peek_empty_n = out_dist_17__empty_n;
  assign krnl_globalSort_L1_L2_5_in_dist2_s_dout = out_dist_17__dout;
  assign krnl_globalSort_L1_L2_5_in_dist2_s_empty_n = out_dist_17__empty_n;
  assign out_dist_17__read = krnl_globalSort_L1_L2_5_in_dist2_s_read;
  assign krnl_globalSort_L1_L2_5_in_id0_peek_dout = out_id_15__dout;
  assign krnl_globalSort_L1_L2_5_in_id0_peek_empty_n = out_id_15__empty_n;
  assign krnl_globalSort_L1_L2_5_in_id0_s_dout = out_id_15__dout;
  assign krnl_globalSort_L1_L2_5_in_id0_s_empty_n = out_id_15__empty_n;
  assign out_id_15__read = krnl_globalSort_L1_L2_5_in_id0_s_read;
  assign krnl_globalSort_L1_L2_5_in_id1_peek_dout = out_id_16__dout;
  assign krnl_globalSort_L1_L2_5_in_id1_peek_empty_n = out_id_16__empty_n;
  assign krnl_globalSort_L1_L2_5_in_id1_s_dout = out_id_16__dout;
  assign krnl_globalSort_L1_L2_5_in_id1_s_empty_n = out_id_16__empty_n;
  assign out_id_16__read = krnl_globalSort_L1_L2_5_in_id1_s_read;
  assign krnl_globalSort_L1_L2_5_in_id2_peek_dout = out_id_17__dout;
  assign krnl_globalSort_L1_L2_5_in_id2_peek_empty_n = out_id_17__empty_n;
  assign krnl_globalSort_L1_L2_5_in_id2_s_dout = out_id_17__dout;
  assign krnl_globalSort_L1_L2_5_in_id2_s_empty_n = out_id_17__empty_n;
  assign out_id_17__read = krnl_globalSort_L1_L2_5_in_id2_s_read;
  assign L1_out_dist_5__din = krnl_globalSort_L1_L2_5_out_dist_din;
  assign krnl_globalSort_L1_L2_5_out_dist_full_n = L1_out_dist_5__full_n;
  assign L1_out_dist_5__write = krnl_globalSort_L1_L2_5_out_dist_write;
  assign L1_out_id_5__din = krnl_globalSort_L1_L2_5_out_id_din;
  assign krnl_globalSort_L1_L2_5_out_id_full_n = L1_out_id_5__full_n;
  assign L1_out_id_5__write = krnl_globalSort_L1_L2_5_out_id_write;
  assign krnl_globalSort_L1_L2_6_ap_clk = ap_clk;
  assign krnl_globalSort_L1_L2_6__ap_done = krnl_globalSort_L1_L2_6_ap_done;
  assign krnl_globalSort_L1_L2_6__ap_idle = krnl_globalSort_L1_L2_6_ap_idle;
  assign krnl_globalSort_L1_L2_6__ap_ready = krnl_globalSort_L1_L2_6_ap_ready;
  assign krnl_globalSort_L1_L2_6_ap_rst_n = ap_rst_n;
  assign krnl_globalSort_L1_L2_6_ap_start = krnl_globalSort_L1_L2_6__ap_start;
  assign krnl_globalSort_L1_L2_6_in_dist0_peek_dout = out_dist_18__dout;
  assign krnl_globalSort_L1_L2_6_in_dist0_peek_empty_n = out_dist_18__empty_n;
  assign krnl_globalSort_L1_L2_6_in_dist0_s_dout = out_dist_18__dout;
  assign krnl_globalSort_L1_L2_6_in_dist0_s_empty_n = out_dist_18__empty_n;
  assign out_dist_18__read = krnl_globalSort_L1_L2_6_in_dist0_s_read;
  assign krnl_globalSort_L1_L2_6_in_dist1_peek_dout = out_dist_19__dout;
  assign krnl_globalSort_L1_L2_6_in_dist1_peek_empty_n = out_dist_19__empty_n;
  assign krnl_globalSort_L1_L2_6_in_dist1_s_dout = out_dist_19__dout;
  assign krnl_globalSort_L1_L2_6_in_dist1_s_empty_n = out_dist_19__empty_n;
  assign out_dist_19__read = krnl_globalSort_L1_L2_6_in_dist1_s_read;
  assign krnl_globalSort_L1_L2_6_in_dist2_peek_dout = out_dist_20__dout;
  assign krnl_globalSort_L1_L2_6_in_dist2_peek_empty_n = out_dist_20__empty_n;
  assign krnl_globalSort_L1_L2_6_in_dist2_s_dout = out_dist_20__dout;
  assign krnl_globalSort_L1_L2_6_in_dist2_s_empty_n = out_dist_20__empty_n;
  assign out_dist_20__read = krnl_globalSort_L1_L2_6_in_dist2_s_read;
  assign krnl_globalSort_L1_L2_6_in_id0_peek_dout = out_id_18__dout;
  assign krnl_globalSort_L1_L2_6_in_id0_peek_empty_n = out_id_18__empty_n;
  assign krnl_globalSort_L1_L2_6_in_id0_s_dout = out_id_18__dout;
  assign krnl_globalSort_L1_L2_6_in_id0_s_empty_n = out_id_18__empty_n;
  assign out_id_18__read = krnl_globalSort_L1_L2_6_in_id0_s_read;
  assign krnl_globalSort_L1_L2_6_in_id1_peek_dout = out_id_19__dout;
  assign krnl_globalSort_L1_L2_6_in_id1_peek_empty_n = out_id_19__empty_n;
  assign krnl_globalSort_L1_L2_6_in_id1_s_dout = out_id_19__dout;
  assign krnl_globalSort_L1_L2_6_in_id1_s_empty_n = out_id_19__empty_n;
  assign out_id_19__read = krnl_globalSort_L1_L2_6_in_id1_s_read;
  assign krnl_globalSort_L1_L2_6_in_id2_peek_dout = out_id_20__dout;
  assign krnl_globalSort_L1_L2_6_in_id2_peek_empty_n = out_id_20__empty_n;
  assign krnl_globalSort_L1_L2_6_in_id2_s_dout = out_id_20__dout;
  assign krnl_globalSort_L1_L2_6_in_id2_s_empty_n = out_id_20__empty_n;
  assign out_id_20__read = krnl_globalSort_L1_L2_6_in_id2_s_read;
  assign L1_out_dist_6__din = krnl_globalSort_L1_L2_6_out_dist_din;
  assign krnl_globalSort_L1_L2_6_out_dist_full_n = L1_out_dist_6__full_n;
  assign L1_out_dist_6__write = krnl_globalSort_L1_L2_6_out_dist_write;
  assign L1_out_id_6__din = krnl_globalSort_L1_L2_6_out_id_din;
  assign krnl_globalSort_L1_L2_6_out_id_full_n = L1_out_id_6__full_n;
  assign L1_out_id_6__write = krnl_globalSort_L1_L2_6_out_id_write;
  assign krnl_globalSort_L1_L2_7_ap_clk = ap_clk;
  assign krnl_globalSort_L1_L2_7__ap_done = krnl_globalSort_L1_L2_7_ap_done;
  assign krnl_globalSort_L1_L2_7__ap_idle = krnl_globalSort_L1_L2_7_ap_idle;
  assign krnl_globalSort_L1_L2_7__ap_ready = krnl_globalSort_L1_L2_7_ap_ready;
  assign krnl_globalSort_L1_L2_7_ap_rst_n = ap_rst_n;
  assign krnl_globalSort_L1_L2_7_ap_start = krnl_globalSort_L1_L2_7__ap_start;
  assign krnl_globalSort_L1_L2_7_in_dist0_peek_dout = out_dist_21__dout;
  assign krnl_globalSort_L1_L2_7_in_dist0_peek_empty_n = out_dist_21__empty_n;
  assign krnl_globalSort_L1_L2_7_in_dist0_s_dout = out_dist_21__dout;
  assign krnl_globalSort_L1_L2_7_in_dist0_s_empty_n = out_dist_21__empty_n;
  assign out_dist_21__read = krnl_globalSort_L1_L2_7_in_dist0_s_read;
  assign krnl_globalSort_L1_L2_7_in_dist1_peek_dout = out_dist_22__dout;
  assign krnl_globalSort_L1_L2_7_in_dist1_peek_empty_n = out_dist_22__empty_n;
  assign krnl_globalSort_L1_L2_7_in_dist1_s_dout = out_dist_22__dout;
  assign krnl_globalSort_L1_L2_7_in_dist1_s_empty_n = out_dist_22__empty_n;
  assign out_dist_22__read = krnl_globalSort_L1_L2_7_in_dist1_s_read;
  assign krnl_globalSort_L1_L2_7_in_dist2_peek_dout = out_dist_23__dout;
  assign krnl_globalSort_L1_L2_7_in_dist2_peek_empty_n = out_dist_23__empty_n;
  assign krnl_globalSort_L1_L2_7_in_dist2_s_dout = out_dist_23__dout;
  assign krnl_globalSort_L1_L2_7_in_dist2_s_empty_n = out_dist_23__empty_n;
  assign out_dist_23__read = krnl_globalSort_L1_L2_7_in_dist2_s_read;
  assign krnl_globalSort_L1_L2_7_in_id0_peek_dout = out_id_21__dout;
  assign krnl_globalSort_L1_L2_7_in_id0_peek_empty_n = out_id_21__empty_n;
  assign krnl_globalSort_L1_L2_7_in_id0_s_dout = out_id_21__dout;
  assign krnl_globalSort_L1_L2_7_in_id0_s_empty_n = out_id_21__empty_n;
  assign out_id_21__read = krnl_globalSort_L1_L2_7_in_id0_s_read;
  assign krnl_globalSort_L1_L2_7_in_id1_peek_dout = out_id_22__dout;
  assign krnl_globalSort_L1_L2_7_in_id1_peek_empty_n = out_id_22__empty_n;
  assign krnl_globalSort_L1_L2_7_in_id1_s_dout = out_id_22__dout;
  assign krnl_globalSort_L1_L2_7_in_id1_s_empty_n = out_id_22__empty_n;
  assign out_id_22__read = krnl_globalSort_L1_L2_7_in_id1_s_read;
  assign krnl_globalSort_L1_L2_7_in_id2_peek_dout = out_id_23__dout;
  assign krnl_globalSort_L1_L2_7_in_id2_peek_empty_n = out_id_23__empty_n;
  assign krnl_globalSort_L1_L2_7_in_id2_s_dout = out_id_23__dout;
  assign krnl_globalSort_L1_L2_7_in_id2_s_empty_n = out_id_23__empty_n;
  assign out_id_23__read = krnl_globalSort_L1_L2_7_in_id2_s_read;
  assign L1_out_dist_7__din = krnl_globalSort_L1_L2_7_out_dist_din;
  assign krnl_globalSort_L1_L2_7_out_dist_full_n = L1_out_dist_7__full_n;
  assign L1_out_dist_7__write = krnl_globalSort_L1_L2_7_out_dist_write;
  assign L1_out_id_7__din = krnl_globalSort_L1_L2_7_out_id_din;
  assign krnl_globalSort_L1_L2_7_out_id_full_n = L1_out_id_7__full_n;
  assign L1_out_id_7__write = krnl_globalSort_L1_L2_7_out_id_write;
  assign krnl_globalSort_L1_L2_8_ap_clk = ap_clk;
  assign krnl_globalSort_L1_L2_8__ap_done = krnl_globalSort_L1_L2_8_ap_done;
  assign krnl_globalSort_L1_L2_8__ap_idle = krnl_globalSort_L1_L2_8_ap_idle;
  assign krnl_globalSort_L1_L2_8__ap_ready = krnl_globalSort_L1_L2_8_ap_ready;
  assign krnl_globalSort_L1_L2_8_ap_rst_n = ap_rst_n;
  assign krnl_globalSort_L1_L2_8_ap_start = krnl_globalSort_L1_L2_8__ap_start;
  assign krnl_globalSort_L1_L2_8_in_dist0_peek_dout = out_dist_24__dout;
  assign krnl_globalSort_L1_L2_8_in_dist0_peek_empty_n = out_dist_24__empty_n;
  assign krnl_globalSort_L1_L2_8_in_dist0_s_dout = out_dist_24__dout;
  assign krnl_globalSort_L1_L2_8_in_dist0_s_empty_n = out_dist_24__empty_n;
  assign out_dist_24__read = krnl_globalSort_L1_L2_8_in_dist0_s_read;
  assign krnl_globalSort_L1_L2_8_in_dist1_peek_dout = out_dist_25__dout;
  assign krnl_globalSort_L1_L2_8_in_dist1_peek_empty_n = out_dist_25__empty_n;
  assign krnl_globalSort_L1_L2_8_in_dist1_s_dout = out_dist_25__dout;
  assign krnl_globalSort_L1_L2_8_in_dist1_s_empty_n = out_dist_25__empty_n;
  assign out_dist_25__read = krnl_globalSort_L1_L2_8_in_dist1_s_read;
  assign krnl_globalSort_L1_L2_8_in_dist2_peek_dout = out_dist_26__dout;
  assign krnl_globalSort_L1_L2_8_in_dist2_peek_empty_n = out_dist_26__empty_n;
  assign krnl_globalSort_L1_L2_8_in_dist2_s_dout = out_dist_26__dout;
  assign krnl_globalSort_L1_L2_8_in_dist2_s_empty_n = out_dist_26__empty_n;
  assign out_dist_26__read = krnl_globalSort_L1_L2_8_in_dist2_s_read;
  assign krnl_globalSort_L1_L2_8_in_id0_peek_dout = out_id_24__dout;
  assign krnl_globalSort_L1_L2_8_in_id0_peek_empty_n = out_id_24__empty_n;
  assign krnl_globalSort_L1_L2_8_in_id0_s_dout = out_id_24__dout;
  assign krnl_globalSort_L1_L2_8_in_id0_s_empty_n = out_id_24__empty_n;
  assign out_id_24__read = krnl_globalSort_L1_L2_8_in_id0_s_read;
  assign krnl_globalSort_L1_L2_8_in_id1_peek_dout = out_id_25__dout;
  assign krnl_globalSort_L1_L2_8_in_id1_peek_empty_n = out_id_25__empty_n;
  assign krnl_globalSort_L1_L2_8_in_id1_s_dout = out_id_25__dout;
  assign krnl_globalSort_L1_L2_8_in_id1_s_empty_n = out_id_25__empty_n;
  assign out_id_25__read = krnl_globalSort_L1_L2_8_in_id1_s_read;
  assign krnl_globalSort_L1_L2_8_in_id2_peek_dout = out_id_26__dout;
  assign krnl_globalSort_L1_L2_8_in_id2_peek_empty_n = out_id_26__empty_n;
  assign krnl_globalSort_L1_L2_8_in_id2_s_dout = out_id_26__dout;
  assign krnl_globalSort_L1_L2_8_in_id2_s_empty_n = out_id_26__empty_n;
  assign out_id_26__read = krnl_globalSort_L1_L2_8_in_id2_s_read;
  assign L1_out_dist_8__din = krnl_globalSort_L1_L2_8_out_dist_din;
  assign krnl_globalSort_L1_L2_8_out_dist_full_n = L1_out_dist_8__full_n;
  assign L1_out_dist_8__write = krnl_globalSort_L1_L2_8_out_dist_write;
  assign L1_out_id_8__din = krnl_globalSort_L1_L2_8_out_id_din;
  assign krnl_globalSort_L1_L2_8_out_id_full_n = L1_out_id_8__full_n;
  assign L1_out_id_8__write = krnl_globalSort_L1_L2_8_out_id_write;
  assign krnl_globalSort_L1_L2_9_ap_clk = ap_clk;
  assign krnl_globalSort_L1_L2_9__ap_done = krnl_globalSort_L1_L2_9_ap_done;
  assign krnl_globalSort_L1_L2_9__ap_idle = krnl_globalSort_L1_L2_9_ap_idle;
  assign krnl_globalSort_L1_L2_9__ap_ready = krnl_globalSort_L1_L2_9_ap_ready;
  assign krnl_globalSort_L1_L2_9_ap_rst_n = ap_rst_n;
  assign krnl_globalSort_L1_L2_9_ap_start = krnl_globalSort_L1_L2_9__ap_start;
  assign krnl_globalSort_L1_L2_9_in_dist0_peek_dout = out_dist_27__dout;
  assign krnl_globalSort_L1_L2_9_in_dist0_peek_empty_n = out_dist_27__empty_n;
  assign krnl_globalSort_L1_L2_9_in_dist0_s_dout = out_dist_27__dout;
  assign krnl_globalSort_L1_L2_9_in_dist0_s_empty_n = out_dist_27__empty_n;
  assign out_dist_27__read = krnl_globalSort_L1_L2_9_in_dist0_s_read;
  assign krnl_globalSort_L1_L2_9_in_dist1_peek_dout = out_dist_28__dout;
  assign krnl_globalSort_L1_L2_9_in_dist1_peek_empty_n = out_dist_28__empty_n;
  assign krnl_globalSort_L1_L2_9_in_dist1_s_dout = out_dist_28__dout;
  assign krnl_globalSort_L1_L2_9_in_dist1_s_empty_n = out_dist_28__empty_n;
  assign out_dist_28__read = krnl_globalSort_L1_L2_9_in_dist1_s_read;
  assign krnl_globalSort_L1_L2_9_in_dist2_peek_dout = out_dist_29__dout;
  assign krnl_globalSort_L1_L2_9_in_dist2_peek_empty_n = out_dist_29__empty_n;
  assign krnl_globalSort_L1_L2_9_in_dist2_s_dout = out_dist_29__dout;
  assign krnl_globalSort_L1_L2_9_in_dist2_s_empty_n = out_dist_29__empty_n;
  assign out_dist_29__read = krnl_globalSort_L1_L2_9_in_dist2_s_read;
  assign krnl_globalSort_L1_L2_9_in_id0_peek_dout = out_id_27__dout;
  assign krnl_globalSort_L1_L2_9_in_id0_peek_empty_n = out_id_27__empty_n;
  assign krnl_globalSort_L1_L2_9_in_id0_s_dout = out_id_27__dout;
  assign krnl_globalSort_L1_L2_9_in_id0_s_empty_n = out_id_27__empty_n;
  assign out_id_27__read = krnl_globalSort_L1_L2_9_in_id0_s_read;
  assign krnl_globalSort_L1_L2_9_in_id1_peek_dout = out_id_28__dout;
  assign krnl_globalSort_L1_L2_9_in_id1_peek_empty_n = out_id_28__empty_n;
  assign krnl_globalSort_L1_L2_9_in_id1_s_dout = out_id_28__dout;
  assign krnl_globalSort_L1_L2_9_in_id1_s_empty_n = out_id_28__empty_n;
  assign out_id_28__read = krnl_globalSort_L1_L2_9_in_id1_s_read;
  assign krnl_globalSort_L1_L2_9_in_id2_peek_dout = out_id_29__dout;
  assign krnl_globalSort_L1_L2_9_in_id2_peek_empty_n = out_id_29__empty_n;
  assign krnl_globalSort_L1_L2_9_in_id2_s_dout = out_id_29__dout;
  assign krnl_globalSort_L1_L2_9_in_id2_s_empty_n = out_id_29__empty_n;
  assign out_id_29__read = krnl_globalSort_L1_L2_9_in_id2_s_read;
  assign L1_out_dist_9__din = krnl_globalSort_L1_L2_9_out_dist_din;
  assign krnl_globalSort_L1_L2_9_out_dist_full_n = L1_out_dist_9__full_n;
  assign L1_out_dist_9__write = krnl_globalSort_L1_L2_9_out_dist_write;
  assign L1_out_id_9__din = krnl_globalSort_L1_L2_9_out_id_din;
  assign krnl_globalSort_L1_L2_9_out_id_full_n = L1_out_id_9__full_n;
  assign L1_out_id_9__write = krnl_globalSort_L1_L2_9_out_id_write;
  assign krnl_globalSort_L1_L2_10_ap_clk = ap_clk;
  assign krnl_globalSort_L1_L2_10__ap_done = krnl_globalSort_L1_L2_10_ap_done;
  assign krnl_globalSort_L1_L2_10__ap_idle = krnl_globalSort_L1_L2_10_ap_idle;
  assign krnl_globalSort_L1_L2_10__ap_ready = krnl_globalSort_L1_L2_10_ap_ready;
  assign krnl_globalSort_L1_L2_10_ap_rst_n = ap_rst_n;
  assign krnl_globalSort_L1_L2_10_ap_start = krnl_globalSort_L1_L2_10__ap_start;
  assign krnl_globalSort_L1_L2_10_in_dist0_peek_dout = out_dist_30__dout;
  assign krnl_globalSort_L1_L2_10_in_dist0_peek_empty_n = out_dist_30__empty_n;
  assign krnl_globalSort_L1_L2_10_in_dist0_s_dout = out_dist_30__dout;
  assign krnl_globalSort_L1_L2_10_in_dist0_s_empty_n = out_dist_30__empty_n;
  assign out_dist_30__read = krnl_globalSort_L1_L2_10_in_dist0_s_read;
  assign krnl_globalSort_L1_L2_10_in_dist1_peek_dout = out_dist_31__dout;
  assign krnl_globalSort_L1_L2_10_in_dist1_peek_empty_n = out_dist_31__empty_n;
  assign krnl_globalSort_L1_L2_10_in_dist1_s_dout = out_dist_31__dout;
  assign krnl_globalSort_L1_L2_10_in_dist1_s_empty_n = out_dist_31__empty_n;
  assign out_dist_31__read = krnl_globalSort_L1_L2_10_in_dist1_s_read;
  assign krnl_globalSort_L1_L2_10_in_dist2_peek_dout = out_dist_32__dout;
  assign krnl_globalSort_L1_L2_10_in_dist2_peek_empty_n = out_dist_32__empty_n;
  assign krnl_globalSort_L1_L2_10_in_dist2_s_dout = out_dist_32__dout;
  assign krnl_globalSort_L1_L2_10_in_dist2_s_empty_n = out_dist_32__empty_n;
  assign out_dist_32__read = krnl_globalSort_L1_L2_10_in_dist2_s_read;
  assign krnl_globalSort_L1_L2_10_in_id0_peek_dout = out_id_30__dout;
  assign krnl_globalSort_L1_L2_10_in_id0_peek_empty_n = out_id_30__empty_n;
  assign krnl_globalSort_L1_L2_10_in_id0_s_dout = out_id_30__dout;
  assign krnl_globalSort_L1_L2_10_in_id0_s_empty_n = out_id_30__empty_n;
  assign out_id_30__read = krnl_globalSort_L1_L2_10_in_id0_s_read;
  assign krnl_globalSort_L1_L2_10_in_id1_peek_dout = out_id_31__dout;
  assign krnl_globalSort_L1_L2_10_in_id1_peek_empty_n = out_id_31__empty_n;
  assign krnl_globalSort_L1_L2_10_in_id1_s_dout = out_id_31__dout;
  assign krnl_globalSort_L1_L2_10_in_id1_s_empty_n = out_id_31__empty_n;
  assign out_id_31__read = krnl_globalSort_L1_L2_10_in_id1_s_read;
  assign krnl_globalSort_L1_L2_10_in_id2_peek_dout = out_id_32__dout;
  assign krnl_globalSort_L1_L2_10_in_id2_peek_empty_n = out_id_32__empty_n;
  assign krnl_globalSort_L1_L2_10_in_id2_s_dout = out_id_32__dout;
  assign krnl_globalSort_L1_L2_10_in_id2_s_empty_n = out_id_32__empty_n;
  assign out_id_32__read = krnl_globalSort_L1_L2_10_in_id2_s_read;
  assign L1_out_dist_10__din = krnl_globalSort_L1_L2_10_out_dist_din;
  assign krnl_globalSort_L1_L2_10_out_dist_full_n = L1_out_dist_10__full_n;
  assign L1_out_dist_10__write = krnl_globalSort_L1_L2_10_out_dist_write;
  assign L1_out_id_10__din = krnl_globalSort_L1_L2_10_out_id_din;
  assign krnl_globalSort_L1_L2_10_out_id_full_n = L1_out_id_10__full_n;
  assign L1_out_id_10__write = krnl_globalSort_L1_L2_10_out_id_write;
  assign krnl_globalSort_L1_L2_11_ap_clk = ap_clk;
  assign krnl_globalSort_L1_L2_11__ap_done = krnl_globalSort_L1_L2_11_ap_done;
  assign krnl_globalSort_L1_L2_11__ap_idle = krnl_globalSort_L1_L2_11_ap_idle;
  assign krnl_globalSort_L1_L2_11__ap_ready = krnl_globalSort_L1_L2_11_ap_ready;
  assign krnl_globalSort_L1_L2_11_ap_rst_n = ap_rst_n;
  assign krnl_globalSort_L1_L2_11_ap_start = krnl_globalSort_L1_L2_11__ap_start;
  assign krnl_globalSort_L1_L2_11_in_dist0_peek_dout = out_dist_33__dout;
  assign krnl_globalSort_L1_L2_11_in_dist0_peek_empty_n = out_dist_33__empty_n;
  assign krnl_globalSort_L1_L2_11_in_dist0_s_dout = out_dist_33__dout;
  assign krnl_globalSort_L1_L2_11_in_dist0_s_empty_n = out_dist_33__empty_n;
  assign out_dist_33__read = krnl_globalSort_L1_L2_11_in_dist0_s_read;
  assign krnl_globalSort_L1_L2_11_in_dist1_peek_dout = out_dist_34__dout;
  assign krnl_globalSort_L1_L2_11_in_dist1_peek_empty_n = out_dist_34__empty_n;
  assign krnl_globalSort_L1_L2_11_in_dist1_s_dout = out_dist_34__dout;
  assign krnl_globalSort_L1_L2_11_in_dist1_s_empty_n = out_dist_34__empty_n;
  assign out_dist_34__read = krnl_globalSort_L1_L2_11_in_dist1_s_read;
  assign krnl_globalSort_L1_L2_11_in_dist2_peek_dout = out_dist_35__dout;
  assign krnl_globalSort_L1_L2_11_in_dist2_peek_empty_n = out_dist_35__empty_n;
  assign krnl_globalSort_L1_L2_11_in_dist2_s_dout = out_dist_35__dout;
  assign krnl_globalSort_L1_L2_11_in_dist2_s_empty_n = out_dist_35__empty_n;
  assign out_dist_35__read = krnl_globalSort_L1_L2_11_in_dist2_s_read;
  assign krnl_globalSort_L1_L2_11_in_id0_peek_dout = out_id_33__dout;
  assign krnl_globalSort_L1_L2_11_in_id0_peek_empty_n = out_id_33__empty_n;
  assign krnl_globalSort_L1_L2_11_in_id0_s_dout = out_id_33__dout;
  assign krnl_globalSort_L1_L2_11_in_id0_s_empty_n = out_id_33__empty_n;
  assign out_id_33__read = krnl_globalSort_L1_L2_11_in_id0_s_read;
  assign krnl_globalSort_L1_L2_11_in_id1_peek_dout = out_id_34__dout;
  assign krnl_globalSort_L1_L2_11_in_id1_peek_empty_n = out_id_34__empty_n;
  assign krnl_globalSort_L1_L2_11_in_id1_s_dout = out_id_34__dout;
  assign krnl_globalSort_L1_L2_11_in_id1_s_empty_n = out_id_34__empty_n;
  assign out_id_34__read = krnl_globalSort_L1_L2_11_in_id1_s_read;
  assign krnl_globalSort_L1_L2_11_in_id2_peek_dout = out_id_35__dout;
  assign krnl_globalSort_L1_L2_11_in_id2_peek_empty_n = out_id_35__empty_n;
  assign krnl_globalSort_L1_L2_11_in_id2_s_dout = out_id_35__dout;
  assign krnl_globalSort_L1_L2_11_in_id2_s_empty_n = out_id_35__empty_n;
  assign out_id_35__read = krnl_globalSort_L1_L2_11_in_id2_s_read;
  assign L1_out_dist_11__din = krnl_globalSort_L1_L2_11_out_dist_din;
  assign krnl_globalSort_L1_L2_11_out_dist_full_n = L1_out_dist_11__full_n;
  assign L1_out_dist_11__write = krnl_globalSort_L1_L2_11_out_dist_write;
  assign L1_out_id_11__din = krnl_globalSort_L1_L2_11_out_id_din;
  assign krnl_globalSort_L1_L2_11_out_id_full_n = L1_out_id_11__full_n;
  assign L1_out_id_11__write = krnl_globalSort_L1_L2_11_out_id_write;
  assign krnl_globalSort_L1_L2_12_ap_clk = ap_clk;
  assign krnl_globalSort_L1_L2_12__ap_done = krnl_globalSort_L1_L2_12_ap_done;
  assign krnl_globalSort_L1_L2_12__ap_idle = krnl_globalSort_L1_L2_12_ap_idle;
  assign krnl_globalSort_L1_L2_12__ap_ready = krnl_globalSort_L1_L2_12_ap_ready;
  assign krnl_globalSort_L1_L2_12_ap_rst_n = ap_rst_n;
  assign krnl_globalSort_L1_L2_12_ap_start = krnl_globalSort_L1_L2_12__ap_start;
  assign krnl_globalSort_L1_L2_12_in_dist0_peek_dout = out_dist_36__dout;
  assign krnl_globalSort_L1_L2_12_in_dist0_peek_empty_n = out_dist_36__empty_n;
  assign krnl_globalSort_L1_L2_12_in_dist0_s_dout = out_dist_36__dout;
  assign krnl_globalSort_L1_L2_12_in_dist0_s_empty_n = out_dist_36__empty_n;
  assign out_dist_36__read = krnl_globalSort_L1_L2_12_in_dist0_s_read;
  assign krnl_globalSort_L1_L2_12_in_dist1_peek_dout = out_dist_37__dout;
  assign krnl_globalSort_L1_L2_12_in_dist1_peek_empty_n = out_dist_37__empty_n;
  assign krnl_globalSort_L1_L2_12_in_dist1_s_dout = out_dist_37__dout;
  assign krnl_globalSort_L1_L2_12_in_dist1_s_empty_n = out_dist_37__empty_n;
  assign out_dist_37__read = krnl_globalSort_L1_L2_12_in_dist1_s_read;
  assign krnl_globalSort_L1_L2_12_in_dist2_peek_dout = out_dist_38__dout;
  assign krnl_globalSort_L1_L2_12_in_dist2_peek_empty_n = out_dist_38__empty_n;
  assign krnl_globalSort_L1_L2_12_in_dist2_s_dout = out_dist_38__dout;
  assign krnl_globalSort_L1_L2_12_in_dist2_s_empty_n = out_dist_38__empty_n;
  assign out_dist_38__read = krnl_globalSort_L1_L2_12_in_dist2_s_read;
  assign krnl_globalSort_L1_L2_12_in_id0_peek_dout = out_id_36__dout;
  assign krnl_globalSort_L1_L2_12_in_id0_peek_empty_n = out_id_36__empty_n;
  assign krnl_globalSort_L1_L2_12_in_id0_s_dout = out_id_36__dout;
  assign krnl_globalSort_L1_L2_12_in_id0_s_empty_n = out_id_36__empty_n;
  assign out_id_36__read = krnl_globalSort_L1_L2_12_in_id0_s_read;
  assign krnl_globalSort_L1_L2_12_in_id1_peek_dout = out_id_37__dout;
  assign krnl_globalSort_L1_L2_12_in_id1_peek_empty_n = out_id_37__empty_n;
  assign krnl_globalSort_L1_L2_12_in_id1_s_dout = out_id_37__dout;
  assign krnl_globalSort_L1_L2_12_in_id1_s_empty_n = out_id_37__empty_n;
  assign out_id_37__read = krnl_globalSort_L1_L2_12_in_id1_s_read;
  assign krnl_globalSort_L1_L2_12_in_id2_peek_dout = out_id_38__dout;
  assign krnl_globalSort_L1_L2_12_in_id2_peek_empty_n = out_id_38__empty_n;
  assign krnl_globalSort_L1_L2_12_in_id2_s_dout = out_id_38__dout;
  assign krnl_globalSort_L1_L2_12_in_id2_s_empty_n = out_id_38__empty_n;
  assign out_id_38__read = krnl_globalSort_L1_L2_12_in_id2_s_read;
  assign L1_out_dist_12__din = krnl_globalSort_L1_L2_12_out_dist_din;
  assign krnl_globalSort_L1_L2_12_out_dist_full_n = L1_out_dist_12__full_n;
  assign L1_out_dist_12__write = krnl_globalSort_L1_L2_12_out_dist_write;
  assign L1_out_id_12__din = krnl_globalSort_L1_L2_12_out_id_din;
  assign krnl_globalSort_L1_L2_12_out_id_full_n = L1_out_id_12__full_n;
  assign L1_out_id_12__write = krnl_globalSort_L1_L2_12_out_id_write;
  assign krnl_globalSort_L1_L2_13_ap_clk = ap_clk;
  assign krnl_globalSort_L1_L2_13__ap_done = krnl_globalSort_L1_L2_13_ap_done;
  assign krnl_globalSort_L1_L2_13__ap_idle = krnl_globalSort_L1_L2_13_ap_idle;
  assign krnl_globalSort_L1_L2_13__ap_ready = krnl_globalSort_L1_L2_13_ap_ready;
  assign krnl_globalSort_L1_L2_13_ap_rst_n = ap_rst_n;
  assign krnl_globalSort_L1_L2_13_ap_start = krnl_globalSort_L1_L2_13__ap_start;
  assign krnl_globalSort_L1_L2_13_in_dist0_peek_dout = out_dist_39__dout;
  assign krnl_globalSort_L1_L2_13_in_dist0_peek_empty_n = out_dist_39__empty_n;
  assign krnl_globalSort_L1_L2_13_in_dist0_s_dout = out_dist_39__dout;
  assign krnl_globalSort_L1_L2_13_in_dist0_s_empty_n = out_dist_39__empty_n;
  assign out_dist_39__read = krnl_globalSort_L1_L2_13_in_dist0_s_read;
  assign krnl_globalSort_L1_L2_13_in_dist1_peek_dout = out_dist_40__dout;
  assign krnl_globalSort_L1_L2_13_in_dist1_peek_empty_n = out_dist_40__empty_n;
  assign krnl_globalSort_L1_L2_13_in_dist1_s_dout = out_dist_40__dout;
  assign krnl_globalSort_L1_L2_13_in_dist1_s_empty_n = out_dist_40__empty_n;
  assign out_dist_40__read = krnl_globalSort_L1_L2_13_in_dist1_s_read;
  assign krnl_globalSort_L1_L2_13_in_dist2_peek_dout = out_dist_41__dout;
  assign krnl_globalSort_L1_L2_13_in_dist2_peek_empty_n = out_dist_41__empty_n;
  assign krnl_globalSort_L1_L2_13_in_dist2_s_dout = out_dist_41__dout;
  assign krnl_globalSort_L1_L2_13_in_dist2_s_empty_n = out_dist_41__empty_n;
  assign out_dist_41__read = krnl_globalSort_L1_L2_13_in_dist2_s_read;
  assign krnl_globalSort_L1_L2_13_in_id0_peek_dout = out_id_39__dout;
  assign krnl_globalSort_L1_L2_13_in_id0_peek_empty_n = out_id_39__empty_n;
  assign krnl_globalSort_L1_L2_13_in_id0_s_dout = out_id_39__dout;
  assign krnl_globalSort_L1_L2_13_in_id0_s_empty_n = out_id_39__empty_n;
  assign out_id_39__read = krnl_globalSort_L1_L2_13_in_id0_s_read;
  assign krnl_globalSort_L1_L2_13_in_id1_peek_dout = out_id_40__dout;
  assign krnl_globalSort_L1_L2_13_in_id1_peek_empty_n = out_id_40__empty_n;
  assign krnl_globalSort_L1_L2_13_in_id1_s_dout = out_id_40__dout;
  assign krnl_globalSort_L1_L2_13_in_id1_s_empty_n = out_id_40__empty_n;
  assign out_id_40__read = krnl_globalSort_L1_L2_13_in_id1_s_read;
  assign krnl_globalSort_L1_L2_13_in_id2_peek_dout = out_id_41__dout;
  assign krnl_globalSort_L1_L2_13_in_id2_peek_empty_n = out_id_41__empty_n;
  assign krnl_globalSort_L1_L2_13_in_id2_s_dout = out_id_41__dout;
  assign krnl_globalSort_L1_L2_13_in_id2_s_empty_n = out_id_41__empty_n;
  assign out_id_41__read = krnl_globalSort_L1_L2_13_in_id2_s_read;
  assign L1_out_dist_13__din = krnl_globalSort_L1_L2_13_out_dist_din;
  assign krnl_globalSort_L1_L2_13_out_dist_full_n = L1_out_dist_13__full_n;
  assign L1_out_dist_13__write = krnl_globalSort_L1_L2_13_out_dist_write;
  assign L1_out_id_13__din = krnl_globalSort_L1_L2_13_out_id_din;
  assign krnl_globalSort_L1_L2_13_out_id_full_n = L1_out_id_13__full_n;
  assign L1_out_id_13__write = krnl_globalSort_L1_L2_13_out_id_write;
  assign krnl_globalSort_L1_L2_14_ap_clk = ap_clk;
  assign krnl_globalSort_L1_L2_14__ap_done = krnl_globalSort_L1_L2_14_ap_done;
  assign krnl_globalSort_L1_L2_14__ap_idle = krnl_globalSort_L1_L2_14_ap_idle;
  assign krnl_globalSort_L1_L2_14__ap_ready = krnl_globalSort_L1_L2_14_ap_ready;
  assign krnl_globalSort_L1_L2_14_ap_rst_n = ap_rst_n;
  assign krnl_globalSort_L1_L2_14_ap_start = krnl_globalSort_L1_L2_14__ap_start;
  assign krnl_globalSort_L1_L2_14_in_dist0_peek_dout = out_dist_42__dout;
  assign krnl_globalSort_L1_L2_14_in_dist0_peek_empty_n = out_dist_42__empty_n;
  assign krnl_globalSort_L1_L2_14_in_dist0_s_dout = out_dist_42__dout;
  assign krnl_globalSort_L1_L2_14_in_dist0_s_empty_n = out_dist_42__empty_n;
  assign out_dist_42__read = krnl_globalSort_L1_L2_14_in_dist0_s_read;
  assign krnl_globalSort_L1_L2_14_in_dist1_peek_dout = out_dist_43__dout;
  assign krnl_globalSort_L1_L2_14_in_dist1_peek_empty_n = out_dist_43__empty_n;
  assign krnl_globalSort_L1_L2_14_in_dist1_s_dout = out_dist_43__dout;
  assign krnl_globalSort_L1_L2_14_in_dist1_s_empty_n = out_dist_43__empty_n;
  assign out_dist_43__read = krnl_globalSort_L1_L2_14_in_dist1_s_read;
  assign krnl_globalSort_L1_L2_14_in_dist2_peek_dout = out_dist_44__dout;
  assign krnl_globalSort_L1_L2_14_in_dist2_peek_empty_n = out_dist_44__empty_n;
  assign krnl_globalSort_L1_L2_14_in_dist2_s_dout = out_dist_44__dout;
  assign krnl_globalSort_L1_L2_14_in_dist2_s_empty_n = out_dist_44__empty_n;
  assign out_dist_44__read = krnl_globalSort_L1_L2_14_in_dist2_s_read;
  assign krnl_globalSort_L1_L2_14_in_id0_peek_dout = out_id_42__dout;
  assign krnl_globalSort_L1_L2_14_in_id0_peek_empty_n = out_id_42__empty_n;
  assign krnl_globalSort_L1_L2_14_in_id0_s_dout = out_id_42__dout;
  assign krnl_globalSort_L1_L2_14_in_id0_s_empty_n = out_id_42__empty_n;
  assign out_id_42__read = krnl_globalSort_L1_L2_14_in_id0_s_read;
  assign krnl_globalSort_L1_L2_14_in_id1_peek_dout = out_id_43__dout;
  assign krnl_globalSort_L1_L2_14_in_id1_peek_empty_n = out_id_43__empty_n;
  assign krnl_globalSort_L1_L2_14_in_id1_s_dout = out_id_43__dout;
  assign krnl_globalSort_L1_L2_14_in_id1_s_empty_n = out_id_43__empty_n;
  assign out_id_43__read = krnl_globalSort_L1_L2_14_in_id1_s_read;
  assign krnl_globalSort_L1_L2_14_in_id2_peek_dout = out_id_44__dout;
  assign krnl_globalSort_L1_L2_14_in_id2_peek_empty_n = out_id_44__empty_n;
  assign krnl_globalSort_L1_L2_14_in_id2_s_dout = out_id_44__dout;
  assign krnl_globalSort_L1_L2_14_in_id2_s_empty_n = out_id_44__empty_n;
  assign out_id_44__read = krnl_globalSort_L1_L2_14_in_id2_s_read;
  assign L1_out_dist_14__din = krnl_globalSort_L1_L2_14_out_dist_din;
  assign krnl_globalSort_L1_L2_14_out_dist_full_n = L1_out_dist_14__full_n;
  assign L1_out_dist_14__write = krnl_globalSort_L1_L2_14_out_dist_write;
  assign L1_out_id_14__din = krnl_globalSort_L1_L2_14_out_id_din;
  assign krnl_globalSort_L1_L2_14_out_id_full_n = L1_out_id_14__full_n;
  assign L1_out_id_14__write = krnl_globalSort_L1_L2_14_out_id_write;
  assign krnl_globalSort_L1_L2_15_ap_clk = ap_clk;
  assign krnl_globalSort_L1_L2_15__ap_done = krnl_globalSort_L1_L2_15_ap_done;
  assign krnl_globalSort_L1_L2_15__ap_idle = krnl_globalSort_L1_L2_15_ap_idle;
  assign krnl_globalSort_L1_L2_15__ap_ready = krnl_globalSort_L1_L2_15_ap_ready;
  assign krnl_globalSort_L1_L2_15_ap_rst_n = ap_rst_n;
  assign krnl_globalSort_L1_L2_15_ap_start = krnl_globalSort_L1_L2_15__ap_start;
  assign krnl_globalSort_L1_L2_15_in_dist0_peek_dout = out_dist_45__dout;
  assign krnl_globalSort_L1_L2_15_in_dist0_peek_empty_n = out_dist_45__empty_n;
  assign krnl_globalSort_L1_L2_15_in_dist0_s_dout = out_dist_45__dout;
  assign krnl_globalSort_L1_L2_15_in_dist0_s_empty_n = out_dist_45__empty_n;
  assign out_dist_45__read = krnl_globalSort_L1_L2_15_in_dist0_s_read;
  assign krnl_globalSort_L1_L2_15_in_dist1_peek_dout = out_dist_46__dout;
  assign krnl_globalSort_L1_L2_15_in_dist1_peek_empty_n = out_dist_46__empty_n;
  assign krnl_globalSort_L1_L2_15_in_dist1_s_dout = out_dist_46__dout;
  assign krnl_globalSort_L1_L2_15_in_dist1_s_empty_n = out_dist_46__empty_n;
  assign out_dist_46__read = krnl_globalSort_L1_L2_15_in_dist1_s_read;
  assign krnl_globalSort_L1_L2_15_in_dist2_peek_dout = out_dist_47__dout;
  assign krnl_globalSort_L1_L2_15_in_dist2_peek_empty_n = out_dist_47__empty_n;
  assign krnl_globalSort_L1_L2_15_in_dist2_s_dout = out_dist_47__dout;
  assign krnl_globalSort_L1_L2_15_in_dist2_s_empty_n = out_dist_47__empty_n;
  assign out_dist_47__read = krnl_globalSort_L1_L2_15_in_dist2_s_read;
  assign krnl_globalSort_L1_L2_15_in_id0_peek_dout = out_id_45__dout;
  assign krnl_globalSort_L1_L2_15_in_id0_peek_empty_n = out_id_45__empty_n;
  assign krnl_globalSort_L1_L2_15_in_id0_s_dout = out_id_45__dout;
  assign krnl_globalSort_L1_L2_15_in_id0_s_empty_n = out_id_45__empty_n;
  assign out_id_45__read = krnl_globalSort_L1_L2_15_in_id0_s_read;
  assign krnl_globalSort_L1_L2_15_in_id1_peek_dout = out_id_46__dout;
  assign krnl_globalSort_L1_L2_15_in_id1_peek_empty_n = out_id_46__empty_n;
  assign krnl_globalSort_L1_L2_15_in_id1_s_dout = out_id_46__dout;
  assign krnl_globalSort_L1_L2_15_in_id1_s_empty_n = out_id_46__empty_n;
  assign out_id_46__read = krnl_globalSort_L1_L2_15_in_id1_s_read;
  assign krnl_globalSort_L1_L2_15_in_id2_peek_dout = out_id_47__dout;
  assign krnl_globalSort_L1_L2_15_in_id2_peek_empty_n = out_id_47__empty_n;
  assign krnl_globalSort_L1_L2_15_in_id2_s_dout = out_id_47__dout;
  assign krnl_globalSort_L1_L2_15_in_id2_s_empty_n = out_id_47__empty_n;
  assign out_id_47__read = krnl_globalSort_L1_L2_15_in_id2_s_read;
  assign L1_out_dist_15__din = krnl_globalSort_L1_L2_15_out_dist_din;
  assign krnl_globalSort_L1_L2_15_out_dist_full_n = L1_out_dist_15__full_n;
  assign L1_out_dist_15__write = krnl_globalSort_L1_L2_15_out_dist_write;
  assign L1_out_id_15__din = krnl_globalSort_L1_L2_15_out_id_din;
  assign krnl_globalSort_L1_L2_15_out_id_full_n = L1_out_id_15__full_n;
  assign L1_out_id_15__write = krnl_globalSort_L1_L2_15_out_id_write;
  assign krnl_globalSort_L1_L2_16_ap_clk = ap_clk;
  assign krnl_globalSort_L1_L2_16__ap_done = krnl_globalSort_L1_L2_16_ap_done;
  assign krnl_globalSort_L1_L2_16__ap_idle = krnl_globalSort_L1_L2_16_ap_idle;
  assign krnl_globalSort_L1_L2_16__ap_ready = krnl_globalSort_L1_L2_16_ap_ready;
  assign krnl_globalSort_L1_L2_16_ap_rst_n = ap_rst_n;
  assign krnl_globalSort_L1_L2_16_ap_start = krnl_globalSort_L1_L2_16__ap_start;
  assign krnl_globalSort_L1_L2_16_in_dist0_peek_dout = out_dist_48__dout;
  assign krnl_globalSort_L1_L2_16_in_dist0_peek_empty_n = out_dist_48__empty_n;
  assign krnl_globalSort_L1_L2_16_in_dist0_s_dout = out_dist_48__dout;
  assign krnl_globalSort_L1_L2_16_in_dist0_s_empty_n = out_dist_48__empty_n;
  assign out_dist_48__read = krnl_globalSort_L1_L2_16_in_dist0_s_read;
  assign krnl_globalSort_L1_L2_16_in_dist1_peek_dout = out_dist_49__dout;
  assign krnl_globalSort_L1_L2_16_in_dist1_peek_empty_n = out_dist_49__empty_n;
  assign krnl_globalSort_L1_L2_16_in_dist1_s_dout = out_dist_49__dout;
  assign krnl_globalSort_L1_L2_16_in_dist1_s_empty_n = out_dist_49__empty_n;
  assign out_dist_49__read = krnl_globalSort_L1_L2_16_in_dist1_s_read;
  assign krnl_globalSort_L1_L2_16_in_dist2_peek_dout = out_dist_50__dout;
  assign krnl_globalSort_L1_L2_16_in_dist2_peek_empty_n = out_dist_50__empty_n;
  assign krnl_globalSort_L1_L2_16_in_dist2_s_dout = out_dist_50__dout;
  assign krnl_globalSort_L1_L2_16_in_dist2_s_empty_n = out_dist_50__empty_n;
  assign out_dist_50__read = krnl_globalSort_L1_L2_16_in_dist2_s_read;
  assign krnl_globalSort_L1_L2_16_in_id0_peek_dout = out_id_48__dout;
  assign krnl_globalSort_L1_L2_16_in_id0_peek_empty_n = out_id_48__empty_n;
  assign krnl_globalSort_L1_L2_16_in_id0_s_dout = out_id_48__dout;
  assign krnl_globalSort_L1_L2_16_in_id0_s_empty_n = out_id_48__empty_n;
  assign out_id_48__read = krnl_globalSort_L1_L2_16_in_id0_s_read;
  assign krnl_globalSort_L1_L2_16_in_id1_peek_dout = out_id_49__dout;
  assign krnl_globalSort_L1_L2_16_in_id1_peek_empty_n = out_id_49__empty_n;
  assign krnl_globalSort_L1_L2_16_in_id1_s_dout = out_id_49__dout;
  assign krnl_globalSort_L1_L2_16_in_id1_s_empty_n = out_id_49__empty_n;
  assign out_id_49__read = krnl_globalSort_L1_L2_16_in_id1_s_read;
  assign krnl_globalSort_L1_L2_16_in_id2_peek_dout = out_id_50__dout;
  assign krnl_globalSort_L1_L2_16_in_id2_peek_empty_n = out_id_50__empty_n;
  assign krnl_globalSort_L1_L2_16_in_id2_s_dout = out_id_50__dout;
  assign krnl_globalSort_L1_L2_16_in_id2_s_empty_n = out_id_50__empty_n;
  assign out_id_50__read = krnl_globalSort_L1_L2_16_in_id2_s_read;
  assign L1_out_dist_16__din = krnl_globalSort_L1_L2_16_out_dist_din;
  assign krnl_globalSort_L1_L2_16_out_dist_full_n = L1_out_dist_16__full_n;
  assign L1_out_dist_16__write = krnl_globalSort_L1_L2_16_out_dist_write;
  assign L1_out_id_16__din = krnl_globalSort_L1_L2_16_out_id_din;
  assign krnl_globalSort_L1_L2_16_out_id_full_n = L1_out_id_16__full_n;
  assign L1_out_id_16__write = krnl_globalSort_L1_L2_16_out_id_write;
  assign krnl_globalSort_L1_L2_17_ap_clk = ap_clk;
  assign krnl_globalSort_L1_L2_17__ap_done = krnl_globalSort_L1_L2_17_ap_done;
  assign krnl_globalSort_L1_L2_17__ap_idle = krnl_globalSort_L1_L2_17_ap_idle;
  assign krnl_globalSort_L1_L2_17__ap_ready = krnl_globalSort_L1_L2_17_ap_ready;
  assign krnl_globalSort_L1_L2_17_ap_rst_n = ap_rst_n;
  assign krnl_globalSort_L1_L2_17_ap_start = krnl_globalSort_L1_L2_17__ap_start;
  assign krnl_globalSort_L1_L2_17_in_dist0_peek_dout = out_dist_51__dout;
  assign krnl_globalSort_L1_L2_17_in_dist0_peek_empty_n = out_dist_51__empty_n;
  assign krnl_globalSort_L1_L2_17_in_dist0_s_dout = out_dist_51__dout;
  assign krnl_globalSort_L1_L2_17_in_dist0_s_empty_n = out_dist_51__empty_n;
  assign out_dist_51__read = krnl_globalSort_L1_L2_17_in_dist0_s_read;
  assign krnl_globalSort_L1_L2_17_in_dist1_peek_dout = out_dist_52__dout;
  assign krnl_globalSort_L1_L2_17_in_dist1_peek_empty_n = out_dist_52__empty_n;
  assign krnl_globalSort_L1_L2_17_in_dist1_s_dout = out_dist_52__dout;
  assign krnl_globalSort_L1_L2_17_in_dist1_s_empty_n = out_dist_52__empty_n;
  assign out_dist_52__read = krnl_globalSort_L1_L2_17_in_dist1_s_read;
  assign krnl_globalSort_L1_L2_17_in_dist2_peek_dout = out_dist_53__dout;
  assign krnl_globalSort_L1_L2_17_in_dist2_peek_empty_n = out_dist_53__empty_n;
  assign krnl_globalSort_L1_L2_17_in_dist2_s_dout = out_dist_53__dout;
  assign krnl_globalSort_L1_L2_17_in_dist2_s_empty_n = out_dist_53__empty_n;
  assign out_dist_53__read = krnl_globalSort_L1_L2_17_in_dist2_s_read;
  assign krnl_globalSort_L1_L2_17_in_id0_peek_dout = out_id_51__dout;
  assign krnl_globalSort_L1_L2_17_in_id0_peek_empty_n = out_id_51__empty_n;
  assign krnl_globalSort_L1_L2_17_in_id0_s_dout = out_id_51__dout;
  assign krnl_globalSort_L1_L2_17_in_id0_s_empty_n = out_id_51__empty_n;
  assign out_id_51__read = krnl_globalSort_L1_L2_17_in_id0_s_read;
  assign krnl_globalSort_L1_L2_17_in_id1_peek_dout = out_id_52__dout;
  assign krnl_globalSort_L1_L2_17_in_id1_peek_empty_n = out_id_52__empty_n;
  assign krnl_globalSort_L1_L2_17_in_id1_s_dout = out_id_52__dout;
  assign krnl_globalSort_L1_L2_17_in_id1_s_empty_n = out_id_52__empty_n;
  assign out_id_52__read = krnl_globalSort_L1_L2_17_in_id1_s_read;
  assign krnl_globalSort_L1_L2_17_in_id2_peek_dout = out_id_53__dout;
  assign krnl_globalSort_L1_L2_17_in_id2_peek_empty_n = out_id_53__empty_n;
  assign krnl_globalSort_L1_L2_17_in_id2_s_dout = out_id_53__dout;
  assign krnl_globalSort_L1_L2_17_in_id2_s_empty_n = out_id_53__empty_n;
  assign out_id_53__read = krnl_globalSort_L1_L2_17_in_id2_s_read;
  assign L1_out_dist_17__din = krnl_globalSort_L1_L2_17_out_dist_din;
  assign krnl_globalSort_L1_L2_17_out_dist_full_n = L1_out_dist_17__full_n;
  assign L1_out_dist_17__write = krnl_globalSort_L1_L2_17_out_dist_write;
  assign L1_out_id_17__din = krnl_globalSort_L1_L2_17_out_id_din;
  assign krnl_globalSort_L1_L2_17_out_id_full_n = L1_out_id_17__full_n;
  assign L1_out_id_17__write = krnl_globalSort_L1_L2_17_out_id_write;
  assign krnl_globalSort_L1_L2_18_ap_clk = ap_clk;
  assign krnl_globalSort_L1_L2_18__ap_done = krnl_globalSort_L1_L2_18_ap_done;
  assign krnl_globalSort_L1_L2_18__ap_idle = krnl_globalSort_L1_L2_18_ap_idle;
  assign krnl_globalSort_L1_L2_18__ap_ready = krnl_globalSort_L1_L2_18_ap_ready;
  assign krnl_globalSort_L1_L2_18_ap_rst_n = ap_rst_n;
  assign krnl_globalSort_L1_L2_18_ap_start = krnl_globalSort_L1_L2_18__ap_start;
  assign krnl_globalSort_L1_L2_18_in_dist0_peek_dout = L1_out_dist_0__dout;
  assign krnl_globalSort_L1_L2_18_in_dist0_peek_empty_n = L1_out_dist_0__empty_n;
  assign krnl_globalSort_L1_L2_18_in_dist0_s_dout = L1_out_dist_0__dout;
  assign krnl_globalSort_L1_L2_18_in_dist0_s_empty_n = L1_out_dist_0__empty_n;
  assign L1_out_dist_0__read = krnl_globalSort_L1_L2_18_in_dist0_s_read;
  assign krnl_globalSort_L1_L2_18_in_dist1_peek_dout = L1_out_dist_1__dout;
  assign krnl_globalSort_L1_L2_18_in_dist1_peek_empty_n = L1_out_dist_1__empty_n;
  assign krnl_globalSort_L1_L2_18_in_dist1_s_dout = L1_out_dist_1__dout;
  assign krnl_globalSort_L1_L2_18_in_dist1_s_empty_n = L1_out_dist_1__empty_n;
  assign L1_out_dist_1__read = krnl_globalSort_L1_L2_18_in_dist1_s_read;
  assign krnl_globalSort_L1_L2_18_in_dist2_peek_dout = L1_out_dist_2__dout;
  assign krnl_globalSort_L1_L2_18_in_dist2_peek_empty_n = L1_out_dist_2__empty_n;
  assign krnl_globalSort_L1_L2_18_in_dist2_s_dout = L1_out_dist_2__dout;
  assign krnl_globalSort_L1_L2_18_in_dist2_s_empty_n = L1_out_dist_2__empty_n;
  assign L1_out_dist_2__read = krnl_globalSort_L1_L2_18_in_dist2_s_read;
  assign krnl_globalSort_L1_L2_18_in_id0_peek_dout = L1_out_id_0__dout;
  assign krnl_globalSort_L1_L2_18_in_id0_peek_empty_n = L1_out_id_0__empty_n;
  assign krnl_globalSort_L1_L2_18_in_id0_s_dout = L1_out_id_0__dout;
  assign krnl_globalSort_L1_L2_18_in_id0_s_empty_n = L1_out_id_0__empty_n;
  assign L1_out_id_0__read = krnl_globalSort_L1_L2_18_in_id0_s_read;
  assign krnl_globalSort_L1_L2_18_in_id1_peek_dout = L1_out_id_1__dout;
  assign krnl_globalSort_L1_L2_18_in_id1_peek_empty_n = L1_out_id_1__empty_n;
  assign krnl_globalSort_L1_L2_18_in_id1_s_dout = L1_out_id_1__dout;
  assign krnl_globalSort_L1_L2_18_in_id1_s_empty_n = L1_out_id_1__empty_n;
  assign L1_out_id_1__read = krnl_globalSort_L1_L2_18_in_id1_s_read;
  assign krnl_globalSort_L1_L2_18_in_id2_peek_dout = L1_out_id_2__dout;
  assign krnl_globalSort_L1_L2_18_in_id2_peek_empty_n = L1_out_id_2__empty_n;
  assign krnl_globalSort_L1_L2_18_in_id2_s_dout = L1_out_id_2__dout;
  assign krnl_globalSort_L1_L2_18_in_id2_s_empty_n = L1_out_id_2__empty_n;
  assign L1_out_id_2__read = krnl_globalSort_L1_L2_18_in_id2_s_read;
  assign L2_out_dist0__din = krnl_globalSort_L1_L2_18_out_dist_din;
  assign krnl_globalSort_L1_L2_18_out_dist_full_n = L2_out_dist0__full_n;
  assign L2_out_dist0__write = krnl_globalSort_L1_L2_18_out_dist_write;
  assign L2_out_id0__din = krnl_globalSort_L1_L2_18_out_id_din;
  assign krnl_globalSort_L1_L2_18_out_id_full_n = L2_out_id0__full_n;
  assign L2_out_id0__write = krnl_globalSort_L1_L2_18_out_id_write;
  assign krnl_globalSort_L1_L2_19_ap_clk = ap_clk;
  assign krnl_globalSort_L1_L2_19__ap_done = krnl_globalSort_L1_L2_19_ap_done;
  assign krnl_globalSort_L1_L2_19__ap_idle = krnl_globalSort_L1_L2_19_ap_idle;
  assign krnl_globalSort_L1_L2_19__ap_ready = krnl_globalSort_L1_L2_19_ap_ready;
  assign krnl_globalSort_L1_L2_19_ap_rst_n = ap_rst_n;
  assign krnl_globalSort_L1_L2_19_ap_start = krnl_globalSort_L1_L2_19__ap_start;
  assign krnl_globalSort_L1_L2_19_in_dist0_peek_dout = L1_out_dist_3__dout;
  assign krnl_globalSort_L1_L2_19_in_dist0_peek_empty_n = L1_out_dist_3__empty_n;
  assign krnl_globalSort_L1_L2_19_in_dist0_s_dout = L1_out_dist_3__dout;
  assign krnl_globalSort_L1_L2_19_in_dist0_s_empty_n = L1_out_dist_3__empty_n;
  assign L1_out_dist_3__read = krnl_globalSort_L1_L2_19_in_dist0_s_read;
  assign krnl_globalSort_L1_L2_19_in_dist1_peek_dout = L1_out_dist_4__dout;
  assign krnl_globalSort_L1_L2_19_in_dist1_peek_empty_n = L1_out_dist_4__empty_n;
  assign krnl_globalSort_L1_L2_19_in_dist1_s_dout = L1_out_dist_4__dout;
  assign krnl_globalSort_L1_L2_19_in_dist1_s_empty_n = L1_out_dist_4__empty_n;
  assign L1_out_dist_4__read = krnl_globalSort_L1_L2_19_in_dist1_s_read;
  assign krnl_globalSort_L1_L2_19_in_dist2_peek_dout = L1_out_dist_5__dout;
  assign krnl_globalSort_L1_L2_19_in_dist2_peek_empty_n = L1_out_dist_5__empty_n;
  assign krnl_globalSort_L1_L2_19_in_dist2_s_dout = L1_out_dist_5__dout;
  assign krnl_globalSort_L1_L2_19_in_dist2_s_empty_n = L1_out_dist_5__empty_n;
  assign L1_out_dist_5__read = krnl_globalSort_L1_L2_19_in_dist2_s_read;
  assign krnl_globalSort_L1_L2_19_in_id0_peek_dout = L1_out_id_3__dout;
  assign krnl_globalSort_L1_L2_19_in_id0_peek_empty_n = L1_out_id_3__empty_n;
  assign krnl_globalSort_L1_L2_19_in_id0_s_dout = L1_out_id_3__dout;
  assign krnl_globalSort_L1_L2_19_in_id0_s_empty_n = L1_out_id_3__empty_n;
  assign L1_out_id_3__read = krnl_globalSort_L1_L2_19_in_id0_s_read;
  assign krnl_globalSort_L1_L2_19_in_id1_peek_dout = L1_out_id_4__dout;
  assign krnl_globalSort_L1_L2_19_in_id1_peek_empty_n = L1_out_id_4__empty_n;
  assign krnl_globalSort_L1_L2_19_in_id1_s_dout = L1_out_id_4__dout;
  assign krnl_globalSort_L1_L2_19_in_id1_s_empty_n = L1_out_id_4__empty_n;
  assign L1_out_id_4__read = krnl_globalSort_L1_L2_19_in_id1_s_read;
  assign krnl_globalSort_L1_L2_19_in_id2_peek_dout = L1_out_id_5__dout;
  assign krnl_globalSort_L1_L2_19_in_id2_peek_empty_n = L1_out_id_5__empty_n;
  assign krnl_globalSort_L1_L2_19_in_id2_s_dout = L1_out_id_5__dout;
  assign krnl_globalSort_L1_L2_19_in_id2_s_empty_n = L1_out_id_5__empty_n;
  assign L1_out_id_5__read = krnl_globalSort_L1_L2_19_in_id2_s_read;
  assign L2_out_dist1__din = krnl_globalSort_L1_L2_19_out_dist_din;
  assign krnl_globalSort_L1_L2_19_out_dist_full_n = L2_out_dist1__full_n;
  assign L2_out_dist1__write = krnl_globalSort_L1_L2_19_out_dist_write;
  assign L2_out_id1__din = krnl_globalSort_L1_L2_19_out_id_din;
  assign krnl_globalSort_L1_L2_19_out_id_full_n = L2_out_id1__full_n;
  assign L2_out_id1__write = krnl_globalSort_L1_L2_19_out_id_write;
  assign krnl_globalSort_L1_L2_20_ap_clk = ap_clk;
  assign krnl_globalSort_L1_L2_20__ap_done = krnl_globalSort_L1_L2_20_ap_done;
  assign krnl_globalSort_L1_L2_20__ap_idle = krnl_globalSort_L1_L2_20_ap_idle;
  assign krnl_globalSort_L1_L2_20__ap_ready = krnl_globalSort_L1_L2_20_ap_ready;
  assign krnl_globalSort_L1_L2_20_ap_rst_n = ap_rst_n;
  assign krnl_globalSort_L1_L2_20_ap_start = krnl_globalSort_L1_L2_20__ap_start;
  assign krnl_globalSort_L1_L2_20_in_dist0_peek_dout = L1_out_dist_6__dout;
  assign krnl_globalSort_L1_L2_20_in_dist0_peek_empty_n = L1_out_dist_6__empty_n;
  assign krnl_globalSort_L1_L2_20_in_dist0_s_dout = L1_out_dist_6__dout;
  assign krnl_globalSort_L1_L2_20_in_dist0_s_empty_n = L1_out_dist_6__empty_n;
  assign L1_out_dist_6__read = krnl_globalSort_L1_L2_20_in_dist0_s_read;
  assign krnl_globalSort_L1_L2_20_in_dist1_peek_dout = L1_out_dist_7__dout;
  assign krnl_globalSort_L1_L2_20_in_dist1_peek_empty_n = L1_out_dist_7__empty_n;
  assign krnl_globalSort_L1_L2_20_in_dist1_s_dout = L1_out_dist_7__dout;
  assign krnl_globalSort_L1_L2_20_in_dist1_s_empty_n = L1_out_dist_7__empty_n;
  assign L1_out_dist_7__read = krnl_globalSort_L1_L2_20_in_dist1_s_read;
  assign krnl_globalSort_L1_L2_20_in_dist2_peek_dout = L1_out_dist_8__dout;
  assign krnl_globalSort_L1_L2_20_in_dist2_peek_empty_n = L1_out_dist_8__empty_n;
  assign krnl_globalSort_L1_L2_20_in_dist2_s_dout = L1_out_dist_8__dout;
  assign krnl_globalSort_L1_L2_20_in_dist2_s_empty_n = L1_out_dist_8__empty_n;
  assign L1_out_dist_8__read = krnl_globalSort_L1_L2_20_in_dist2_s_read;
  assign krnl_globalSort_L1_L2_20_in_id0_peek_dout = L1_out_id_6__dout;
  assign krnl_globalSort_L1_L2_20_in_id0_peek_empty_n = L1_out_id_6__empty_n;
  assign krnl_globalSort_L1_L2_20_in_id0_s_dout = L1_out_id_6__dout;
  assign krnl_globalSort_L1_L2_20_in_id0_s_empty_n = L1_out_id_6__empty_n;
  assign L1_out_id_6__read = krnl_globalSort_L1_L2_20_in_id0_s_read;
  assign krnl_globalSort_L1_L2_20_in_id1_peek_dout = L1_out_id_7__dout;
  assign krnl_globalSort_L1_L2_20_in_id1_peek_empty_n = L1_out_id_7__empty_n;
  assign krnl_globalSort_L1_L2_20_in_id1_s_dout = L1_out_id_7__dout;
  assign krnl_globalSort_L1_L2_20_in_id1_s_empty_n = L1_out_id_7__empty_n;
  assign L1_out_id_7__read = krnl_globalSort_L1_L2_20_in_id1_s_read;
  assign krnl_globalSort_L1_L2_20_in_id2_peek_dout = L1_out_id_8__dout;
  assign krnl_globalSort_L1_L2_20_in_id2_peek_empty_n = L1_out_id_8__empty_n;
  assign krnl_globalSort_L1_L2_20_in_id2_s_dout = L1_out_id_8__dout;
  assign krnl_globalSort_L1_L2_20_in_id2_s_empty_n = L1_out_id_8__empty_n;
  assign L1_out_id_8__read = krnl_globalSort_L1_L2_20_in_id2_s_read;
  assign L2_out_dist2__din = krnl_globalSort_L1_L2_20_out_dist_din;
  assign krnl_globalSort_L1_L2_20_out_dist_full_n = L2_out_dist2__full_n;
  assign L2_out_dist2__write = krnl_globalSort_L1_L2_20_out_dist_write;
  assign L2_out_id2__din = krnl_globalSort_L1_L2_20_out_id_din;
  assign krnl_globalSort_L1_L2_20_out_id_full_n = L2_out_id2__full_n;
  assign L2_out_id2__write = krnl_globalSort_L1_L2_20_out_id_write;
  assign krnl_globalSort_L1_L2_21_ap_clk = ap_clk;
  assign krnl_globalSort_L1_L2_21__ap_done = krnl_globalSort_L1_L2_21_ap_done;
  assign krnl_globalSort_L1_L2_21__ap_idle = krnl_globalSort_L1_L2_21_ap_idle;
  assign krnl_globalSort_L1_L2_21__ap_ready = krnl_globalSort_L1_L2_21_ap_ready;
  assign krnl_globalSort_L1_L2_21_ap_rst_n = ap_rst_n;
  assign krnl_globalSort_L1_L2_21_ap_start = krnl_globalSort_L1_L2_21__ap_start;
  assign krnl_globalSort_L1_L2_21_in_dist0_peek_dout = L1_out_dist_9__dout;
  assign krnl_globalSort_L1_L2_21_in_dist0_peek_empty_n = L1_out_dist_9__empty_n;
  assign krnl_globalSort_L1_L2_21_in_dist0_s_dout = L1_out_dist_9__dout;
  assign krnl_globalSort_L1_L2_21_in_dist0_s_empty_n = L1_out_dist_9__empty_n;
  assign L1_out_dist_9__read = krnl_globalSort_L1_L2_21_in_dist0_s_read;
  assign krnl_globalSort_L1_L2_21_in_dist1_peek_dout = L1_out_dist_10__dout;
  assign krnl_globalSort_L1_L2_21_in_dist1_peek_empty_n = L1_out_dist_10__empty_n;
  assign krnl_globalSort_L1_L2_21_in_dist1_s_dout = L1_out_dist_10__dout;
  assign krnl_globalSort_L1_L2_21_in_dist1_s_empty_n = L1_out_dist_10__empty_n;
  assign L1_out_dist_10__read = krnl_globalSort_L1_L2_21_in_dist1_s_read;
  assign krnl_globalSort_L1_L2_21_in_dist2_peek_dout = L1_out_dist_11__dout;
  assign krnl_globalSort_L1_L2_21_in_dist2_peek_empty_n = L1_out_dist_11__empty_n;
  assign krnl_globalSort_L1_L2_21_in_dist2_s_dout = L1_out_dist_11__dout;
  assign krnl_globalSort_L1_L2_21_in_dist2_s_empty_n = L1_out_dist_11__empty_n;
  assign L1_out_dist_11__read = krnl_globalSort_L1_L2_21_in_dist2_s_read;
  assign krnl_globalSort_L1_L2_21_in_id0_peek_dout = L1_out_id_9__dout;
  assign krnl_globalSort_L1_L2_21_in_id0_peek_empty_n = L1_out_id_9__empty_n;
  assign krnl_globalSort_L1_L2_21_in_id0_s_dout = L1_out_id_9__dout;
  assign krnl_globalSort_L1_L2_21_in_id0_s_empty_n = L1_out_id_9__empty_n;
  assign L1_out_id_9__read = krnl_globalSort_L1_L2_21_in_id0_s_read;
  assign krnl_globalSort_L1_L2_21_in_id1_peek_dout = L1_out_id_10__dout;
  assign krnl_globalSort_L1_L2_21_in_id1_peek_empty_n = L1_out_id_10__empty_n;
  assign krnl_globalSort_L1_L2_21_in_id1_s_dout = L1_out_id_10__dout;
  assign krnl_globalSort_L1_L2_21_in_id1_s_empty_n = L1_out_id_10__empty_n;
  assign L1_out_id_10__read = krnl_globalSort_L1_L2_21_in_id1_s_read;
  assign krnl_globalSort_L1_L2_21_in_id2_peek_dout = L1_out_id_11__dout;
  assign krnl_globalSort_L1_L2_21_in_id2_peek_empty_n = L1_out_id_11__empty_n;
  assign krnl_globalSort_L1_L2_21_in_id2_s_dout = L1_out_id_11__dout;
  assign krnl_globalSort_L1_L2_21_in_id2_s_empty_n = L1_out_id_11__empty_n;
  assign L1_out_id_11__read = krnl_globalSort_L1_L2_21_in_id2_s_read;
  assign L2_out_dist3__din = krnl_globalSort_L1_L2_21_out_dist_din;
  assign krnl_globalSort_L1_L2_21_out_dist_full_n = L2_out_dist3__full_n;
  assign L2_out_dist3__write = krnl_globalSort_L1_L2_21_out_dist_write;
  assign L2_out_id3__din = krnl_globalSort_L1_L2_21_out_id_din;
  assign krnl_globalSort_L1_L2_21_out_id_full_n = L2_out_id3__full_n;
  assign L2_out_id3__write = krnl_globalSort_L1_L2_21_out_id_write;
  assign krnl_globalSort_L1_L2_22_ap_clk = ap_clk;
  assign krnl_globalSort_L1_L2_22__ap_done = krnl_globalSort_L1_L2_22_ap_done;
  assign krnl_globalSort_L1_L2_22__ap_idle = krnl_globalSort_L1_L2_22_ap_idle;
  assign krnl_globalSort_L1_L2_22__ap_ready = krnl_globalSort_L1_L2_22_ap_ready;
  assign krnl_globalSort_L1_L2_22_ap_rst_n = ap_rst_n;
  assign krnl_globalSort_L1_L2_22_ap_start = krnl_globalSort_L1_L2_22__ap_start;
  assign krnl_globalSort_L1_L2_22_in_dist0_peek_dout = L1_out_dist_12__dout;
  assign krnl_globalSort_L1_L2_22_in_dist0_peek_empty_n = L1_out_dist_12__empty_n;
  assign krnl_globalSort_L1_L2_22_in_dist0_s_dout = L1_out_dist_12__dout;
  assign krnl_globalSort_L1_L2_22_in_dist0_s_empty_n = L1_out_dist_12__empty_n;
  assign L1_out_dist_12__read = krnl_globalSort_L1_L2_22_in_dist0_s_read;
  assign krnl_globalSort_L1_L2_22_in_dist1_peek_dout = L1_out_dist_13__dout;
  assign krnl_globalSort_L1_L2_22_in_dist1_peek_empty_n = L1_out_dist_13__empty_n;
  assign krnl_globalSort_L1_L2_22_in_dist1_s_dout = L1_out_dist_13__dout;
  assign krnl_globalSort_L1_L2_22_in_dist1_s_empty_n = L1_out_dist_13__empty_n;
  assign L1_out_dist_13__read = krnl_globalSort_L1_L2_22_in_dist1_s_read;
  assign krnl_globalSort_L1_L2_22_in_dist2_peek_dout = L1_out_dist_14__dout;
  assign krnl_globalSort_L1_L2_22_in_dist2_peek_empty_n = L1_out_dist_14__empty_n;
  assign krnl_globalSort_L1_L2_22_in_dist2_s_dout = L1_out_dist_14__dout;
  assign krnl_globalSort_L1_L2_22_in_dist2_s_empty_n = L1_out_dist_14__empty_n;
  assign L1_out_dist_14__read = krnl_globalSort_L1_L2_22_in_dist2_s_read;
  assign krnl_globalSort_L1_L2_22_in_id0_peek_dout = L1_out_id_12__dout;
  assign krnl_globalSort_L1_L2_22_in_id0_peek_empty_n = L1_out_id_12__empty_n;
  assign krnl_globalSort_L1_L2_22_in_id0_s_dout = L1_out_id_12__dout;
  assign krnl_globalSort_L1_L2_22_in_id0_s_empty_n = L1_out_id_12__empty_n;
  assign L1_out_id_12__read = krnl_globalSort_L1_L2_22_in_id0_s_read;
  assign krnl_globalSort_L1_L2_22_in_id1_peek_dout = L1_out_id_13__dout;
  assign krnl_globalSort_L1_L2_22_in_id1_peek_empty_n = L1_out_id_13__empty_n;
  assign krnl_globalSort_L1_L2_22_in_id1_s_dout = L1_out_id_13__dout;
  assign krnl_globalSort_L1_L2_22_in_id1_s_empty_n = L1_out_id_13__empty_n;
  assign L1_out_id_13__read = krnl_globalSort_L1_L2_22_in_id1_s_read;
  assign krnl_globalSort_L1_L2_22_in_id2_peek_dout = L1_out_id_14__dout;
  assign krnl_globalSort_L1_L2_22_in_id2_peek_empty_n = L1_out_id_14__empty_n;
  assign krnl_globalSort_L1_L2_22_in_id2_s_dout = L1_out_id_14__dout;
  assign krnl_globalSort_L1_L2_22_in_id2_s_empty_n = L1_out_id_14__empty_n;
  assign L1_out_id_14__read = krnl_globalSort_L1_L2_22_in_id2_s_read;
  assign L2_out_dist4__din = krnl_globalSort_L1_L2_22_out_dist_din;
  assign krnl_globalSort_L1_L2_22_out_dist_full_n = L2_out_dist4__full_n;
  assign L2_out_dist4__write = krnl_globalSort_L1_L2_22_out_dist_write;
  assign L2_out_id4__din = krnl_globalSort_L1_L2_22_out_id_din;
  assign krnl_globalSort_L1_L2_22_out_id_full_n = L2_out_id4__full_n;
  assign L2_out_id4__write = krnl_globalSort_L1_L2_22_out_id_write;
  assign krnl_globalSort_L1_L2_23_ap_clk = ap_clk;
  assign krnl_globalSort_L1_L2_23__ap_done = krnl_globalSort_L1_L2_23_ap_done;
  assign krnl_globalSort_L1_L2_23__ap_idle = krnl_globalSort_L1_L2_23_ap_idle;
  assign krnl_globalSort_L1_L2_23__ap_ready = krnl_globalSort_L1_L2_23_ap_ready;
  assign krnl_globalSort_L1_L2_23_ap_rst_n = ap_rst_n;
  assign krnl_globalSort_L1_L2_23_ap_start = krnl_globalSort_L1_L2_23__ap_start;
  assign krnl_globalSort_L1_L2_23_in_dist0_peek_dout = L1_out_dist_15__dout;
  assign krnl_globalSort_L1_L2_23_in_dist0_peek_empty_n = L1_out_dist_15__empty_n;
  assign krnl_globalSort_L1_L2_23_in_dist0_s_dout = L1_out_dist_15__dout;
  assign krnl_globalSort_L1_L2_23_in_dist0_s_empty_n = L1_out_dist_15__empty_n;
  assign L1_out_dist_15__read = krnl_globalSort_L1_L2_23_in_dist0_s_read;
  assign krnl_globalSort_L1_L2_23_in_dist1_peek_dout = L1_out_dist_16__dout;
  assign krnl_globalSort_L1_L2_23_in_dist1_peek_empty_n = L1_out_dist_16__empty_n;
  assign krnl_globalSort_L1_L2_23_in_dist1_s_dout = L1_out_dist_16__dout;
  assign krnl_globalSort_L1_L2_23_in_dist1_s_empty_n = L1_out_dist_16__empty_n;
  assign L1_out_dist_16__read = krnl_globalSort_L1_L2_23_in_dist1_s_read;
  assign krnl_globalSort_L1_L2_23_in_dist2_peek_dout = L1_out_dist_17__dout;
  assign krnl_globalSort_L1_L2_23_in_dist2_peek_empty_n = L1_out_dist_17__empty_n;
  assign krnl_globalSort_L1_L2_23_in_dist2_s_dout = L1_out_dist_17__dout;
  assign krnl_globalSort_L1_L2_23_in_dist2_s_empty_n = L1_out_dist_17__empty_n;
  assign L1_out_dist_17__read = krnl_globalSort_L1_L2_23_in_dist2_s_read;
  assign krnl_globalSort_L1_L2_23_in_id0_peek_dout = L1_out_id_15__dout;
  assign krnl_globalSort_L1_L2_23_in_id0_peek_empty_n = L1_out_id_15__empty_n;
  assign krnl_globalSort_L1_L2_23_in_id0_s_dout = L1_out_id_15__dout;
  assign krnl_globalSort_L1_L2_23_in_id0_s_empty_n = L1_out_id_15__empty_n;
  assign L1_out_id_15__read = krnl_globalSort_L1_L2_23_in_id0_s_read;
  assign krnl_globalSort_L1_L2_23_in_id1_peek_dout = L1_out_id_16__dout;
  assign krnl_globalSort_L1_L2_23_in_id1_peek_empty_n = L1_out_id_16__empty_n;
  assign krnl_globalSort_L1_L2_23_in_id1_s_dout = L1_out_id_16__dout;
  assign krnl_globalSort_L1_L2_23_in_id1_s_empty_n = L1_out_id_16__empty_n;
  assign L1_out_id_16__read = krnl_globalSort_L1_L2_23_in_id1_s_read;
  assign krnl_globalSort_L1_L2_23_in_id2_peek_dout = L1_out_id_17__dout;
  assign krnl_globalSort_L1_L2_23_in_id2_peek_empty_n = L1_out_id_17__empty_n;
  assign krnl_globalSort_L1_L2_23_in_id2_s_dout = L1_out_id_17__dout;
  assign krnl_globalSort_L1_L2_23_in_id2_s_empty_n = L1_out_id_17__empty_n;
  assign L1_out_id_17__read = krnl_globalSort_L1_L2_23_in_id2_s_read;
  assign L2_out_dist5__din = krnl_globalSort_L1_L2_23_out_dist_din;
  assign krnl_globalSort_L1_L2_23_out_dist_full_n = L2_out_dist5__full_n;
  assign L2_out_dist5__write = krnl_globalSort_L1_L2_23_out_dist_write;
  assign L2_out_id5__din = krnl_globalSort_L1_L2_23_out_id_din;
  assign krnl_globalSort_L1_L2_23_out_id_full_n = L2_out_id5__full_n;
  assign L2_out_id5__write = krnl_globalSort_L1_L2_23_out_id_write;
  assign krnl_globalSort_L1_L2_24_ap_clk = ap_clk;
  assign krnl_globalSort_L1_L2_24__ap_done = krnl_globalSort_L1_L2_24_ap_done;
  assign krnl_globalSort_L1_L2_24__ap_idle = krnl_globalSort_L1_L2_24_ap_idle;
  assign krnl_globalSort_L1_L2_24__ap_ready = krnl_globalSort_L1_L2_24_ap_ready;
  assign krnl_globalSort_L1_L2_24_ap_rst_n = ap_rst_n;
  assign krnl_globalSort_L1_L2_24_ap_start = krnl_globalSort_L1_L2_24__ap_start;
  assign krnl_globalSort_L1_L2_24_in_dist0_peek_dout = L2_out_dist0__dout;
  assign krnl_globalSort_L1_L2_24_in_dist0_peek_empty_n = L2_out_dist0__empty_n;
  assign krnl_globalSort_L1_L2_24_in_dist0_s_dout = L2_out_dist0__dout;
  assign krnl_globalSort_L1_L2_24_in_dist0_s_empty_n = L2_out_dist0__empty_n;
  assign L2_out_dist0__read = krnl_globalSort_L1_L2_24_in_dist0_s_read;
  assign krnl_globalSort_L1_L2_24_in_dist1_peek_dout = L2_out_dist1__dout;
  assign krnl_globalSort_L1_L2_24_in_dist1_peek_empty_n = L2_out_dist1__empty_n;
  assign krnl_globalSort_L1_L2_24_in_dist1_s_dout = L2_out_dist1__dout;
  assign krnl_globalSort_L1_L2_24_in_dist1_s_empty_n = L2_out_dist1__empty_n;
  assign L2_out_dist1__read = krnl_globalSort_L1_L2_24_in_dist1_s_read;
  assign krnl_globalSort_L1_L2_24_in_dist2_peek_dout = L2_out_dist2__dout;
  assign krnl_globalSort_L1_L2_24_in_dist2_peek_empty_n = L2_out_dist2__empty_n;
  assign krnl_globalSort_L1_L2_24_in_dist2_s_dout = L2_out_dist2__dout;
  assign krnl_globalSort_L1_L2_24_in_dist2_s_empty_n = L2_out_dist2__empty_n;
  assign L2_out_dist2__read = krnl_globalSort_L1_L2_24_in_dist2_s_read;
  assign krnl_globalSort_L1_L2_24_in_id0_peek_dout = L2_out_id0__dout;
  assign krnl_globalSort_L1_L2_24_in_id0_peek_empty_n = L2_out_id0__empty_n;
  assign krnl_globalSort_L1_L2_24_in_id0_s_dout = L2_out_id0__dout;
  assign krnl_globalSort_L1_L2_24_in_id0_s_empty_n = L2_out_id0__empty_n;
  assign L2_out_id0__read = krnl_globalSort_L1_L2_24_in_id0_s_read;
  assign krnl_globalSort_L1_L2_24_in_id1_peek_dout = L2_out_id1__dout;
  assign krnl_globalSort_L1_L2_24_in_id1_peek_empty_n = L2_out_id1__empty_n;
  assign krnl_globalSort_L1_L2_24_in_id1_s_dout = L2_out_id1__dout;
  assign krnl_globalSort_L1_L2_24_in_id1_s_empty_n = L2_out_id1__empty_n;
  assign L2_out_id1__read = krnl_globalSort_L1_L2_24_in_id1_s_read;
  assign krnl_globalSort_L1_L2_24_in_id2_peek_dout = L2_out_id2__dout;
  assign krnl_globalSort_L1_L2_24_in_id2_peek_empty_n = L2_out_id2__empty_n;
  assign krnl_globalSort_L1_L2_24_in_id2_s_dout = L2_out_id2__dout;
  assign krnl_globalSort_L1_L2_24_in_id2_s_empty_n = L2_out_id2__empty_n;
  assign L2_out_id2__read = krnl_globalSort_L1_L2_24_in_id2_s_read;
  assign L3_out_dist0__din = krnl_globalSort_L1_L2_24_out_dist_din;
  assign krnl_globalSort_L1_L2_24_out_dist_full_n = L3_out_dist0__full_n;
  assign L3_out_dist0__write = krnl_globalSort_L1_L2_24_out_dist_write;
  assign L3_out_id0__din = krnl_globalSort_L1_L2_24_out_id_din;
  assign krnl_globalSort_L1_L2_24_out_id_full_n = L3_out_id0__full_n;
  assign L3_out_id0__write = krnl_globalSort_L1_L2_24_out_id_write;
  assign krnl_globalSort_L1_L2_25_ap_clk = ap_clk;
  assign krnl_globalSort_L1_L2_25__ap_done = krnl_globalSort_L1_L2_25_ap_done;
  assign krnl_globalSort_L1_L2_25__ap_idle = krnl_globalSort_L1_L2_25_ap_idle;
  assign krnl_globalSort_L1_L2_25__ap_ready = krnl_globalSort_L1_L2_25_ap_ready;
  assign krnl_globalSort_L1_L2_25_ap_rst_n = ap_rst_n;
  assign krnl_globalSort_L1_L2_25_ap_start = krnl_globalSort_L1_L2_25__ap_start;
  assign krnl_globalSort_L1_L2_25_in_dist0_peek_dout = L2_out_dist3__dout;
  assign krnl_globalSort_L1_L2_25_in_dist0_peek_empty_n = L2_out_dist3__empty_n;
  assign krnl_globalSort_L1_L2_25_in_dist0_s_dout = L2_out_dist3__dout;
  assign krnl_globalSort_L1_L2_25_in_dist0_s_empty_n = L2_out_dist3__empty_n;
  assign L2_out_dist3__read = krnl_globalSort_L1_L2_25_in_dist0_s_read;
  assign krnl_globalSort_L1_L2_25_in_dist1_peek_dout = L2_out_dist4__dout;
  assign krnl_globalSort_L1_L2_25_in_dist1_peek_empty_n = L2_out_dist4__empty_n;
  assign krnl_globalSort_L1_L2_25_in_dist1_s_dout = L2_out_dist4__dout;
  assign krnl_globalSort_L1_L2_25_in_dist1_s_empty_n = L2_out_dist4__empty_n;
  assign L2_out_dist4__read = krnl_globalSort_L1_L2_25_in_dist1_s_read;
  assign krnl_globalSort_L1_L2_25_in_dist2_peek_dout = L2_out_dist5__dout;
  assign krnl_globalSort_L1_L2_25_in_dist2_peek_empty_n = L2_out_dist5__empty_n;
  assign krnl_globalSort_L1_L2_25_in_dist2_s_dout = L2_out_dist5__dout;
  assign krnl_globalSort_L1_L2_25_in_dist2_s_empty_n = L2_out_dist5__empty_n;
  assign L2_out_dist5__read = krnl_globalSort_L1_L2_25_in_dist2_s_read;
  assign krnl_globalSort_L1_L2_25_in_id0_peek_dout = L2_out_id3__dout;
  assign krnl_globalSort_L1_L2_25_in_id0_peek_empty_n = L2_out_id3__empty_n;
  assign krnl_globalSort_L1_L2_25_in_id0_s_dout = L2_out_id3__dout;
  assign krnl_globalSort_L1_L2_25_in_id0_s_empty_n = L2_out_id3__empty_n;
  assign L2_out_id3__read = krnl_globalSort_L1_L2_25_in_id0_s_read;
  assign krnl_globalSort_L1_L2_25_in_id1_peek_dout = L2_out_id4__dout;
  assign krnl_globalSort_L1_L2_25_in_id1_peek_empty_n = L2_out_id4__empty_n;
  assign krnl_globalSort_L1_L2_25_in_id1_s_dout = L2_out_id4__dout;
  assign krnl_globalSort_L1_L2_25_in_id1_s_empty_n = L2_out_id4__empty_n;
  assign L2_out_id4__read = krnl_globalSort_L1_L2_25_in_id1_s_read;
  assign krnl_globalSort_L1_L2_25_in_id2_peek_dout = L2_out_id5__dout;
  assign krnl_globalSort_L1_L2_25_in_id2_peek_empty_n = L2_out_id5__empty_n;
  assign krnl_globalSort_L1_L2_25_in_id2_s_dout = L2_out_id5__dout;
  assign krnl_globalSort_L1_L2_25_in_id2_s_empty_n = L2_out_id5__empty_n;
  assign L2_out_id5__read = krnl_globalSort_L1_L2_25_in_id2_s_read;
  assign L3_out_dist1__din = krnl_globalSort_L1_L2_25_out_dist_din;
  assign krnl_globalSort_L1_L2_25_out_dist_full_n = L3_out_dist1__full_n;
  assign L3_out_dist1__write = krnl_globalSort_L1_L2_25_out_dist_write;
  assign L3_out_id1__din = krnl_globalSort_L1_L2_25_out_id_din;
  assign krnl_globalSort_L1_L2_25_out_id_full_n = L3_out_id1__full_n;
  assign L3_out_id1__write = krnl_globalSort_L1_L2_25_out_id_write;
  assign krnl_globalSort_L3_0_ap_clk = ap_clk;
  assign krnl_globalSort_L3_0__ap_done = krnl_globalSort_L3_0_ap_done;
  assign krnl_globalSort_L3_0__ap_idle = krnl_globalSort_L3_0_ap_idle;
  assign krnl_globalSort_L3_0__ap_ready = krnl_globalSort_L3_0_ap_ready;
  assign krnl_globalSort_L3_0_ap_rst_n = ap_rst_n;
  assign krnl_globalSort_L3_0_ap_start = krnl_globalSort_L3_0__ap_start;
  assign krnl_globalSort_L3_0_in_dist0_peek_dout = L3_out_dist0__dout;
  assign krnl_globalSort_L3_0_in_dist0_peek_empty_n = L3_out_dist0__empty_n;
  assign krnl_globalSort_L3_0_in_dist0_s_dout = L3_out_dist0__dout;
  assign krnl_globalSort_L3_0_in_dist0_s_empty_n = L3_out_dist0__empty_n;
  assign L3_out_dist0__read = krnl_globalSort_L3_0_in_dist0_s_read;
  assign krnl_globalSort_L3_0_in_dist1_peek_dout = L3_out_dist1__dout;
  assign krnl_globalSort_L3_0_in_dist1_peek_empty_n = L3_out_dist1__empty_n;
  assign krnl_globalSort_L3_0_in_dist1_s_dout = L3_out_dist1__dout;
  assign krnl_globalSort_L3_0_in_dist1_s_empty_n = L3_out_dist1__empty_n;
  assign L3_out_dist1__read = krnl_globalSort_L3_0_in_dist1_s_read;
  assign krnl_globalSort_L3_0_in_id0_peek_dout = L3_out_id0__dout;
  assign krnl_globalSort_L3_0_in_id0_peek_empty_n = L3_out_id0__empty_n;
  assign krnl_globalSort_L3_0_in_id0_s_dout = L3_out_id0__dout;
  assign krnl_globalSort_L3_0_in_id0_s_empty_n = L3_out_id0__empty_n;
  assign L3_out_id0__read = krnl_globalSort_L3_0_in_id0_s_read;
  assign krnl_globalSort_L3_0_in_id1_peek_dout = L3_out_id1__dout;
  assign krnl_globalSort_L3_0_in_id1_peek_empty_n = L3_out_id1__empty_n;
  assign krnl_globalSort_L3_0_in_id1_s_dout = L3_out_id1__dout;
  assign krnl_globalSort_L3_0_in_id1_s_empty_n = L3_out_id1__empty_n;
  assign L3_out_id1__read = krnl_globalSort_L3_0_in_id1_s_read;
  assign krnl_globalSort_L3_0_output_knnDist_read_addr_offset = krnl_globalSort_L3_0___L4_out_dist__q0;
  assign L4_out_dist_read_addr__din = krnl_globalSort_L3_0_output_knnDist_read_addr_s_din;
  assign krnl_globalSort_L3_0_output_knnDist_read_addr_s_full_n = L4_out_dist_read_addr__full_n;
  assign L4_out_dist_read_addr__write = krnl_globalSort_L3_0_output_knnDist_read_addr_s_write;
  assign krnl_globalSort_L3_0_output_knnDist_read_data_peek_dout = { 1'b0 , L4_out_dist_read_data__dout };
  assign krnl_globalSort_L3_0_output_knnDist_read_data_peek_empty_n = L4_out_dist_read_data__empty_n;
  assign krnl_globalSort_L3_0_output_knnDist_read_data_s_dout = { 1'b0 , L4_out_dist_read_data__dout };
  assign krnl_globalSort_L3_0_output_knnDist_read_data_s_empty_n = L4_out_dist_read_data__empty_n;
  assign L4_out_dist_read_data__read = krnl_globalSort_L3_0_output_knnDist_read_data_s_read;
  assign krnl_globalSort_L3_0_output_knnDist_write_addr_offset = krnl_globalSort_L3_0___L4_out_dist__q0;
  assign L4_out_dist_write_addr__din = krnl_globalSort_L3_0_output_knnDist_write_addr_s_din;
  assign krnl_globalSort_L3_0_output_knnDist_write_addr_s_full_n = L4_out_dist_write_addr__full_n;
  assign L4_out_dist_write_addr__write = krnl_globalSort_L3_0_output_knnDist_write_addr_s_write;
  assign L4_out_dist_write_data__din = krnl_globalSort_L3_0_output_knnDist_write_data_din;
  assign krnl_globalSort_L3_0_output_knnDist_write_data_full_n = L4_out_dist_write_data__full_n;
  assign L4_out_dist_write_data__write = krnl_globalSort_L3_0_output_knnDist_write_data_write;
  assign krnl_globalSort_L3_0_output_knnDist_write_resp_peek_dout = { 1'b0 , L4_out_dist_write_resp__dout };
  assign krnl_globalSort_L3_0_output_knnDist_write_resp_peek_empty_n = L4_out_dist_write_resp__empty_n;
  assign krnl_globalSort_L3_0_output_knnDist_write_resp_s_dout = { 1'b0 , L4_out_dist_write_resp__dout };
  assign krnl_globalSort_L3_0_output_knnDist_write_resp_s_empty_n = L4_out_dist_write_resp__empty_n;
  assign L4_out_dist_write_resp__read = krnl_globalSort_L3_0_output_knnDist_write_resp_s_read;
  assign krnl_globalSort_L3_0_output_knnId_read_addr_offset = krnl_globalSort_L3_0___L4_out_id__q0;
  assign L4_out_id_read_addr__din = krnl_globalSort_L3_0_output_knnId_read_addr_s_din;
  assign krnl_globalSort_L3_0_output_knnId_read_addr_s_full_n = L4_out_id_read_addr__full_n;
  assign L4_out_id_read_addr__write = krnl_globalSort_L3_0_output_knnId_read_addr_s_write;
  assign krnl_globalSort_L3_0_output_knnId_read_data_peek_dout = { 1'b0 , L4_out_id_read_data__dout };
  assign krnl_globalSort_L3_0_output_knnId_read_data_peek_empty_n = L4_out_id_read_data__empty_n;
  assign krnl_globalSort_L3_0_output_knnId_read_data_s_dout = { 1'b0 , L4_out_id_read_data__dout };
  assign krnl_globalSort_L3_0_output_knnId_read_data_s_empty_n = L4_out_id_read_data__empty_n;
  assign L4_out_id_read_data__read = krnl_globalSort_L3_0_output_knnId_read_data_s_read;
  assign krnl_globalSort_L3_0_output_knnId_write_addr_offset = krnl_globalSort_L3_0___L4_out_id__q0;
  assign L4_out_id_write_addr__din = krnl_globalSort_L3_0_output_knnId_write_addr_s_din;
  assign krnl_globalSort_L3_0_output_knnId_write_addr_s_full_n = L4_out_id_write_addr__full_n;
  assign L4_out_id_write_addr__write = krnl_globalSort_L3_0_output_knnId_write_addr_s_write;
  assign L4_out_id_write_data__din = krnl_globalSort_L3_0_output_knnId_write_data_din;
  assign krnl_globalSort_L3_0_output_knnId_write_data_full_n = L4_out_id_write_data__full_n;
  assign L4_out_id_write_data__write = krnl_globalSort_L3_0_output_knnId_write_data_write;
  assign krnl_globalSort_L3_0_output_knnId_write_resp_peek_dout = { 1'b0 , L4_out_id_write_resp__dout };
  assign krnl_globalSort_L3_0_output_knnId_write_resp_peek_empty_n = L4_out_id_write_resp__empty_n;
  assign krnl_globalSort_L3_0_output_knnId_write_resp_s_dout = { 1'b0 , L4_out_id_write_resp__dout };
  assign krnl_globalSort_L3_0_output_knnId_write_resp_s_empty_n = L4_out_id_write_resp__empty_n;
  assign L4_out_id_write_resp__read = krnl_globalSort_L3_0_output_knnId_write_resp_s_read;
  assign krnl_partialKnn_wrapper_0_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_0_0__ap_done = krnl_partialKnn_wrapper_0_0_ap_done;
  assign krnl_partialKnn_wrapper_0_0__ap_idle = krnl_partialKnn_wrapper_0_0_ap_idle;
  assign krnl_partialKnn_wrapper_0_0__ap_ready = krnl_partialKnn_wrapper_0_0_ap_ready;
  assign krnl_partialKnn_wrapper_0_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_0_0_ap_start = krnl_partialKnn_wrapper_0_0__ap_start;
  assign out_dist_0__din = krnl_partialKnn_wrapper_0_0_out_dist_din;
  assign krnl_partialKnn_wrapper_0_0_out_dist_full_n = out_dist_0__full_n;
  assign out_dist_0__write = krnl_partialKnn_wrapper_0_0_out_dist_write;
  assign out_id_0__din = krnl_partialKnn_wrapper_0_0_out_id_din;
  assign krnl_partialKnn_wrapper_0_0_out_id_full_n = out_id_0__full_n;
  assign out_id_0__write = krnl_partialKnn_wrapper_0_0_out_id_write;
  assign krnl_partialKnn_wrapper_0_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_0_0___in_0__q0;
  assign in_0_read_addr__din = krnl_partialKnn_wrapper_0_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_0_0_searchSpace_0_read_addr_s_full_n = in_0_read_addr__full_n;
  assign in_0_read_addr__write = krnl_partialKnn_wrapper_0_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_0_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_0_read_data__dout };
  assign krnl_partialKnn_wrapper_0_0_searchSpace_0_read_data_peek_empty_n = in_0_read_data__empty_n;
  assign krnl_partialKnn_wrapper_0_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_0_read_data__dout };
  assign krnl_partialKnn_wrapper_0_0_searchSpace_0_read_data_s_empty_n = in_0_read_data__empty_n;
  assign in_0_read_data__read = krnl_partialKnn_wrapper_0_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_0_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_0_0___in_0__q0;
  assign in_0_write_addr__din = krnl_partialKnn_wrapper_0_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_0_0_searchSpace_0_write_addr_s_full_n = in_0_write_addr__full_n;
  assign in_0_write_addr__write = krnl_partialKnn_wrapper_0_0_searchSpace_0_write_addr_s_write;
  assign in_0_write_data__din = krnl_partialKnn_wrapper_0_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_0_0_searchSpace_0_write_data_full_n = in_0_write_data__full_n;
  assign in_0_write_data__write = krnl_partialKnn_wrapper_0_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_0_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_0_write_resp__dout };
  assign krnl_partialKnn_wrapper_0_0_searchSpace_write_resp_peek_empty_n = in_0_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_0_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_0_write_resp__dout };
  assign krnl_partialKnn_wrapper_0_0_searchSpace_0_write_resp_s_empty_n = in_0_write_resp__empty_n;
  assign in_0_write_resp__read = krnl_partialKnn_wrapper_0_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_0_0_start_id_0 = 64'd0;
  assign krnl_partialKnn_wrapper_1_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_1_0__ap_done = krnl_partialKnn_wrapper_1_0_ap_done;
  assign krnl_partialKnn_wrapper_1_0__ap_idle = krnl_partialKnn_wrapper_1_0_ap_idle;
  assign krnl_partialKnn_wrapper_1_0__ap_ready = krnl_partialKnn_wrapper_1_0_ap_ready;
  assign krnl_partialKnn_wrapper_1_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_1_0_ap_start = krnl_partialKnn_wrapper_1_0__ap_start;
  assign out_dist_1__din = krnl_partialKnn_wrapper_1_0_out_dist_din;
  assign krnl_partialKnn_wrapper_1_0_out_dist_full_n = out_dist_1__full_n;
  assign out_dist_1__write = krnl_partialKnn_wrapper_1_0_out_dist_write;
  assign out_id_1__din = krnl_partialKnn_wrapper_1_0_out_id_din;
  assign krnl_partialKnn_wrapper_1_0_out_id_full_n = out_id_1__full_n;
  assign out_id_1__write = krnl_partialKnn_wrapper_1_0_out_id_write;
  assign krnl_partialKnn_wrapper_1_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_1_0___in_1__q0;
  assign in_1_read_addr__din = krnl_partialKnn_wrapper_1_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_1_0_searchSpace_0_read_addr_s_full_n = in_1_read_addr__full_n;
  assign in_1_read_addr__write = krnl_partialKnn_wrapper_1_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_1_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_1_read_data__dout };
  assign krnl_partialKnn_wrapper_1_0_searchSpace_0_read_data_peek_empty_n = in_1_read_data__empty_n;
  assign krnl_partialKnn_wrapper_1_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_1_read_data__dout };
  assign krnl_partialKnn_wrapper_1_0_searchSpace_0_read_data_s_empty_n = in_1_read_data__empty_n;
  assign in_1_read_data__read = krnl_partialKnn_wrapper_1_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_1_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_1_0___in_1__q0;
  assign in_1_write_addr__din = krnl_partialKnn_wrapper_1_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_1_0_searchSpace_0_write_addr_s_full_n = in_1_write_addr__full_n;
  assign in_1_write_addr__write = krnl_partialKnn_wrapper_1_0_searchSpace_0_write_addr_s_write;
  assign in_1_write_data__din = krnl_partialKnn_wrapper_1_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_1_0_searchSpace_0_write_data_full_n = in_1_write_data__full_n;
  assign in_1_write_data__write = krnl_partialKnn_wrapper_1_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_1_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_1_write_resp__dout };
  assign krnl_partialKnn_wrapper_1_0_searchSpace_write_resp_peek_empty_n = in_1_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_1_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_1_write_resp__dout };
  assign krnl_partialKnn_wrapper_1_0_searchSpace_0_write_resp_s_empty_n = in_1_write_resp__empty_n;
  assign in_1_write_resp__read = krnl_partialKnn_wrapper_1_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_1_0_start_id_0 = 64'd8192;
  assign krnl_partialKnn_wrapper_10_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_10_0__ap_done = krnl_partialKnn_wrapper_10_0_ap_done;
  assign krnl_partialKnn_wrapper_10_0__ap_idle = krnl_partialKnn_wrapper_10_0_ap_idle;
  assign krnl_partialKnn_wrapper_10_0__ap_ready = krnl_partialKnn_wrapper_10_0_ap_ready;
  assign krnl_partialKnn_wrapper_10_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_10_0_ap_start = krnl_partialKnn_wrapper_10_0__ap_start;
  assign out_dist_10__din = krnl_partialKnn_wrapper_10_0_out_dist_din;
  assign krnl_partialKnn_wrapper_10_0_out_dist_full_n = out_dist_10__full_n;
  assign out_dist_10__write = krnl_partialKnn_wrapper_10_0_out_dist_write;
  assign out_id_10__din = krnl_partialKnn_wrapper_10_0_out_id_din;
  assign krnl_partialKnn_wrapper_10_0_out_id_full_n = out_id_10__full_n;
  assign out_id_10__write = krnl_partialKnn_wrapper_10_0_out_id_write;
  assign krnl_partialKnn_wrapper_10_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_10_0___in_10__q0;
  assign in_10_read_addr__din = krnl_partialKnn_wrapper_10_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_10_0_searchSpace_0_read_addr_s_full_n = in_10_read_addr__full_n;
  assign in_10_read_addr__write = krnl_partialKnn_wrapper_10_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_10_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_10_read_data__dout };
  assign krnl_partialKnn_wrapper_10_0_searchSpace_read_data_peek_empty_n = in_10_read_data__empty_n;
  assign krnl_partialKnn_wrapper_10_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_10_read_data__dout };
  assign krnl_partialKnn_wrapper_10_0_searchSpace_0_read_data_s_empty_n = in_10_read_data__empty_n;
  assign in_10_read_data__read = krnl_partialKnn_wrapper_10_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_10_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_10_0___in_10__q0;
  assign in_10_write_addr__din = krnl_partialKnn_wrapper_10_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_10_0_searchSpace_0_write_addr_s_full_n = in_10_write_addr__full_n;
  assign in_10_write_addr__write = krnl_partialKnn_wrapper_10_0_searchSpace_0_write_addr_s_write;
  assign in_10_write_data__din = krnl_partialKnn_wrapper_10_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_10_0_searchSpace_0_write_data_full_n = in_10_write_data__full_n;
  assign in_10_write_data__write = krnl_partialKnn_wrapper_10_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_10_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_10_write_resp__dout };
  assign krnl_partialKnn_wrapper_10_0_searchSpace_write_resp_peek_empty_n = in_10_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_10_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_10_write_resp__dout };
  assign krnl_partialKnn_wrapper_10_0_searchSpace_0_write_resp_s_empty_n = in_10_write_resp__empty_n;
  assign in_10_write_resp__read = krnl_partialKnn_wrapper_10_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_10_0_start_id_0 = 64'd81920;
  assign krnl_partialKnn_wrapper_11_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_11_0__ap_done = krnl_partialKnn_wrapper_11_0_ap_done;
  assign krnl_partialKnn_wrapper_11_0__ap_idle = krnl_partialKnn_wrapper_11_0_ap_idle;
  assign krnl_partialKnn_wrapper_11_0__ap_ready = krnl_partialKnn_wrapper_11_0_ap_ready;
  assign krnl_partialKnn_wrapper_11_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_11_0_ap_start = krnl_partialKnn_wrapper_11_0__ap_start;
  assign out_dist_11__din = krnl_partialKnn_wrapper_11_0_out_dist_din;
  assign krnl_partialKnn_wrapper_11_0_out_dist_full_n = out_dist_11__full_n;
  assign out_dist_11__write = krnl_partialKnn_wrapper_11_0_out_dist_write;
  assign out_id_11__din = krnl_partialKnn_wrapper_11_0_out_id_din;
  assign krnl_partialKnn_wrapper_11_0_out_id_full_n = out_id_11__full_n;
  assign out_id_11__write = krnl_partialKnn_wrapper_11_0_out_id_write;
  assign krnl_partialKnn_wrapper_11_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_11_0___in_11__q0;
  assign in_11_read_addr__din = krnl_partialKnn_wrapper_11_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_11_0_searchSpace_0_read_addr_s_full_n = in_11_read_addr__full_n;
  assign in_11_read_addr__write = krnl_partialKnn_wrapper_11_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_11_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_11_read_data__dout };
  assign krnl_partialKnn_wrapper_11_0_searchSpace_read_data_peek_empty_n = in_11_read_data__empty_n;
  assign krnl_partialKnn_wrapper_11_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_11_read_data__dout };
  assign krnl_partialKnn_wrapper_11_0_searchSpace_0_read_data_s_empty_n = in_11_read_data__empty_n;
  assign in_11_read_data__read = krnl_partialKnn_wrapper_11_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_11_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_11_0___in_11__q0;
  assign in_11_write_addr__din = krnl_partialKnn_wrapper_11_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_11_0_searchSpace_0_write_addr_s_full_n = in_11_write_addr__full_n;
  assign in_11_write_addr__write = krnl_partialKnn_wrapper_11_0_searchSpace_0_write_addr_s_write;
  assign in_11_write_data__din = krnl_partialKnn_wrapper_11_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_11_0_searchSpace_0_write_data_full_n = in_11_write_data__full_n;
  assign in_11_write_data__write = krnl_partialKnn_wrapper_11_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_11_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_11_write_resp__dout };
  assign krnl_partialKnn_wrapper_11_0_searchSpace_write_resp_peek_empty_n = in_11_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_11_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_11_write_resp__dout };
  assign krnl_partialKnn_wrapper_11_0_searchSpace_0_write_resp_s_empty_n = in_11_write_resp__empty_n;
  assign in_11_write_resp__read = krnl_partialKnn_wrapper_11_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_11_0_start_id_0 = 64'd90112;
  assign krnl_partialKnn_wrapper_12_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_12_0__ap_done = krnl_partialKnn_wrapper_12_0_ap_done;
  assign krnl_partialKnn_wrapper_12_0__ap_idle = krnl_partialKnn_wrapper_12_0_ap_idle;
  assign krnl_partialKnn_wrapper_12_0__ap_ready = krnl_partialKnn_wrapper_12_0_ap_ready;
  assign krnl_partialKnn_wrapper_12_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_12_0_ap_start = krnl_partialKnn_wrapper_12_0__ap_start;
  assign out_dist_12__din = krnl_partialKnn_wrapper_12_0_out_dist_din;
  assign krnl_partialKnn_wrapper_12_0_out_dist_full_n = out_dist_12__full_n;
  assign out_dist_12__write = krnl_partialKnn_wrapper_12_0_out_dist_write;
  assign out_id_12__din = krnl_partialKnn_wrapper_12_0_out_id_din;
  assign krnl_partialKnn_wrapper_12_0_out_id_full_n = out_id_12__full_n;
  assign out_id_12__write = krnl_partialKnn_wrapper_12_0_out_id_write;
  assign krnl_partialKnn_wrapper_12_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_12_0___in_12__q0;
  assign in_12_read_addr__din = krnl_partialKnn_wrapper_12_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_12_0_searchSpace_0_read_addr_s_full_n = in_12_read_addr__full_n;
  assign in_12_read_addr__write = krnl_partialKnn_wrapper_12_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_12_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_12_read_data__dout };
  assign krnl_partialKnn_wrapper_12_0_searchSpace_read_data_peek_empty_n = in_12_read_data__empty_n;
  assign krnl_partialKnn_wrapper_12_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_12_read_data__dout };
  assign krnl_partialKnn_wrapper_12_0_searchSpace_0_read_data_s_empty_n = in_12_read_data__empty_n;
  assign in_12_read_data__read = krnl_partialKnn_wrapper_12_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_12_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_12_0___in_12__q0;
  assign in_12_write_addr__din = krnl_partialKnn_wrapper_12_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_12_0_searchSpace_0_write_addr_s_full_n = in_12_write_addr__full_n;
  assign in_12_write_addr__write = krnl_partialKnn_wrapper_12_0_searchSpace_0_write_addr_s_write;
  assign in_12_write_data__din = krnl_partialKnn_wrapper_12_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_12_0_searchSpace_0_write_data_full_n = in_12_write_data__full_n;
  assign in_12_write_data__write = krnl_partialKnn_wrapper_12_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_12_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_12_write_resp__dout };
  assign krnl_partialKnn_wrapper_12_0_searchSpace_write_resp_peek_empty_n = in_12_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_12_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_12_write_resp__dout };
  assign krnl_partialKnn_wrapper_12_0_searchSpace_0_write_resp_s_empty_n = in_12_write_resp__empty_n;
  assign in_12_write_resp__read = krnl_partialKnn_wrapper_12_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_12_0_start_id_0 = 64'd98304;
  assign krnl_partialKnn_wrapper_13_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_13_0__ap_done = krnl_partialKnn_wrapper_13_0_ap_done;
  assign krnl_partialKnn_wrapper_13_0__ap_idle = krnl_partialKnn_wrapper_13_0_ap_idle;
  assign krnl_partialKnn_wrapper_13_0__ap_ready = krnl_partialKnn_wrapper_13_0_ap_ready;
  assign krnl_partialKnn_wrapper_13_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_13_0_ap_start = krnl_partialKnn_wrapper_13_0__ap_start;
  assign out_dist_13__din = krnl_partialKnn_wrapper_13_0_out_dist_din;
  assign krnl_partialKnn_wrapper_13_0_out_dist_full_n = out_dist_13__full_n;
  assign out_dist_13__write = krnl_partialKnn_wrapper_13_0_out_dist_write;
  assign out_id_13__din = krnl_partialKnn_wrapper_13_0_out_id_din;
  assign krnl_partialKnn_wrapper_13_0_out_id_full_n = out_id_13__full_n;
  assign out_id_13__write = krnl_partialKnn_wrapper_13_0_out_id_write;
  assign krnl_partialKnn_wrapper_13_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_13_0___in_13__q0;
  assign in_13_read_addr__din = krnl_partialKnn_wrapper_13_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_13_0_searchSpace_0_read_addr_s_full_n = in_13_read_addr__full_n;
  assign in_13_read_addr__write = krnl_partialKnn_wrapper_13_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_13_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_13_read_data__dout };
  assign krnl_partialKnn_wrapper_13_0_searchSpace_read_data_peek_empty_n = in_13_read_data__empty_n;
  assign krnl_partialKnn_wrapper_13_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_13_read_data__dout };
  assign krnl_partialKnn_wrapper_13_0_searchSpace_0_read_data_s_empty_n = in_13_read_data__empty_n;
  assign in_13_read_data__read = krnl_partialKnn_wrapper_13_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_13_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_13_0___in_13__q0;
  assign in_13_write_addr__din = krnl_partialKnn_wrapper_13_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_13_0_searchSpace_0_write_addr_s_full_n = in_13_write_addr__full_n;
  assign in_13_write_addr__write = krnl_partialKnn_wrapper_13_0_searchSpace_0_write_addr_s_write;
  assign in_13_write_data__din = krnl_partialKnn_wrapper_13_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_13_0_searchSpace_0_write_data_full_n = in_13_write_data__full_n;
  assign in_13_write_data__write = krnl_partialKnn_wrapper_13_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_13_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_13_write_resp__dout };
  assign krnl_partialKnn_wrapper_13_0_searchSpace_write_resp_peek_empty_n = in_13_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_13_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_13_write_resp__dout };
  assign krnl_partialKnn_wrapper_13_0_searchSpace_0_write_resp_s_empty_n = in_13_write_resp__empty_n;
  assign in_13_write_resp__read = krnl_partialKnn_wrapper_13_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_13_0_start_id_0 = 64'd106496;
  assign krnl_partialKnn_wrapper_14_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_14_0__ap_done = krnl_partialKnn_wrapper_14_0_ap_done;
  assign krnl_partialKnn_wrapper_14_0__ap_idle = krnl_partialKnn_wrapper_14_0_ap_idle;
  assign krnl_partialKnn_wrapper_14_0__ap_ready = krnl_partialKnn_wrapper_14_0_ap_ready;
  assign krnl_partialKnn_wrapper_14_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_14_0_ap_start = krnl_partialKnn_wrapper_14_0__ap_start;
  assign out_dist_14__din = krnl_partialKnn_wrapper_14_0_out_dist_din;
  assign krnl_partialKnn_wrapper_14_0_out_dist_full_n = out_dist_14__full_n;
  assign out_dist_14__write = krnl_partialKnn_wrapper_14_0_out_dist_write;
  assign out_id_14__din = krnl_partialKnn_wrapper_14_0_out_id_din;
  assign krnl_partialKnn_wrapper_14_0_out_id_full_n = out_id_14__full_n;
  assign out_id_14__write = krnl_partialKnn_wrapper_14_0_out_id_write;
  assign krnl_partialKnn_wrapper_14_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_14_0___in_14__q0;
  assign in_14_read_addr__din = krnl_partialKnn_wrapper_14_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_14_0_searchSpace_0_read_addr_s_full_n = in_14_read_addr__full_n;
  assign in_14_read_addr__write = krnl_partialKnn_wrapper_14_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_14_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_14_read_data__dout };
  assign krnl_partialKnn_wrapper_14_0_searchSpace_read_data_peek_empty_n = in_14_read_data__empty_n;
  assign krnl_partialKnn_wrapper_14_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_14_read_data__dout };
  assign krnl_partialKnn_wrapper_14_0_searchSpace_0_read_data_s_empty_n = in_14_read_data__empty_n;
  assign in_14_read_data__read = krnl_partialKnn_wrapper_14_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_14_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_14_0___in_14__q0;
  assign in_14_write_addr__din = krnl_partialKnn_wrapper_14_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_14_0_searchSpace_0_write_addr_s_full_n = in_14_write_addr__full_n;
  assign in_14_write_addr__write = krnl_partialKnn_wrapper_14_0_searchSpace_0_write_addr_s_write;
  assign in_14_write_data__din = krnl_partialKnn_wrapper_14_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_14_0_searchSpace_0_write_data_full_n = in_14_write_data__full_n;
  assign in_14_write_data__write = krnl_partialKnn_wrapper_14_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_14_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_14_write_resp__dout };
  assign krnl_partialKnn_wrapper_14_0_searchSpace_write_resp_peek_empty_n = in_14_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_14_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_14_write_resp__dout };
  assign krnl_partialKnn_wrapper_14_0_searchSpace_0_write_resp_s_empty_n = in_14_write_resp__empty_n;
  assign in_14_write_resp__read = krnl_partialKnn_wrapper_14_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_14_0_start_id_0 = 64'd114688;
  assign krnl_partialKnn_wrapper_15_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_15_0__ap_done = krnl_partialKnn_wrapper_15_0_ap_done;
  assign krnl_partialKnn_wrapper_15_0__ap_idle = krnl_partialKnn_wrapper_15_0_ap_idle;
  assign krnl_partialKnn_wrapper_15_0__ap_ready = krnl_partialKnn_wrapper_15_0_ap_ready;
  assign krnl_partialKnn_wrapper_15_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_15_0_ap_start = krnl_partialKnn_wrapper_15_0__ap_start;
  assign out_dist_15__din = krnl_partialKnn_wrapper_15_0_out_dist_din;
  assign krnl_partialKnn_wrapper_15_0_out_dist_full_n = out_dist_15__full_n;
  assign out_dist_15__write = krnl_partialKnn_wrapper_15_0_out_dist_write;
  assign out_id_15__din = krnl_partialKnn_wrapper_15_0_out_id_din;
  assign krnl_partialKnn_wrapper_15_0_out_id_full_n = out_id_15__full_n;
  assign out_id_15__write = krnl_partialKnn_wrapper_15_0_out_id_write;
  assign krnl_partialKnn_wrapper_15_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_15_0___in_15__q0;
  assign in_15_read_addr__din = krnl_partialKnn_wrapper_15_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_15_0_searchSpace_0_read_addr_s_full_n = in_15_read_addr__full_n;
  assign in_15_read_addr__write = krnl_partialKnn_wrapper_15_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_15_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_15_read_data__dout };
  assign krnl_partialKnn_wrapper_15_0_searchSpace_read_data_peek_empty_n = in_15_read_data__empty_n;
  assign krnl_partialKnn_wrapper_15_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_15_read_data__dout };
  assign krnl_partialKnn_wrapper_15_0_searchSpace_0_read_data_s_empty_n = in_15_read_data__empty_n;
  assign in_15_read_data__read = krnl_partialKnn_wrapper_15_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_15_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_15_0___in_15__q0;
  assign in_15_write_addr__din = krnl_partialKnn_wrapper_15_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_15_0_searchSpace_0_write_addr_s_full_n = in_15_write_addr__full_n;
  assign in_15_write_addr__write = krnl_partialKnn_wrapper_15_0_searchSpace_0_write_addr_s_write;
  assign in_15_write_data__din = krnl_partialKnn_wrapper_15_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_15_0_searchSpace_0_write_data_full_n = in_15_write_data__full_n;
  assign in_15_write_data__write = krnl_partialKnn_wrapper_15_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_15_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_15_write_resp__dout };
  assign krnl_partialKnn_wrapper_15_0_searchSpace_write_resp_peek_empty_n = in_15_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_15_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_15_write_resp__dout };
  assign krnl_partialKnn_wrapper_15_0_searchSpace_0_write_resp_s_empty_n = in_15_write_resp__empty_n;
  assign in_15_write_resp__read = krnl_partialKnn_wrapper_15_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_15_0_start_id_0 = 64'd122880;
  assign krnl_partialKnn_wrapper_16_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_16_0__ap_done = krnl_partialKnn_wrapper_16_0_ap_done;
  assign krnl_partialKnn_wrapper_16_0__ap_idle = krnl_partialKnn_wrapper_16_0_ap_idle;
  assign krnl_partialKnn_wrapper_16_0__ap_ready = krnl_partialKnn_wrapper_16_0_ap_ready;
  assign krnl_partialKnn_wrapper_16_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_16_0_ap_start = krnl_partialKnn_wrapper_16_0__ap_start;
  assign out_dist_16__din = krnl_partialKnn_wrapper_16_0_out_dist_din;
  assign krnl_partialKnn_wrapper_16_0_out_dist_full_n = out_dist_16__full_n;
  assign out_dist_16__write = krnl_partialKnn_wrapper_16_0_out_dist_write;
  assign out_id_16__din = krnl_partialKnn_wrapper_16_0_out_id_din;
  assign krnl_partialKnn_wrapper_16_0_out_id_full_n = out_id_16__full_n;
  assign out_id_16__write = krnl_partialKnn_wrapper_16_0_out_id_write;
  assign krnl_partialKnn_wrapper_16_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_16_0___in_16__q0;
  assign in_16_read_addr__din = krnl_partialKnn_wrapper_16_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_16_0_searchSpace_0_read_addr_s_full_n = in_16_read_addr__full_n;
  assign in_16_read_addr__write = krnl_partialKnn_wrapper_16_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_16_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_16_read_data__dout };
  assign krnl_partialKnn_wrapper_16_0_searchSpace_read_data_peek_empty_n = in_16_read_data__empty_n;
  assign krnl_partialKnn_wrapper_16_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_16_read_data__dout };
  assign krnl_partialKnn_wrapper_16_0_searchSpace_0_read_data_s_empty_n = in_16_read_data__empty_n;
  assign in_16_read_data__read = krnl_partialKnn_wrapper_16_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_16_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_16_0___in_16__q0;
  assign in_16_write_addr__din = krnl_partialKnn_wrapper_16_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_16_0_searchSpace_0_write_addr_s_full_n = in_16_write_addr__full_n;
  assign in_16_write_addr__write = krnl_partialKnn_wrapper_16_0_searchSpace_0_write_addr_s_write;
  assign in_16_write_data__din = krnl_partialKnn_wrapper_16_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_16_0_searchSpace_0_write_data_full_n = in_16_write_data__full_n;
  assign in_16_write_data__write = krnl_partialKnn_wrapper_16_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_16_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_16_write_resp__dout };
  assign krnl_partialKnn_wrapper_16_0_searchSpace_write_resp_peek_empty_n = in_16_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_16_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_16_write_resp__dout };
  assign krnl_partialKnn_wrapper_16_0_searchSpace_0_write_resp_s_empty_n = in_16_write_resp__empty_n;
  assign in_16_write_resp__read = krnl_partialKnn_wrapper_16_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_16_0_start_id_0 = 64'd131072;
  assign krnl_partialKnn_wrapper_17_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_17_0__ap_done = krnl_partialKnn_wrapper_17_0_ap_done;
  assign krnl_partialKnn_wrapper_17_0__ap_idle = krnl_partialKnn_wrapper_17_0_ap_idle;
  assign krnl_partialKnn_wrapper_17_0__ap_ready = krnl_partialKnn_wrapper_17_0_ap_ready;
  assign krnl_partialKnn_wrapper_17_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_17_0_ap_start = krnl_partialKnn_wrapper_17_0__ap_start;
  assign out_dist_17__din = krnl_partialKnn_wrapper_17_0_out_dist_din;
  assign krnl_partialKnn_wrapper_17_0_out_dist_full_n = out_dist_17__full_n;
  assign out_dist_17__write = krnl_partialKnn_wrapper_17_0_out_dist_write;
  assign out_id_17__din = krnl_partialKnn_wrapper_17_0_out_id_din;
  assign krnl_partialKnn_wrapper_17_0_out_id_full_n = out_id_17__full_n;
  assign out_id_17__write = krnl_partialKnn_wrapper_17_0_out_id_write;
  assign krnl_partialKnn_wrapper_17_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_17_0___in_17__q0;
  assign in_17_read_addr__din = krnl_partialKnn_wrapper_17_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_17_0_searchSpace_0_read_addr_s_full_n = in_17_read_addr__full_n;
  assign in_17_read_addr__write = krnl_partialKnn_wrapper_17_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_17_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_17_read_data__dout };
  assign krnl_partialKnn_wrapper_17_0_searchSpace_read_data_peek_empty_n = in_17_read_data__empty_n;
  assign krnl_partialKnn_wrapper_17_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_17_read_data__dout };
  assign krnl_partialKnn_wrapper_17_0_searchSpace_0_read_data_s_empty_n = in_17_read_data__empty_n;
  assign in_17_read_data__read = krnl_partialKnn_wrapper_17_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_17_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_17_0___in_17__q0;
  assign in_17_write_addr__din = krnl_partialKnn_wrapper_17_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_17_0_searchSpace_0_write_addr_s_full_n = in_17_write_addr__full_n;
  assign in_17_write_addr__write = krnl_partialKnn_wrapper_17_0_searchSpace_0_write_addr_s_write;
  assign in_17_write_data__din = krnl_partialKnn_wrapper_17_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_17_0_searchSpace_0_write_data_full_n = in_17_write_data__full_n;
  assign in_17_write_data__write = krnl_partialKnn_wrapper_17_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_17_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_17_write_resp__dout };
  assign krnl_partialKnn_wrapper_17_0_searchSpace_write_resp_peek_empty_n = in_17_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_17_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_17_write_resp__dout };
  assign krnl_partialKnn_wrapper_17_0_searchSpace_0_write_resp_s_empty_n = in_17_write_resp__empty_n;
  assign in_17_write_resp__read = krnl_partialKnn_wrapper_17_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_17_0_start_id_0 = 64'd139264;
  assign krnl_partialKnn_wrapper_18_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_18_0__ap_done = krnl_partialKnn_wrapper_18_0_ap_done;
  assign krnl_partialKnn_wrapper_18_0__ap_idle = krnl_partialKnn_wrapper_18_0_ap_idle;
  assign krnl_partialKnn_wrapper_18_0__ap_ready = krnl_partialKnn_wrapper_18_0_ap_ready;
  assign krnl_partialKnn_wrapper_18_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_18_0_ap_start = krnl_partialKnn_wrapper_18_0__ap_start;
  assign out_dist_18__din = krnl_partialKnn_wrapper_18_0_out_dist_din;
  assign krnl_partialKnn_wrapper_18_0_out_dist_full_n = out_dist_18__full_n;
  assign out_dist_18__write = krnl_partialKnn_wrapper_18_0_out_dist_write;
  assign out_id_18__din = krnl_partialKnn_wrapper_18_0_out_id_din;
  assign krnl_partialKnn_wrapper_18_0_out_id_full_n = out_id_18__full_n;
  assign out_id_18__write = krnl_partialKnn_wrapper_18_0_out_id_write;
  assign krnl_partialKnn_wrapper_18_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_18_0___in_18__q0;
  assign in_18_read_addr__din = krnl_partialKnn_wrapper_18_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_18_0_searchSpace_0_read_addr_s_full_n = in_18_read_addr__full_n;
  assign in_18_read_addr__write = krnl_partialKnn_wrapper_18_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_18_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_18_read_data__dout };
  assign krnl_partialKnn_wrapper_18_0_searchSpace_read_data_peek_empty_n = in_18_read_data__empty_n;
  assign krnl_partialKnn_wrapper_18_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_18_read_data__dout };
  assign krnl_partialKnn_wrapper_18_0_searchSpace_0_read_data_s_empty_n = in_18_read_data__empty_n;
  assign in_18_read_data__read = krnl_partialKnn_wrapper_18_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_18_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_18_0___in_18__q0;
  assign in_18_write_addr__din = krnl_partialKnn_wrapper_18_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_18_0_searchSpace_0_write_addr_s_full_n = in_18_write_addr__full_n;
  assign in_18_write_addr__write = krnl_partialKnn_wrapper_18_0_searchSpace_0_write_addr_s_write;
  assign in_18_write_data__din = krnl_partialKnn_wrapper_18_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_18_0_searchSpace_0_write_data_full_n = in_18_write_data__full_n;
  assign in_18_write_data__write = krnl_partialKnn_wrapper_18_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_18_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_18_write_resp__dout };
  assign krnl_partialKnn_wrapper_18_0_searchSpace_write_resp_peek_empty_n = in_18_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_18_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_18_write_resp__dout };
  assign krnl_partialKnn_wrapper_18_0_searchSpace_0_write_resp_s_empty_n = in_18_write_resp__empty_n;
  assign in_18_write_resp__read = krnl_partialKnn_wrapper_18_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_18_0_start_id_0 = 64'd147456;
  assign krnl_partialKnn_wrapper_19_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_19_0__ap_done = krnl_partialKnn_wrapper_19_0_ap_done;
  assign krnl_partialKnn_wrapper_19_0__ap_idle = krnl_partialKnn_wrapper_19_0_ap_idle;
  assign krnl_partialKnn_wrapper_19_0__ap_ready = krnl_partialKnn_wrapper_19_0_ap_ready;
  assign krnl_partialKnn_wrapper_19_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_19_0_ap_start = krnl_partialKnn_wrapper_19_0__ap_start;
  assign out_dist_19__din = krnl_partialKnn_wrapper_19_0_out_dist_din;
  assign krnl_partialKnn_wrapper_19_0_out_dist_full_n = out_dist_19__full_n;
  assign out_dist_19__write = krnl_partialKnn_wrapper_19_0_out_dist_write;
  assign out_id_19__din = krnl_partialKnn_wrapper_19_0_out_id_din;
  assign krnl_partialKnn_wrapper_19_0_out_id_full_n = out_id_19__full_n;
  assign out_id_19__write = krnl_partialKnn_wrapper_19_0_out_id_write;
  assign krnl_partialKnn_wrapper_19_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_19_0___in_19__q0;
  assign in_19_read_addr__din = krnl_partialKnn_wrapper_19_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_19_0_searchSpace_0_read_addr_s_full_n = in_19_read_addr__full_n;
  assign in_19_read_addr__write = krnl_partialKnn_wrapper_19_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_19_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_19_read_data__dout };
  assign krnl_partialKnn_wrapper_19_0_searchSpace_read_data_peek_empty_n = in_19_read_data__empty_n;
  assign krnl_partialKnn_wrapper_19_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_19_read_data__dout };
  assign krnl_partialKnn_wrapper_19_0_searchSpace_0_read_data_s_empty_n = in_19_read_data__empty_n;
  assign in_19_read_data__read = krnl_partialKnn_wrapper_19_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_19_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_19_0___in_19__q0;
  assign in_19_write_addr__din = krnl_partialKnn_wrapper_19_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_19_0_searchSpace_0_write_addr_s_full_n = in_19_write_addr__full_n;
  assign in_19_write_addr__write = krnl_partialKnn_wrapper_19_0_searchSpace_0_write_addr_s_write;
  assign in_19_write_data__din = krnl_partialKnn_wrapper_19_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_19_0_searchSpace_0_write_data_full_n = in_19_write_data__full_n;
  assign in_19_write_data__write = krnl_partialKnn_wrapper_19_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_19_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_19_write_resp__dout };
  assign krnl_partialKnn_wrapper_19_0_searchSpace_write_resp_peek_empty_n = in_19_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_19_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_19_write_resp__dout };
  assign krnl_partialKnn_wrapper_19_0_searchSpace_0_write_resp_s_empty_n = in_19_write_resp__empty_n;
  assign in_19_write_resp__read = krnl_partialKnn_wrapper_19_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_19_0_start_id_0 = 64'd155648;
  assign krnl_partialKnn_wrapper_2_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_2_0__ap_done = krnl_partialKnn_wrapper_2_0_ap_done;
  assign krnl_partialKnn_wrapper_2_0__ap_idle = krnl_partialKnn_wrapper_2_0_ap_idle;
  assign krnl_partialKnn_wrapper_2_0__ap_ready = krnl_partialKnn_wrapper_2_0_ap_ready;
  assign krnl_partialKnn_wrapper_2_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_2_0_ap_start = krnl_partialKnn_wrapper_2_0__ap_start;
  assign out_dist_2__din = krnl_partialKnn_wrapper_2_0_out_dist_din;
  assign krnl_partialKnn_wrapper_2_0_out_dist_full_n = out_dist_2__full_n;
  assign out_dist_2__write = krnl_partialKnn_wrapper_2_0_out_dist_write;
  assign out_id_2__din = krnl_partialKnn_wrapper_2_0_out_id_din;
  assign krnl_partialKnn_wrapper_2_0_out_id_full_n = out_id_2__full_n;
  assign out_id_2__write = krnl_partialKnn_wrapper_2_0_out_id_write;
  assign krnl_partialKnn_wrapper_2_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_2_0___in_2__q0;
  assign in_2_read_addr__din = krnl_partialKnn_wrapper_2_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_2_0_searchSpace_0_read_addr_s_full_n = in_2_read_addr__full_n;
  assign in_2_read_addr__write = krnl_partialKnn_wrapper_2_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_2_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_2_read_data__dout };
  assign krnl_partialKnn_wrapper_2_0_searchSpace_0_read_data_peek_empty_n = in_2_read_data__empty_n;
  assign krnl_partialKnn_wrapper_2_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_2_read_data__dout };
  assign krnl_partialKnn_wrapper_2_0_searchSpace_0_read_data_s_empty_n = in_2_read_data__empty_n;
  assign in_2_read_data__read = krnl_partialKnn_wrapper_2_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_2_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_2_0___in_2__q0;
  assign in_2_write_addr__din = krnl_partialKnn_wrapper_2_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_2_0_searchSpace_0_write_addr_s_full_n = in_2_write_addr__full_n;
  assign in_2_write_addr__write = krnl_partialKnn_wrapper_2_0_searchSpace_0_write_addr_s_write;
  assign in_2_write_data__din = krnl_partialKnn_wrapper_2_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_2_0_searchSpace_0_write_data_full_n = in_2_write_data__full_n;
  assign in_2_write_data__write = krnl_partialKnn_wrapper_2_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_2_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_2_write_resp__dout };
  assign krnl_partialKnn_wrapper_2_0_searchSpace_write_resp_peek_empty_n = in_2_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_2_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_2_write_resp__dout };
  assign krnl_partialKnn_wrapper_2_0_searchSpace_0_write_resp_s_empty_n = in_2_write_resp__empty_n;
  assign in_2_write_resp__read = krnl_partialKnn_wrapper_2_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_2_0_start_id_0 = 64'd16384;
  assign krnl_partialKnn_wrapper_20_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_20_0__ap_done = krnl_partialKnn_wrapper_20_0_ap_done;
  assign krnl_partialKnn_wrapper_20_0__ap_idle = krnl_partialKnn_wrapper_20_0_ap_idle;
  assign krnl_partialKnn_wrapper_20_0__ap_ready = krnl_partialKnn_wrapper_20_0_ap_ready;
  assign krnl_partialKnn_wrapper_20_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_20_0_ap_start = krnl_partialKnn_wrapper_20_0__ap_start;
  assign out_dist_20__din = krnl_partialKnn_wrapper_20_0_out_dist_din;
  assign krnl_partialKnn_wrapper_20_0_out_dist_full_n = out_dist_20__full_n;
  assign out_dist_20__write = krnl_partialKnn_wrapper_20_0_out_dist_write;
  assign out_id_20__din = krnl_partialKnn_wrapper_20_0_out_id_din;
  assign krnl_partialKnn_wrapper_20_0_out_id_full_n = out_id_20__full_n;
  assign out_id_20__write = krnl_partialKnn_wrapper_20_0_out_id_write;
  assign krnl_partialKnn_wrapper_20_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_20_0___in_20__q0;
  assign in_20_read_addr__din = krnl_partialKnn_wrapper_20_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_20_0_searchSpace_0_read_addr_s_full_n = in_20_read_addr__full_n;
  assign in_20_read_addr__write = krnl_partialKnn_wrapper_20_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_20_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_20_read_data__dout };
  assign krnl_partialKnn_wrapper_20_0_searchSpace_read_data_peek_empty_n = in_20_read_data__empty_n;
  assign krnl_partialKnn_wrapper_20_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_20_read_data__dout };
  assign krnl_partialKnn_wrapper_20_0_searchSpace_0_read_data_s_empty_n = in_20_read_data__empty_n;
  assign in_20_read_data__read = krnl_partialKnn_wrapper_20_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_20_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_20_0___in_20__q0;
  assign in_20_write_addr__din = krnl_partialKnn_wrapper_20_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_20_0_searchSpace_0_write_addr_s_full_n = in_20_write_addr__full_n;
  assign in_20_write_addr__write = krnl_partialKnn_wrapper_20_0_searchSpace_0_write_addr_s_write;
  assign in_20_write_data__din = krnl_partialKnn_wrapper_20_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_20_0_searchSpace_0_write_data_full_n = in_20_write_data__full_n;
  assign in_20_write_data__write = krnl_partialKnn_wrapper_20_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_20_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_20_write_resp__dout };
  assign krnl_partialKnn_wrapper_20_0_searchSpace_write_resp_peek_empty_n = in_20_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_20_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_20_write_resp__dout };
  assign krnl_partialKnn_wrapper_20_0_searchSpace_0_write_resp_s_empty_n = in_20_write_resp__empty_n;
  assign in_20_write_resp__read = krnl_partialKnn_wrapper_20_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_20_0_start_id_0 = 64'd163840;
  assign krnl_partialKnn_wrapper_21_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_21_0__ap_done = krnl_partialKnn_wrapper_21_0_ap_done;
  assign krnl_partialKnn_wrapper_21_0__ap_idle = krnl_partialKnn_wrapper_21_0_ap_idle;
  assign krnl_partialKnn_wrapper_21_0__ap_ready = krnl_partialKnn_wrapper_21_0_ap_ready;
  assign krnl_partialKnn_wrapper_21_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_21_0_ap_start = krnl_partialKnn_wrapper_21_0__ap_start;
  assign out_dist_21__din = krnl_partialKnn_wrapper_21_0_out_dist_din;
  assign krnl_partialKnn_wrapper_21_0_out_dist_full_n = out_dist_21__full_n;
  assign out_dist_21__write = krnl_partialKnn_wrapper_21_0_out_dist_write;
  assign out_id_21__din = krnl_partialKnn_wrapper_21_0_out_id_din;
  assign krnl_partialKnn_wrapper_21_0_out_id_full_n = out_id_21__full_n;
  assign out_id_21__write = krnl_partialKnn_wrapper_21_0_out_id_write;
  assign krnl_partialKnn_wrapper_21_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_21_0___in_21__q0;
  assign in_21_read_addr__din = krnl_partialKnn_wrapper_21_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_21_0_searchSpace_0_read_addr_s_full_n = in_21_read_addr__full_n;
  assign in_21_read_addr__write = krnl_partialKnn_wrapper_21_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_21_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_21_read_data__dout };
  assign krnl_partialKnn_wrapper_21_0_searchSpace_read_data_peek_empty_n = in_21_read_data__empty_n;
  assign krnl_partialKnn_wrapper_21_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_21_read_data__dout };
  assign krnl_partialKnn_wrapper_21_0_searchSpace_0_read_data_s_empty_n = in_21_read_data__empty_n;
  assign in_21_read_data__read = krnl_partialKnn_wrapper_21_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_21_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_21_0___in_21__q0;
  assign in_21_write_addr__din = krnl_partialKnn_wrapper_21_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_21_0_searchSpace_0_write_addr_s_full_n = in_21_write_addr__full_n;
  assign in_21_write_addr__write = krnl_partialKnn_wrapper_21_0_searchSpace_0_write_addr_s_write;
  assign in_21_write_data__din = krnl_partialKnn_wrapper_21_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_21_0_searchSpace_0_write_data_full_n = in_21_write_data__full_n;
  assign in_21_write_data__write = krnl_partialKnn_wrapper_21_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_21_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_21_write_resp__dout };
  assign krnl_partialKnn_wrapper_21_0_searchSpace_write_resp_peek_empty_n = in_21_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_21_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_21_write_resp__dout };
  assign krnl_partialKnn_wrapper_21_0_searchSpace_0_write_resp_s_empty_n = in_21_write_resp__empty_n;
  assign in_21_write_resp__read = krnl_partialKnn_wrapper_21_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_21_0_start_id_0 = 64'd172032;
  assign krnl_partialKnn_wrapper_22_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_22_0__ap_done = krnl_partialKnn_wrapper_22_0_ap_done;
  assign krnl_partialKnn_wrapper_22_0__ap_idle = krnl_partialKnn_wrapper_22_0_ap_idle;
  assign krnl_partialKnn_wrapper_22_0__ap_ready = krnl_partialKnn_wrapper_22_0_ap_ready;
  assign krnl_partialKnn_wrapper_22_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_22_0_ap_start = krnl_partialKnn_wrapper_22_0__ap_start;
  assign out_dist_22__din = krnl_partialKnn_wrapper_22_0_out_dist_din;
  assign krnl_partialKnn_wrapper_22_0_out_dist_full_n = out_dist_22__full_n;
  assign out_dist_22__write = krnl_partialKnn_wrapper_22_0_out_dist_write;
  assign out_id_22__din = krnl_partialKnn_wrapper_22_0_out_id_din;
  assign krnl_partialKnn_wrapper_22_0_out_id_full_n = out_id_22__full_n;
  assign out_id_22__write = krnl_partialKnn_wrapper_22_0_out_id_write;
  assign krnl_partialKnn_wrapper_22_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_22_0___in_22__q0;
  assign in_22_read_addr__din = krnl_partialKnn_wrapper_22_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_22_0_searchSpace_0_read_addr_s_full_n = in_22_read_addr__full_n;
  assign in_22_read_addr__write = krnl_partialKnn_wrapper_22_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_22_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_22_read_data__dout };
  assign krnl_partialKnn_wrapper_22_0_searchSpace_read_data_peek_empty_n = in_22_read_data__empty_n;
  assign krnl_partialKnn_wrapper_22_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_22_read_data__dout };
  assign krnl_partialKnn_wrapper_22_0_searchSpace_0_read_data_s_empty_n = in_22_read_data__empty_n;
  assign in_22_read_data__read = krnl_partialKnn_wrapper_22_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_22_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_22_0___in_22__q0;
  assign in_22_write_addr__din = krnl_partialKnn_wrapper_22_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_22_0_searchSpace_0_write_addr_s_full_n = in_22_write_addr__full_n;
  assign in_22_write_addr__write = krnl_partialKnn_wrapper_22_0_searchSpace_0_write_addr_s_write;
  assign in_22_write_data__din = krnl_partialKnn_wrapper_22_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_22_0_searchSpace_0_write_data_full_n = in_22_write_data__full_n;
  assign in_22_write_data__write = krnl_partialKnn_wrapper_22_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_22_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_22_write_resp__dout };
  assign krnl_partialKnn_wrapper_22_0_searchSpace_write_resp_peek_empty_n = in_22_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_22_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_22_write_resp__dout };
  assign krnl_partialKnn_wrapper_22_0_searchSpace_0_write_resp_s_empty_n = in_22_write_resp__empty_n;
  assign in_22_write_resp__read = krnl_partialKnn_wrapper_22_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_22_0_start_id_0 = 64'd180224;
  assign krnl_partialKnn_wrapper_23_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_23_0__ap_done = krnl_partialKnn_wrapper_23_0_ap_done;
  assign krnl_partialKnn_wrapper_23_0__ap_idle = krnl_partialKnn_wrapper_23_0_ap_idle;
  assign krnl_partialKnn_wrapper_23_0__ap_ready = krnl_partialKnn_wrapper_23_0_ap_ready;
  assign krnl_partialKnn_wrapper_23_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_23_0_ap_start = krnl_partialKnn_wrapper_23_0__ap_start;
  assign out_dist_23__din = krnl_partialKnn_wrapper_23_0_out_dist_din;
  assign krnl_partialKnn_wrapper_23_0_out_dist_full_n = out_dist_23__full_n;
  assign out_dist_23__write = krnl_partialKnn_wrapper_23_0_out_dist_write;
  assign out_id_23__din = krnl_partialKnn_wrapper_23_0_out_id_din;
  assign krnl_partialKnn_wrapper_23_0_out_id_full_n = out_id_23__full_n;
  assign out_id_23__write = krnl_partialKnn_wrapper_23_0_out_id_write;
  assign krnl_partialKnn_wrapper_23_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_23_0___in_23__q0;
  assign in_23_read_addr__din = krnl_partialKnn_wrapper_23_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_23_0_searchSpace_0_read_addr_s_full_n = in_23_read_addr__full_n;
  assign in_23_read_addr__write = krnl_partialKnn_wrapper_23_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_23_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_23_read_data__dout };
  assign krnl_partialKnn_wrapper_23_0_searchSpace_read_data_peek_empty_n = in_23_read_data__empty_n;
  assign krnl_partialKnn_wrapper_23_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_23_read_data__dout };
  assign krnl_partialKnn_wrapper_23_0_searchSpace_0_read_data_s_empty_n = in_23_read_data__empty_n;
  assign in_23_read_data__read = krnl_partialKnn_wrapper_23_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_23_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_23_0___in_23__q0;
  assign in_23_write_addr__din = krnl_partialKnn_wrapper_23_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_23_0_searchSpace_0_write_addr_s_full_n = in_23_write_addr__full_n;
  assign in_23_write_addr__write = krnl_partialKnn_wrapper_23_0_searchSpace_0_write_addr_s_write;
  assign in_23_write_data__din = krnl_partialKnn_wrapper_23_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_23_0_searchSpace_0_write_data_full_n = in_23_write_data__full_n;
  assign in_23_write_data__write = krnl_partialKnn_wrapper_23_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_23_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_23_write_resp__dout };
  assign krnl_partialKnn_wrapper_23_0_searchSpace_write_resp_peek_empty_n = in_23_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_23_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_23_write_resp__dout };
  assign krnl_partialKnn_wrapper_23_0_searchSpace_0_write_resp_s_empty_n = in_23_write_resp__empty_n;
  assign in_23_write_resp__read = krnl_partialKnn_wrapper_23_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_23_0_start_id_0 = 64'd188416;
  assign krnl_partialKnn_wrapper_24_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_24_0__ap_done = krnl_partialKnn_wrapper_24_0_ap_done;
  assign krnl_partialKnn_wrapper_24_0__ap_idle = krnl_partialKnn_wrapper_24_0_ap_idle;
  assign krnl_partialKnn_wrapper_24_0__ap_ready = krnl_partialKnn_wrapper_24_0_ap_ready;
  assign krnl_partialKnn_wrapper_24_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_24_0_ap_start = krnl_partialKnn_wrapper_24_0__ap_start;
  assign out_dist_24__din = krnl_partialKnn_wrapper_24_0_out_dist_din;
  assign krnl_partialKnn_wrapper_24_0_out_dist_full_n = out_dist_24__full_n;
  assign out_dist_24__write = krnl_partialKnn_wrapper_24_0_out_dist_write;
  assign out_id_24__din = krnl_partialKnn_wrapper_24_0_out_id_din;
  assign krnl_partialKnn_wrapper_24_0_out_id_full_n = out_id_24__full_n;
  assign out_id_24__write = krnl_partialKnn_wrapper_24_0_out_id_write;
  assign krnl_partialKnn_wrapper_24_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_24_0___in_24__q0;
  assign in_24_read_addr__din = krnl_partialKnn_wrapper_24_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_24_0_searchSpace_0_read_addr_s_full_n = in_24_read_addr__full_n;
  assign in_24_read_addr__write = krnl_partialKnn_wrapper_24_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_24_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_24_read_data__dout };
  assign krnl_partialKnn_wrapper_24_0_searchSpace_read_data_peek_empty_n = in_24_read_data__empty_n;
  assign krnl_partialKnn_wrapper_24_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_24_read_data__dout };
  assign krnl_partialKnn_wrapper_24_0_searchSpace_0_read_data_s_empty_n = in_24_read_data__empty_n;
  assign in_24_read_data__read = krnl_partialKnn_wrapper_24_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_24_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_24_0___in_24__q0;
  assign in_24_write_addr__din = krnl_partialKnn_wrapper_24_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_24_0_searchSpace_0_write_addr_s_full_n = in_24_write_addr__full_n;
  assign in_24_write_addr__write = krnl_partialKnn_wrapper_24_0_searchSpace_0_write_addr_s_write;
  assign in_24_write_data__din = krnl_partialKnn_wrapper_24_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_24_0_searchSpace_0_write_data_full_n = in_24_write_data__full_n;
  assign in_24_write_data__write = krnl_partialKnn_wrapper_24_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_24_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_24_write_resp__dout };
  assign krnl_partialKnn_wrapper_24_0_searchSpace_write_resp_peek_empty_n = in_24_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_24_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_24_write_resp__dout };
  assign krnl_partialKnn_wrapper_24_0_searchSpace_0_write_resp_s_empty_n = in_24_write_resp__empty_n;
  assign in_24_write_resp__read = krnl_partialKnn_wrapper_24_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_24_0_start_id_0 = 64'd196608;
  assign krnl_partialKnn_wrapper_25_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_25_0__ap_done = krnl_partialKnn_wrapper_25_0_ap_done;
  assign krnl_partialKnn_wrapper_25_0__ap_idle = krnl_partialKnn_wrapper_25_0_ap_idle;
  assign krnl_partialKnn_wrapper_25_0__ap_ready = krnl_partialKnn_wrapper_25_0_ap_ready;
  assign krnl_partialKnn_wrapper_25_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_25_0_ap_start = krnl_partialKnn_wrapper_25_0__ap_start;
  assign out_dist_25__din = krnl_partialKnn_wrapper_25_0_out_dist_din;
  assign krnl_partialKnn_wrapper_25_0_out_dist_full_n = out_dist_25__full_n;
  assign out_dist_25__write = krnl_partialKnn_wrapper_25_0_out_dist_write;
  assign out_id_25__din = krnl_partialKnn_wrapper_25_0_out_id_din;
  assign krnl_partialKnn_wrapper_25_0_out_id_full_n = out_id_25__full_n;
  assign out_id_25__write = krnl_partialKnn_wrapper_25_0_out_id_write;
  assign krnl_partialKnn_wrapper_25_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_25_0___in_25__q0;
  assign in_25_read_addr__din = krnl_partialKnn_wrapper_25_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_25_0_searchSpace_0_read_addr_s_full_n = in_25_read_addr__full_n;
  assign in_25_read_addr__write = krnl_partialKnn_wrapper_25_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_25_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_25_read_data__dout };
  assign krnl_partialKnn_wrapper_25_0_searchSpace_read_data_peek_empty_n = in_25_read_data__empty_n;
  assign krnl_partialKnn_wrapper_25_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_25_read_data__dout };
  assign krnl_partialKnn_wrapper_25_0_searchSpace_0_read_data_s_empty_n = in_25_read_data__empty_n;
  assign in_25_read_data__read = krnl_partialKnn_wrapper_25_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_25_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_25_0___in_25__q0;
  assign in_25_write_addr__din = krnl_partialKnn_wrapper_25_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_25_0_searchSpace_0_write_addr_s_full_n = in_25_write_addr__full_n;
  assign in_25_write_addr__write = krnl_partialKnn_wrapper_25_0_searchSpace_0_write_addr_s_write;
  assign in_25_write_data__din = krnl_partialKnn_wrapper_25_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_25_0_searchSpace_0_write_data_full_n = in_25_write_data__full_n;
  assign in_25_write_data__write = krnl_partialKnn_wrapper_25_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_25_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_25_write_resp__dout };
  assign krnl_partialKnn_wrapper_25_0_searchSpace_write_resp_peek_empty_n = in_25_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_25_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_25_write_resp__dout };
  assign krnl_partialKnn_wrapper_25_0_searchSpace_0_write_resp_s_empty_n = in_25_write_resp__empty_n;
  assign in_25_write_resp__read = krnl_partialKnn_wrapper_25_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_25_0_start_id_0 = 64'd204800;
  assign krnl_partialKnn_wrapper_26_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_26_0__ap_done = krnl_partialKnn_wrapper_26_0_ap_done;
  assign krnl_partialKnn_wrapper_26_0__ap_idle = krnl_partialKnn_wrapper_26_0_ap_idle;
  assign krnl_partialKnn_wrapper_26_0__ap_ready = krnl_partialKnn_wrapper_26_0_ap_ready;
  assign krnl_partialKnn_wrapper_26_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_26_0_ap_start = krnl_partialKnn_wrapper_26_0__ap_start;
  assign out_dist_26__din = krnl_partialKnn_wrapper_26_0_out_dist_din;
  assign krnl_partialKnn_wrapper_26_0_out_dist_full_n = out_dist_26__full_n;
  assign out_dist_26__write = krnl_partialKnn_wrapper_26_0_out_dist_write;
  assign out_id_26__din = krnl_partialKnn_wrapper_26_0_out_id_din;
  assign krnl_partialKnn_wrapper_26_0_out_id_full_n = out_id_26__full_n;
  assign out_id_26__write = krnl_partialKnn_wrapper_26_0_out_id_write;
  assign krnl_partialKnn_wrapper_26_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_26_0___in_26__q0;
  assign in_26_read_addr__din = krnl_partialKnn_wrapper_26_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_26_0_searchSpace_0_read_addr_s_full_n = in_26_read_addr__full_n;
  assign in_26_read_addr__write = krnl_partialKnn_wrapper_26_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_26_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_26_read_data__dout };
  assign krnl_partialKnn_wrapper_26_0_searchSpace_read_data_peek_empty_n = in_26_read_data__empty_n;
  assign krnl_partialKnn_wrapper_26_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_26_read_data__dout };
  assign krnl_partialKnn_wrapper_26_0_searchSpace_0_read_data_s_empty_n = in_26_read_data__empty_n;
  assign in_26_read_data__read = krnl_partialKnn_wrapper_26_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_26_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_26_0___in_26__q0;
  assign in_26_write_addr__din = krnl_partialKnn_wrapper_26_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_26_0_searchSpace_0_write_addr_s_full_n = in_26_write_addr__full_n;
  assign in_26_write_addr__write = krnl_partialKnn_wrapper_26_0_searchSpace_0_write_addr_s_write;
  assign in_26_write_data__din = krnl_partialKnn_wrapper_26_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_26_0_searchSpace_0_write_data_full_n = in_26_write_data__full_n;
  assign in_26_write_data__write = krnl_partialKnn_wrapper_26_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_26_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_26_write_resp__dout };
  assign krnl_partialKnn_wrapper_26_0_searchSpace_write_resp_peek_empty_n = in_26_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_26_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_26_write_resp__dout };
  assign krnl_partialKnn_wrapper_26_0_searchSpace_0_write_resp_s_empty_n = in_26_write_resp__empty_n;
  assign in_26_write_resp__read = krnl_partialKnn_wrapper_26_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_26_0_start_id_0 = 64'd212992;
  assign krnl_partialKnn_wrapper_27_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_27_0__ap_done = krnl_partialKnn_wrapper_27_0_ap_done;
  assign krnl_partialKnn_wrapper_27_0__ap_idle = krnl_partialKnn_wrapper_27_0_ap_idle;
  assign krnl_partialKnn_wrapper_27_0__ap_ready = krnl_partialKnn_wrapper_27_0_ap_ready;
  assign krnl_partialKnn_wrapper_27_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_27_0_ap_start = krnl_partialKnn_wrapper_27_0__ap_start;
  assign out_dist_27__din = krnl_partialKnn_wrapper_27_0_out_dist_din;
  assign krnl_partialKnn_wrapper_27_0_out_dist_full_n = out_dist_27__full_n;
  assign out_dist_27__write = krnl_partialKnn_wrapper_27_0_out_dist_write;
  assign out_id_27__din = krnl_partialKnn_wrapper_27_0_out_id_din;
  assign krnl_partialKnn_wrapper_27_0_out_id_full_n = out_id_27__full_n;
  assign out_id_27__write = krnl_partialKnn_wrapper_27_0_out_id_write;
  assign krnl_partialKnn_wrapper_27_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_27_0___in_27__q0;
  assign in_27_read_addr__din = krnl_partialKnn_wrapper_27_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_27_0_searchSpace_0_read_addr_s_full_n = in_27_read_addr__full_n;
  assign in_27_read_addr__write = krnl_partialKnn_wrapper_27_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_27_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_27_read_data__dout };
  assign krnl_partialKnn_wrapper_27_0_searchSpace_read_data_peek_empty_n = in_27_read_data__empty_n;
  assign krnl_partialKnn_wrapper_27_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_27_read_data__dout };
  assign krnl_partialKnn_wrapper_27_0_searchSpace_0_read_data_s_empty_n = in_27_read_data__empty_n;
  assign in_27_read_data__read = krnl_partialKnn_wrapper_27_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_27_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_27_0___in_27__q0;
  assign in_27_write_addr__din = krnl_partialKnn_wrapper_27_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_27_0_searchSpace_0_write_addr_s_full_n = in_27_write_addr__full_n;
  assign in_27_write_addr__write = krnl_partialKnn_wrapper_27_0_searchSpace_0_write_addr_s_write;
  assign in_27_write_data__din = krnl_partialKnn_wrapper_27_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_27_0_searchSpace_0_write_data_full_n = in_27_write_data__full_n;
  assign in_27_write_data__write = krnl_partialKnn_wrapper_27_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_27_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_27_write_resp__dout };
  assign krnl_partialKnn_wrapper_27_0_searchSpace_write_resp_peek_empty_n = in_27_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_27_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_27_write_resp__dout };
  assign krnl_partialKnn_wrapper_27_0_searchSpace_0_write_resp_s_empty_n = in_27_write_resp__empty_n;
  assign in_27_write_resp__read = krnl_partialKnn_wrapper_27_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_27_0_start_id_0 = 64'd221184;
  assign krnl_partialKnn_wrapper_28_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_28_0__ap_done = krnl_partialKnn_wrapper_28_0_ap_done;
  assign krnl_partialKnn_wrapper_28_0__ap_idle = krnl_partialKnn_wrapper_28_0_ap_idle;
  assign krnl_partialKnn_wrapper_28_0__ap_ready = krnl_partialKnn_wrapper_28_0_ap_ready;
  assign krnl_partialKnn_wrapper_28_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_28_0_ap_start = krnl_partialKnn_wrapper_28_0__ap_start;
  assign out_dist_28__din = krnl_partialKnn_wrapper_28_0_out_dist_din;
  assign krnl_partialKnn_wrapper_28_0_out_dist_full_n = out_dist_28__full_n;
  assign out_dist_28__write = krnl_partialKnn_wrapper_28_0_out_dist_write;
  assign out_id_28__din = krnl_partialKnn_wrapper_28_0_out_id_din;
  assign krnl_partialKnn_wrapper_28_0_out_id_full_n = out_id_28__full_n;
  assign out_id_28__write = krnl_partialKnn_wrapper_28_0_out_id_write;
  assign krnl_partialKnn_wrapper_28_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_28_0___in_28__q0;
  assign in_28_read_addr__din = krnl_partialKnn_wrapper_28_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_28_0_searchSpace_0_read_addr_s_full_n = in_28_read_addr__full_n;
  assign in_28_read_addr__write = krnl_partialKnn_wrapper_28_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_28_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_28_read_data__dout };
  assign krnl_partialKnn_wrapper_28_0_searchSpace_read_data_peek_empty_n = in_28_read_data__empty_n;
  assign krnl_partialKnn_wrapper_28_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_28_read_data__dout };
  assign krnl_partialKnn_wrapper_28_0_searchSpace_0_read_data_s_empty_n = in_28_read_data__empty_n;
  assign in_28_read_data__read = krnl_partialKnn_wrapper_28_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_28_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_28_0___in_28__q0;
  assign in_28_write_addr__din = krnl_partialKnn_wrapper_28_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_28_0_searchSpace_0_write_addr_s_full_n = in_28_write_addr__full_n;
  assign in_28_write_addr__write = krnl_partialKnn_wrapper_28_0_searchSpace_0_write_addr_s_write;
  assign in_28_write_data__din = krnl_partialKnn_wrapper_28_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_28_0_searchSpace_0_write_data_full_n = in_28_write_data__full_n;
  assign in_28_write_data__write = krnl_partialKnn_wrapper_28_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_28_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_28_write_resp__dout };
  assign krnl_partialKnn_wrapper_28_0_searchSpace_write_resp_peek_empty_n = in_28_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_28_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_28_write_resp__dout };
  assign krnl_partialKnn_wrapper_28_0_searchSpace_0_write_resp_s_empty_n = in_28_write_resp__empty_n;
  assign in_28_write_resp__read = krnl_partialKnn_wrapper_28_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_28_0_start_id_0 = 64'd229376;
  assign krnl_partialKnn_wrapper_29_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_29_0__ap_done = krnl_partialKnn_wrapper_29_0_ap_done;
  assign krnl_partialKnn_wrapper_29_0__ap_idle = krnl_partialKnn_wrapper_29_0_ap_idle;
  assign krnl_partialKnn_wrapper_29_0__ap_ready = krnl_partialKnn_wrapper_29_0_ap_ready;
  assign krnl_partialKnn_wrapper_29_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_29_0_ap_start = krnl_partialKnn_wrapper_29_0__ap_start;
  assign out_dist_29__din = krnl_partialKnn_wrapper_29_0_out_dist_din;
  assign krnl_partialKnn_wrapper_29_0_out_dist_full_n = out_dist_29__full_n;
  assign out_dist_29__write = krnl_partialKnn_wrapper_29_0_out_dist_write;
  assign out_id_29__din = krnl_partialKnn_wrapper_29_0_out_id_din;
  assign krnl_partialKnn_wrapper_29_0_out_id_full_n = out_id_29__full_n;
  assign out_id_29__write = krnl_partialKnn_wrapper_29_0_out_id_write;
  assign krnl_partialKnn_wrapper_29_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_29_0___in_29__q0;
  assign in_29_read_addr__din = krnl_partialKnn_wrapper_29_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_29_0_searchSpace_0_read_addr_s_full_n = in_29_read_addr__full_n;
  assign in_29_read_addr__write = krnl_partialKnn_wrapper_29_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_29_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_29_read_data__dout };
  assign krnl_partialKnn_wrapper_29_0_searchSpace_read_data_peek_empty_n = in_29_read_data__empty_n;
  assign krnl_partialKnn_wrapper_29_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_29_read_data__dout };
  assign krnl_partialKnn_wrapper_29_0_searchSpace_0_read_data_s_empty_n = in_29_read_data__empty_n;
  assign in_29_read_data__read = krnl_partialKnn_wrapper_29_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_29_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_29_0___in_29__q0;
  assign in_29_write_addr__din = krnl_partialKnn_wrapper_29_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_29_0_searchSpace_0_write_addr_s_full_n = in_29_write_addr__full_n;
  assign in_29_write_addr__write = krnl_partialKnn_wrapper_29_0_searchSpace_0_write_addr_s_write;
  assign in_29_write_data__din = krnl_partialKnn_wrapper_29_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_29_0_searchSpace_0_write_data_full_n = in_29_write_data__full_n;
  assign in_29_write_data__write = krnl_partialKnn_wrapper_29_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_29_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_29_write_resp__dout };
  assign krnl_partialKnn_wrapper_29_0_searchSpace_write_resp_peek_empty_n = in_29_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_29_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_29_write_resp__dout };
  assign krnl_partialKnn_wrapper_29_0_searchSpace_0_write_resp_s_empty_n = in_29_write_resp__empty_n;
  assign in_29_write_resp__read = krnl_partialKnn_wrapper_29_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_29_0_start_id_0 = 64'd237568;
  assign krnl_partialKnn_wrapper_3_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_3_0__ap_done = krnl_partialKnn_wrapper_3_0_ap_done;
  assign krnl_partialKnn_wrapper_3_0__ap_idle = krnl_partialKnn_wrapper_3_0_ap_idle;
  assign krnl_partialKnn_wrapper_3_0__ap_ready = krnl_partialKnn_wrapper_3_0_ap_ready;
  assign krnl_partialKnn_wrapper_3_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_3_0_ap_start = krnl_partialKnn_wrapper_3_0__ap_start;
  assign out_dist_3__din = krnl_partialKnn_wrapper_3_0_out_dist_din;
  assign krnl_partialKnn_wrapper_3_0_out_dist_full_n = out_dist_3__full_n;
  assign out_dist_3__write = krnl_partialKnn_wrapper_3_0_out_dist_write;
  assign out_id_3__din = krnl_partialKnn_wrapper_3_0_out_id_din;
  assign krnl_partialKnn_wrapper_3_0_out_id_full_n = out_id_3__full_n;
  assign out_id_3__write = krnl_partialKnn_wrapper_3_0_out_id_write;
  assign krnl_partialKnn_wrapper_3_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_3_0___in_3__q0;
  assign in_3_read_addr__din = krnl_partialKnn_wrapper_3_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_3_0_searchSpace_0_read_addr_s_full_n = in_3_read_addr__full_n;
  assign in_3_read_addr__write = krnl_partialKnn_wrapper_3_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_3_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_3_read_data__dout };
  assign krnl_partialKnn_wrapper_3_0_searchSpace_0_read_data_peek_empty_n = in_3_read_data__empty_n;
  assign krnl_partialKnn_wrapper_3_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_3_read_data__dout };
  assign krnl_partialKnn_wrapper_3_0_searchSpace_0_read_data_s_empty_n = in_3_read_data__empty_n;
  assign in_3_read_data__read = krnl_partialKnn_wrapper_3_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_3_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_3_0___in_3__q0;
  assign in_3_write_addr__din = krnl_partialKnn_wrapper_3_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_3_0_searchSpace_0_write_addr_s_full_n = in_3_write_addr__full_n;
  assign in_3_write_addr__write = krnl_partialKnn_wrapper_3_0_searchSpace_0_write_addr_s_write;
  assign in_3_write_data__din = krnl_partialKnn_wrapper_3_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_3_0_searchSpace_0_write_data_full_n = in_3_write_data__full_n;
  assign in_3_write_data__write = krnl_partialKnn_wrapper_3_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_3_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_3_write_resp__dout };
  assign krnl_partialKnn_wrapper_3_0_searchSpace_write_resp_peek_empty_n = in_3_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_3_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_3_write_resp__dout };
  assign krnl_partialKnn_wrapper_3_0_searchSpace_0_write_resp_s_empty_n = in_3_write_resp__empty_n;
  assign in_3_write_resp__read = krnl_partialKnn_wrapper_3_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_3_0_start_id_0 = 64'd24576;
  assign krnl_partialKnn_wrapper_30_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_30_0__ap_done = krnl_partialKnn_wrapper_30_0_ap_done;
  assign krnl_partialKnn_wrapper_30_0__ap_idle = krnl_partialKnn_wrapper_30_0_ap_idle;
  assign krnl_partialKnn_wrapper_30_0__ap_ready = krnl_partialKnn_wrapper_30_0_ap_ready;
  assign krnl_partialKnn_wrapper_30_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_30_0_ap_start = krnl_partialKnn_wrapper_30_0__ap_start;
  assign out_dist_30__din = krnl_partialKnn_wrapper_30_0_out_dist_din;
  assign krnl_partialKnn_wrapper_30_0_out_dist_full_n = out_dist_30__full_n;
  assign out_dist_30__write = krnl_partialKnn_wrapper_30_0_out_dist_write;
  assign out_id_30__din = krnl_partialKnn_wrapper_30_0_out_id_din;
  assign krnl_partialKnn_wrapper_30_0_out_id_full_n = out_id_30__full_n;
  assign out_id_30__write = krnl_partialKnn_wrapper_30_0_out_id_write;
  assign krnl_partialKnn_wrapper_30_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_30_0___in_30__q0;
  assign in_30_read_addr__din = krnl_partialKnn_wrapper_30_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_30_0_searchSpace_0_read_addr_s_full_n = in_30_read_addr__full_n;
  assign in_30_read_addr__write = krnl_partialKnn_wrapper_30_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_30_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_30_read_data__dout };
  assign krnl_partialKnn_wrapper_30_0_searchSpace_read_data_peek_empty_n = in_30_read_data__empty_n;
  assign krnl_partialKnn_wrapper_30_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_30_read_data__dout };
  assign krnl_partialKnn_wrapper_30_0_searchSpace_0_read_data_s_empty_n = in_30_read_data__empty_n;
  assign in_30_read_data__read = krnl_partialKnn_wrapper_30_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_30_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_30_0___in_30__q0;
  assign in_30_write_addr__din = krnl_partialKnn_wrapper_30_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_30_0_searchSpace_0_write_addr_s_full_n = in_30_write_addr__full_n;
  assign in_30_write_addr__write = krnl_partialKnn_wrapper_30_0_searchSpace_0_write_addr_s_write;
  assign in_30_write_data__din = krnl_partialKnn_wrapper_30_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_30_0_searchSpace_0_write_data_full_n = in_30_write_data__full_n;
  assign in_30_write_data__write = krnl_partialKnn_wrapper_30_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_30_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_30_write_resp__dout };
  assign krnl_partialKnn_wrapper_30_0_searchSpace_write_resp_peek_empty_n = in_30_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_30_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_30_write_resp__dout };
  assign krnl_partialKnn_wrapper_30_0_searchSpace_0_write_resp_s_empty_n = in_30_write_resp__empty_n;
  assign in_30_write_resp__read = krnl_partialKnn_wrapper_30_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_30_0_start_id_0 = 64'd245760;
  assign krnl_partialKnn_wrapper_31_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_31_0__ap_done = krnl_partialKnn_wrapper_31_0_ap_done;
  assign krnl_partialKnn_wrapper_31_0__ap_idle = krnl_partialKnn_wrapper_31_0_ap_idle;
  assign krnl_partialKnn_wrapper_31_0__ap_ready = krnl_partialKnn_wrapper_31_0_ap_ready;
  assign krnl_partialKnn_wrapper_31_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_31_0_ap_start = krnl_partialKnn_wrapper_31_0__ap_start;
  assign out_dist_31__din = krnl_partialKnn_wrapper_31_0_out_dist_din;
  assign krnl_partialKnn_wrapper_31_0_out_dist_full_n = out_dist_31__full_n;
  assign out_dist_31__write = krnl_partialKnn_wrapper_31_0_out_dist_write;
  assign out_id_31__din = krnl_partialKnn_wrapper_31_0_out_id_din;
  assign krnl_partialKnn_wrapper_31_0_out_id_full_n = out_id_31__full_n;
  assign out_id_31__write = krnl_partialKnn_wrapper_31_0_out_id_write;
  assign krnl_partialKnn_wrapper_31_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_31_0___in_31__q0;
  assign in_31_read_addr__din = krnl_partialKnn_wrapper_31_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_31_0_searchSpace_0_read_addr_s_full_n = in_31_read_addr__full_n;
  assign in_31_read_addr__write = krnl_partialKnn_wrapper_31_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_31_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_31_read_data__dout };
  assign krnl_partialKnn_wrapper_31_0_searchSpace_read_data_peek_empty_n = in_31_read_data__empty_n;
  assign krnl_partialKnn_wrapper_31_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_31_read_data__dout };
  assign krnl_partialKnn_wrapper_31_0_searchSpace_0_read_data_s_empty_n = in_31_read_data__empty_n;
  assign in_31_read_data__read = krnl_partialKnn_wrapper_31_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_31_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_31_0___in_31__q0;
  assign in_31_write_addr__din = krnl_partialKnn_wrapper_31_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_31_0_searchSpace_0_write_addr_s_full_n = in_31_write_addr__full_n;
  assign in_31_write_addr__write = krnl_partialKnn_wrapper_31_0_searchSpace_0_write_addr_s_write;
  assign in_31_write_data__din = krnl_partialKnn_wrapper_31_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_31_0_searchSpace_0_write_data_full_n = in_31_write_data__full_n;
  assign in_31_write_data__write = krnl_partialKnn_wrapper_31_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_31_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_31_write_resp__dout };
  assign krnl_partialKnn_wrapper_31_0_searchSpace_write_resp_peek_empty_n = in_31_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_31_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_31_write_resp__dout };
  assign krnl_partialKnn_wrapper_31_0_searchSpace_0_write_resp_s_empty_n = in_31_write_resp__empty_n;
  assign in_31_write_resp__read = krnl_partialKnn_wrapper_31_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_31_0_start_id_0 = 64'd253952;
  assign krnl_partialKnn_wrapper_32_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_32_0__ap_done = krnl_partialKnn_wrapper_32_0_ap_done;
  assign krnl_partialKnn_wrapper_32_0__ap_idle = krnl_partialKnn_wrapper_32_0_ap_idle;
  assign krnl_partialKnn_wrapper_32_0__ap_ready = krnl_partialKnn_wrapper_32_0_ap_ready;
  assign krnl_partialKnn_wrapper_32_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_32_0_ap_start = krnl_partialKnn_wrapper_32_0__ap_start;
  assign out_dist_32__din = krnl_partialKnn_wrapper_32_0_out_dist_din;
  assign krnl_partialKnn_wrapper_32_0_out_dist_full_n = out_dist_32__full_n;
  assign out_dist_32__write = krnl_partialKnn_wrapper_32_0_out_dist_write;
  assign out_id_32__din = krnl_partialKnn_wrapper_32_0_out_id_din;
  assign krnl_partialKnn_wrapper_32_0_out_id_full_n = out_id_32__full_n;
  assign out_id_32__write = krnl_partialKnn_wrapper_32_0_out_id_write;
  assign krnl_partialKnn_wrapper_32_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_32_0___in_32__q0;
  assign in_32_read_addr__din = krnl_partialKnn_wrapper_32_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_32_0_searchSpace_0_read_addr_s_full_n = in_32_read_addr__full_n;
  assign in_32_read_addr__write = krnl_partialKnn_wrapper_32_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_32_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_32_read_data__dout };
  assign krnl_partialKnn_wrapper_32_0_searchSpace_read_data_peek_empty_n = in_32_read_data__empty_n;
  assign krnl_partialKnn_wrapper_32_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_32_read_data__dout };
  assign krnl_partialKnn_wrapper_32_0_searchSpace_0_read_data_s_empty_n = in_32_read_data__empty_n;
  assign in_32_read_data__read = krnl_partialKnn_wrapper_32_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_32_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_32_0___in_32__q0;
  assign in_32_write_addr__din = krnl_partialKnn_wrapper_32_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_32_0_searchSpace_0_write_addr_s_full_n = in_32_write_addr__full_n;
  assign in_32_write_addr__write = krnl_partialKnn_wrapper_32_0_searchSpace_0_write_addr_s_write;
  assign in_32_write_data__din = krnl_partialKnn_wrapper_32_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_32_0_searchSpace_0_write_data_full_n = in_32_write_data__full_n;
  assign in_32_write_data__write = krnl_partialKnn_wrapper_32_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_32_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_32_write_resp__dout };
  assign krnl_partialKnn_wrapper_32_0_searchSpace_write_resp_peek_empty_n = in_32_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_32_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_32_write_resp__dout };
  assign krnl_partialKnn_wrapper_32_0_searchSpace_0_write_resp_s_empty_n = in_32_write_resp__empty_n;
  assign in_32_write_resp__read = krnl_partialKnn_wrapper_32_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_32_0_start_id_0 = 64'd262144;
  assign krnl_partialKnn_wrapper_33_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_33_0__ap_done = krnl_partialKnn_wrapper_33_0_ap_done;
  assign krnl_partialKnn_wrapper_33_0__ap_idle = krnl_partialKnn_wrapper_33_0_ap_idle;
  assign krnl_partialKnn_wrapper_33_0__ap_ready = krnl_partialKnn_wrapper_33_0_ap_ready;
  assign krnl_partialKnn_wrapper_33_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_33_0_ap_start = krnl_partialKnn_wrapper_33_0__ap_start;
  assign out_dist_33__din = krnl_partialKnn_wrapper_33_0_out_dist_din;
  assign krnl_partialKnn_wrapper_33_0_out_dist_full_n = out_dist_33__full_n;
  assign out_dist_33__write = krnl_partialKnn_wrapper_33_0_out_dist_write;
  assign out_id_33__din = krnl_partialKnn_wrapper_33_0_out_id_din;
  assign krnl_partialKnn_wrapper_33_0_out_id_full_n = out_id_33__full_n;
  assign out_id_33__write = krnl_partialKnn_wrapper_33_0_out_id_write;
  assign krnl_partialKnn_wrapper_33_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_33_0___in_33__q0;
  assign in_33_read_addr__din = krnl_partialKnn_wrapper_33_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_33_0_searchSpace_0_read_addr_s_full_n = in_33_read_addr__full_n;
  assign in_33_read_addr__write = krnl_partialKnn_wrapper_33_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_33_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_33_read_data__dout };
  assign krnl_partialKnn_wrapper_33_0_searchSpace_read_data_peek_empty_n = in_33_read_data__empty_n;
  assign krnl_partialKnn_wrapper_33_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_33_read_data__dout };
  assign krnl_partialKnn_wrapper_33_0_searchSpace_0_read_data_s_empty_n = in_33_read_data__empty_n;
  assign in_33_read_data__read = krnl_partialKnn_wrapper_33_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_33_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_33_0___in_33__q0;
  assign in_33_write_addr__din = krnl_partialKnn_wrapper_33_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_33_0_searchSpace_0_write_addr_s_full_n = in_33_write_addr__full_n;
  assign in_33_write_addr__write = krnl_partialKnn_wrapper_33_0_searchSpace_0_write_addr_s_write;
  assign in_33_write_data__din = krnl_partialKnn_wrapper_33_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_33_0_searchSpace_0_write_data_full_n = in_33_write_data__full_n;
  assign in_33_write_data__write = krnl_partialKnn_wrapper_33_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_33_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_33_write_resp__dout };
  assign krnl_partialKnn_wrapper_33_0_searchSpace_write_resp_peek_empty_n = in_33_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_33_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_33_write_resp__dout };
  assign krnl_partialKnn_wrapper_33_0_searchSpace_0_write_resp_s_empty_n = in_33_write_resp__empty_n;
  assign in_33_write_resp__read = krnl_partialKnn_wrapper_33_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_33_0_start_id_0 = 64'd270336;
  assign krnl_partialKnn_wrapper_34_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_34_0__ap_done = krnl_partialKnn_wrapper_34_0_ap_done;
  assign krnl_partialKnn_wrapper_34_0__ap_idle = krnl_partialKnn_wrapper_34_0_ap_idle;
  assign krnl_partialKnn_wrapper_34_0__ap_ready = krnl_partialKnn_wrapper_34_0_ap_ready;
  assign krnl_partialKnn_wrapper_34_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_34_0_ap_start = krnl_partialKnn_wrapper_34_0__ap_start;
  assign out_dist_34__din = krnl_partialKnn_wrapper_34_0_out_dist_din;
  assign krnl_partialKnn_wrapper_34_0_out_dist_full_n = out_dist_34__full_n;
  assign out_dist_34__write = krnl_partialKnn_wrapper_34_0_out_dist_write;
  assign out_id_34__din = krnl_partialKnn_wrapper_34_0_out_id_din;
  assign krnl_partialKnn_wrapper_34_0_out_id_full_n = out_id_34__full_n;
  assign out_id_34__write = krnl_partialKnn_wrapper_34_0_out_id_write;
  assign krnl_partialKnn_wrapper_34_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_34_0___in_34__q0;
  assign in_34_read_addr__din = krnl_partialKnn_wrapper_34_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_34_0_searchSpace_0_read_addr_s_full_n = in_34_read_addr__full_n;
  assign in_34_read_addr__write = krnl_partialKnn_wrapper_34_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_34_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_34_read_data__dout };
  assign krnl_partialKnn_wrapper_34_0_searchSpace_read_data_peek_empty_n = in_34_read_data__empty_n;
  assign krnl_partialKnn_wrapper_34_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_34_read_data__dout };
  assign krnl_partialKnn_wrapper_34_0_searchSpace_0_read_data_s_empty_n = in_34_read_data__empty_n;
  assign in_34_read_data__read = krnl_partialKnn_wrapper_34_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_34_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_34_0___in_34__q0;
  assign in_34_write_addr__din = krnl_partialKnn_wrapper_34_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_34_0_searchSpace_0_write_addr_s_full_n = in_34_write_addr__full_n;
  assign in_34_write_addr__write = krnl_partialKnn_wrapper_34_0_searchSpace_0_write_addr_s_write;
  assign in_34_write_data__din = krnl_partialKnn_wrapper_34_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_34_0_searchSpace_0_write_data_full_n = in_34_write_data__full_n;
  assign in_34_write_data__write = krnl_partialKnn_wrapper_34_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_34_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_34_write_resp__dout };
  assign krnl_partialKnn_wrapper_34_0_searchSpace_write_resp_peek_empty_n = in_34_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_34_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_34_write_resp__dout };
  assign krnl_partialKnn_wrapper_34_0_searchSpace_0_write_resp_s_empty_n = in_34_write_resp__empty_n;
  assign in_34_write_resp__read = krnl_partialKnn_wrapper_34_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_34_0_start_id_0 = 64'd278528;
  assign krnl_partialKnn_wrapper_35_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_35_0__ap_done = krnl_partialKnn_wrapper_35_0_ap_done;
  assign krnl_partialKnn_wrapper_35_0__ap_idle = krnl_partialKnn_wrapper_35_0_ap_idle;
  assign krnl_partialKnn_wrapper_35_0__ap_ready = krnl_partialKnn_wrapper_35_0_ap_ready;
  assign krnl_partialKnn_wrapper_35_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_35_0_ap_start = krnl_partialKnn_wrapper_35_0__ap_start;
  assign out_dist_35__din = krnl_partialKnn_wrapper_35_0_out_dist_din;
  assign krnl_partialKnn_wrapper_35_0_out_dist_full_n = out_dist_35__full_n;
  assign out_dist_35__write = krnl_partialKnn_wrapper_35_0_out_dist_write;
  assign out_id_35__din = krnl_partialKnn_wrapper_35_0_out_id_din;
  assign krnl_partialKnn_wrapper_35_0_out_id_full_n = out_id_35__full_n;
  assign out_id_35__write = krnl_partialKnn_wrapper_35_0_out_id_write;
  assign krnl_partialKnn_wrapper_35_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_35_0___in_35__q0;
  assign in_35_read_addr__din = krnl_partialKnn_wrapper_35_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_35_0_searchSpace_0_read_addr_s_full_n = in_35_read_addr__full_n;
  assign in_35_read_addr__write = krnl_partialKnn_wrapper_35_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_35_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_35_read_data__dout };
  assign krnl_partialKnn_wrapper_35_0_searchSpace_read_data_peek_empty_n = in_35_read_data__empty_n;
  assign krnl_partialKnn_wrapper_35_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_35_read_data__dout };
  assign krnl_partialKnn_wrapper_35_0_searchSpace_0_read_data_s_empty_n = in_35_read_data__empty_n;
  assign in_35_read_data__read = krnl_partialKnn_wrapper_35_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_35_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_35_0___in_35__q0;
  assign in_35_write_addr__din = krnl_partialKnn_wrapper_35_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_35_0_searchSpace_0_write_addr_s_full_n = in_35_write_addr__full_n;
  assign in_35_write_addr__write = krnl_partialKnn_wrapper_35_0_searchSpace_0_write_addr_s_write;
  assign in_35_write_data__din = krnl_partialKnn_wrapper_35_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_35_0_searchSpace_0_write_data_full_n = in_35_write_data__full_n;
  assign in_35_write_data__write = krnl_partialKnn_wrapper_35_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_35_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_35_write_resp__dout };
  assign krnl_partialKnn_wrapper_35_0_searchSpace_write_resp_peek_empty_n = in_35_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_35_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_35_write_resp__dout };
  assign krnl_partialKnn_wrapper_35_0_searchSpace_0_write_resp_s_empty_n = in_35_write_resp__empty_n;
  assign in_35_write_resp__read = krnl_partialKnn_wrapper_35_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_35_0_start_id_0 = 64'd286720;
  assign krnl_partialKnn_wrapper_36_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_36_0__ap_done = krnl_partialKnn_wrapper_36_0_ap_done;
  assign krnl_partialKnn_wrapper_36_0__ap_idle = krnl_partialKnn_wrapper_36_0_ap_idle;
  assign krnl_partialKnn_wrapper_36_0__ap_ready = krnl_partialKnn_wrapper_36_0_ap_ready;
  assign krnl_partialKnn_wrapper_36_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_36_0_ap_start = krnl_partialKnn_wrapper_36_0__ap_start;
  assign out_dist_36__din = krnl_partialKnn_wrapper_36_0_out_dist_din;
  assign krnl_partialKnn_wrapper_36_0_out_dist_full_n = out_dist_36__full_n;
  assign out_dist_36__write = krnl_partialKnn_wrapper_36_0_out_dist_write;
  assign out_id_36__din = krnl_partialKnn_wrapper_36_0_out_id_din;
  assign krnl_partialKnn_wrapper_36_0_out_id_full_n = out_id_36__full_n;
  assign out_id_36__write = krnl_partialKnn_wrapper_36_0_out_id_write;
  assign krnl_partialKnn_wrapper_36_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_36_0___in_36__q0;
  assign in_36_read_addr__din = krnl_partialKnn_wrapper_36_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_36_0_searchSpace_0_read_addr_s_full_n = in_36_read_addr__full_n;
  assign in_36_read_addr__write = krnl_partialKnn_wrapper_36_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_36_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_36_read_data__dout };
  assign krnl_partialKnn_wrapper_36_0_searchSpace_read_data_peek_empty_n = in_36_read_data__empty_n;
  assign krnl_partialKnn_wrapper_36_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_36_read_data__dout };
  assign krnl_partialKnn_wrapper_36_0_searchSpace_0_read_data_s_empty_n = in_36_read_data__empty_n;
  assign in_36_read_data__read = krnl_partialKnn_wrapper_36_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_36_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_36_0___in_36__q0;
  assign in_36_write_addr__din = krnl_partialKnn_wrapper_36_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_36_0_searchSpace_0_write_addr_s_full_n = in_36_write_addr__full_n;
  assign in_36_write_addr__write = krnl_partialKnn_wrapper_36_0_searchSpace_0_write_addr_s_write;
  assign in_36_write_data__din = krnl_partialKnn_wrapper_36_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_36_0_searchSpace_0_write_data_full_n = in_36_write_data__full_n;
  assign in_36_write_data__write = krnl_partialKnn_wrapper_36_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_36_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_36_write_resp__dout };
  assign krnl_partialKnn_wrapper_36_0_searchSpace_write_resp_peek_empty_n = in_36_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_36_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_36_write_resp__dout };
  assign krnl_partialKnn_wrapper_36_0_searchSpace_0_write_resp_s_empty_n = in_36_write_resp__empty_n;
  assign in_36_write_resp__read = krnl_partialKnn_wrapper_36_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_36_0_start_id_0 = 64'd294912;
  assign krnl_partialKnn_wrapper_37_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_37_0__ap_done = krnl_partialKnn_wrapper_37_0_ap_done;
  assign krnl_partialKnn_wrapper_37_0__ap_idle = krnl_partialKnn_wrapper_37_0_ap_idle;
  assign krnl_partialKnn_wrapper_37_0__ap_ready = krnl_partialKnn_wrapper_37_0_ap_ready;
  assign krnl_partialKnn_wrapper_37_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_37_0_ap_start = krnl_partialKnn_wrapper_37_0__ap_start;
  assign out_dist_37__din = krnl_partialKnn_wrapper_37_0_out_dist_din;
  assign krnl_partialKnn_wrapper_37_0_out_dist_full_n = out_dist_37__full_n;
  assign out_dist_37__write = krnl_partialKnn_wrapper_37_0_out_dist_write;
  assign out_id_37__din = krnl_partialKnn_wrapper_37_0_out_id_din;
  assign krnl_partialKnn_wrapper_37_0_out_id_full_n = out_id_37__full_n;
  assign out_id_37__write = krnl_partialKnn_wrapper_37_0_out_id_write;
  assign krnl_partialKnn_wrapper_37_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_37_0___in_37__q0;
  assign in_37_read_addr__din = krnl_partialKnn_wrapper_37_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_37_0_searchSpace_0_read_addr_s_full_n = in_37_read_addr__full_n;
  assign in_37_read_addr__write = krnl_partialKnn_wrapper_37_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_37_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_37_read_data__dout };
  assign krnl_partialKnn_wrapper_37_0_searchSpace_read_data_peek_empty_n = in_37_read_data__empty_n;
  assign krnl_partialKnn_wrapper_37_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_37_read_data__dout };
  assign krnl_partialKnn_wrapper_37_0_searchSpace_0_read_data_s_empty_n = in_37_read_data__empty_n;
  assign in_37_read_data__read = krnl_partialKnn_wrapper_37_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_37_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_37_0___in_37__q0;
  assign in_37_write_addr__din = krnl_partialKnn_wrapper_37_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_37_0_searchSpace_0_write_addr_s_full_n = in_37_write_addr__full_n;
  assign in_37_write_addr__write = krnl_partialKnn_wrapper_37_0_searchSpace_0_write_addr_s_write;
  assign in_37_write_data__din = krnl_partialKnn_wrapper_37_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_37_0_searchSpace_0_write_data_full_n = in_37_write_data__full_n;
  assign in_37_write_data__write = krnl_partialKnn_wrapper_37_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_37_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_37_write_resp__dout };
  assign krnl_partialKnn_wrapper_37_0_searchSpace_write_resp_peek_empty_n = in_37_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_37_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_37_write_resp__dout };
  assign krnl_partialKnn_wrapper_37_0_searchSpace_0_write_resp_s_empty_n = in_37_write_resp__empty_n;
  assign in_37_write_resp__read = krnl_partialKnn_wrapper_37_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_37_0_start_id_0 = 64'd303104;
  assign krnl_partialKnn_wrapper_38_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_38_0__ap_done = krnl_partialKnn_wrapper_38_0_ap_done;
  assign krnl_partialKnn_wrapper_38_0__ap_idle = krnl_partialKnn_wrapper_38_0_ap_idle;
  assign krnl_partialKnn_wrapper_38_0__ap_ready = krnl_partialKnn_wrapper_38_0_ap_ready;
  assign krnl_partialKnn_wrapper_38_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_38_0_ap_start = krnl_partialKnn_wrapper_38_0__ap_start;
  assign out_dist_38__din = krnl_partialKnn_wrapper_38_0_out_dist_din;
  assign krnl_partialKnn_wrapper_38_0_out_dist_full_n = out_dist_38__full_n;
  assign out_dist_38__write = krnl_partialKnn_wrapper_38_0_out_dist_write;
  assign out_id_38__din = krnl_partialKnn_wrapper_38_0_out_id_din;
  assign krnl_partialKnn_wrapper_38_0_out_id_full_n = out_id_38__full_n;
  assign out_id_38__write = krnl_partialKnn_wrapper_38_0_out_id_write;
  assign krnl_partialKnn_wrapper_38_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_38_0___in_38__q0;
  assign in_38_read_addr__din = krnl_partialKnn_wrapper_38_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_38_0_searchSpace_0_read_addr_s_full_n = in_38_read_addr__full_n;
  assign in_38_read_addr__write = krnl_partialKnn_wrapper_38_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_38_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_38_read_data__dout };
  assign krnl_partialKnn_wrapper_38_0_searchSpace_read_data_peek_empty_n = in_38_read_data__empty_n;
  assign krnl_partialKnn_wrapper_38_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_38_read_data__dout };
  assign krnl_partialKnn_wrapper_38_0_searchSpace_0_read_data_s_empty_n = in_38_read_data__empty_n;
  assign in_38_read_data__read = krnl_partialKnn_wrapper_38_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_38_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_38_0___in_38__q0;
  assign in_38_write_addr__din = krnl_partialKnn_wrapper_38_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_38_0_searchSpace_0_write_addr_s_full_n = in_38_write_addr__full_n;
  assign in_38_write_addr__write = krnl_partialKnn_wrapper_38_0_searchSpace_0_write_addr_s_write;
  assign in_38_write_data__din = krnl_partialKnn_wrapper_38_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_38_0_searchSpace_0_write_data_full_n = in_38_write_data__full_n;
  assign in_38_write_data__write = krnl_partialKnn_wrapper_38_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_38_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_38_write_resp__dout };
  assign krnl_partialKnn_wrapper_38_0_searchSpace_write_resp_peek_empty_n = in_38_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_38_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_38_write_resp__dout };
  assign krnl_partialKnn_wrapper_38_0_searchSpace_0_write_resp_s_empty_n = in_38_write_resp__empty_n;
  assign in_38_write_resp__read = krnl_partialKnn_wrapper_38_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_38_0_start_id_0 = 64'd311296;
  assign krnl_partialKnn_wrapper_39_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_39_0__ap_done = krnl_partialKnn_wrapper_39_0_ap_done;
  assign krnl_partialKnn_wrapper_39_0__ap_idle = krnl_partialKnn_wrapper_39_0_ap_idle;
  assign krnl_partialKnn_wrapper_39_0__ap_ready = krnl_partialKnn_wrapper_39_0_ap_ready;
  assign krnl_partialKnn_wrapper_39_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_39_0_ap_start = krnl_partialKnn_wrapper_39_0__ap_start;
  assign out_dist_39__din = krnl_partialKnn_wrapper_39_0_out_dist_din;
  assign krnl_partialKnn_wrapper_39_0_out_dist_full_n = out_dist_39__full_n;
  assign out_dist_39__write = krnl_partialKnn_wrapper_39_0_out_dist_write;
  assign out_id_39__din = krnl_partialKnn_wrapper_39_0_out_id_din;
  assign krnl_partialKnn_wrapper_39_0_out_id_full_n = out_id_39__full_n;
  assign out_id_39__write = krnl_partialKnn_wrapper_39_0_out_id_write;
  assign krnl_partialKnn_wrapper_39_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_39_0___in_39__q0;
  assign in_39_read_addr__din = krnl_partialKnn_wrapper_39_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_39_0_searchSpace_0_read_addr_s_full_n = in_39_read_addr__full_n;
  assign in_39_read_addr__write = krnl_partialKnn_wrapper_39_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_39_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_39_read_data__dout };
  assign krnl_partialKnn_wrapper_39_0_searchSpace_read_data_peek_empty_n = in_39_read_data__empty_n;
  assign krnl_partialKnn_wrapper_39_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_39_read_data__dout };
  assign krnl_partialKnn_wrapper_39_0_searchSpace_0_read_data_s_empty_n = in_39_read_data__empty_n;
  assign in_39_read_data__read = krnl_partialKnn_wrapper_39_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_39_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_39_0___in_39__q0;
  assign in_39_write_addr__din = krnl_partialKnn_wrapper_39_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_39_0_searchSpace_0_write_addr_s_full_n = in_39_write_addr__full_n;
  assign in_39_write_addr__write = krnl_partialKnn_wrapper_39_0_searchSpace_0_write_addr_s_write;
  assign in_39_write_data__din = krnl_partialKnn_wrapper_39_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_39_0_searchSpace_0_write_data_full_n = in_39_write_data__full_n;
  assign in_39_write_data__write = krnl_partialKnn_wrapper_39_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_39_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_39_write_resp__dout };
  assign krnl_partialKnn_wrapper_39_0_searchSpace_write_resp_peek_empty_n = in_39_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_39_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_39_write_resp__dout };
  assign krnl_partialKnn_wrapper_39_0_searchSpace_0_write_resp_s_empty_n = in_39_write_resp__empty_n;
  assign in_39_write_resp__read = krnl_partialKnn_wrapper_39_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_39_0_start_id_0 = 64'd319488;
  assign krnl_partialKnn_wrapper_4_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_4_0__ap_done = krnl_partialKnn_wrapper_4_0_ap_done;
  assign krnl_partialKnn_wrapper_4_0__ap_idle = krnl_partialKnn_wrapper_4_0_ap_idle;
  assign krnl_partialKnn_wrapper_4_0__ap_ready = krnl_partialKnn_wrapper_4_0_ap_ready;
  assign krnl_partialKnn_wrapper_4_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_4_0_ap_start = krnl_partialKnn_wrapper_4_0__ap_start;
  assign out_dist_4__din = krnl_partialKnn_wrapper_4_0_out_dist_din;
  assign krnl_partialKnn_wrapper_4_0_out_dist_full_n = out_dist_4__full_n;
  assign out_dist_4__write = krnl_partialKnn_wrapper_4_0_out_dist_write;
  assign out_id_4__din = krnl_partialKnn_wrapper_4_0_out_id_din;
  assign krnl_partialKnn_wrapper_4_0_out_id_full_n = out_id_4__full_n;
  assign out_id_4__write = krnl_partialKnn_wrapper_4_0_out_id_write;
  assign krnl_partialKnn_wrapper_4_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_4_0___in_4__q0;
  assign in_4_read_addr__din = krnl_partialKnn_wrapper_4_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_4_0_searchSpace_0_read_addr_s_full_n = in_4_read_addr__full_n;
  assign in_4_read_addr__write = krnl_partialKnn_wrapper_4_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_4_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_4_read_data__dout };
  assign krnl_partialKnn_wrapper_4_0_searchSpace_0_read_data_peek_empty_n = in_4_read_data__empty_n;
  assign krnl_partialKnn_wrapper_4_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_4_read_data__dout };
  assign krnl_partialKnn_wrapper_4_0_searchSpace_0_read_data_s_empty_n = in_4_read_data__empty_n;
  assign in_4_read_data__read = krnl_partialKnn_wrapper_4_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_4_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_4_0___in_4__q0;
  assign in_4_write_addr__din = krnl_partialKnn_wrapper_4_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_4_0_searchSpace_0_write_addr_s_full_n = in_4_write_addr__full_n;
  assign in_4_write_addr__write = krnl_partialKnn_wrapper_4_0_searchSpace_0_write_addr_s_write;
  assign in_4_write_data__din = krnl_partialKnn_wrapper_4_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_4_0_searchSpace_0_write_data_full_n = in_4_write_data__full_n;
  assign in_4_write_data__write = krnl_partialKnn_wrapper_4_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_4_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_4_write_resp__dout };
  assign krnl_partialKnn_wrapper_4_0_searchSpace_write_resp_peek_empty_n = in_4_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_4_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_4_write_resp__dout };
  assign krnl_partialKnn_wrapper_4_0_searchSpace_0_write_resp_s_empty_n = in_4_write_resp__empty_n;
  assign in_4_write_resp__read = krnl_partialKnn_wrapper_4_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_4_0_start_id_0 = 64'd32768;
  assign krnl_partialKnn_wrapper_40_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_40_0__ap_done = krnl_partialKnn_wrapper_40_0_ap_done;
  assign krnl_partialKnn_wrapper_40_0__ap_idle = krnl_partialKnn_wrapper_40_0_ap_idle;
  assign krnl_partialKnn_wrapper_40_0__ap_ready = krnl_partialKnn_wrapper_40_0_ap_ready;
  assign krnl_partialKnn_wrapper_40_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_40_0_ap_start = krnl_partialKnn_wrapper_40_0__ap_start;
  assign out_dist_40__din = krnl_partialKnn_wrapper_40_0_out_dist_din;
  assign krnl_partialKnn_wrapper_40_0_out_dist_full_n = out_dist_40__full_n;
  assign out_dist_40__write = krnl_partialKnn_wrapper_40_0_out_dist_write;
  assign out_id_40__din = krnl_partialKnn_wrapper_40_0_out_id_din;
  assign krnl_partialKnn_wrapper_40_0_out_id_full_n = out_id_40__full_n;
  assign out_id_40__write = krnl_partialKnn_wrapper_40_0_out_id_write;
  assign krnl_partialKnn_wrapper_40_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_40_0___in_40__q0;
  assign in_40_read_addr__din = krnl_partialKnn_wrapper_40_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_40_0_searchSpace_0_read_addr_s_full_n = in_40_read_addr__full_n;
  assign in_40_read_addr__write = krnl_partialKnn_wrapper_40_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_40_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_40_read_data__dout };
  assign krnl_partialKnn_wrapper_40_0_searchSpace_read_data_peek_empty_n = in_40_read_data__empty_n;
  assign krnl_partialKnn_wrapper_40_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_40_read_data__dout };
  assign krnl_partialKnn_wrapper_40_0_searchSpace_0_read_data_s_empty_n = in_40_read_data__empty_n;
  assign in_40_read_data__read = krnl_partialKnn_wrapper_40_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_40_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_40_0___in_40__q0;
  assign in_40_write_addr__din = krnl_partialKnn_wrapper_40_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_40_0_searchSpace_0_write_addr_s_full_n = in_40_write_addr__full_n;
  assign in_40_write_addr__write = krnl_partialKnn_wrapper_40_0_searchSpace_0_write_addr_s_write;
  assign in_40_write_data__din = krnl_partialKnn_wrapper_40_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_40_0_searchSpace_0_write_data_full_n = in_40_write_data__full_n;
  assign in_40_write_data__write = krnl_partialKnn_wrapper_40_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_40_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_40_write_resp__dout };
  assign krnl_partialKnn_wrapper_40_0_searchSpace_write_resp_peek_empty_n = in_40_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_40_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_40_write_resp__dout };
  assign krnl_partialKnn_wrapper_40_0_searchSpace_0_write_resp_s_empty_n = in_40_write_resp__empty_n;
  assign in_40_write_resp__read = krnl_partialKnn_wrapper_40_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_40_0_start_id_0 = 64'd327680;
  assign krnl_partialKnn_wrapper_41_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_41_0__ap_done = krnl_partialKnn_wrapper_41_0_ap_done;
  assign krnl_partialKnn_wrapper_41_0__ap_idle = krnl_partialKnn_wrapper_41_0_ap_idle;
  assign krnl_partialKnn_wrapper_41_0__ap_ready = krnl_partialKnn_wrapper_41_0_ap_ready;
  assign krnl_partialKnn_wrapper_41_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_41_0_ap_start = krnl_partialKnn_wrapper_41_0__ap_start;
  assign out_dist_41__din = krnl_partialKnn_wrapper_41_0_out_dist_din;
  assign krnl_partialKnn_wrapper_41_0_out_dist_full_n = out_dist_41__full_n;
  assign out_dist_41__write = krnl_partialKnn_wrapper_41_0_out_dist_write;
  assign out_id_41__din = krnl_partialKnn_wrapper_41_0_out_id_din;
  assign krnl_partialKnn_wrapper_41_0_out_id_full_n = out_id_41__full_n;
  assign out_id_41__write = krnl_partialKnn_wrapper_41_0_out_id_write;
  assign krnl_partialKnn_wrapper_41_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_41_0___in_41__q0;
  assign in_41_read_addr__din = krnl_partialKnn_wrapper_41_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_41_0_searchSpace_0_read_addr_s_full_n = in_41_read_addr__full_n;
  assign in_41_read_addr__write = krnl_partialKnn_wrapper_41_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_41_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_41_read_data__dout };
  assign krnl_partialKnn_wrapper_41_0_searchSpace_read_data_peek_empty_n = in_41_read_data__empty_n;
  assign krnl_partialKnn_wrapper_41_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_41_read_data__dout };
  assign krnl_partialKnn_wrapper_41_0_searchSpace_0_read_data_s_empty_n = in_41_read_data__empty_n;
  assign in_41_read_data__read = krnl_partialKnn_wrapper_41_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_41_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_41_0___in_41__q0;
  assign in_41_write_addr__din = krnl_partialKnn_wrapper_41_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_41_0_searchSpace_0_write_addr_s_full_n = in_41_write_addr__full_n;
  assign in_41_write_addr__write = krnl_partialKnn_wrapper_41_0_searchSpace_0_write_addr_s_write;
  assign in_41_write_data__din = krnl_partialKnn_wrapper_41_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_41_0_searchSpace_0_write_data_full_n = in_41_write_data__full_n;
  assign in_41_write_data__write = krnl_partialKnn_wrapper_41_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_41_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_41_write_resp__dout };
  assign krnl_partialKnn_wrapper_41_0_searchSpace_write_resp_peek_empty_n = in_41_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_41_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_41_write_resp__dout };
  assign krnl_partialKnn_wrapper_41_0_searchSpace_0_write_resp_s_empty_n = in_41_write_resp__empty_n;
  assign in_41_write_resp__read = krnl_partialKnn_wrapper_41_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_41_0_start_id_0 = 64'd335872;
  assign krnl_partialKnn_wrapper_42_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_42_0__ap_done = krnl_partialKnn_wrapper_42_0_ap_done;
  assign krnl_partialKnn_wrapper_42_0__ap_idle = krnl_partialKnn_wrapper_42_0_ap_idle;
  assign krnl_partialKnn_wrapper_42_0__ap_ready = krnl_partialKnn_wrapper_42_0_ap_ready;
  assign krnl_partialKnn_wrapper_42_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_42_0_ap_start = krnl_partialKnn_wrapper_42_0__ap_start;
  assign out_dist_42__din = krnl_partialKnn_wrapper_42_0_out_dist_din;
  assign krnl_partialKnn_wrapper_42_0_out_dist_full_n = out_dist_42__full_n;
  assign out_dist_42__write = krnl_partialKnn_wrapper_42_0_out_dist_write;
  assign out_id_42__din = krnl_partialKnn_wrapper_42_0_out_id_din;
  assign krnl_partialKnn_wrapper_42_0_out_id_full_n = out_id_42__full_n;
  assign out_id_42__write = krnl_partialKnn_wrapper_42_0_out_id_write;
  assign krnl_partialKnn_wrapper_42_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_42_0___in_42__q0;
  assign in_42_read_addr__din = krnl_partialKnn_wrapper_42_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_42_0_searchSpace_0_read_addr_s_full_n = in_42_read_addr__full_n;
  assign in_42_read_addr__write = krnl_partialKnn_wrapper_42_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_42_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_42_read_data__dout };
  assign krnl_partialKnn_wrapper_42_0_searchSpace_read_data_peek_empty_n = in_42_read_data__empty_n;
  assign krnl_partialKnn_wrapper_42_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_42_read_data__dout };
  assign krnl_partialKnn_wrapper_42_0_searchSpace_0_read_data_s_empty_n = in_42_read_data__empty_n;
  assign in_42_read_data__read = krnl_partialKnn_wrapper_42_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_42_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_42_0___in_42__q0;
  assign in_42_write_addr__din = krnl_partialKnn_wrapper_42_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_42_0_searchSpace_0_write_addr_s_full_n = in_42_write_addr__full_n;
  assign in_42_write_addr__write = krnl_partialKnn_wrapper_42_0_searchSpace_0_write_addr_s_write;
  assign in_42_write_data__din = krnl_partialKnn_wrapper_42_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_42_0_searchSpace_0_write_data_full_n = in_42_write_data__full_n;
  assign in_42_write_data__write = krnl_partialKnn_wrapper_42_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_42_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_42_write_resp__dout };
  assign krnl_partialKnn_wrapper_42_0_searchSpace_write_resp_peek_empty_n = in_42_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_42_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_42_write_resp__dout };
  assign krnl_partialKnn_wrapper_42_0_searchSpace_0_write_resp_s_empty_n = in_42_write_resp__empty_n;
  assign in_42_write_resp__read = krnl_partialKnn_wrapper_42_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_42_0_start_id_0 = 64'd344064;
  assign krnl_partialKnn_wrapper_43_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_43_0__ap_done = krnl_partialKnn_wrapper_43_0_ap_done;
  assign krnl_partialKnn_wrapper_43_0__ap_idle = krnl_partialKnn_wrapper_43_0_ap_idle;
  assign krnl_partialKnn_wrapper_43_0__ap_ready = krnl_partialKnn_wrapper_43_0_ap_ready;
  assign krnl_partialKnn_wrapper_43_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_43_0_ap_start = krnl_partialKnn_wrapper_43_0__ap_start;
  assign out_dist_43__din = krnl_partialKnn_wrapper_43_0_out_dist_din;
  assign krnl_partialKnn_wrapper_43_0_out_dist_full_n = out_dist_43__full_n;
  assign out_dist_43__write = krnl_partialKnn_wrapper_43_0_out_dist_write;
  assign out_id_43__din = krnl_partialKnn_wrapper_43_0_out_id_din;
  assign krnl_partialKnn_wrapper_43_0_out_id_full_n = out_id_43__full_n;
  assign out_id_43__write = krnl_partialKnn_wrapper_43_0_out_id_write;
  assign krnl_partialKnn_wrapper_43_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_43_0___in_43__q0;
  assign in_43_read_addr__din = krnl_partialKnn_wrapper_43_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_43_0_searchSpace_0_read_addr_s_full_n = in_43_read_addr__full_n;
  assign in_43_read_addr__write = krnl_partialKnn_wrapper_43_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_43_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_43_read_data__dout };
  assign krnl_partialKnn_wrapper_43_0_searchSpace_read_data_peek_empty_n = in_43_read_data__empty_n;
  assign krnl_partialKnn_wrapper_43_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_43_read_data__dout };
  assign krnl_partialKnn_wrapper_43_0_searchSpace_0_read_data_s_empty_n = in_43_read_data__empty_n;
  assign in_43_read_data__read = krnl_partialKnn_wrapper_43_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_43_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_43_0___in_43__q0;
  assign in_43_write_addr__din = krnl_partialKnn_wrapper_43_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_43_0_searchSpace_0_write_addr_s_full_n = in_43_write_addr__full_n;
  assign in_43_write_addr__write = krnl_partialKnn_wrapper_43_0_searchSpace_0_write_addr_s_write;
  assign in_43_write_data__din = krnl_partialKnn_wrapper_43_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_43_0_searchSpace_0_write_data_full_n = in_43_write_data__full_n;
  assign in_43_write_data__write = krnl_partialKnn_wrapper_43_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_43_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_43_write_resp__dout };
  assign krnl_partialKnn_wrapper_43_0_searchSpace_write_resp_peek_empty_n = in_43_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_43_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_43_write_resp__dout };
  assign krnl_partialKnn_wrapper_43_0_searchSpace_0_write_resp_s_empty_n = in_43_write_resp__empty_n;
  assign in_43_write_resp__read = krnl_partialKnn_wrapper_43_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_43_0_start_id_0 = 64'd352256;
  assign krnl_partialKnn_wrapper_44_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_44_0__ap_done = krnl_partialKnn_wrapper_44_0_ap_done;
  assign krnl_partialKnn_wrapper_44_0__ap_idle = krnl_partialKnn_wrapper_44_0_ap_idle;
  assign krnl_partialKnn_wrapper_44_0__ap_ready = krnl_partialKnn_wrapper_44_0_ap_ready;
  assign krnl_partialKnn_wrapper_44_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_44_0_ap_start = krnl_partialKnn_wrapper_44_0__ap_start;
  assign out_dist_44__din = krnl_partialKnn_wrapper_44_0_out_dist_din;
  assign krnl_partialKnn_wrapper_44_0_out_dist_full_n = out_dist_44__full_n;
  assign out_dist_44__write = krnl_partialKnn_wrapper_44_0_out_dist_write;
  assign out_id_44__din = krnl_partialKnn_wrapper_44_0_out_id_din;
  assign krnl_partialKnn_wrapper_44_0_out_id_full_n = out_id_44__full_n;
  assign out_id_44__write = krnl_partialKnn_wrapper_44_0_out_id_write;
  assign krnl_partialKnn_wrapper_44_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_44_0___in_44__q0;
  assign in_44_read_addr__din = krnl_partialKnn_wrapper_44_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_44_0_searchSpace_0_read_addr_s_full_n = in_44_read_addr__full_n;
  assign in_44_read_addr__write = krnl_partialKnn_wrapper_44_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_44_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_44_read_data__dout };
  assign krnl_partialKnn_wrapper_44_0_searchSpace_read_data_peek_empty_n = in_44_read_data__empty_n;
  assign krnl_partialKnn_wrapper_44_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_44_read_data__dout };
  assign krnl_partialKnn_wrapper_44_0_searchSpace_0_read_data_s_empty_n = in_44_read_data__empty_n;
  assign in_44_read_data__read = krnl_partialKnn_wrapper_44_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_44_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_44_0___in_44__q0;
  assign in_44_write_addr__din = krnl_partialKnn_wrapper_44_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_44_0_searchSpace_0_write_addr_s_full_n = in_44_write_addr__full_n;
  assign in_44_write_addr__write = krnl_partialKnn_wrapper_44_0_searchSpace_0_write_addr_s_write;
  assign in_44_write_data__din = krnl_partialKnn_wrapper_44_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_44_0_searchSpace_0_write_data_full_n = in_44_write_data__full_n;
  assign in_44_write_data__write = krnl_partialKnn_wrapper_44_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_44_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_44_write_resp__dout };
  assign krnl_partialKnn_wrapper_44_0_searchSpace_write_resp_peek_empty_n = in_44_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_44_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_44_write_resp__dout };
  assign krnl_partialKnn_wrapper_44_0_searchSpace_0_write_resp_s_empty_n = in_44_write_resp__empty_n;
  assign in_44_write_resp__read = krnl_partialKnn_wrapper_44_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_44_0_start_id_0 = 64'd360448;
  assign krnl_partialKnn_wrapper_45_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_45_0__ap_done = krnl_partialKnn_wrapper_45_0_ap_done;
  assign krnl_partialKnn_wrapper_45_0__ap_idle = krnl_partialKnn_wrapper_45_0_ap_idle;
  assign krnl_partialKnn_wrapper_45_0__ap_ready = krnl_partialKnn_wrapper_45_0_ap_ready;
  assign krnl_partialKnn_wrapper_45_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_45_0_ap_start = krnl_partialKnn_wrapper_45_0__ap_start;
  assign out_dist_45__din = krnl_partialKnn_wrapper_45_0_out_dist_din;
  assign krnl_partialKnn_wrapper_45_0_out_dist_full_n = out_dist_45__full_n;
  assign out_dist_45__write = krnl_partialKnn_wrapper_45_0_out_dist_write;
  assign out_id_45__din = krnl_partialKnn_wrapper_45_0_out_id_din;
  assign krnl_partialKnn_wrapper_45_0_out_id_full_n = out_id_45__full_n;
  assign out_id_45__write = krnl_partialKnn_wrapper_45_0_out_id_write;
  assign krnl_partialKnn_wrapper_45_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_45_0___in_45__q0;
  assign in_45_read_addr__din = krnl_partialKnn_wrapper_45_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_45_0_searchSpace_0_read_addr_s_full_n = in_45_read_addr__full_n;
  assign in_45_read_addr__write = krnl_partialKnn_wrapper_45_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_45_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_45_read_data__dout };
  assign krnl_partialKnn_wrapper_45_0_searchSpace_read_data_peek_empty_n = in_45_read_data__empty_n;
  assign krnl_partialKnn_wrapper_45_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_45_read_data__dout };
  assign krnl_partialKnn_wrapper_45_0_searchSpace_0_read_data_s_empty_n = in_45_read_data__empty_n;
  assign in_45_read_data__read = krnl_partialKnn_wrapper_45_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_45_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_45_0___in_45__q0;
  assign in_45_write_addr__din = krnl_partialKnn_wrapper_45_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_45_0_searchSpace_0_write_addr_s_full_n = in_45_write_addr__full_n;
  assign in_45_write_addr__write = krnl_partialKnn_wrapper_45_0_searchSpace_0_write_addr_s_write;
  assign in_45_write_data__din = krnl_partialKnn_wrapper_45_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_45_0_searchSpace_0_write_data_full_n = in_45_write_data__full_n;
  assign in_45_write_data__write = krnl_partialKnn_wrapper_45_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_45_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_45_write_resp__dout };
  assign krnl_partialKnn_wrapper_45_0_searchSpace_write_resp_peek_empty_n = in_45_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_45_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_45_write_resp__dout };
  assign krnl_partialKnn_wrapper_45_0_searchSpace_0_write_resp_s_empty_n = in_45_write_resp__empty_n;
  assign in_45_write_resp__read = krnl_partialKnn_wrapper_45_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_45_0_start_id_0 = 64'd368640;
  assign krnl_partialKnn_wrapper_46_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_46_0__ap_done = krnl_partialKnn_wrapper_46_0_ap_done;
  assign krnl_partialKnn_wrapper_46_0__ap_idle = krnl_partialKnn_wrapper_46_0_ap_idle;
  assign krnl_partialKnn_wrapper_46_0__ap_ready = krnl_partialKnn_wrapper_46_0_ap_ready;
  assign krnl_partialKnn_wrapper_46_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_46_0_ap_start = krnl_partialKnn_wrapper_46_0__ap_start;
  assign out_dist_46__din = krnl_partialKnn_wrapper_46_0_out_dist_din;
  assign krnl_partialKnn_wrapper_46_0_out_dist_full_n = out_dist_46__full_n;
  assign out_dist_46__write = krnl_partialKnn_wrapper_46_0_out_dist_write;
  assign out_id_46__din = krnl_partialKnn_wrapper_46_0_out_id_din;
  assign krnl_partialKnn_wrapper_46_0_out_id_full_n = out_id_46__full_n;
  assign out_id_46__write = krnl_partialKnn_wrapper_46_0_out_id_write;
  assign krnl_partialKnn_wrapper_46_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_46_0___in_46__q0;
  assign in_46_read_addr__din = krnl_partialKnn_wrapper_46_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_46_0_searchSpace_0_read_addr_s_full_n = in_46_read_addr__full_n;
  assign in_46_read_addr__write = krnl_partialKnn_wrapper_46_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_46_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_46_read_data__dout };
  assign krnl_partialKnn_wrapper_46_0_searchSpace_read_data_peek_empty_n = in_46_read_data__empty_n;
  assign krnl_partialKnn_wrapper_46_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_46_read_data__dout };
  assign krnl_partialKnn_wrapper_46_0_searchSpace_0_read_data_s_empty_n = in_46_read_data__empty_n;
  assign in_46_read_data__read = krnl_partialKnn_wrapper_46_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_46_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_46_0___in_46__q0;
  assign in_46_write_addr__din = krnl_partialKnn_wrapper_46_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_46_0_searchSpace_0_write_addr_s_full_n = in_46_write_addr__full_n;
  assign in_46_write_addr__write = krnl_partialKnn_wrapper_46_0_searchSpace_0_write_addr_s_write;
  assign in_46_write_data__din = krnl_partialKnn_wrapper_46_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_46_0_searchSpace_0_write_data_full_n = in_46_write_data__full_n;
  assign in_46_write_data__write = krnl_partialKnn_wrapper_46_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_46_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_46_write_resp__dout };
  assign krnl_partialKnn_wrapper_46_0_searchSpace_write_resp_peek_empty_n = in_46_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_46_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_46_write_resp__dout };
  assign krnl_partialKnn_wrapper_46_0_searchSpace_0_write_resp_s_empty_n = in_46_write_resp__empty_n;
  assign in_46_write_resp__read = krnl_partialKnn_wrapper_46_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_46_0_start_id_0 = 64'd376832;
  assign krnl_partialKnn_wrapper_47_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_47_0__ap_done = krnl_partialKnn_wrapper_47_0_ap_done;
  assign krnl_partialKnn_wrapper_47_0__ap_idle = krnl_partialKnn_wrapper_47_0_ap_idle;
  assign krnl_partialKnn_wrapper_47_0__ap_ready = krnl_partialKnn_wrapper_47_0_ap_ready;
  assign krnl_partialKnn_wrapper_47_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_47_0_ap_start = krnl_partialKnn_wrapper_47_0__ap_start;
  assign out_dist_47__din = krnl_partialKnn_wrapper_47_0_out_dist_din;
  assign krnl_partialKnn_wrapper_47_0_out_dist_full_n = out_dist_47__full_n;
  assign out_dist_47__write = krnl_partialKnn_wrapper_47_0_out_dist_write;
  assign out_id_47__din = krnl_partialKnn_wrapper_47_0_out_id_din;
  assign krnl_partialKnn_wrapper_47_0_out_id_full_n = out_id_47__full_n;
  assign out_id_47__write = krnl_partialKnn_wrapper_47_0_out_id_write;
  assign krnl_partialKnn_wrapper_47_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_47_0___in_47__q0;
  assign in_47_read_addr__din = krnl_partialKnn_wrapper_47_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_47_0_searchSpace_0_read_addr_s_full_n = in_47_read_addr__full_n;
  assign in_47_read_addr__write = krnl_partialKnn_wrapper_47_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_47_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_47_read_data__dout };
  assign krnl_partialKnn_wrapper_47_0_searchSpace_read_data_peek_empty_n = in_47_read_data__empty_n;
  assign krnl_partialKnn_wrapper_47_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_47_read_data__dout };
  assign krnl_partialKnn_wrapper_47_0_searchSpace_0_read_data_s_empty_n = in_47_read_data__empty_n;
  assign in_47_read_data__read = krnl_partialKnn_wrapper_47_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_47_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_47_0___in_47__q0;
  assign in_47_write_addr__din = krnl_partialKnn_wrapper_47_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_47_0_searchSpace_0_write_addr_s_full_n = in_47_write_addr__full_n;
  assign in_47_write_addr__write = krnl_partialKnn_wrapper_47_0_searchSpace_0_write_addr_s_write;
  assign in_47_write_data__din = krnl_partialKnn_wrapper_47_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_47_0_searchSpace_0_write_data_full_n = in_47_write_data__full_n;
  assign in_47_write_data__write = krnl_partialKnn_wrapper_47_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_47_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_47_write_resp__dout };
  assign krnl_partialKnn_wrapper_47_0_searchSpace_write_resp_peek_empty_n = in_47_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_47_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_47_write_resp__dout };
  assign krnl_partialKnn_wrapper_47_0_searchSpace_0_write_resp_s_empty_n = in_47_write_resp__empty_n;
  assign in_47_write_resp__read = krnl_partialKnn_wrapper_47_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_47_0_start_id_0 = 64'd385024;
  assign krnl_partialKnn_wrapper_48_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_48_0__ap_done = krnl_partialKnn_wrapper_48_0_ap_done;
  assign krnl_partialKnn_wrapper_48_0__ap_idle = krnl_partialKnn_wrapper_48_0_ap_idle;
  assign krnl_partialKnn_wrapper_48_0__ap_ready = krnl_partialKnn_wrapper_48_0_ap_ready;
  assign krnl_partialKnn_wrapper_48_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_48_0_ap_start = krnl_partialKnn_wrapper_48_0__ap_start;
  assign out_dist_48__din = krnl_partialKnn_wrapper_48_0_out_dist_din;
  assign krnl_partialKnn_wrapper_48_0_out_dist_full_n = out_dist_48__full_n;
  assign out_dist_48__write = krnl_partialKnn_wrapper_48_0_out_dist_write;
  assign out_id_48__din = krnl_partialKnn_wrapper_48_0_out_id_din;
  assign krnl_partialKnn_wrapper_48_0_out_id_full_n = out_id_48__full_n;
  assign out_id_48__write = krnl_partialKnn_wrapper_48_0_out_id_write;
  assign krnl_partialKnn_wrapper_48_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_48_0___in_48__q0;
  assign in_48_read_addr__din = krnl_partialKnn_wrapper_48_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_48_0_searchSpace_0_read_addr_s_full_n = in_48_read_addr__full_n;
  assign in_48_read_addr__write = krnl_partialKnn_wrapper_48_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_48_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_48_read_data__dout };
  assign krnl_partialKnn_wrapper_48_0_searchSpace_read_data_peek_empty_n = in_48_read_data__empty_n;
  assign krnl_partialKnn_wrapper_48_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_48_read_data__dout };
  assign krnl_partialKnn_wrapper_48_0_searchSpace_0_read_data_s_empty_n = in_48_read_data__empty_n;
  assign in_48_read_data__read = krnl_partialKnn_wrapper_48_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_48_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_48_0___in_48__q0;
  assign in_48_write_addr__din = krnl_partialKnn_wrapper_48_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_48_0_searchSpace_0_write_addr_s_full_n = in_48_write_addr__full_n;
  assign in_48_write_addr__write = krnl_partialKnn_wrapper_48_0_searchSpace_0_write_addr_s_write;
  assign in_48_write_data__din = krnl_partialKnn_wrapper_48_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_48_0_searchSpace_0_write_data_full_n = in_48_write_data__full_n;
  assign in_48_write_data__write = krnl_partialKnn_wrapper_48_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_48_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_48_write_resp__dout };
  assign krnl_partialKnn_wrapper_48_0_searchSpace_write_resp_peek_empty_n = in_48_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_48_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_48_write_resp__dout };
  assign krnl_partialKnn_wrapper_48_0_searchSpace_0_write_resp_s_empty_n = in_48_write_resp__empty_n;
  assign in_48_write_resp__read = krnl_partialKnn_wrapper_48_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_48_0_start_id_0 = 64'd393216;
  assign krnl_partialKnn_wrapper_49_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_49_0__ap_done = krnl_partialKnn_wrapper_49_0_ap_done;
  assign krnl_partialKnn_wrapper_49_0__ap_idle = krnl_partialKnn_wrapper_49_0_ap_idle;
  assign krnl_partialKnn_wrapper_49_0__ap_ready = krnl_partialKnn_wrapper_49_0_ap_ready;
  assign krnl_partialKnn_wrapper_49_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_49_0_ap_start = krnl_partialKnn_wrapper_49_0__ap_start;
  assign out_dist_49__din = krnl_partialKnn_wrapper_49_0_out_dist_din;
  assign krnl_partialKnn_wrapper_49_0_out_dist_full_n = out_dist_49__full_n;
  assign out_dist_49__write = krnl_partialKnn_wrapper_49_0_out_dist_write;
  assign out_id_49__din = krnl_partialKnn_wrapper_49_0_out_id_din;
  assign krnl_partialKnn_wrapper_49_0_out_id_full_n = out_id_49__full_n;
  assign out_id_49__write = krnl_partialKnn_wrapper_49_0_out_id_write;
  assign krnl_partialKnn_wrapper_49_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_49_0___in_49__q0;
  assign in_49_read_addr__din = krnl_partialKnn_wrapper_49_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_49_0_searchSpace_0_read_addr_s_full_n = in_49_read_addr__full_n;
  assign in_49_read_addr__write = krnl_partialKnn_wrapper_49_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_49_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_49_read_data__dout };
  assign krnl_partialKnn_wrapper_49_0_searchSpace_read_data_peek_empty_n = in_49_read_data__empty_n;
  assign krnl_partialKnn_wrapper_49_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_49_read_data__dout };
  assign krnl_partialKnn_wrapper_49_0_searchSpace_0_read_data_s_empty_n = in_49_read_data__empty_n;
  assign in_49_read_data__read = krnl_partialKnn_wrapper_49_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_49_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_49_0___in_49__q0;
  assign in_49_write_addr__din = krnl_partialKnn_wrapper_49_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_49_0_searchSpace_0_write_addr_s_full_n = in_49_write_addr__full_n;
  assign in_49_write_addr__write = krnl_partialKnn_wrapper_49_0_searchSpace_0_write_addr_s_write;
  assign in_49_write_data__din = krnl_partialKnn_wrapper_49_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_49_0_searchSpace_0_write_data_full_n = in_49_write_data__full_n;
  assign in_49_write_data__write = krnl_partialKnn_wrapper_49_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_49_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_49_write_resp__dout };
  assign krnl_partialKnn_wrapper_49_0_searchSpace_write_resp_peek_empty_n = in_49_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_49_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_49_write_resp__dout };
  assign krnl_partialKnn_wrapper_49_0_searchSpace_0_write_resp_s_empty_n = in_49_write_resp__empty_n;
  assign in_49_write_resp__read = krnl_partialKnn_wrapper_49_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_49_0_start_id_0 = 64'd401408;
  assign krnl_partialKnn_wrapper_5_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_5_0__ap_done = krnl_partialKnn_wrapper_5_0_ap_done;
  assign krnl_partialKnn_wrapper_5_0__ap_idle = krnl_partialKnn_wrapper_5_0_ap_idle;
  assign krnl_partialKnn_wrapper_5_0__ap_ready = krnl_partialKnn_wrapper_5_0_ap_ready;
  assign krnl_partialKnn_wrapper_5_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_5_0_ap_start = krnl_partialKnn_wrapper_5_0__ap_start;
  assign out_dist_5__din = krnl_partialKnn_wrapper_5_0_out_dist_din;
  assign krnl_partialKnn_wrapper_5_0_out_dist_full_n = out_dist_5__full_n;
  assign out_dist_5__write = krnl_partialKnn_wrapper_5_0_out_dist_write;
  assign out_id_5__din = krnl_partialKnn_wrapper_5_0_out_id_din;
  assign krnl_partialKnn_wrapper_5_0_out_id_full_n = out_id_5__full_n;
  assign out_id_5__write = krnl_partialKnn_wrapper_5_0_out_id_write;
  assign krnl_partialKnn_wrapper_5_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_5_0___in_5__q0;
  assign in_5_read_addr__din = krnl_partialKnn_wrapper_5_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_5_0_searchSpace_0_read_addr_s_full_n = in_5_read_addr__full_n;
  assign in_5_read_addr__write = krnl_partialKnn_wrapper_5_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_5_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_5_read_data__dout };
  assign krnl_partialKnn_wrapper_5_0_searchSpace_0_read_data_peek_empty_n = in_5_read_data__empty_n;
  assign krnl_partialKnn_wrapper_5_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_5_read_data__dout };
  assign krnl_partialKnn_wrapper_5_0_searchSpace_0_read_data_s_empty_n = in_5_read_data__empty_n;
  assign in_5_read_data__read = krnl_partialKnn_wrapper_5_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_5_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_5_0___in_5__q0;
  assign in_5_write_addr__din = krnl_partialKnn_wrapper_5_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_5_0_searchSpace_0_write_addr_s_full_n = in_5_write_addr__full_n;
  assign in_5_write_addr__write = krnl_partialKnn_wrapper_5_0_searchSpace_0_write_addr_s_write;
  assign in_5_write_data__din = krnl_partialKnn_wrapper_5_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_5_0_searchSpace_0_write_data_full_n = in_5_write_data__full_n;
  assign in_5_write_data__write = krnl_partialKnn_wrapper_5_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_5_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_5_write_resp__dout };
  assign krnl_partialKnn_wrapper_5_0_searchSpace_write_resp_peek_empty_n = in_5_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_5_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_5_write_resp__dout };
  assign krnl_partialKnn_wrapper_5_0_searchSpace_0_write_resp_s_empty_n = in_5_write_resp__empty_n;
  assign in_5_write_resp__read = krnl_partialKnn_wrapper_5_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_5_0_start_id_0 = 64'd40960;
  assign krnl_partialKnn_wrapper_50_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_50_0__ap_done = krnl_partialKnn_wrapper_50_0_ap_done;
  assign krnl_partialKnn_wrapper_50_0__ap_idle = krnl_partialKnn_wrapper_50_0_ap_idle;
  assign krnl_partialKnn_wrapper_50_0__ap_ready = krnl_partialKnn_wrapper_50_0_ap_ready;
  assign krnl_partialKnn_wrapper_50_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_50_0_ap_start = krnl_partialKnn_wrapper_50_0__ap_start;
  assign out_dist_50__din = krnl_partialKnn_wrapper_50_0_out_dist_din;
  assign krnl_partialKnn_wrapper_50_0_out_dist_full_n = out_dist_50__full_n;
  assign out_dist_50__write = krnl_partialKnn_wrapper_50_0_out_dist_write;
  assign out_id_50__din = krnl_partialKnn_wrapper_50_0_out_id_din;
  assign krnl_partialKnn_wrapper_50_0_out_id_full_n = out_id_50__full_n;
  assign out_id_50__write = krnl_partialKnn_wrapper_50_0_out_id_write;
  assign krnl_partialKnn_wrapper_50_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_50_0___in_50__q0;
  assign in_50_read_addr__din = krnl_partialKnn_wrapper_50_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_50_0_searchSpace_0_read_addr_s_full_n = in_50_read_addr__full_n;
  assign in_50_read_addr__write = krnl_partialKnn_wrapper_50_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_50_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_50_read_data__dout };
  assign krnl_partialKnn_wrapper_50_0_searchSpace_read_data_peek_empty_n = in_50_read_data__empty_n;
  assign krnl_partialKnn_wrapper_50_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_50_read_data__dout };
  assign krnl_partialKnn_wrapper_50_0_searchSpace_0_read_data_s_empty_n = in_50_read_data__empty_n;
  assign in_50_read_data__read = krnl_partialKnn_wrapper_50_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_50_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_50_0___in_50__q0;
  assign in_50_write_addr__din = krnl_partialKnn_wrapper_50_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_50_0_searchSpace_0_write_addr_s_full_n = in_50_write_addr__full_n;
  assign in_50_write_addr__write = krnl_partialKnn_wrapper_50_0_searchSpace_0_write_addr_s_write;
  assign in_50_write_data__din = krnl_partialKnn_wrapper_50_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_50_0_searchSpace_0_write_data_full_n = in_50_write_data__full_n;
  assign in_50_write_data__write = krnl_partialKnn_wrapper_50_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_50_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_50_write_resp__dout };
  assign krnl_partialKnn_wrapper_50_0_searchSpace_write_resp_peek_empty_n = in_50_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_50_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_50_write_resp__dout };
  assign krnl_partialKnn_wrapper_50_0_searchSpace_0_write_resp_s_empty_n = in_50_write_resp__empty_n;
  assign in_50_write_resp__read = krnl_partialKnn_wrapper_50_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_50_0_start_id_0 = 64'd409600;
  assign krnl_partialKnn_wrapper_51_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_51_0__ap_done = krnl_partialKnn_wrapper_51_0_ap_done;
  assign krnl_partialKnn_wrapper_51_0__ap_idle = krnl_partialKnn_wrapper_51_0_ap_idle;
  assign krnl_partialKnn_wrapper_51_0__ap_ready = krnl_partialKnn_wrapper_51_0_ap_ready;
  assign krnl_partialKnn_wrapper_51_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_51_0_ap_start = krnl_partialKnn_wrapper_51_0__ap_start;
  assign out_dist_51__din = krnl_partialKnn_wrapper_51_0_out_dist_din;
  assign krnl_partialKnn_wrapper_51_0_out_dist_full_n = out_dist_51__full_n;
  assign out_dist_51__write = krnl_partialKnn_wrapper_51_0_out_dist_write;
  assign out_id_51__din = krnl_partialKnn_wrapper_51_0_out_id_din;
  assign krnl_partialKnn_wrapper_51_0_out_id_full_n = out_id_51__full_n;
  assign out_id_51__write = krnl_partialKnn_wrapper_51_0_out_id_write;
  assign krnl_partialKnn_wrapper_51_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_51_0___in_51__q0;
  assign in_51_read_addr__din = krnl_partialKnn_wrapper_51_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_51_0_searchSpace_0_read_addr_s_full_n = in_51_read_addr__full_n;
  assign in_51_read_addr__write = krnl_partialKnn_wrapper_51_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_51_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_51_read_data__dout };
  assign krnl_partialKnn_wrapper_51_0_searchSpace_read_data_peek_empty_n = in_51_read_data__empty_n;
  assign krnl_partialKnn_wrapper_51_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_51_read_data__dout };
  assign krnl_partialKnn_wrapper_51_0_searchSpace_0_read_data_s_empty_n = in_51_read_data__empty_n;
  assign in_51_read_data__read = krnl_partialKnn_wrapper_51_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_51_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_51_0___in_51__q0;
  assign in_51_write_addr__din = krnl_partialKnn_wrapper_51_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_51_0_searchSpace_0_write_addr_s_full_n = in_51_write_addr__full_n;
  assign in_51_write_addr__write = krnl_partialKnn_wrapper_51_0_searchSpace_0_write_addr_s_write;
  assign in_51_write_data__din = krnl_partialKnn_wrapper_51_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_51_0_searchSpace_0_write_data_full_n = in_51_write_data__full_n;
  assign in_51_write_data__write = krnl_partialKnn_wrapper_51_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_51_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_51_write_resp__dout };
  assign krnl_partialKnn_wrapper_51_0_searchSpace_write_resp_peek_empty_n = in_51_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_51_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_51_write_resp__dout };
  assign krnl_partialKnn_wrapper_51_0_searchSpace_0_write_resp_s_empty_n = in_51_write_resp__empty_n;
  assign in_51_write_resp__read = krnl_partialKnn_wrapper_51_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_51_0_start_id_0 = 64'd417792;
  assign krnl_partialKnn_wrapper_52_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_52_0__ap_done = krnl_partialKnn_wrapper_52_0_ap_done;
  assign krnl_partialKnn_wrapper_52_0__ap_idle = krnl_partialKnn_wrapper_52_0_ap_idle;
  assign krnl_partialKnn_wrapper_52_0__ap_ready = krnl_partialKnn_wrapper_52_0_ap_ready;
  assign krnl_partialKnn_wrapper_52_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_52_0_ap_start = krnl_partialKnn_wrapper_52_0__ap_start;
  assign out_dist_52__din = krnl_partialKnn_wrapper_52_0_out_dist_din;
  assign krnl_partialKnn_wrapper_52_0_out_dist_full_n = out_dist_52__full_n;
  assign out_dist_52__write = krnl_partialKnn_wrapper_52_0_out_dist_write;
  assign out_id_52__din = krnl_partialKnn_wrapper_52_0_out_id_din;
  assign krnl_partialKnn_wrapper_52_0_out_id_full_n = out_id_52__full_n;
  assign out_id_52__write = krnl_partialKnn_wrapper_52_0_out_id_write;
  assign krnl_partialKnn_wrapper_52_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_52_0___in_52__q0;
  assign in_52_read_addr__din = krnl_partialKnn_wrapper_52_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_52_0_searchSpace_0_read_addr_s_full_n = in_52_read_addr__full_n;
  assign in_52_read_addr__write = krnl_partialKnn_wrapper_52_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_52_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_52_read_data__dout };
  assign krnl_partialKnn_wrapper_52_0_searchSpace_read_data_peek_empty_n = in_52_read_data__empty_n;
  assign krnl_partialKnn_wrapper_52_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_52_read_data__dout };
  assign krnl_partialKnn_wrapper_52_0_searchSpace_0_read_data_s_empty_n = in_52_read_data__empty_n;
  assign in_52_read_data__read = krnl_partialKnn_wrapper_52_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_52_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_52_0___in_52__q0;
  assign in_52_write_addr__din = krnl_partialKnn_wrapper_52_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_52_0_searchSpace_0_write_addr_s_full_n = in_52_write_addr__full_n;
  assign in_52_write_addr__write = krnl_partialKnn_wrapper_52_0_searchSpace_0_write_addr_s_write;
  assign in_52_write_data__din = krnl_partialKnn_wrapper_52_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_52_0_searchSpace_0_write_data_full_n = in_52_write_data__full_n;
  assign in_52_write_data__write = krnl_partialKnn_wrapper_52_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_52_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_52_write_resp__dout };
  assign krnl_partialKnn_wrapper_52_0_searchSpace_write_resp_peek_empty_n = in_52_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_52_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_52_write_resp__dout };
  assign krnl_partialKnn_wrapper_52_0_searchSpace_0_write_resp_s_empty_n = in_52_write_resp__empty_n;
  assign in_52_write_resp__read = krnl_partialKnn_wrapper_52_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_52_0_start_id_0 = 64'd425984;
  assign krnl_partialKnn_wrapper_53_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_53_0__ap_done = krnl_partialKnn_wrapper_53_0_ap_done;
  assign krnl_partialKnn_wrapper_53_0__ap_idle = krnl_partialKnn_wrapper_53_0_ap_idle;
  assign krnl_partialKnn_wrapper_53_0__ap_ready = krnl_partialKnn_wrapper_53_0_ap_ready;
  assign krnl_partialKnn_wrapper_53_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_53_0_ap_start = krnl_partialKnn_wrapper_53_0__ap_start;
  assign out_dist_53__din = krnl_partialKnn_wrapper_53_0_out_dist_din;
  assign krnl_partialKnn_wrapper_53_0_out_dist_full_n = out_dist_53__full_n;
  assign out_dist_53__write = krnl_partialKnn_wrapper_53_0_out_dist_write;
  assign out_id_53__din = krnl_partialKnn_wrapper_53_0_out_id_din;
  assign krnl_partialKnn_wrapper_53_0_out_id_full_n = out_id_53__full_n;
  assign out_id_53__write = krnl_partialKnn_wrapper_53_0_out_id_write;
  assign krnl_partialKnn_wrapper_53_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_53_0___in_53__q0;
  assign in_53_read_addr__din = krnl_partialKnn_wrapper_53_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_53_0_searchSpace_0_read_addr_s_full_n = in_53_read_addr__full_n;
  assign in_53_read_addr__write = krnl_partialKnn_wrapper_53_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_53_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_53_read_data__dout };
  assign krnl_partialKnn_wrapper_53_0_searchSpace_read_data_peek_empty_n = in_53_read_data__empty_n;
  assign krnl_partialKnn_wrapper_53_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_53_read_data__dout };
  assign krnl_partialKnn_wrapper_53_0_searchSpace_0_read_data_s_empty_n = in_53_read_data__empty_n;
  assign in_53_read_data__read = krnl_partialKnn_wrapper_53_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_53_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_53_0___in_53__q0;
  assign in_53_write_addr__din = krnl_partialKnn_wrapper_53_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_53_0_searchSpace_0_write_addr_s_full_n = in_53_write_addr__full_n;
  assign in_53_write_addr__write = krnl_partialKnn_wrapper_53_0_searchSpace_0_write_addr_s_write;
  assign in_53_write_data__din = krnl_partialKnn_wrapper_53_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_53_0_searchSpace_0_write_data_full_n = in_53_write_data__full_n;
  assign in_53_write_data__write = krnl_partialKnn_wrapper_53_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_53_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_53_write_resp__dout };
  assign krnl_partialKnn_wrapper_53_0_searchSpace_write_resp_peek_empty_n = in_53_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_53_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_53_write_resp__dout };
  assign krnl_partialKnn_wrapper_53_0_searchSpace_0_write_resp_s_empty_n = in_53_write_resp__empty_n;
  assign in_53_write_resp__read = krnl_partialKnn_wrapper_53_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_53_0_start_id_0 = 64'd434176;
  assign krnl_partialKnn_wrapper_6_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_6_0__ap_done = krnl_partialKnn_wrapper_6_0_ap_done;
  assign krnl_partialKnn_wrapper_6_0__ap_idle = krnl_partialKnn_wrapper_6_0_ap_idle;
  assign krnl_partialKnn_wrapper_6_0__ap_ready = krnl_partialKnn_wrapper_6_0_ap_ready;
  assign krnl_partialKnn_wrapper_6_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_6_0_ap_start = krnl_partialKnn_wrapper_6_0__ap_start;
  assign out_dist_6__din = krnl_partialKnn_wrapper_6_0_out_dist_din;
  assign krnl_partialKnn_wrapper_6_0_out_dist_full_n = out_dist_6__full_n;
  assign out_dist_6__write = krnl_partialKnn_wrapper_6_0_out_dist_write;
  assign out_id_6__din = krnl_partialKnn_wrapper_6_0_out_id_din;
  assign krnl_partialKnn_wrapper_6_0_out_id_full_n = out_id_6__full_n;
  assign out_id_6__write = krnl_partialKnn_wrapper_6_0_out_id_write;
  assign krnl_partialKnn_wrapper_6_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_6_0___in_6__q0;
  assign in_6_read_addr__din = krnl_partialKnn_wrapper_6_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_6_0_searchSpace_0_read_addr_s_full_n = in_6_read_addr__full_n;
  assign in_6_read_addr__write = krnl_partialKnn_wrapper_6_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_6_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_6_read_data__dout };
  assign krnl_partialKnn_wrapper_6_0_searchSpace_0_read_data_peek_empty_n = in_6_read_data__empty_n;
  assign krnl_partialKnn_wrapper_6_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_6_read_data__dout };
  assign krnl_partialKnn_wrapper_6_0_searchSpace_0_read_data_s_empty_n = in_6_read_data__empty_n;
  assign in_6_read_data__read = krnl_partialKnn_wrapper_6_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_6_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_6_0___in_6__q0;
  assign in_6_write_addr__din = krnl_partialKnn_wrapper_6_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_6_0_searchSpace_0_write_addr_s_full_n = in_6_write_addr__full_n;
  assign in_6_write_addr__write = krnl_partialKnn_wrapper_6_0_searchSpace_0_write_addr_s_write;
  assign in_6_write_data__din = krnl_partialKnn_wrapper_6_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_6_0_searchSpace_0_write_data_full_n = in_6_write_data__full_n;
  assign in_6_write_data__write = krnl_partialKnn_wrapper_6_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_6_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_6_write_resp__dout };
  assign krnl_partialKnn_wrapper_6_0_searchSpace_write_resp_peek_empty_n = in_6_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_6_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_6_write_resp__dout };
  assign krnl_partialKnn_wrapper_6_0_searchSpace_0_write_resp_s_empty_n = in_6_write_resp__empty_n;
  assign in_6_write_resp__read = krnl_partialKnn_wrapper_6_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_6_0_start_id_0 = 64'd49152;
  assign krnl_partialKnn_wrapper_7_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_7_0__ap_done = krnl_partialKnn_wrapper_7_0_ap_done;
  assign krnl_partialKnn_wrapper_7_0__ap_idle = krnl_partialKnn_wrapper_7_0_ap_idle;
  assign krnl_partialKnn_wrapper_7_0__ap_ready = krnl_partialKnn_wrapper_7_0_ap_ready;
  assign krnl_partialKnn_wrapper_7_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_7_0_ap_start = krnl_partialKnn_wrapper_7_0__ap_start;
  assign out_dist_7__din = krnl_partialKnn_wrapper_7_0_out_dist_din;
  assign krnl_partialKnn_wrapper_7_0_out_dist_full_n = out_dist_7__full_n;
  assign out_dist_7__write = krnl_partialKnn_wrapper_7_0_out_dist_write;
  assign out_id_7__din = krnl_partialKnn_wrapper_7_0_out_id_din;
  assign krnl_partialKnn_wrapper_7_0_out_id_full_n = out_id_7__full_n;
  assign out_id_7__write = krnl_partialKnn_wrapper_7_0_out_id_write;
  assign krnl_partialKnn_wrapper_7_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_7_0___in_7__q0;
  assign in_7_read_addr__din = krnl_partialKnn_wrapper_7_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_7_0_searchSpace_0_read_addr_s_full_n = in_7_read_addr__full_n;
  assign in_7_read_addr__write = krnl_partialKnn_wrapper_7_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_7_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_7_read_data__dout };
  assign krnl_partialKnn_wrapper_7_0_searchSpace_0_read_data_peek_empty_n = in_7_read_data__empty_n;
  assign krnl_partialKnn_wrapper_7_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_7_read_data__dout };
  assign krnl_partialKnn_wrapper_7_0_searchSpace_0_read_data_s_empty_n = in_7_read_data__empty_n;
  assign in_7_read_data__read = krnl_partialKnn_wrapper_7_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_7_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_7_0___in_7__q0;
  assign in_7_write_addr__din = krnl_partialKnn_wrapper_7_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_7_0_searchSpace_0_write_addr_s_full_n = in_7_write_addr__full_n;
  assign in_7_write_addr__write = krnl_partialKnn_wrapper_7_0_searchSpace_0_write_addr_s_write;
  assign in_7_write_data__din = krnl_partialKnn_wrapper_7_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_7_0_searchSpace_0_write_data_full_n = in_7_write_data__full_n;
  assign in_7_write_data__write = krnl_partialKnn_wrapper_7_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_7_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_7_write_resp__dout };
  assign krnl_partialKnn_wrapper_7_0_searchSpace_write_resp_peek_empty_n = in_7_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_7_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_7_write_resp__dout };
  assign krnl_partialKnn_wrapper_7_0_searchSpace_0_write_resp_s_empty_n = in_7_write_resp__empty_n;
  assign in_7_write_resp__read = krnl_partialKnn_wrapper_7_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_7_0_start_id_0 = 64'd57344;
  assign krnl_partialKnn_wrapper_8_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_8_0__ap_done = krnl_partialKnn_wrapper_8_0_ap_done;
  assign krnl_partialKnn_wrapper_8_0__ap_idle = krnl_partialKnn_wrapper_8_0_ap_idle;
  assign krnl_partialKnn_wrapper_8_0__ap_ready = krnl_partialKnn_wrapper_8_0_ap_ready;
  assign krnl_partialKnn_wrapper_8_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_8_0_ap_start = krnl_partialKnn_wrapper_8_0__ap_start;
  assign out_dist_8__din = krnl_partialKnn_wrapper_8_0_out_dist_din;
  assign krnl_partialKnn_wrapper_8_0_out_dist_full_n = out_dist_8__full_n;
  assign out_dist_8__write = krnl_partialKnn_wrapper_8_0_out_dist_write;
  assign out_id_8__din = krnl_partialKnn_wrapper_8_0_out_id_din;
  assign krnl_partialKnn_wrapper_8_0_out_id_full_n = out_id_8__full_n;
  assign out_id_8__write = krnl_partialKnn_wrapper_8_0_out_id_write;
  assign krnl_partialKnn_wrapper_8_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_8_0___in_8__q0;
  assign in_8_read_addr__din = krnl_partialKnn_wrapper_8_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_8_0_searchSpace_0_read_addr_s_full_n = in_8_read_addr__full_n;
  assign in_8_read_addr__write = krnl_partialKnn_wrapper_8_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_8_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_8_read_data__dout };
  assign krnl_partialKnn_wrapper_8_0_searchSpace_0_read_data_peek_empty_n = in_8_read_data__empty_n;
  assign krnl_partialKnn_wrapper_8_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_8_read_data__dout };
  assign krnl_partialKnn_wrapper_8_0_searchSpace_0_read_data_s_empty_n = in_8_read_data__empty_n;
  assign in_8_read_data__read = krnl_partialKnn_wrapper_8_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_8_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_8_0___in_8__q0;
  assign in_8_write_addr__din = krnl_partialKnn_wrapper_8_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_8_0_searchSpace_0_write_addr_s_full_n = in_8_write_addr__full_n;
  assign in_8_write_addr__write = krnl_partialKnn_wrapper_8_0_searchSpace_0_write_addr_s_write;
  assign in_8_write_data__din = krnl_partialKnn_wrapper_8_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_8_0_searchSpace_0_write_data_full_n = in_8_write_data__full_n;
  assign in_8_write_data__write = krnl_partialKnn_wrapper_8_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_8_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_8_write_resp__dout };
  assign krnl_partialKnn_wrapper_8_0_searchSpace_write_resp_peek_empty_n = in_8_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_8_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_8_write_resp__dout };
  assign krnl_partialKnn_wrapper_8_0_searchSpace_0_write_resp_s_empty_n = in_8_write_resp__empty_n;
  assign in_8_write_resp__read = krnl_partialKnn_wrapper_8_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_8_0_start_id_0 = 64'd65536;
  assign krnl_partialKnn_wrapper_9_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_9_0__ap_done = krnl_partialKnn_wrapper_9_0_ap_done;
  assign krnl_partialKnn_wrapper_9_0__ap_idle = krnl_partialKnn_wrapper_9_0_ap_idle;
  assign krnl_partialKnn_wrapper_9_0__ap_ready = krnl_partialKnn_wrapper_9_0_ap_ready;
  assign krnl_partialKnn_wrapper_9_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_9_0_ap_start = krnl_partialKnn_wrapper_9_0__ap_start;
  assign out_dist_9__din = krnl_partialKnn_wrapper_9_0_out_dist_din;
  assign krnl_partialKnn_wrapper_9_0_out_dist_full_n = out_dist_9__full_n;
  assign out_dist_9__write = krnl_partialKnn_wrapper_9_0_out_dist_write;
  assign out_id_9__din = krnl_partialKnn_wrapper_9_0_out_id_din;
  assign krnl_partialKnn_wrapper_9_0_out_id_full_n = out_id_9__full_n;
  assign out_id_9__write = krnl_partialKnn_wrapper_9_0_out_id_write;
  assign krnl_partialKnn_wrapper_9_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_9_0___in_9__q0;
  assign in_9_read_addr__din = krnl_partialKnn_wrapper_9_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_9_0_searchSpace_0_read_addr_s_full_n = in_9_read_addr__full_n;
  assign in_9_read_addr__write = krnl_partialKnn_wrapper_9_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_9_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_9_read_data__dout };
  assign krnl_partialKnn_wrapper_9_0_searchSpace_0_read_data_peek_empty_n = in_9_read_data__empty_n;
  assign krnl_partialKnn_wrapper_9_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_9_read_data__dout };
  assign krnl_partialKnn_wrapper_9_0_searchSpace_0_read_data_s_empty_n = in_9_read_data__empty_n;
  assign in_9_read_data__read = krnl_partialKnn_wrapper_9_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_9_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_9_0___in_9__q0;
  assign in_9_write_addr__din = krnl_partialKnn_wrapper_9_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_9_0_searchSpace_0_write_addr_s_full_n = in_9_write_addr__full_n;
  assign in_9_write_addr__write = krnl_partialKnn_wrapper_9_0_searchSpace_0_write_addr_s_write;
  assign in_9_write_data__din = krnl_partialKnn_wrapper_9_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_9_0_searchSpace_0_write_data_full_n = in_9_write_data__full_n;
  assign in_9_write_data__write = krnl_partialKnn_wrapper_9_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_9_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_9_write_resp__dout };
  assign krnl_partialKnn_wrapper_9_0_searchSpace_write_resp_peek_empty_n = in_9_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_9_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_9_write_resp__dout };
  assign krnl_partialKnn_wrapper_9_0_searchSpace_0_write_resp_s_empty_n = in_9_write_resp__empty_n;
  assign in_9_write_resp__read = krnl_partialKnn_wrapper_9_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_9_0_start_id_0 = 64'd73728;
  assign L4_out_dist__m_axi_clk = ap_clk;
  assign m_axi_L4_out_dist_ARADDR = L4_out_dist__m_axi_m_axi_ARADDR;
  assign m_axi_L4_out_dist_ARBURST = L4_out_dist__m_axi_m_axi_ARBURST;
  assign m_axi_L4_out_dist_ARCACHE = L4_out_dist__m_axi_m_axi_ARCACHE;
  assign m_axi_L4_out_dist_ARID = L4_out_dist__m_axi_m_axi_ARID;
  assign m_axi_L4_out_dist_ARLEN = L4_out_dist__m_axi_m_axi_ARLEN;
  assign m_axi_L4_out_dist_ARLOCK = L4_out_dist__m_axi_m_axi_ARLOCK;
  assign m_axi_L4_out_dist_ARPROT = L4_out_dist__m_axi_m_axi_ARPROT;
  assign m_axi_L4_out_dist_ARQOS = L4_out_dist__m_axi_m_axi_ARQOS;
  assign L4_out_dist__m_axi_m_axi_ARREADY = m_axi_L4_out_dist_ARREADY;
  assign m_axi_L4_out_dist_ARSIZE = L4_out_dist__m_axi_m_axi_ARSIZE;
  assign m_axi_L4_out_dist_ARVALID = L4_out_dist__m_axi_m_axi_ARVALID;
  assign m_axi_L4_out_dist_AWADDR = L4_out_dist__m_axi_m_axi_AWADDR;
  assign m_axi_L4_out_dist_AWBURST = L4_out_dist__m_axi_m_axi_AWBURST;
  assign m_axi_L4_out_dist_AWCACHE = L4_out_dist__m_axi_m_axi_AWCACHE;
  assign m_axi_L4_out_dist_AWID = L4_out_dist__m_axi_m_axi_AWID;
  assign m_axi_L4_out_dist_AWLEN = L4_out_dist__m_axi_m_axi_AWLEN;
  assign m_axi_L4_out_dist_AWLOCK = L4_out_dist__m_axi_m_axi_AWLOCK;
  assign m_axi_L4_out_dist_AWPROT = L4_out_dist__m_axi_m_axi_AWPROT;
  assign m_axi_L4_out_dist_AWQOS = L4_out_dist__m_axi_m_axi_AWQOS;
  assign L4_out_dist__m_axi_m_axi_AWREADY = m_axi_L4_out_dist_AWREADY;
  assign m_axi_L4_out_dist_AWSIZE = L4_out_dist__m_axi_m_axi_AWSIZE;
  assign m_axi_L4_out_dist_AWVALID = L4_out_dist__m_axi_m_axi_AWVALID;
  assign L4_out_dist__m_axi_m_axi_BID = m_axi_L4_out_dist_BID;
  assign m_axi_L4_out_dist_BREADY = L4_out_dist__m_axi_m_axi_BREADY;
  assign L4_out_dist__m_axi_m_axi_BRESP = m_axi_L4_out_dist_BRESP;
  assign L4_out_dist__m_axi_m_axi_BVALID = m_axi_L4_out_dist_BVALID;
  assign L4_out_dist__m_axi_m_axi_RDATA = m_axi_L4_out_dist_RDATA;
  assign L4_out_dist__m_axi_m_axi_RID = m_axi_L4_out_dist_RID;
  assign L4_out_dist__m_axi_m_axi_RLAST = m_axi_L4_out_dist_RLAST;
  assign m_axi_L4_out_dist_RREADY = L4_out_dist__m_axi_m_axi_RREADY;
  assign L4_out_dist__m_axi_m_axi_RRESP = m_axi_L4_out_dist_RRESP;
  assign L4_out_dist__m_axi_m_axi_RVALID = m_axi_L4_out_dist_RVALID;
  assign m_axi_L4_out_dist_WDATA = L4_out_dist__m_axi_m_axi_WDATA;
  assign m_axi_L4_out_dist_WLAST = L4_out_dist__m_axi_m_axi_WLAST;
  assign L4_out_dist__m_axi_m_axi_WREADY = m_axi_L4_out_dist_WREADY;
  assign m_axi_L4_out_dist_WSTRB = L4_out_dist__m_axi_m_axi_WSTRB;
  assign m_axi_L4_out_dist_WVALID = L4_out_dist__m_axi_m_axi_WVALID;
  assign L4_out_dist__m_axi_read_addr_din = L4_out_dist_read_addr__din;
  assign L4_out_dist_read_addr__full_n = L4_out_dist__m_axi_read_addr_full_n;
  assign L4_out_dist__m_axi_read_addr_write = L4_out_dist_read_addr__write;
  assign L4_out_dist_read_data__dout = L4_out_dist__m_axi_read_data_dout;
  assign L4_out_dist_read_data__empty_n = L4_out_dist__m_axi_read_data_empty_n;
  assign L4_out_dist__m_axi_read_data_read = L4_out_dist_read_data__read;
  assign L4_out_dist__m_axi_rst = ~ ap_rst_n;
  assign L4_out_dist__m_axi_write_addr_din = L4_out_dist_write_addr__din;
  assign L4_out_dist_write_addr__full_n = L4_out_dist__m_axi_write_addr_full_n;
  assign L4_out_dist__m_axi_write_addr_write = L4_out_dist_write_addr__write;
  assign L4_out_dist__m_axi_write_data_din = L4_out_dist_write_data__din;
  assign L4_out_dist_write_data__full_n = L4_out_dist__m_axi_write_data_full_n;
  assign L4_out_dist__m_axi_write_data_write = L4_out_dist_write_data__write;
  assign L4_out_dist_write_resp__dout = L4_out_dist__m_axi_write_resp_dout;
  assign L4_out_dist_write_resp__empty_n = L4_out_dist__m_axi_write_resp_empty_n;
  assign L4_out_dist__m_axi_write_resp_read = L4_out_dist_write_resp__read;
  assign L4_out_id__m_axi_clk = ap_clk;
  assign m_axi_L4_out_id_ARADDR = L4_out_id__m_axi_m_axi_ARADDR;
  assign m_axi_L4_out_id_ARBURST = L4_out_id__m_axi_m_axi_ARBURST;
  assign m_axi_L4_out_id_ARCACHE = L4_out_id__m_axi_m_axi_ARCACHE;
  assign m_axi_L4_out_id_ARID = L4_out_id__m_axi_m_axi_ARID;
  assign m_axi_L4_out_id_ARLEN = L4_out_id__m_axi_m_axi_ARLEN;
  assign m_axi_L4_out_id_ARLOCK = L4_out_id__m_axi_m_axi_ARLOCK;
  assign m_axi_L4_out_id_ARPROT = L4_out_id__m_axi_m_axi_ARPROT;
  assign m_axi_L4_out_id_ARQOS = L4_out_id__m_axi_m_axi_ARQOS;
  assign L4_out_id__m_axi_m_axi_ARREADY = m_axi_L4_out_id_ARREADY;
  assign m_axi_L4_out_id_ARSIZE = L4_out_id__m_axi_m_axi_ARSIZE;
  assign m_axi_L4_out_id_ARVALID = L4_out_id__m_axi_m_axi_ARVALID;
  assign m_axi_L4_out_id_AWADDR = L4_out_id__m_axi_m_axi_AWADDR;
  assign m_axi_L4_out_id_AWBURST = L4_out_id__m_axi_m_axi_AWBURST;
  assign m_axi_L4_out_id_AWCACHE = L4_out_id__m_axi_m_axi_AWCACHE;
  assign m_axi_L4_out_id_AWID = L4_out_id__m_axi_m_axi_AWID;
  assign m_axi_L4_out_id_AWLEN = L4_out_id__m_axi_m_axi_AWLEN;
  assign m_axi_L4_out_id_AWLOCK = L4_out_id__m_axi_m_axi_AWLOCK;
  assign m_axi_L4_out_id_AWPROT = L4_out_id__m_axi_m_axi_AWPROT;
  assign m_axi_L4_out_id_AWQOS = L4_out_id__m_axi_m_axi_AWQOS;
  assign L4_out_id__m_axi_m_axi_AWREADY = m_axi_L4_out_id_AWREADY;
  assign m_axi_L4_out_id_AWSIZE = L4_out_id__m_axi_m_axi_AWSIZE;
  assign m_axi_L4_out_id_AWVALID = L4_out_id__m_axi_m_axi_AWVALID;
  assign L4_out_id__m_axi_m_axi_BID = m_axi_L4_out_id_BID;
  assign m_axi_L4_out_id_BREADY = L4_out_id__m_axi_m_axi_BREADY;
  assign L4_out_id__m_axi_m_axi_BRESP = m_axi_L4_out_id_BRESP;
  assign L4_out_id__m_axi_m_axi_BVALID = m_axi_L4_out_id_BVALID;
  assign L4_out_id__m_axi_m_axi_RDATA = m_axi_L4_out_id_RDATA;
  assign L4_out_id__m_axi_m_axi_RID = m_axi_L4_out_id_RID;
  assign L4_out_id__m_axi_m_axi_RLAST = m_axi_L4_out_id_RLAST;
  assign m_axi_L4_out_id_RREADY = L4_out_id__m_axi_m_axi_RREADY;
  assign L4_out_id__m_axi_m_axi_RRESP = m_axi_L4_out_id_RRESP;
  assign L4_out_id__m_axi_m_axi_RVALID = m_axi_L4_out_id_RVALID;
  assign m_axi_L4_out_id_WDATA = L4_out_id__m_axi_m_axi_WDATA;
  assign m_axi_L4_out_id_WLAST = L4_out_id__m_axi_m_axi_WLAST;
  assign L4_out_id__m_axi_m_axi_WREADY = m_axi_L4_out_id_WREADY;
  assign m_axi_L4_out_id_WSTRB = L4_out_id__m_axi_m_axi_WSTRB;
  assign m_axi_L4_out_id_WVALID = L4_out_id__m_axi_m_axi_WVALID;
  assign L4_out_id__m_axi_read_addr_din = L4_out_id_read_addr__din;
  assign L4_out_id_read_addr__full_n = L4_out_id__m_axi_read_addr_full_n;
  assign L4_out_id__m_axi_read_addr_write = L4_out_id_read_addr__write;
  assign L4_out_id_read_data__dout = L4_out_id__m_axi_read_data_dout;
  assign L4_out_id_read_data__empty_n = L4_out_id__m_axi_read_data_empty_n;
  assign L4_out_id__m_axi_read_data_read = L4_out_id_read_data__read;
  assign L4_out_id__m_axi_rst = ~ ap_rst_n;
  assign L4_out_id__m_axi_write_addr_din = L4_out_id_write_addr__din;
  assign L4_out_id_write_addr__full_n = L4_out_id__m_axi_write_addr_full_n;
  assign L4_out_id__m_axi_write_addr_write = L4_out_id_write_addr__write;
  assign L4_out_id__m_axi_write_data_din = L4_out_id_write_data__din;
  assign L4_out_id_write_data__full_n = L4_out_id__m_axi_write_data_full_n;
  assign L4_out_id__m_axi_write_data_write = L4_out_id_write_data__write;
  assign L4_out_id_write_resp__dout = L4_out_id__m_axi_write_resp_dout;
  assign L4_out_id_write_resp__empty_n = L4_out_id__m_axi_write_resp_empty_n;
  assign L4_out_id__m_axi_write_resp_read = L4_out_id_write_resp__read;
  assign in_0__m_axi_clk = ap_clk;
  assign m_axi_in_0_ARADDR = in_0__m_axi_m_axi_ARADDR;
  assign m_axi_in_0_ARBURST = in_0__m_axi_m_axi_ARBURST;
  assign m_axi_in_0_ARCACHE = in_0__m_axi_m_axi_ARCACHE;
  assign m_axi_in_0_ARID = in_0__m_axi_m_axi_ARID;
  assign m_axi_in_0_ARLEN = in_0__m_axi_m_axi_ARLEN;
  assign m_axi_in_0_ARLOCK = in_0__m_axi_m_axi_ARLOCK;
  assign m_axi_in_0_ARPROT = in_0__m_axi_m_axi_ARPROT;
  assign m_axi_in_0_ARQOS = in_0__m_axi_m_axi_ARQOS;
  assign in_0__m_axi_m_axi_ARREADY = m_axi_in_0_ARREADY;
  assign m_axi_in_0_ARSIZE = in_0__m_axi_m_axi_ARSIZE;
  assign m_axi_in_0_ARVALID = in_0__m_axi_m_axi_ARVALID;
  assign m_axi_in_0_AWADDR = in_0__m_axi_m_axi_AWADDR;
  assign m_axi_in_0_AWBURST = in_0__m_axi_m_axi_AWBURST;
  assign m_axi_in_0_AWCACHE = in_0__m_axi_m_axi_AWCACHE;
  assign m_axi_in_0_AWID = in_0__m_axi_m_axi_AWID;
  assign m_axi_in_0_AWLEN = in_0__m_axi_m_axi_AWLEN;
  assign m_axi_in_0_AWLOCK = in_0__m_axi_m_axi_AWLOCK;
  assign m_axi_in_0_AWPROT = in_0__m_axi_m_axi_AWPROT;
  assign m_axi_in_0_AWQOS = in_0__m_axi_m_axi_AWQOS;
  assign in_0__m_axi_m_axi_AWREADY = m_axi_in_0_AWREADY;
  assign m_axi_in_0_AWSIZE = in_0__m_axi_m_axi_AWSIZE;
  assign m_axi_in_0_AWVALID = in_0__m_axi_m_axi_AWVALID;
  assign in_0__m_axi_m_axi_BID = m_axi_in_0_BID;
  assign m_axi_in_0_BREADY = in_0__m_axi_m_axi_BREADY;
  assign in_0__m_axi_m_axi_BRESP = m_axi_in_0_BRESP;
  assign in_0__m_axi_m_axi_BVALID = m_axi_in_0_BVALID;
  assign in_0__m_axi_m_axi_RDATA = m_axi_in_0_RDATA;
  assign in_0__m_axi_m_axi_RID = m_axi_in_0_RID;
  assign in_0__m_axi_m_axi_RLAST = m_axi_in_0_RLAST;
  assign m_axi_in_0_RREADY = in_0__m_axi_m_axi_RREADY;
  assign in_0__m_axi_m_axi_RRESP = m_axi_in_0_RRESP;
  assign in_0__m_axi_m_axi_RVALID = m_axi_in_0_RVALID;
  assign m_axi_in_0_WDATA = in_0__m_axi_m_axi_WDATA;
  assign m_axi_in_0_WLAST = in_0__m_axi_m_axi_WLAST;
  assign in_0__m_axi_m_axi_WREADY = m_axi_in_0_WREADY;
  assign m_axi_in_0_WSTRB = in_0__m_axi_m_axi_WSTRB;
  assign m_axi_in_0_WVALID = in_0__m_axi_m_axi_WVALID;
  assign in_0__m_axi_read_addr_din = in_0_read_addr__din;
  assign in_0_read_addr__full_n = in_0__m_axi_read_addr_full_n;
  assign in_0__m_axi_read_addr_write = in_0_read_addr__write;
  assign in_0_read_data__dout = in_0__m_axi_read_data_dout;
  assign in_0_read_data__empty_n = in_0__m_axi_read_data_empty_n;
  assign in_0__m_axi_read_data_read = in_0_read_data__read;
  assign in_0__m_axi_rst = ~ ap_rst_n;
  assign in_0__m_axi_write_addr_din = in_0_write_addr__din;
  assign in_0_write_addr__full_n = in_0__m_axi_write_addr_full_n;
  assign in_0__m_axi_write_addr_write = in_0_write_addr__write;
  assign in_0__m_axi_write_data_din = in_0_write_data__din;
  assign in_0_write_data__full_n = in_0__m_axi_write_data_full_n;
  assign in_0__m_axi_write_data_write = in_0_write_data__write;
  assign in_0_write_resp__dout = in_0__m_axi_write_resp_dout;
  assign in_0_write_resp__empty_n = in_0__m_axi_write_resp_empty_n;
  assign in_0__m_axi_write_resp_read = in_0_write_resp__read;
  assign in_1__m_axi_clk = ap_clk;
  assign m_axi_in_1_ARADDR = in_1__m_axi_m_axi_ARADDR;
  assign m_axi_in_1_ARBURST = in_1__m_axi_m_axi_ARBURST;
  assign m_axi_in_1_ARCACHE = in_1__m_axi_m_axi_ARCACHE;
  assign m_axi_in_1_ARID = in_1__m_axi_m_axi_ARID;
  assign m_axi_in_1_ARLEN = in_1__m_axi_m_axi_ARLEN;
  assign m_axi_in_1_ARLOCK = in_1__m_axi_m_axi_ARLOCK;
  assign m_axi_in_1_ARPROT = in_1__m_axi_m_axi_ARPROT;
  assign m_axi_in_1_ARQOS = in_1__m_axi_m_axi_ARQOS;
  assign in_1__m_axi_m_axi_ARREADY = m_axi_in_1_ARREADY;
  assign m_axi_in_1_ARSIZE = in_1__m_axi_m_axi_ARSIZE;
  assign m_axi_in_1_ARVALID = in_1__m_axi_m_axi_ARVALID;
  assign m_axi_in_1_AWADDR = in_1__m_axi_m_axi_AWADDR;
  assign m_axi_in_1_AWBURST = in_1__m_axi_m_axi_AWBURST;
  assign m_axi_in_1_AWCACHE = in_1__m_axi_m_axi_AWCACHE;
  assign m_axi_in_1_AWID = in_1__m_axi_m_axi_AWID;
  assign m_axi_in_1_AWLEN = in_1__m_axi_m_axi_AWLEN;
  assign m_axi_in_1_AWLOCK = in_1__m_axi_m_axi_AWLOCK;
  assign m_axi_in_1_AWPROT = in_1__m_axi_m_axi_AWPROT;
  assign m_axi_in_1_AWQOS = in_1__m_axi_m_axi_AWQOS;
  assign in_1__m_axi_m_axi_AWREADY = m_axi_in_1_AWREADY;
  assign m_axi_in_1_AWSIZE = in_1__m_axi_m_axi_AWSIZE;
  assign m_axi_in_1_AWVALID = in_1__m_axi_m_axi_AWVALID;
  assign in_1__m_axi_m_axi_BID = m_axi_in_1_BID;
  assign m_axi_in_1_BREADY = in_1__m_axi_m_axi_BREADY;
  assign in_1__m_axi_m_axi_BRESP = m_axi_in_1_BRESP;
  assign in_1__m_axi_m_axi_BVALID = m_axi_in_1_BVALID;
  assign in_1__m_axi_m_axi_RDATA = m_axi_in_1_RDATA;
  assign in_1__m_axi_m_axi_RID = m_axi_in_1_RID;
  assign in_1__m_axi_m_axi_RLAST = m_axi_in_1_RLAST;
  assign m_axi_in_1_RREADY = in_1__m_axi_m_axi_RREADY;
  assign in_1__m_axi_m_axi_RRESP = m_axi_in_1_RRESP;
  assign in_1__m_axi_m_axi_RVALID = m_axi_in_1_RVALID;
  assign m_axi_in_1_WDATA = in_1__m_axi_m_axi_WDATA;
  assign m_axi_in_1_WLAST = in_1__m_axi_m_axi_WLAST;
  assign in_1__m_axi_m_axi_WREADY = m_axi_in_1_WREADY;
  assign m_axi_in_1_WSTRB = in_1__m_axi_m_axi_WSTRB;
  assign m_axi_in_1_WVALID = in_1__m_axi_m_axi_WVALID;
  assign in_1__m_axi_read_addr_din = in_1_read_addr__din;
  assign in_1_read_addr__full_n = in_1__m_axi_read_addr_full_n;
  assign in_1__m_axi_read_addr_write = in_1_read_addr__write;
  assign in_1_read_data__dout = in_1__m_axi_read_data_dout;
  assign in_1_read_data__empty_n = in_1__m_axi_read_data_empty_n;
  assign in_1__m_axi_read_data_read = in_1_read_data__read;
  assign in_1__m_axi_rst = ~ ap_rst_n;
  assign in_1__m_axi_write_addr_din = in_1_write_addr__din;
  assign in_1_write_addr__full_n = in_1__m_axi_write_addr_full_n;
  assign in_1__m_axi_write_addr_write = in_1_write_addr__write;
  assign in_1__m_axi_write_data_din = in_1_write_data__din;
  assign in_1_write_data__full_n = in_1__m_axi_write_data_full_n;
  assign in_1__m_axi_write_data_write = in_1_write_data__write;
  assign in_1_write_resp__dout = in_1__m_axi_write_resp_dout;
  assign in_1_write_resp__empty_n = in_1__m_axi_write_resp_empty_n;
  assign in_1__m_axi_write_resp_read = in_1_write_resp__read;
  assign in_10__m_axi_clk = ap_clk;
  assign m_axi_in_10_ARADDR = in_10__m_axi_m_axi_ARADDR;
  assign m_axi_in_10_ARBURST = in_10__m_axi_m_axi_ARBURST;
  assign m_axi_in_10_ARCACHE = in_10__m_axi_m_axi_ARCACHE;
  assign m_axi_in_10_ARID = in_10__m_axi_m_axi_ARID;
  assign m_axi_in_10_ARLEN = in_10__m_axi_m_axi_ARLEN;
  assign m_axi_in_10_ARLOCK = in_10__m_axi_m_axi_ARLOCK;
  assign m_axi_in_10_ARPROT = in_10__m_axi_m_axi_ARPROT;
  assign m_axi_in_10_ARQOS = in_10__m_axi_m_axi_ARQOS;
  assign in_10__m_axi_m_axi_ARREADY = m_axi_in_10_ARREADY;
  assign m_axi_in_10_ARSIZE = in_10__m_axi_m_axi_ARSIZE;
  assign m_axi_in_10_ARVALID = in_10__m_axi_m_axi_ARVALID;
  assign m_axi_in_10_AWADDR = in_10__m_axi_m_axi_AWADDR;
  assign m_axi_in_10_AWBURST = in_10__m_axi_m_axi_AWBURST;
  assign m_axi_in_10_AWCACHE = in_10__m_axi_m_axi_AWCACHE;
  assign m_axi_in_10_AWID = in_10__m_axi_m_axi_AWID;
  assign m_axi_in_10_AWLEN = in_10__m_axi_m_axi_AWLEN;
  assign m_axi_in_10_AWLOCK = in_10__m_axi_m_axi_AWLOCK;
  assign m_axi_in_10_AWPROT = in_10__m_axi_m_axi_AWPROT;
  assign m_axi_in_10_AWQOS = in_10__m_axi_m_axi_AWQOS;
  assign in_10__m_axi_m_axi_AWREADY = m_axi_in_10_AWREADY;
  assign m_axi_in_10_AWSIZE = in_10__m_axi_m_axi_AWSIZE;
  assign m_axi_in_10_AWVALID = in_10__m_axi_m_axi_AWVALID;
  assign in_10__m_axi_m_axi_BID = m_axi_in_10_BID;
  assign m_axi_in_10_BREADY = in_10__m_axi_m_axi_BREADY;
  assign in_10__m_axi_m_axi_BRESP = m_axi_in_10_BRESP;
  assign in_10__m_axi_m_axi_BVALID = m_axi_in_10_BVALID;
  assign in_10__m_axi_m_axi_RDATA = m_axi_in_10_RDATA;
  assign in_10__m_axi_m_axi_RID = m_axi_in_10_RID;
  assign in_10__m_axi_m_axi_RLAST = m_axi_in_10_RLAST;
  assign m_axi_in_10_RREADY = in_10__m_axi_m_axi_RREADY;
  assign in_10__m_axi_m_axi_RRESP = m_axi_in_10_RRESP;
  assign in_10__m_axi_m_axi_RVALID = m_axi_in_10_RVALID;
  assign m_axi_in_10_WDATA = in_10__m_axi_m_axi_WDATA;
  assign m_axi_in_10_WLAST = in_10__m_axi_m_axi_WLAST;
  assign in_10__m_axi_m_axi_WREADY = m_axi_in_10_WREADY;
  assign m_axi_in_10_WSTRB = in_10__m_axi_m_axi_WSTRB;
  assign m_axi_in_10_WVALID = in_10__m_axi_m_axi_WVALID;
  assign in_10__m_axi_read_addr_din = in_10_read_addr__din;
  assign in_10_read_addr__full_n = in_10__m_axi_read_addr_full_n;
  assign in_10__m_axi_read_addr_write = in_10_read_addr__write;
  assign in_10_read_data__dout = in_10__m_axi_read_data_dout;
  assign in_10_read_data__empty_n = in_10__m_axi_read_data_empty_n;
  assign in_10__m_axi_read_data_read = in_10_read_data__read;
  assign in_10__m_axi_rst = ~ ap_rst_n;
  assign in_10__m_axi_write_addr_din = in_10_write_addr__din;
  assign in_10_write_addr__full_n = in_10__m_axi_write_addr_full_n;
  assign in_10__m_axi_write_addr_write = in_10_write_addr__write;
  assign in_10__m_axi_write_data_din = in_10_write_data__din;
  assign in_10_write_data__full_n = in_10__m_axi_write_data_full_n;
  assign in_10__m_axi_write_data_write = in_10_write_data__write;
  assign in_10_write_resp__dout = in_10__m_axi_write_resp_dout;
  assign in_10_write_resp__empty_n = in_10__m_axi_write_resp_empty_n;
  assign in_10__m_axi_write_resp_read = in_10_write_resp__read;
  assign in_11__m_axi_clk = ap_clk;
  assign m_axi_in_11_ARADDR = in_11__m_axi_m_axi_ARADDR;
  assign m_axi_in_11_ARBURST = in_11__m_axi_m_axi_ARBURST;
  assign m_axi_in_11_ARCACHE = in_11__m_axi_m_axi_ARCACHE;
  assign m_axi_in_11_ARID = in_11__m_axi_m_axi_ARID;
  assign m_axi_in_11_ARLEN = in_11__m_axi_m_axi_ARLEN;
  assign m_axi_in_11_ARLOCK = in_11__m_axi_m_axi_ARLOCK;
  assign m_axi_in_11_ARPROT = in_11__m_axi_m_axi_ARPROT;
  assign m_axi_in_11_ARQOS = in_11__m_axi_m_axi_ARQOS;
  assign in_11__m_axi_m_axi_ARREADY = m_axi_in_11_ARREADY;
  assign m_axi_in_11_ARSIZE = in_11__m_axi_m_axi_ARSIZE;
  assign m_axi_in_11_ARVALID = in_11__m_axi_m_axi_ARVALID;
  assign m_axi_in_11_AWADDR = in_11__m_axi_m_axi_AWADDR;
  assign m_axi_in_11_AWBURST = in_11__m_axi_m_axi_AWBURST;
  assign m_axi_in_11_AWCACHE = in_11__m_axi_m_axi_AWCACHE;
  assign m_axi_in_11_AWID = in_11__m_axi_m_axi_AWID;
  assign m_axi_in_11_AWLEN = in_11__m_axi_m_axi_AWLEN;
  assign m_axi_in_11_AWLOCK = in_11__m_axi_m_axi_AWLOCK;
  assign m_axi_in_11_AWPROT = in_11__m_axi_m_axi_AWPROT;
  assign m_axi_in_11_AWQOS = in_11__m_axi_m_axi_AWQOS;
  assign in_11__m_axi_m_axi_AWREADY = m_axi_in_11_AWREADY;
  assign m_axi_in_11_AWSIZE = in_11__m_axi_m_axi_AWSIZE;
  assign m_axi_in_11_AWVALID = in_11__m_axi_m_axi_AWVALID;
  assign in_11__m_axi_m_axi_BID = m_axi_in_11_BID;
  assign m_axi_in_11_BREADY = in_11__m_axi_m_axi_BREADY;
  assign in_11__m_axi_m_axi_BRESP = m_axi_in_11_BRESP;
  assign in_11__m_axi_m_axi_BVALID = m_axi_in_11_BVALID;
  assign in_11__m_axi_m_axi_RDATA = m_axi_in_11_RDATA;
  assign in_11__m_axi_m_axi_RID = m_axi_in_11_RID;
  assign in_11__m_axi_m_axi_RLAST = m_axi_in_11_RLAST;
  assign m_axi_in_11_RREADY = in_11__m_axi_m_axi_RREADY;
  assign in_11__m_axi_m_axi_RRESP = m_axi_in_11_RRESP;
  assign in_11__m_axi_m_axi_RVALID = m_axi_in_11_RVALID;
  assign m_axi_in_11_WDATA = in_11__m_axi_m_axi_WDATA;
  assign m_axi_in_11_WLAST = in_11__m_axi_m_axi_WLAST;
  assign in_11__m_axi_m_axi_WREADY = m_axi_in_11_WREADY;
  assign m_axi_in_11_WSTRB = in_11__m_axi_m_axi_WSTRB;
  assign m_axi_in_11_WVALID = in_11__m_axi_m_axi_WVALID;
  assign in_11__m_axi_read_addr_din = in_11_read_addr__din;
  assign in_11_read_addr__full_n = in_11__m_axi_read_addr_full_n;
  assign in_11__m_axi_read_addr_write = in_11_read_addr__write;
  assign in_11_read_data__dout = in_11__m_axi_read_data_dout;
  assign in_11_read_data__empty_n = in_11__m_axi_read_data_empty_n;
  assign in_11__m_axi_read_data_read = in_11_read_data__read;
  assign in_11__m_axi_rst = ~ ap_rst_n;
  assign in_11__m_axi_write_addr_din = in_11_write_addr__din;
  assign in_11_write_addr__full_n = in_11__m_axi_write_addr_full_n;
  assign in_11__m_axi_write_addr_write = in_11_write_addr__write;
  assign in_11__m_axi_write_data_din = in_11_write_data__din;
  assign in_11_write_data__full_n = in_11__m_axi_write_data_full_n;
  assign in_11__m_axi_write_data_write = in_11_write_data__write;
  assign in_11_write_resp__dout = in_11__m_axi_write_resp_dout;
  assign in_11_write_resp__empty_n = in_11__m_axi_write_resp_empty_n;
  assign in_11__m_axi_write_resp_read = in_11_write_resp__read;
  assign in_12__m_axi_clk = ap_clk;
  assign m_axi_in_12_ARADDR = in_12__m_axi_m_axi_ARADDR;
  assign m_axi_in_12_ARBURST = in_12__m_axi_m_axi_ARBURST;
  assign m_axi_in_12_ARCACHE = in_12__m_axi_m_axi_ARCACHE;
  assign m_axi_in_12_ARID = in_12__m_axi_m_axi_ARID;
  assign m_axi_in_12_ARLEN = in_12__m_axi_m_axi_ARLEN;
  assign m_axi_in_12_ARLOCK = in_12__m_axi_m_axi_ARLOCK;
  assign m_axi_in_12_ARPROT = in_12__m_axi_m_axi_ARPROT;
  assign m_axi_in_12_ARQOS = in_12__m_axi_m_axi_ARQOS;
  assign in_12__m_axi_m_axi_ARREADY = m_axi_in_12_ARREADY;
  assign m_axi_in_12_ARSIZE = in_12__m_axi_m_axi_ARSIZE;
  assign m_axi_in_12_ARVALID = in_12__m_axi_m_axi_ARVALID;
  assign m_axi_in_12_AWADDR = in_12__m_axi_m_axi_AWADDR;
  assign m_axi_in_12_AWBURST = in_12__m_axi_m_axi_AWBURST;
  assign m_axi_in_12_AWCACHE = in_12__m_axi_m_axi_AWCACHE;
  assign m_axi_in_12_AWID = in_12__m_axi_m_axi_AWID;
  assign m_axi_in_12_AWLEN = in_12__m_axi_m_axi_AWLEN;
  assign m_axi_in_12_AWLOCK = in_12__m_axi_m_axi_AWLOCK;
  assign m_axi_in_12_AWPROT = in_12__m_axi_m_axi_AWPROT;
  assign m_axi_in_12_AWQOS = in_12__m_axi_m_axi_AWQOS;
  assign in_12__m_axi_m_axi_AWREADY = m_axi_in_12_AWREADY;
  assign m_axi_in_12_AWSIZE = in_12__m_axi_m_axi_AWSIZE;
  assign m_axi_in_12_AWVALID = in_12__m_axi_m_axi_AWVALID;
  assign in_12__m_axi_m_axi_BID = m_axi_in_12_BID;
  assign m_axi_in_12_BREADY = in_12__m_axi_m_axi_BREADY;
  assign in_12__m_axi_m_axi_BRESP = m_axi_in_12_BRESP;
  assign in_12__m_axi_m_axi_BVALID = m_axi_in_12_BVALID;
  assign in_12__m_axi_m_axi_RDATA = m_axi_in_12_RDATA;
  assign in_12__m_axi_m_axi_RID = m_axi_in_12_RID;
  assign in_12__m_axi_m_axi_RLAST = m_axi_in_12_RLAST;
  assign m_axi_in_12_RREADY = in_12__m_axi_m_axi_RREADY;
  assign in_12__m_axi_m_axi_RRESP = m_axi_in_12_RRESP;
  assign in_12__m_axi_m_axi_RVALID = m_axi_in_12_RVALID;
  assign m_axi_in_12_WDATA = in_12__m_axi_m_axi_WDATA;
  assign m_axi_in_12_WLAST = in_12__m_axi_m_axi_WLAST;
  assign in_12__m_axi_m_axi_WREADY = m_axi_in_12_WREADY;
  assign m_axi_in_12_WSTRB = in_12__m_axi_m_axi_WSTRB;
  assign m_axi_in_12_WVALID = in_12__m_axi_m_axi_WVALID;
  assign in_12__m_axi_read_addr_din = in_12_read_addr__din;
  assign in_12_read_addr__full_n = in_12__m_axi_read_addr_full_n;
  assign in_12__m_axi_read_addr_write = in_12_read_addr__write;
  assign in_12_read_data__dout = in_12__m_axi_read_data_dout;
  assign in_12_read_data__empty_n = in_12__m_axi_read_data_empty_n;
  assign in_12__m_axi_read_data_read = in_12_read_data__read;
  assign in_12__m_axi_rst = ~ ap_rst_n;
  assign in_12__m_axi_write_addr_din = in_12_write_addr__din;
  assign in_12_write_addr__full_n = in_12__m_axi_write_addr_full_n;
  assign in_12__m_axi_write_addr_write = in_12_write_addr__write;
  assign in_12__m_axi_write_data_din = in_12_write_data__din;
  assign in_12_write_data__full_n = in_12__m_axi_write_data_full_n;
  assign in_12__m_axi_write_data_write = in_12_write_data__write;
  assign in_12_write_resp__dout = in_12__m_axi_write_resp_dout;
  assign in_12_write_resp__empty_n = in_12__m_axi_write_resp_empty_n;
  assign in_12__m_axi_write_resp_read = in_12_write_resp__read;
  assign in_13__m_axi_clk = ap_clk;
  assign m_axi_in_13_ARADDR = in_13__m_axi_m_axi_ARADDR;
  assign m_axi_in_13_ARBURST = in_13__m_axi_m_axi_ARBURST;
  assign m_axi_in_13_ARCACHE = in_13__m_axi_m_axi_ARCACHE;
  assign m_axi_in_13_ARID = in_13__m_axi_m_axi_ARID;
  assign m_axi_in_13_ARLEN = in_13__m_axi_m_axi_ARLEN;
  assign m_axi_in_13_ARLOCK = in_13__m_axi_m_axi_ARLOCK;
  assign m_axi_in_13_ARPROT = in_13__m_axi_m_axi_ARPROT;
  assign m_axi_in_13_ARQOS = in_13__m_axi_m_axi_ARQOS;
  assign in_13__m_axi_m_axi_ARREADY = m_axi_in_13_ARREADY;
  assign m_axi_in_13_ARSIZE = in_13__m_axi_m_axi_ARSIZE;
  assign m_axi_in_13_ARVALID = in_13__m_axi_m_axi_ARVALID;
  assign m_axi_in_13_AWADDR = in_13__m_axi_m_axi_AWADDR;
  assign m_axi_in_13_AWBURST = in_13__m_axi_m_axi_AWBURST;
  assign m_axi_in_13_AWCACHE = in_13__m_axi_m_axi_AWCACHE;
  assign m_axi_in_13_AWID = in_13__m_axi_m_axi_AWID;
  assign m_axi_in_13_AWLEN = in_13__m_axi_m_axi_AWLEN;
  assign m_axi_in_13_AWLOCK = in_13__m_axi_m_axi_AWLOCK;
  assign m_axi_in_13_AWPROT = in_13__m_axi_m_axi_AWPROT;
  assign m_axi_in_13_AWQOS = in_13__m_axi_m_axi_AWQOS;
  assign in_13__m_axi_m_axi_AWREADY = m_axi_in_13_AWREADY;
  assign m_axi_in_13_AWSIZE = in_13__m_axi_m_axi_AWSIZE;
  assign m_axi_in_13_AWVALID = in_13__m_axi_m_axi_AWVALID;
  assign in_13__m_axi_m_axi_BID = m_axi_in_13_BID;
  assign m_axi_in_13_BREADY = in_13__m_axi_m_axi_BREADY;
  assign in_13__m_axi_m_axi_BRESP = m_axi_in_13_BRESP;
  assign in_13__m_axi_m_axi_BVALID = m_axi_in_13_BVALID;
  assign in_13__m_axi_m_axi_RDATA = m_axi_in_13_RDATA;
  assign in_13__m_axi_m_axi_RID = m_axi_in_13_RID;
  assign in_13__m_axi_m_axi_RLAST = m_axi_in_13_RLAST;
  assign m_axi_in_13_RREADY = in_13__m_axi_m_axi_RREADY;
  assign in_13__m_axi_m_axi_RRESP = m_axi_in_13_RRESP;
  assign in_13__m_axi_m_axi_RVALID = m_axi_in_13_RVALID;
  assign m_axi_in_13_WDATA = in_13__m_axi_m_axi_WDATA;
  assign m_axi_in_13_WLAST = in_13__m_axi_m_axi_WLAST;
  assign in_13__m_axi_m_axi_WREADY = m_axi_in_13_WREADY;
  assign m_axi_in_13_WSTRB = in_13__m_axi_m_axi_WSTRB;
  assign m_axi_in_13_WVALID = in_13__m_axi_m_axi_WVALID;
  assign in_13__m_axi_read_addr_din = in_13_read_addr__din;
  assign in_13_read_addr__full_n = in_13__m_axi_read_addr_full_n;
  assign in_13__m_axi_read_addr_write = in_13_read_addr__write;
  assign in_13_read_data__dout = in_13__m_axi_read_data_dout;
  assign in_13_read_data__empty_n = in_13__m_axi_read_data_empty_n;
  assign in_13__m_axi_read_data_read = in_13_read_data__read;
  assign in_13__m_axi_rst = ~ ap_rst_n;
  assign in_13__m_axi_write_addr_din = in_13_write_addr__din;
  assign in_13_write_addr__full_n = in_13__m_axi_write_addr_full_n;
  assign in_13__m_axi_write_addr_write = in_13_write_addr__write;
  assign in_13__m_axi_write_data_din = in_13_write_data__din;
  assign in_13_write_data__full_n = in_13__m_axi_write_data_full_n;
  assign in_13__m_axi_write_data_write = in_13_write_data__write;
  assign in_13_write_resp__dout = in_13__m_axi_write_resp_dout;
  assign in_13_write_resp__empty_n = in_13__m_axi_write_resp_empty_n;
  assign in_13__m_axi_write_resp_read = in_13_write_resp__read;
  assign in_14__m_axi_clk = ap_clk;
  assign m_axi_in_14_ARADDR = in_14__m_axi_m_axi_ARADDR;
  assign m_axi_in_14_ARBURST = in_14__m_axi_m_axi_ARBURST;
  assign m_axi_in_14_ARCACHE = in_14__m_axi_m_axi_ARCACHE;
  assign m_axi_in_14_ARID = in_14__m_axi_m_axi_ARID;
  assign m_axi_in_14_ARLEN = in_14__m_axi_m_axi_ARLEN;
  assign m_axi_in_14_ARLOCK = in_14__m_axi_m_axi_ARLOCK;
  assign m_axi_in_14_ARPROT = in_14__m_axi_m_axi_ARPROT;
  assign m_axi_in_14_ARQOS = in_14__m_axi_m_axi_ARQOS;
  assign in_14__m_axi_m_axi_ARREADY = m_axi_in_14_ARREADY;
  assign m_axi_in_14_ARSIZE = in_14__m_axi_m_axi_ARSIZE;
  assign m_axi_in_14_ARVALID = in_14__m_axi_m_axi_ARVALID;
  assign m_axi_in_14_AWADDR = in_14__m_axi_m_axi_AWADDR;
  assign m_axi_in_14_AWBURST = in_14__m_axi_m_axi_AWBURST;
  assign m_axi_in_14_AWCACHE = in_14__m_axi_m_axi_AWCACHE;
  assign m_axi_in_14_AWID = in_14__m_axi_m_axi_AWID;
  assign m_axi_in_14_AWLEN = in_14__m_axi_m_axi_AWLEN;
  assign m_axi_in_14_AWLOCK = in_14__m_axi_m_axi_AWLOCK;
  assign m_axi_in_14_AWPROT = in_14__m_axi_m_axi_AWPROT;
  assign m_axi_in_14_AWQOS = in_14__m_axi_m_axi_AWQOS;
  assign in_14__m_axi_m_axi_AWREADY = m_axi_in_14_AWREADY;
  assign m_axi_in_14_AWSIZE = in_14__m_axi_m_axi_AWSIZE;
  assign m_axi_in_14_AWVALID = in_14__m_axi_m_axi_AWVALID;
  assign in_14__m_axi_m_axi_BID = m_axi_in_14_BID;
  assign m_axi_in_14_BREADY = in_14__m_axi_m_axi_BREADY;
  assign in_14__m_axi_m_axi_BRESP = m_axi_in_14_BRESP;
  assign in_14__m_axi_m_axi_BVALID = m_axi_in_14_BVALID;
  assign in_14__m_axi_m_axi_RDATA = m_axi_in_14_RDATA;
  assign in_14__m_axi_m_axi_RID = m_axi_in_14_RID;
  assign in_14__m_axi_m_axi_RLAST = m_axi_in_14_RLAST;
  assign m_axi_in_14_RREADY = in_14__m_axi_m_axi_RREADY;
  assign in_14__m_axi_m_axi_RRESP = m_axi_in_14_RRESP;
  assign in_14__m_axi_m_axi_RVALID = m_axi_in_14_RVALID;
  assign m_axi_in_14_WDATA = in_14__m_axi_m_axi_WDATA;
  assign m_axi_in_14_WLAST = in_14__m_axi_m_axi_WLAST;
  assign in_14__m_axi_m_axi_WREADY = m_axi_in_14_WREADY;
  assign m_axi_in_14_WSTRB = in_14__m_axi_m_axi_WSTRB;
  assign m_axi_in_14_WVALID = in_14__m_axi_m_axi_WVALID;
  assign in_14__m_axi_read_addr_din = in_14_read_addr__din;
  assign in_14_read_addr__full_n = in_14__m_axi_read_addr_full_n;
  assign in_14__m_axi_read_addr_write = in_14_read_addr__write;
  assign in_14_read_data__dout = in_14__m_axi_read_data_dout;
  assign in_14_read_data__empty_n = in_14__m_axi_read_data_empty_n;
  assign in_14__m_axi_read_data_read = in_14_read_data__read;
  assign in_14__m_axi_rst = ~ ap_rst_n;
  assign in_14__m_axi_write_addr_din = in_14_write_addr__din;
  assign in_14_write_addr__full_n = in_14__m_axi_write_addr_full_n;
  assign in_14__m_axi_write_addr_write = in_14_write_addr__write;
  assign in_14__m_axi_write_data_din = in_14_write_data__din;
  assign in_14_write_data__full_n = in_14__m_axi_write_data_full_n;
  assign in_14__m_axi_write_data_write = in_14_write_data__write;
  assign in_14_write_resp__dout = in_14__m_axi_write_resp_dout;
  assign in_14_write_resp__empty_n = in_14__m_axi_write_resp_empty_n;
  assign in_14__m_axi_write_resp_read = in_14_write_resp__read;
  assign in_15__m_axi_clk = ap_clk;
  assign m_axi_in_15_ARADDR = in_15__m_axi_m_axi_ARADDR;
  assign m_axi_in_15_ARBURST = in_15__m_axi_m_axi_ARBURST;
  assign m_axi_in_15_ARCACHE = in_15__m_axi_m_axi_ARCACHE;
  assign m_axi_in_15_ARID = in_15__m_axi_m_axi_ARID;
  assign m_axi_in_15_ARLEN = in_15__m_axi_m_axi_ARLEN;
  assign m_axi_in_15_ARLOCK = in_15__m_axi_m_axi_ARLOCK;
  assign m_axi_in_15_ARPROT = in_15__m_axi_m_axi_ARPROT;
  assign m_axi_in_15_ARQOS = in_15__m_axi_m_axi_ARQOS;
  assign in_15__m_axi_m_axi_ARREADY = m_axi_in_15_ARREADY;
  assign m_axi_in_15_ARSIZE = in_15__m_axi_m_axi_ARSIZE;
  assign m_axi_in_15_ARVALID = in_15__m_axi_m_axi_ARVALID;
  assign m_axi_in_15_AWADDR = in_15__m_axi_m_axi_AWADDR;
  assign m_axi_in_15_AWBURST = in_15__m_axi_m_axi_AWBURST;
  assign m_axi_in_15_AWCACHE = in_15__m_axi_m_axi_AWCACHE;
  assign m_axi_in_15_AWID = in_15__m_axi_m_axi_AWID;
  assign m_axi_in_15_AWLEN = in_15__m_axi_m_axi_AWLEN;
  assign m_axi_in_15_AWLOCK = in_15__m_axi_m_axi_AWLOCK;
  assign m_axi_in_15_AWPROT = in_15__m_axi_m_axi_AWPROT;
  assign m_axi_in_15_AWQOS = in_15__m_axi_m_axi_AWQOS;
  assign in_15__m_axi_m_axi_AWREADY = m_axi_in_15_AWREADY;
  assign m_axi_in_15_AWSIZE = in_15__m_axi_m_axi_AWSIZE;
  assign m_axi_in_15_AWVALID = in_15__m_axi_m_axi_AWVALID;
  assign in_15__m_axi_m_axi_BID = m_axi_in_15_BID;
  assign m_axi_in_15_BREADY = in_15__m_axi_m_axi_BREADY;
  assign in_15__m_axi_m_axi_BRESP = m_axi_in_15_BRESP;
  assign in_15__m_axi_m_axi_BVALID = m_axi_in_15_BVALID;
  assign in_15__m_axi_m_axi_RDATA = m_axi_in_15_RDATA;
  assign in_15__m_axi_m_axi_RID = m_axi_in_15_RID;
  assign in_15__m_axi_m_axi_RLAST = m_axi_in_15_RLAST;
  assign m_axi_in_15_RREADY = in_15__m_axi_m_axi_RREADY;
  assign in_15__m_axi_m_axi_RRESP = m_axi_in_15_RRESP;
  assign in_15__m_axi_m_axi_RVALID = m_axi_in_15_RVALID;
  assign m_axi_in_15_WDATA = in_15__m_axi_m_axi_WDATA;
  assign m_axi_in_15_WLAST = in_15__m_axi_m_axi_WLAST;
  assign in_15__m_axi_m_axi_WREADY = m_axi_in_15_WREADY;
  assign m_axi_in_15_WSTRB = in_15__m_axi_m_axi_WSTRB;
  assign m_axi_in_15_WVALID = in_15__m_axi_m_axi_WVALID;
  assign in_15__m_axi_read_addr_din = in_15_read_addr__din;
  assign in_15_read_addr__full_n = in_15__m_axi_read_addr_full_n;
  assign in_15__m_axi_read_addr_write = in_15_read_addr__write;
  assign in_15_read_data__dout = in_15__m_axi_read_data_dout;
  assign in_15_read_data__empty_n = in_15__m_axi_read_data_empty_n;
  assign in_15__m_axi_read_data_read = in_15_read_data__read;
  assign in_15__m_axi_rst = ~ ap_rst_n;
  assign in_15__m_axi_write_addr_din = in_15_write_addr__din;
  assign in_15_write_addr__full_n = in_15__m_axi_write_addr_full_n;
  assign in_15__m_axi_write_addr_write = in_15_write_addr__write;
  assign in_15__m_axi_write_data_din = in_15_write_data__din;
  assign in_15_write_data__full_n = in_15__m_axi_write_data_full_n;
  assign in_15__m_axi_write_data_write = in_15_write_data__write;
  assign in_15_write_resp__dout = in_15__m_axi_write_resp_dout;
  assign in_15_write_resp__empty_n = in_15__m_axi_write_resp_empty_n;
  assign in_15__m_axi_write_resp_read = in_15_write_resp__read;
  assign in_16__m_axi_clk = ap_clk;
  assign m_axi_in_16_ARADDR = in_16__m_axi_m_axi_ARADDR;
  assign m_axi_in_16_ARBURST = in_16__m_axi_m_axi_ARBURST;
  assign m_axi_in_16_ARCACHE = in_16__m_axi_m_axi_ARCACHE;
  assign m_axi_in_16_ARID = in_16__m_axi_m_axi_ARID;
  assign m_axi_in_16_ARLEN = in_16__m_axi_m_axi_ARLEN;
  assign m_axi_in_16_ARLOCK = in_16__m_axi_m_axi_ARLOCK;
  assign m_axi_in_16_ARPROT = in_16__m_axi_m_axi_ARPROT;
  assign m_axi_in_16_ARQOS = in_16__m_axi_m_axi_ARQOS;
  assign in_16__m_axi_m_axi_ARREADY = m_axi_in_16_ARREADY;
  assign m_axi_in_16_ARSIZE = in_16__m_axi_m_axi_ARSIZE;
  assign m_axi_in_16_ARVALID = in_16__m_axi_m_axi_ARVALID;
  assign m_axi_in_16_AWADDR = in_16__m_axi_m_axi_AWADDR;
  assign m_axi_in_16_AWBURST = in_16__m_axi_m_axi_AWBURST;
  assign m_axi_in_16_AWCACHE = in_16__m_axi_m_axi_AWCACHE;
  assign m_axi_in_16_AWID = in_16__m_axi_m_axi_AWID;
  assign m_axi_in_16_AWLEN = in_16__m_axi_m_axi_AWLEN;
  assign m_axi_in_16_AWLOCK = in_16__m_axi_m_axi_AWLOCK;
  assign m_axi_in_16_AWPROT = in_16__m_axi_m_axi_AWPROT;
  assign m_axi_in_16_AWQOS = in_16__m_axi_m_axi_AWQOS;
  assign in_16__m_axi_m_axi_AWREADY = m_axi_in_16_AWREADY;
  assign m_axi_in_16_AWSIZE = in_16__m_axi_m_axi_AWSIZE;
  assign m_axi_in_16_AWVALID = in_16__m_axi_m_axi_AWVALID;
  assign in_16__m_axi_m_axi_BID = m_axi_in_16_BID;
  assign m_axi_in_16_BREADY = in_16__m_axi_m_axi_BREADY;
  assign in_16__m_axi_m_axi_BRESP = m_axi_in_16_BRESP;
  assign in_16__m_axi_m_axi_BVALID = m_axi_in_16_BVALID;
  assign in_16__m_axi_m_axi_RDATA = m_axi_in_16_RDATA;
  assign in_16__m_axi_m_axi_RID = m_axi_in_16_RID;
  assign in_16__m_axi_m_axi_RLAST = m_axi_in_16_RLAST;
  assign m_axi_in_16_RREADY = in_16__m_axi_m_axi_RREADY;
  assign in_16__m_axi_m_axi_RRESP = m_axi_in_16_RRESP;
  assign in_16__m_axi_m_axi_RVALID = m_axi_in_16_RVALID;
  assign m_axi_in_16_WDATA = in_16__m_axi_m_axi_WDATA;
  assign m_axi_in_16_WLAST = in_16__m_axi_m_axi_WLAST;
  assign in_16__m_axi_m_axi_WREADY = m_axi_in_16_WREADY;
  assign m_axi_in_16_WSTRB = in_16__m_axi_m_axi_WSTRB;
  assign m_axi_in_16_WVALID = in_16__m_axi_m_axi_WVALID;
  assign in_16__m_axi_read_addr_din = in_16_read_addr__din;
  assign in_16_read_addr__full_n = in_16__m_axi_read_addr_full_n;
  assign in_16__m_axi_read_addr_write = in_16_read_addr__write;
  assign in_16_read_data__dout = in_16__m_axi_read_data_dout;
  assign in_16_read_data__empty_n = in_16__m_axi_read_data_empty_n;
  assign in_16__m_axi_read_data_read = in_16_read_data__read;
  assign in_16__m_axi_rst = ~ ap_rst_n;
  assign in_16__m_axi_write_addr_din = in_16_write_addr__din;
  assign in_16_write_addr__full_n = in_16__m_axi_write_addr_full_n;
  assign in_16__m_axi_write_addr_write = in_16_write_addr__write;
  assign in_16__m_axi_write_data_din = in_16_write_data__din;
  assign in_16_write_data__full_n = in_16__m_axi_write_data_full_n;
  assign in_16__m_axi_write_data_write = in_16_write_data__write;
  assign in_16_write_resp__dout = in_16__m_axi_write_resp_dout;
  assign in_16_write_resp__empty_n = in_16__m_axi_write_resp_empty_n;
  assign in_16__m_axi_write_resp_read = in_16_write_resp__read;
  assign in_17__m_axi_clk = ap_clk;
  assign m_axi_in_17_ARADDR = in_17__m_axi_m_axi_ARADDR;
  assign m_axi_in_17_ARBURST = in_17__m_axi_m_axi_ARBURST;
  assign m_axi_in_17_ARCACHE = in_17__m_axi_m_axi_ARCACHE;
  assign m_axi_in_17_ARID = in_17__m_axi_m_axi_ARID;
  assign m_axi_in_17_ARLEN = in_17__m_axi_m_axi_ARLEN;
  assign m_axi_in_17_ARLOCK = in_17__m_axi_m_axi_ARLOCK;
  assign m_axi_in_17_ARPROT = in_17__m_axi_m_axi_ARPROT;
  assign m_axi_in_17_ARQOS = in_17__m_axi_m_axi_ARQOS;
  assign in_17__m_axi_m_axi_ARREADY = m_axi_in_17_ARREADY;
  assign m_axi_in_17_ARSIZE = in_17__m_axi_m_axi_ARSIZE;
  assign m_axi_in_17_ARVALID = in_17__m_axi_m_axi_ARVALID;
  assign m_axi_in_17_AWADDR = in_17__m_axi_m_axi_AWADDR;
  assign m_axi_in_17_AWBURST = in_17__m_axi_m_axi_AWBURST;
  assign m_axi_in_17_AWCACHE = in_17__m_axi_m_axi_AWCACHE;
  assign m_axi_in_17_AWID = in_17__m_axi_m_axi_AWID;
  assign m_axi_in_17_AWLEN = in_17__m_axi_m_axi_AWLEN;
  assign m_axi_in_17_AWLOCK = in_17__m_axi_m_axi_AWLOCK;
  assign m_axi_in_17_AWPROT = in_17__m_axi_m_axi_AWPROT;
  assign m_axi_in_17_AWQOS = in_17__m_axi_m_axi_AWQOS;
  assign in_17__m_axi_m_axi_AWREADY = m_axi_in_17_AWREADY;
  assign m_axi_in_17_AWSIZE = in_17__m_axi_m_axi_AWSIZE;
  assign m_axi_in_17_AWVALID = in_17__m_axi_m_axi_AWVALID;
  assign in_17__m_axi_m_axi_BID = m_axi_in_17_BID;
  assign m_axi_in_17_BREADY = in_17__m_axi_m_axi_BREADY;
  assign in_17__m_axi_m_axi_BRESP = m_axi_in_17_BRESP;
  assign in_17__m_axi_m_axi_BVALID = m_axi_in_17_BVALID;
  assign in_17__m_axi_m_axi_RDATA = m_axi_in_17_RDATA;
  assign in_17__m_axi_m_axi_RID = m_axi_in_17_RID;
  assign in_17__m_axi_m_axi_RLAST = m_axi_in_17_RLAST;
  assign m_axi_in_17_RREADY = in_17__m_axi_m_axi_RREADY;
  assign in_17__m_axi_m_axi_RRESP = m_axi_in_17_RRESP;
  assign in_17__m_axi_m_axi_RVALID = m_axi_in_17_RVALID;
  assign m_axi_in_17_WDATA = in_17__m_axi_m_axi_WDATA;
  assign m_axi_in_17_WLAST = in_17__m_axi_m_axi_WLAST;
  assign in_17__m_axi_m_axi_WREADY = m_axi_in_17_WREADY;
  assign m_axi_in_17_WSTRB = in_17__m_axi_m_axi_WSTRB;
  assign m_axi_in_17_WVALID = in_17__m_axi_m_axi_WVALID;
  assign in_17__m_axi_read_addr_din = in_17_read_addr__din;
  assign in_17_read_addr__full_n = in_17__m_axi_read_addr_full_n;
  assign in_17__m_axi_read_addr_write = in_17_read_addr__write;
  assign in_17_read_data__dout = in_17__m_axi_read_data_dout;
  assign in_17_read_data__empty_n = in_17__m_axi_read_data_empty_n;
  assign in_17__m_axi_read_data_read = in_17_read_data__read;
  assign in_17__m_axi_rst = ~ ap_rst_n;
  assign in_17__m_axi_write_addr_din = in_17_write_addr__din;
  assign in_17_write_addr__full_n = in_17__m_axi_write_addr_full_n;
  assign in_17__m_axi_write_addr_write = in_17_write_addr__write;
  assign in_17__m_axi_write_data_din = in_17_write_data__din;
  assign in_17_write_data__full_n = in_17__m_axi_write_data_full_n;
  assign in_17__m_axi_write_data_write = in_17_write_data__write;
  assign in_17_write_resp__dout = in_17__m_axi_write_resp_dout;
  assign in_17_write_resp__empty_n = in_17__m_axi_write_resp_empty_n;
  assign in_17__m_axi_write_resp_read = in_17_write_resp__read;
  assign in_18__m_axi_clk = ap_clk;
  assign m_axi_in_18_ARADDR = in_18__m_axi_m_axi_ARADDR;
  assign m_axi_in_18_ARBURST = in_18__m_axi_m_axi_ARBURST;
  assign m_axi_in_18_ARCACHE = in_18__m_axi_m_axi_ARCACHE;
  assign m_axi_in_18_ARID = in_18__m_axi_m_axi_ARID;
  assign m_axi_in_18_ARLEN = in_18__m_axi_m_axi_ARLEN;
  assign m_axi_in_18_ARLOCK = in_18__m_axi_m_axi_ARLOCK;
  assign m_axi_in_18_ARPROT = in_18__m_axi_m_axi_ARPROT;
  assign m_axi_in_18_ARQOS = in_18__m_axi_m_axi_ARQOS;
  assign in_18__m_axi_m_axi_ARREADY = m_axi_in_18_ARREADY;
  assign m_axi_in_18_ARSIZE = in_18__m_axi_m_axi_ARSIZE;
  assign m_axi_in_18_ARVALID = in_18__m_axi_m_axi_ARVALID;
  assign m_axi_in_18_AWADDR = in_18__m_axi_m_axi_AWADDR;
  assign m_axi_in_18_AWBURST = in_18__m_axi_m_axi_AWBURST;
  assign m_axi_in_18_AWCACHE = in_18__m_axi_m_axi_AWCACHE;
  assign m_axi_in_18_AWID = in_18__m_axi_m_axi_AWID;
  assign m_axi_in_18_AWLEN = in_18__m_axi_m_axi_AWLEN;
  assign m_axi_in_18_AWLOCK = in_18__m_axi_m_axi_AWLOCK;
  assign m_axi_in_18_AWPROT = in_18__m_axi_m_axi_AWPROT;
  assign m_axi_in_18_AWQOS = in_18__m_axi_m_axi_AWQOS;
  assign in_18__m_axi_m_axi_AWREADY = m_axi_in_18_AWREADY;
  assign m_axi_in_18_AWSIZE = in_18__m_axi_m_axi_AWSIZE;
  assign m_axi_in_18_AWVALID = in_18__m_axi_m_axi_AWVALID;
  assign in_18__m_axi_m_axi_BID = m_axi_in_18_BID;
  assign m_axi_in_18_BREADY = in_18__m_axi_m_axi_BREADY;
  assign in_18__m_axi_m_axi_BRESP = m_axi_in_18_BRESP;
  assign in_18__m_axi_m_axi_BVALID = m_axi_in_18_BVALID;
  assign in_18__m_axi_m_axi_RDATA = m_axi_in_18_RDATA;
  assign in_18__m_axi_m_axi_RID = m_axi_in_18_RID;
  assign in_18__m_axi_m_axi_RLAST = m_axi_in_18_RLAST;
  assign m_axi_in_18_RREADY = in_18__m_axi_m_axi_RREADY;
  assign in_18__m_axi_m_axi_RRESP = m_axi_in_18_RRESP;
  assign in_18__m_axi_m_axi_RVALID = m_axi_in_18_RVALID;
  assign m_axi_in_18_WDATA = in_18__m_axi_m_axi_WDATA;
  assign m_axi_in_18_WLAST = in_18__m_axi_m_axi_WLAST;
  assign in_18__m_axi_m_axi_WREADY = m_axi_in_18_WREADY;
  assign m_axi_in_18_WSTRB = in_18__m_axi_m_axi_WSTRB;
  assign m_axi_in_18_WVALID = in_18__m_axi_m_axi_WVALID;
  assign in_18__m_axi_read_addr_din = in_18_read_addr__din;
  assign in_18_read_addr__full_n = in_18__m_axi_read_addr_full_n;
  assign in_18__m_axi_read_addr_write = in_18_read_addr__write;
  assign in_18_read_data__dout = in_18__m_axi_read_data_dout;
  assign in_18_read_data__empty_n = in_18__m_axi_read_data_empty_n;
  assign in_18__m_axi_read_data_read = in_18_read_data__read;
  assign in_18__m_axi_rst = ~ ap_rst_n;
  assign in_18__m_axi_write_addr_din = in_18_write_addr__din;
  assign in_18_write_addr__full_n = in_18__m_axi_write_addr_full_n;
  assign in_18__m_axi_write_addr_write = in_18_write_addr__write;
  assign in_18__m_axi_write_data_din = in_18_write_data__din;
  assign in_18_write_data__full_n = in_18__m_axi_write_data_full_n;
  assign in_18__m_axi_write_data_write = in_18_write_data__write;
  assign in_18_write_resp__dout = in_18__m_axi_write_resp_dout;
  assign in_18_write_resp__empty_n = in_18__m_axi_write_resp_empty_n;
  assign in_18__m_axi_write_resp_read = in_18_write_resp__read;
  assign in_19__m_axi_clk = ap_clk;
  assign m_axi_in_19_ARADDR = in_19__m_axi_m_axi_ARADDR;
  assign m_axi_in_19_ARBURST = in_19__m_axi_m_axi_ARBURST;
  assign m_axi_in_19_ARCACHE = in_19__m_axi_m_axi_ARCACHE;
  assign m_axi_in_19_ARID = in_19__m_axi_m_axi_ARID;
  assign m_axi_in_19_ARLEN = in_19__m_axi_m_axi_ARLEN;
  assign m_axi_in_19_ARLOCK = in_19__m_axi_m_axi_ARLOCK;
  assign m_axi_in_19_ARPROT = in_19__m_axi_m_axi_ARPROT;
  assign m_axi_in_19_ARQOS = in_19__m_axi_m_axi_ARQOS;
  assign in_19__m_axi_m_axi_ARREADY = m_axi_in_19_ARREADY;
  assign m_axi_in_19_ARSIZE = in_19__m_axi_m_axi_ARSIZE;
  assign m_axi_in_19_ARVALID = in_19__m_axi_m_axi_ARVALID;
  assign m_axi_in_19_AWADDR = in_19__m_axi_m_axi_AWADDR;
  assign m_axi_in_19_AWBURST = in_19__m_axi_m_axi_AWBURST;
  assign m_axi_in_19_AWCACHE = in_19__m_axi_m_axi_AWCACHE;
  assign m_axi_in_19_AWID = in_19__m_axi_m_axi_AWID;
  assign m_axi_in_19_AWLEN = in_19__m_axi_m_axi_AWLEN;
  assign m_axi_in_19_AWLOCK = in_19__m_axi_m_axi_AWLOCK;
  assign m_axi_in_19_AWPROT = in_19__m_axi_m_axi_AWPROT;
  assign m_axi_in_19_AWQOS = in_19__m_axi_m_axi_AWQOS;
  assign in_19__m_axi_m_axi_AWREADY = m_axi_in_19_AWREADY;
  assign m_axi_in_19_AWSIZE = in_19__m_axi_m_axi_AWSIZE;
  assign m_axi_in_19_AWVALID = in_19__m_axi_m_axi_AWVALID;
  assign in_19__m_axi_m_axi_BID = m_axi_in_19_BID;
  assign m_axi_in_19_BREADY = in_19__m_axi_m_axi_BREADY;
  assign in_19__m_axi_m_axi_BRESP = m_axi_in_19_BRESP;
  assign in_19__m_axi_m_axi_BVALID = m_axi_in_19_BVALID;
  assign in_19__m_axi_m_axi_RDATA = m_axi_in_19_RDATA;
  assign in_19__m_axi_m_axi_RID = m_axi_in_19_RID;
  assign in_19__m_axi_m_axi_RLAST = m_axi_in_19_RLAST;
  assign m_axi_in_19_RREADY = in_19__m_axi_m_axi_RREADY;
  assign in_19__m_axi_m_axi_RRESP = m_axi_in_19_RRESP;
  assign in_19__m_axi_m_axi_RVALID = m_axi_in_19_RVALID;
  assign m_axi_in_19_WDATA = in_19__m_axi_m_axi_WDATA;
  assign m_axi_in_19_WLAST = in_19__m_axi_m_axi_WLAST;
  assign in_19__m_axi_m_axi_WREADY = m_axi_in_19_WREADY;
  assign m_axi_in_19_WSTRB = in_19__m_axi_m_axi_WSTRB;
  assign m_axi_in_19_WVALID = in_19__m_axi_m_axi_WVALID;
  assign in_19__m_axi_read_addr_din = in_19_read_addr__din;
  assign in_19_read_addr__full_n = in_19__m_axi_read_addr_full_n;
  assign in_19__m_axi_read_addr_write = in_19_read_addr__write;
  assign in_19_read_data__dout = in_19__m_axi_read_data_dout;
  assign in_19_read_data__empty_n = in_19__m_axi_read_data_empty_n;
  assign in_19__m_axi_read_data_read = in_19_read_data__read;
  assign in_19__m_axi_rst = ~ ap_rst_n;
  assign in_19__m_axi_write_addr_din = in_19_write_addr__din;
  assign in_19_write_addr__full_n = in_19__m_axi_write_addr_full_n;
  assign in_19__m_axi_write_addr_write = in_19_write_addr__write;
  assign in_19__m_axi_write_data_din = in_19_write_data__din;
  assign in_19_write_data__full_n = in_19__m_axi_write_data_full_n;
  assign in_19__m_axi_write_data_write = in_19_write_data__write;
  assign in_19_write_resp__dout = in_19__m_axi_write_resp_dout;
  assign in_19_write_resp__empty_n = in_19__m_axi_write_resp_empty_n;
  assign in_19__m_axi_write_resp_read = in_19_write_resp__read;
  assign in_2__m_axi_clk = ap_clk;
  assign m_axi_in_2_ARADDR = in_2__m_axi_m_axi_ARADDR;
  assign m_axi_in_2_ARBURST = in_2__m_axi_m_axi_ARBURST;
  assign m_axi_in_2_ARCACHE = in_2__m_axi_m_axi_ARCACHE;
  assign m_axi_in_2_ARID = in_2__m_axi_m_axi_ARID;
  assign m_axi_in_2_ARLEN = in_2__m_axi_m_axi_ARLEN;
  assign m_axi_in_2_ARLOCK = in_2__m_axi_m_axi_ARLOCK;
  assign m_axi_in_2_ARPROT = in_2__m_axi_m_axi_ARPROT;
  assign m_axi_in_2_ARQOS = in_2__m_axi_m_axi_ARQOS;
  assign in_2__m_axi_m_axi_ARREADY = m_axi_in_2_ARREADY;
  assign m_axi_in_2_ARSIZE = in_2__m_axi_m_axi_ARSIZE;
  assign m_axi_in_2_ARVALID = in_2__m_axi_m_axi_ARVALID;
  assign m_axi_in_2_AWADDR = in_2__m_axi_m_axi_AWADDR;
  assign m_axi_in_2_AWBURST = in_2__m_axi_m_axi_AWBURST;
  assign m_axi_in_2_AWCACHE = in_2__m_axi_m_axi_AWCACHE;
  assign m_axi_in_2_AWID = in_2__m_axi_m_axi_AWID;
  assign m_axi_in_2_AWLEN = in_2__m_axi_m_axi_AWLEN;
  assign m_axi_in_2_AWLOCK = in_2__m_axi_m_axi_AWLOCK;
  assign m_axi_in_2_AWPROT = in_2__m_axi_m_axi_AWPROT;
  assign m_axi_in_2_AWQOS = in_2__m_axi_m_axi_AWQOS;
  assign in_2__m_axi_m_axi_AWREADY = m_axi_in_2_AWREADY;
  assign m_axi_in_2_AWSIZE = in_2__m_axi_m_axi_AWSIZE;
  assign m_axi_in_2_AWVALID = in_2__m_axi_m_axi_AWVALID;
  assign in_2__m_axi_m_axi_BID = m_axi_in_2_BID;
  assign m_axi_in_2_BREADY = in_2__m_axi_m_axi_BREADY;
  assign in_2__m_axi_m_axi_BRESP = m_axi_in_2_BRESP;
  assign in_2__m_axi_m_axi_BVALID = m_axi_in_2_BVALID;
  assign in_2__m_axi_m_axi_RDATA = m_axi_in_2_RDATA;
  assign in_2__m_axi_m_axi_RID = m_axi_in_2_RID;
  assign in_2__m_axi_m_axi_RLAST = m_axi_in_2_RLAST;
  assign m_axi_in_2_RREADY = in_2__m_axi_m_axi_RREADY;
  assign in_2__m_axi_m_axi_RRESP = m_axi_in_2_RRESP;
  assign in_2__m_axi_m_axi_RVALID = m_axi_in_2_RVALID;
  assign m_axi_in_2_WDATA = in_2__m_axi_m_axi_WDATA;
  assign m_axi_in_2_WLAST = in_2__m_axi_m_axi_WLAST;
  assign in_2__m_axi_m_axi_WREADY = m_axi_in_2_WREADY;
  assign m_axi_in_2_WSTRB = in_2__m_axi_m_axi_WSTRB;
  assign m_axi_in_2_WVALID = in_2__m_axi_m_axi_WVALID;
  assign in_2__m_axi_read_addr_din = in_2_read_addr__din;
  assign in_2_read_addr__full_n = in_2__m_axi_read_addr_full_n;
  assign in_2__m_axi_read_addr_write = in_2_read_addr__write;
  assign in_2_read_data__dout = in_2__m_axi_read_data_dout;
  assign in_2_read_data__empty_n = in_2__m_axi_read_data_empty_n;
  assign in_2__m_axi_read_data_read = in_2_read_data__read;
  assign in_2__m_axi_rst = ~ ap_rst_n;
  assign in_2__m_axi_write_addr_din = in_2_write_addr__din;
  assign in_2_write_addr__full_n = in_2__m_axi_write_addr_full_n;
  assign in_2__m_axi_write_addr_write = in_2_write_addr__write;
  assign in_2__m_axi_write_data_din = in_2_write_data__din;
  assign in_2_write_data__full_n = in_2__m_axi_write_data_full_n;
  assign in_2__m_axi_write_data_write = in_2_write_data__write;
  assign in_2_write_resp__dout = in_2__m_axi_write_resp_dout;
  assign in_2_write_resp__empty_n = in_2__m_axi_write_resp_empty_n;
  assign in_2__m_axi_write_resp_read = in_2_write_resp__read;
  assign in_20__m_axi_clk = ap_clk;
  assign m_axi_in_20_ARADDR = in_20__m_axi_m_axi_ARADDR;
  assign m_axi_in_20_ARBURST = in_20__m_axi_m_axi_ARBURST;
  assign m_axi_in_20_ARCACHE = in_20__m_axi_m_axi_ARCACHE;
  assign m_axi_in_20_ARID = in_20__m_axi_m_axi_ARID;
  assign m_axi_in_20_ARLEN = in_20__m_axi_m_axi_ARLEN;
  assign m_axi_in_20_ARLOCK = in_20__m_axi_m_axi_ARLOCK;
  assign m_axi_in_20_ARPROT = in_20__m_axi_m_axi_ARPROT;
  assign m_axi_in_20_ARQOS = in_20__m_axi_m_axi_ARQOS;
  assign in_20__m_axi_m_axi_ARREADY = m_axi_in_20_ARREADY;
  assign m_axi_in_20_ARSIZE = in_20__m_axi_m_axi_ARSIZE;
  assign m_axi_in_20_ARVALID = in_20__m_axi_m_axi_ARVALID;
  assign m_axi_in_20_AWADDR = in_20__m_axi_m_axi_AWADDR;
  assign m_axi_in_20_AWBURST = in_20__m_axi_m_axi_AWBURST;
  assign m_axi_in_20_AWCACHE = in_20__m_axi_m_axi_AWCACHE;
  assign m_axi_in_20_AWID = in_20__m_axi_m_axi_AWID;
  assign m_axi_in_20_AWLEN = in_20__m_axi_m_axi_AWLEN;
  assign m_axi_in_20_AWLOCK = in_20__m_axi_m_axi_AWLOCK;
  assign m_axi_in_20_AWPROT = in_20__m_axi_m_axi_AWPROT;
  assign m_axi_in_20_AWQOS = in_20__m_axi_m_axi_AWQOS;
  assign in_20__m_axi_m_axi_AWREADY = m_axi_in_20_AWREADY;
  assign m_axi_in_20_AWSIZE = in_20__m_axi_m_axi_AWSIZE;
  assign m_axi_in_20_AWVALID = in_20__m_axi_m_axi_AWVALID;
  assign in_20__m_axi_m_axi_BID = m_axi_in_20_BID;
  assign m_axi_in_20_BREADY = in_20__m_axi_m_axi_BREADY;
  assign in_20__m_axi_m_axi_BRESP = m_axi_in_20_BRESP;
  assign in_20__m_axi_m_axi_BVALID = m_axi_in_20_BVALID;
  assign in_20__m_axi_m_axi_RDATA = m_axi_in_20_RDATA;
  assign in_20__m_axi_m_axi_RID = m_axi_in_20_RID;
  assign in_20__m_axi_m_axi_RLAST = m_axi_in_20_RLAST;
  assign m_axi_in_20_RREADY = in_20__m_axi_m_axi_RREADY;
  assign in_20__m_axi_m_axi_RRESP = m_axi_in_20_RRESP;
  assign in_20__m_axi_m_axi_RVALID = m_axi_in_20_RVALID;
  assign m_axi_in_20_WDATA = in_20__m_axi_m_axi_WDATA;
  assign m_axi_in_20_WLAST = in_20__m_axi_m_axi_WLAST;
  assign in_20__m_axi_m_axi_WREADY = m_axi_in_20_WREADY;
  assign m_axi_in_20_WSTRB = in_20__m_axi_m_axi_WSTRB;
  assign m_axi_in_20_WVALID = in_20__m_axi_m_axi_WVALID;
  assign in_20__m_axi_read_addr_din = in_20_read_addr__din;
  assign in_20_read_addr__full_n = in_20__m_axi_read_addr_full_n;
  assign in_20__m_axi_read_addr_write = in_20_read_addr__write;
  assign in_20_read_data__dout = in_20__m_axi_read_data_dout;
  assign in_20_read_data__empty_n = in_20__m_axi_read_data_empty_n;
  assign in_20__m_axi_read_data_read = in_20_read_data__read;
  assign in_20__m_axi_rst = ~ ap_rst_n;
  assign in_20__m_axi_write_addr_din = in_20_write_addr__din;
  assign in_20_write_addr__full_n = in_20__m_axi_write_addr_full_n;
  assign in_20__m_axi_write_addr_write = in_20_write_addr__write;
  assign in_20__m_axi_write_data_din = in_20_write_data__din;
  assign in_20_write_data__full_n = in_20__m_axi_write_data_full_n;
  assign in_20__m_axi_write_data_write = in_20_write_data__write;
  assign in_20_write_resp__dout = in_20__m_axi_write_resp_dout;
  assign in_20_write_resp__empty_n = in_20__m_axi_write_resp_empty_n;
  assign in_20__m_axi_write_resp_read = in_20_write_resp__read;
  assign in_21__m_axi_clk = ap_clk;
  assign m_axi_in_21_ARADDR = in_21__m_axi_m_axi_ARADDR;
  assign m_axi_in_21_ARBURST = in_21__m_axi_m_axi_ARBURST;
  assign m_axi_in_21_ARCACHE = in_21__m_axi_m_axi_ARCACHE;
  assign m_axi_in_21_ARID = in_21__m_axi_m_axi_ARID;
  assign m_axi_in_21_ARLEN = in_21__m_axi_m_axi_ARLEN;
  assign m_axi_in_21_ARLOCK = in_21__m_axi_m_axi_ARLOCK;
  assign m_axi_in_21_ARPROT = in_21__m_axi_m_axi_ARPROT;
  assign m_axi_in_21_ARQOS = in_21__m_axi_m_axi_ARQOS;
  assign in_21__m_axi_m_axi_ARREADY = m_axi_in_21_ARREADY;
  assign m_axi_in_21_ARSIZE = in_21__m_axi_m_axi_ARSIZE;
  assign m_axi_in_21_ARVALID = in_21__m_axi_m_axi_ARVALID;
  assign m_axi_in_21_AWADDR = in_21__m_axi_m_axi_AWADDR;
  assign m_axi_in_21_AWBURST = in_21__m_axi_m_axi_AWBURST;
  assign m_axi_in_21_AWCACHE = in_21__m_axi_m_axi_AWCACHE;
  assign m_axi_in_21_AWID = in_21__m_axi_m_axi_AWID;
  assign m_axi_in_21_AWLEN = in_21__m_axi_m_axi_AWLEN;
  assign m_axi_in_21_AWLOCK = in_21__m_axi_m_axi_AWLOCK;
  assign m_axi_in_21_AWPROT = in_21__m_axi_m_axi_AWPROT;
  assign m_axi_in_21_AWQOS = in_21__m_axi_m_axi_AWQOS;
  assign in_21__m_axi_m_axi_AWREADY = m_axi_in_21_AWREADY;
  assign m_axi_in_21_AWSIZE = in_21__m_axi_m_axi_AWSIZE;
  assign m_axi_in_21_AWVALID = in_21__m_axi_m_axi_AWVALID;
  assign in_21__m_axi_m_axi_BID = m_axi_in_21_BID;
  assign m_axi_in_21_BREADY = in_21__m_axi_m_axi_BREADY;
  assign in_21__m_axi_m_axi_BRESP = m_axi_in_21_BRESP;
  assign in_21__m_axi_m_axi_BVALID = m_axi_in_21_BVALID;
  assign in_21__m_axi_m_axi_RDATA = m_axi_in_21_RDATA;
  assign in_21__m_axi_m_axi_RID = m_axi_in_21_RID;
  assign in_21__m_axi_m_axi_RLAST = m_axi_in_21_RLAST;
  assign m_axi_in_21_RREADY = in_21__m_axi_m_axi_RREADY;
  assign in_21__m_axi_m_axi_RRESP = m_axi_in_21_RRESP;
  assign in_21__m_axi_m_axi_RVALID = m_axi_in_21_RVALID;
  assign m_axi_in_21_WDATA = in_21__m_axi_m_axi_WDATA;
  assign m_axi_in_21_WLAST = in_21__m_axi_m_axi_WLAST;
  assign in_21__m_axi_m_axi_WREADY = m_axi_in_21_WREADY;
  assign m_axi_in_21_WSTRB = in_21__m_axi_m_axi_WSTRB;
  assign m_axi_in_21_WVALID = in_21__m_axi_m_axi_WVALID;
  assign in_21__m_axi_read_addr_din = in_21_read_addr__din;
  assign in_21_read_addr__full_n = in_21__m_axi_read_addr_full_n;
  assign in_21__m_axi_read_addr_write = in_21_read_addr__write;
  assign in_21_read_data__dout = in_21__m_axi_read_data_dout;
  assign in_21_read_data__empty_n = in_21__m_axi_read_data_empty_n;
  assign in_21__m_axi_read_data_read = in_21_read_data__read;
  assign in_21__m_axi_rst = ~ ap_rst_n;
  assign in_21__m_axi_write_addr_din = in_21_write_addr__din;
  assign in_21_write_addr__full_n = in_21__m_axi_write_addr_full_n;
  assign in_21__m_axi_write_addr_write = in_21_write_addr__write;
  assign in_21__m_axi_write_data_din = in_21_write_data__din;
  assign in_21_write_data__full_n = in_21__m_axi_write_data_full_n;
  assign in_21__m_axi_write_data_write = in_21_write_data__write;
  assign in_21_write_resp__dout = in_21__m_axi_write_resp_dout;
  assign in_21_write_resp__empty_n = in_21__m_axi_write_resp_empty_n;
  assign in_21__m_axi_write_resp_read = in_21_write_resp__read;
  assign in_22__m_axi_clk = ap_clk;
  assign m_axi_in_22_ARADDR = in_22__m_axi_m_axi_ARADDR;
  assign m_axi_in_22_ARBURST = in_22__m_axi_m_axi_ARBURST;
  assign m_axi_in_22_ARCACHE = in_22__m_axi_m_axi_ARCACHE;
  assign m_axi_in_22_ARID = in_22__m_axi_m_axi_ARID;
  assign m_axi_in_22_ARLEN = in_22__m_axi_m_axi_ARLEN;
  assign m_axi_in_22_ARLOCK = in_22__m_axi_m_axi_ARLOCK;
  assign m_axi_in_22_ARPROT = in_22__m_axi_m_axi_ARPROT;
  assign m_axi_in_22_ARQOS = in_22__m_axi_m_axi_ARQOS;
  assign in_22__m_axi_m_axi_ARREADY = m_axi_in_22_ARREADY;
  assign m_axi_in_22_ARSIZE = in_22__m_axi_m_axi_ARSIZE;
  assign m_axi_in_22_ARVALID = in_22__m_axi_m_axi_ARVALID;
  assign m_axi_in_22_AWADDR = in_22__m_axi_m_axi_AWADDR;
  assign m_axi_in_22_AWBURST = in_22__m_axi_m_axi_AWBURST;
  assign m_axi_in_22_AWCACHE = in_22__m_axi_m_axi_AWCACHE;
  assign m_axi_in_22_AWID = in_22__m_axi_m_axi_AWID;
  assign m_axi_in_22_AWLEN = in_22__m_axi_m_axi_AWLEN;
  assign m_axi_in_22_AWLOCK = in_22__m_axi_m_axi_AWLOCK;
  assign m_axi_in_22_AWPROT = in_22__m_axi_m_axi_AWPROT;
  assign m_axi_in_22_AWQOS = in_22__m_axi_m_axi_AWQOS;
  assign in_22__m_axi_m_axi_AWREADY = m_axi_in_22_AWREADY;
  assign m_axi_in_22_AWSIZE = in_22__m_axi_m_axi_AWSIZE;
  assign m_axi_in_22_AWVALID = in_22__m_axi_m_axi_AWVALID;
  assign in_22__m_axi_m_axi_BID = m_axi_in_22_BID;
  assign m_axi_in_22_BREADY = in_22__m_axi_m_axi_BREADY;
  assign in_22__m_axi_m_axi_BRESP = m_axi_in_22_BRESP;
  assign in_22__m_axi_m_axi_BVALID = m_axi_in_22_BVALID;
  assign in_22__m_axi_m_axi_RDATA = m_axi_in_22_RDATA;
  assign in_22__m_axi_m_axi_RID = m_axi_in_22_RID;
  assign in_22__m_axi_m_axi_RLAST = m_axi_in_22_RLAST;
  assign m_axi_in_22_RREADY = in_22__m_axi_m_axi_RREADY;
  assign in_22__m_axi_m_axi_RRESP = m_axi_in_22_RRESP;
  assign in_22__m_axi_m_axi_RVALID = m_axi_in_22_RVALID;
  assign m_axi_in_22_WDATA = in_22__m_axi_m_axi_WDATA;
  assign m_axi_in_22_WLAST = in_22__m_axi_m_axi_WLAST;
  assign in_22__m_axi_m_axi_WREADY = m_axi_in_22_WREADY;
  assign m_axi_in_22_WSTRB = in_22__m_axi_m_axi_WSTRB;
  assign m_axi_in_22_WVALID = in_22__m_axi_m_axi_WVALID;
  assign in_22__m_axi_read_addr_din = in_22_read_addr__din;
  assign in_22_read_addr__full_n = in_22__m_axi_read_addr_full_n;
  assign in_22__m_axi_read_addr_write = in_22_read_addr__write;
  assign in_22_read_data__dout = in_22__m_axi_read_data_dout;
  assign in_22_read_data__empty_n = in_22__m_axi_read_data_empty_n;
  assign in_22__m_axi_read_data_read = in_22_read_data__read;
  assign in_22__m_axi_rst = ~ ap_rst_n;
  assign in_22__m_axi_write_addr_din = in_22_write_addr__din;
  assign in_22_write_addr__full_n = in_22__m_axi_write_addr_full_n;
  assign in_22__m_axi_write_addr_write = in_22_write_addr__write;
  assign in_22__m_axi_write_data_din = in_22_write_data__din;
  assign in_22_write_data__full_n = in_22__m_axi_write_data_full_n;
  assign in_22__m_axi_write_data_write = in_22_write_data__write;
  assign in_22_write_resp__dout = in_22__m_axi_write_resp_dout;
  assign in_22_write_resp__empty_n = in_22__m_axi_write_resp_empty_n;
  assign in_22__m_axi_write_resp_read = in_22_write_resp__read;
  assign in_23__m_axi_clk = ap_clk;
  assign m_axi_in_23_ARADDR = in_23__m_axi_m_axi_ARADDR;
  assign m_axi_in_23_ARBURST = in_23__m_axi_m_axi_ARBURST;
  assign m_axi_in_23_ARCACHE = in_23__m_axi_m_axi_ARCACHE;
  assign m_axi_in_23_ARID = in_23__m_axi_m_axi_ARID;
  assign m_axi_in_23_ARLEN = in_23__m_axi_m_axi_ARLEN;
  assign m_axi_in_23_ARLOCK = in_23__m_axi_m_axi_ARLOCK;
  assign m_axi_in_23_ARPROT = in_23__m_axi_m_axi_ARPROT;
  assign m_axi_in_23_ARQOS = in_23__m_axi_m_axi_ARQOS;
  assign in_23__m_axi_m_axi_ARREADY = m_axi_in_23_ARREADY;
  assign m_axi_in_23_ARSIZE = in_23__m_axi_m_axi_ARSIZE;
  assign m_axi_in_23_ARVALID = in_23__m_axi_m_axi_ARVALID;
  assign m_axi_in_23_AWADDR = in_23__m_axi_m_axi_AWADDR;
  assign m_axi_in_23_AWBURST = in_23__m_axi_m_axi_AWBURST;
  assign m_axi_in_23_AWCACHE = in_23__m_axi_m_axi_AWCACHE;
  assign m_axi_in_23_AWID = in_23__m_axi_m_axi_AWID;
  assign m_axi_in_23_AWLEN = in_23__m_axi_m_axi_AWLEN;
  assign m_axi_in_23_AWLOCK = in_23__m_axi_m_axi_AWLOCK;
  assign m_axi_in_23_AWPROT = in_23__m_axi_m_axi_AWPROT;
  assign m_axi_in_23_AWQOS = in_23__m_axi_m_axi_AWQOS;
  assign in_23__m_axi_m_axi_AWREADY = m_axi_in_23_AWREADY;
  assign m_axi_in_23_AWSIZE = in_23__m_axi_m_axi_AWSIZE;
  assign m_axi_in_23_AWVALID = in_23__m_axi_m_axi_AWVALID;
  assign in_23__m_axi_m_axi_BID = m_axi_in_23_BID;
  assign m_axi_in_23_BREADY = in_23__m_axi_m_axi_BREADY;
  assign in_23__m_axi_m_axi_BRESP = m_axi_in_23_BRESP;
  assign in_23__m_axi_m_axi_BVALID = m_axi_in_23_BVALID;
  assign in_23__m_axi_m_axi_RDATA = m_axi_in_23_RDATA;
  assign in_23__m_axi_m_axi_RID = m_axi_in_23_RID;
  assign in_23__m_axi_m_axi_RLAST = m_axi_in_23_RLAST;
  assign m_axi_in_23_RREADY = in_23__m_axi_m_axi_RREADY;
  assign in_23__m_axi_m_axi_RRESP = m_axi_in_23_RRESP;
  assign in_23__m_axi_m_axi_RVALID = m_axi_in_23_RVALID;
  assign m_axi_in_23_WDATA = in_23__m_axi_m_axi_WDATA;
  assign m_axi_in_23_WLAST = in_23__m_axi_m_axi_WLAST;
  assign in_23__m_axi_m_axi_WREADY = m_axi_in_23_WREADY;
  assign m_axi_in_23_WSTRB = in_23__m_axi_m_axi_WSTRB;
  assign m_axi_in_23_WVALID = in_23__m_axi_m_axi_WVALID;
  assign in_23__m_axi_read_addr_din = in_23_read_addr__din;
  assign in_23_read_addr__full_n = in_23__m_axi_read_addr_full_n;
  assign in_23__m_axi_read_addr_write = in_23_read_addr__write;
  assign in_23_read_data__dout = in_23__m_axi_read_data_dout;
  assign in_23_read_data__empty_n = in_23__m_axi_read_data_empty_n;
  assign in_23__m_axi_read_data_read = in_23_read_data__read;
  assign in_23__m_axi_rst = ~ ap_rst_n;
  assign in_23__m_axi_write_addr_din = in_23_write_addr__din;
  assign in_23_write_addr__full_n = in_23__m_axi_write_addr_full_n;
  assign in_23__m_axi_write_addr_write = in_23_write_addr__write;
  assign in_23__m_axi_write_data_din = in_23_write_data__din;
  assign in_23_write_data__full_n = in_23__m_axi_write_data_full_n;
  assign in_23__m_axi_write_data_write = in_23_write_data__write;
  assign in_23_write_resp__dout = in_23__m_axi_write_resp_dout;
  assign in_23_write_resp__empty_n = in_23__m_axi_write_resp_empty_n;
  assign in_23__m_axi_write_resp_read = in_23_write_resp__read;
  assign in_24__m_axi_clk = ap_clk;
  assign m_axi_in_24_ARADDR = in_24__m_axi_m_axi_ARADDR;
  assign m_axi_in_24_ARBURST = in_24__m_axi_m_axi_ARBURST;
  assign m_axi_in_24_ARCACHE = in_24__m_axi_m_axi_ARCACHE;
  assign m_axi_in_24_ARID = in_24__m_axi_m_axi_ARID;
  assign m_axi_in_24_ARLEN = in_24__m_axi_m_axi_ARLEN;
  assign m_axi_in_24_ARLOCK = in_24__m_axi_m_axi_ARLOCK;
  assign m_axi_in_24_ARPROT = in_24__m_axi_m_axi_ARPROT;
  assign m_axi_in_24_ARQOS = in_24__m_axi_m_axi_ARQOS;
  assign in_24__m_axi_m_axi_ARREADY = m_axi_in_24_ARREADY;
  assign m_axi_in_24_ARSIZE = in_24__m_axi_m_axi_ARSIZE;
  assign m_axi_in_24_ARVALID = in_24__m_axi_m_axi_ARVALID;
  assign m_axi_in_24_AWADDR = in_24__m_axi_m_axi_AWADDR;
  assign m_axi_in_24_AWBURST = in_24__m_axi_m_axi_AWBURST;
  assign m_axi_in_24_AWCACHE = in_24__m_axi_m_axi_AWCACHE;
  assign m_axi_in_24_AWID = in_24__m_axi_m_axi_AWID;
  assign m_axi_in_24_AWLEN = in_24__m_axi_m_axi_AWLEN;
  assign m_axi_in_24_AWLOCK = in_24__m_axi_m_axi_AWLOCK;
  assign m_axi_in_24_AWPROT = in_24__m_axi_m_axi_AWPROT;
  assign m_axi_in_24_AWQOS = in_24__m_axi_m_axi_AWQOS;
  assign in_24__m_axi_m_axi_AWREADY = m_axi_in_24_AWREADY;
  assign m_axi_in_24_AWSIZE = in_24__m_axi_m_axi_AWSIZE;
  assign m_axi_in_24_AWVALID = in_24__m_axi_m_axi_AWVALID;
  assign in_24__m_axi_m_axi_BID = m_axi_in_24_BID;
  assign m_axi_in_24_BREADY = in_24__m_axi_m_axi_BREADY;
  assign in_24__m_axi_m_axi_BRESP = m_axi_in_24_BRESP;
  assign in_24__m_axi_m_axi_BVALID = m_axi_in_24_BVALID;
  assign in_24__m_axi_m_axi_RDATA = m_axi_in_24_RDATA;
  assign in_24__m_axi_m_axi_RID = m_axi_in_24_RID;
  assign in_24__m_axi_m_axi_RLAST = m_axi_in_24_RLAST;
  assign m_axi_in_24_RREADY = in_24__m_axi_m_axi_RREADY;
  assign in_24__m_axi_m_axi_RRESP = m_axi_in_24_RRESP;
  assign in_24__m_axi_m_axi_RVALID = m_axi_in_24_RVALID;
  assign m_axi_in_24_WDATA = in_24__m_axi_m_axi_WDATA;
  assign m_axi_in_24_WLAST = in_24__m_axi_m_axi_WLAST;
  assign in_24__m_axi_m_axi_WREADY = m_axi_in_24_WREADY;
  assign m_axi_in_24_WSTRB = in_24__m_axi_m_axi_WSTRB;
  assign m_axi_in_24_WVALID = in_24__m_axi_m_axi_WVALID;
  assign in_24__m_axi_read_addr_din = in_24_read_addr__din;
  assign in_24_read_addr__full_n = in_24__m_axi_read_addr_full_n;
  assign in_24__m_axi_read_addr_write = in_24_read_addr__write;
  assign in_24_read_data__dout = in_24__m_axi_read_data_dout;
  assign in_24_read_data__empty_n = in_24__m_axi_read_data_empty_n;
  assign in_24__m_axi_read_data_read = in_24_read_data__read;
  assign in_24__m_axi_rst = ~ ap_rst_n;
  assign in_24__m_axi_write_addr_din = in_24_write_addr__din;
  assign in_24_write_addr__full_n = in_24__m_axi_write_addr_full_n;
  assign in_24__m_axi_write_addr_write = in_24_write_addr__write;
  assign in_24__m_axi_write_data_din = in_24_write_data__din;
  assign in_24_write_data__full_n = in_24__m_axi_write_data_full_n;
  assign in_24__m_axi_write_data_write = in_24_write_data__write;
  assign in_24_write_resp__dout = in_24__m_axi_write_resp_dout;
  assign in_24_write_resp__empty_n = in_24__m_axi_write_resp_empty_n;
  assign in_24__m_axi_write_resp_read = in_24_write_resp__read;
  assign in_25__m_axi_clk = ap_clk;
  assign m_axi_in_25_ARADDR = in_25__m_axi_m_axi_ARADDR;
  assign m_axi_in_25_ARBURST = in_25__m_axi_m_axi_ARBURST;
  assign m_axi_in_25_ARCACHE = in_25__m_axi_m_axi_ARCACHE;
  assign m_axi_in_25_ARID = in_25__m_axi_m_axi_ARID;
  assign m_axi_in_25_ARLEN = in_25__m_axi_m_axi_ARLEN;
  assign m_axi_in_25_ARLOCK = in_25__m_axi_m_axi_ARLOCK;
  assign m_axi_in_25_ARPROT = in_25__m_axi_m_axi_ARPROT;
  assign m_axi_in_25_ARQOS = in_25__m_axi_m_axi_ARQOS;
  assign in_25__m_axi_m_axi_ARREADY = m_axi_in_25_ARREADY;
  assign m_axi_in_25_ARSIZE = in_25__m_axi_m_axi_ARSIZE;
  assign m_axi_in_25_ARVALID = in_25__m_axi_m_axi_ARVALID;
  assign m_axi_in_25_AWADDR = in_25__m_axi_m_axi_AWADDR;
  assign m_axi_in_25_AWBURST = in_25__m_axi_m_axi_AWBURST;
  assign m_axi_in_25_AWCACHE = in_25__m_axi_m_axi_AWCACHE;
  assign m_axi_in_25_AWID = in_25__m_axi_m_axi_AWID;
  assign m_axi_in_25_AWLEN = in_25__m_axi_m_axi_AWLEN;
  assign m_axi_in_25_AWLOCK = in_25__m_axi_m_axi_AWLOCK;
  assign m_axi_in_25_AWPROT = in_25__m_axi_m_axi_AWPROT;
  assign m_axi_in_25_AWQOS = in_25__m_axi_m_axi_AWQOS;
  assign in_25__m_axi_m_axi_AWREADY = m_axi_in_25_AWREADY;
  assign m_axi_in_25_AWSIZE = in_25__m_axi_m_axi_AWSIZE;
  assign m_axi_in_25_AWVALID = in_25__m_axi_m_axi_AWVALID;
  assign in_25__m_axi_m_axi_BID = m_axi_in_25_BID;
  assign m_axi_in_25_BREADY = in_25__m_axi_m_axi_BREADY;
  assign in_25__m_axi_m_axi_BRESP = m_axi_in_25_BRESP;
  assign in_25__m_axi_m_axi_BVALID = m_axi_in_25_BVALID;
  assign in_25__m_axi_m_axi_RDATA = m_axi_in_25_RDATA;
  assign in_25__m_axi_m_axi_RID = m_axi_in_25_RID;
  assign in_25__m_axi_m_axi_RLAST = m_axi_in_25_RLAST;
  assign m_axi_in_25_RREADY = in_25__m_axi_m_axi_RREADY;
  assign in_25__m_axi_m_axi_RRESP = m_axi_in_25_RRESP;
  assign in_25__m_axi_m_axi_RVALID = m_axi_in_25_RVALID;
  assign m_axi_in_25_WDATA = in_25__m_axi_m_axi_WDATA;
  assign m_axi_in_25_WLAST = in_25__m_axi_m_axi_WLAST;
  assign in_25__m_axi_m_axi_WREADY = m_axi_in_25_WREADY;
  assign m_axi_in_25_WSTRB = in_25__m_axi_m_axi_WSTRB;
  assign m_axi_in_25_WVALID = in_25__m_axi_m_axi_WVALID;
  assign in_25__m_axi_read_addr_din = in_25_read_addr__din;
  assign in_25_read_addr__full_n = in_25__m_axi_read_addr_full_n;
  assign in_25__m_axi_read_addr_write = in_25_read_addr__write;
  assign in_25_read_data__dout = in_25__m_axi_read_data_dout;
  assign in_25_read_data__empty_n = in_25__m_axi_read_data_empty_n;
  assign in_25__m_axi_read_data_read = in_25_read_data__read;
  assign in_25__m_axi_rst = ~ ap_rst_n;
  assign in_25__m_axi_write_addr_din = in_25_write_addr__din;
  assign in_25_write_addr__full_n = in_25__m_axi_write_addr_full_n;
  assign in_25__m_axi_write_addr_write = in_25_write_addr__write;
  assign in_25__m_axi_write_data_din = in_25_write_data__din;
  assign in_25_write_data__full_n = in_25__m_axi_write_data_full_n;
  assign in_25__m_axi_write_data_write = in_25_write_data__write;
  assign in_25_write_resp__dout = in_25__m_axi_write_resp_dout;
  assign in_25_write_resp__empty_n = in_25__m_axi_write_resp_empty_n;
  assign in_25__m_axi_write_resp_read = in_25_write_resp__read;
  assign in_26__m_axi_clk = ap_clk;
  assign m_axi_in_26_ARADDR = in_26__m_axi_m_axi_ARADDR;
  assign m_axi_in_26_ARBURST = in_26__m_axi_m_axi_ARBURST;
  assign m_axi_in_26_ARCACHE = in_26__m_axi_m_axi_ARCACHE;
  assign m_axi_in_26_ARID = in_26__m_axi_m_axi_ARID;
  assign m_axi_in_26_ARLEN = in_26__m_axi_m_axi_ARLEN;
  assign m_axi_in_26_ARLOCK = in_26__m_axi_m_axi_ARLOCK;
  assign m_axi_in_26_ARPROT = in_26__m_axi_m_axi_ARPROT;
  assign m_axi_in_26_ARQOS = in_26__m_axi_m_axi_ARQOS;
  assign in_26__m_axi_m_axi_ARREADY = m_axi_in_26_ARREADY;
  assign m_axi_in_26_ARSIZE = in_26__m_axi_m_axi_ARSIZE;
  assign m_axi_in_26_ARVALID = in_26__m_axi_m_axi_ARVALID;
  assign m_axi_in_26_AWADDR = in_26__m_axi_m_axi_AWADDR;
  assign m_axi_in_26_AWBURST = in_26__m_axi_m_axi_AWBURST;
  assign m_axi_in_26_AWCACHE = in_26__m_axi_m_axi_AWCACHE;
  assign m_axi_in_26_AWID = in_26__m_axi_m_axi_AWID;
  assign m_axi_in_26_AWLEN = in_26__m_axi_m_axi_AWLEN;
  assign m_axi_in_26_AWLOCK = in_26__m_axi_m_axi_AWLOCK;
  assign m_axi_in_26_AWPROT = in_26__m_axi_m_axi_AWPROT;
  assign m_axi_in_26_AWQOS = in_26__m_axi_m_axi_AWQOS;
  assign in_26__m_axi_m_axi_AWREADY = m_axi_in_26_AWREADY;
  assign m_axi_in_26_AWSIZE = in_26__m_axi_m_axi_AWSIZE;
  assign m_axi_in_26_AWVALID = in_26__m_axi_m_axi_AWVALID;
  assign in_26__m_axi_m_axi_BID = m_axi_in_26_BID;
  assign m_axi_in_26_BREADY = in_26__m_axi_m_axi_BREADY;
  assign in_26__m_axi_m_axi_BRESP = m_axi_in_26_BRESP;
  assign in_26__m_axi_m_axi_BVALID = m_axi_in_26_BVALID;
  assign in_26__m_axi_m_axi_RDATA = m_axi_in_26_RDATA;
  assign in_26__m_axi_m_axi_RID = m_axi_in_26_RID;
  assign in_26__m_axi_m_axi_RLAST = m_axi_in_26_RLAST;
  assign m_axi_in_26_RREADY = in_26__m_axi_m_axi_RREADY;
  assign in_26__m_axi_m_axi_RRESP = m_axi_in_26_RRESP;
  assign in_26__m_axi_m_axi_RVALID = m_axi_in_26_RVALID;
  assign m_axi_in_26_WDATA = in_26__m_axi_m_axi_WDATA;
  assign m_axi_in_26_WLAST = in_26__m_axi_m_axi_WLAST;
  assign in_26__m_axi_m_axi_WREADY = m_axi_in_26_WREADY;
  assign m_axi_in_26_WSTRB = in_26__m_axi_m_axi_WSTRB;
  assign m_axi_in_26_WVALID = in_26__m_axi_m_axi_WVALID;
  assign in_26__m_axi_read_addr_din = in_26_read_addr__din;
  assign in_26_read_addr__full_n = in_26__m_axi_read_addr_full_n;
  assign in_26__m_axi_read_addr_write = in_26_read_addr__write;
  assign in_26_read_data__dout = in_26__m_axi_read_data_dout;
  assign in_26_read_data__empty_n = in_26__m_axi_read_data_empty_n;
  assign in_26__m_axi_read_data_read = in_26_read_data__read;
  assign in_26__m_axi_rst = ~ ap_rst_n;
  assign in_26__m_axi_write_addr_din = in_26_write_addr__din;
  assign in_26_write_addr__full_n = in_26__m_axi_write_addr_full_n;
  assign in_26__m_axi_write_addr_write = in_26_write_addr__write;
  assign in_26__m_axi_write_data_din = in_26_write_data__din;
  assign in_26_write_data__full_n = in_26__m_axi_write_data_full_n;
  assign in_26__m_axi_write_data_write = in_26_write_data__write;
  assign in_26_write_resp__dout = in_26__m_axi_write_resp_dout;
  assign in_26_write_resp__empty_n = in_26__m_axi_write_resp_empty_n;
  assign in_26__m_axi_write_resp_read = in_26_write_resp__read;
  assign in_27__m_axi_clk = ap_clk;
  assign m_axi_in_27_ARADDR = in_27__m_axi_m_axi_ARADDR;
  assign m_axi_in_27_ARBURST = in_27__m_axi_m_axi_ARBURST;
  assign m_axi_in_27_ARCACHE = in_27__m_axi_m_axi_ARCACHE;
  assign m_axi_in_27_ARID = in_27__m_axi_m_axi_ARID;
  assign m_axi_in_27_ARLEN = in_27__m_axi_m_axi_ARLEN;
  assign m_axi_in_27_ARLOCK = in_27__m_axi_m_axi_ARLOCK;
  assign m_axi_in_27_ARPROT = in_27__m_axi_m_axi_ARPROT;
  assign m_axi_in_27_ARQOS = in_27__m_axi_m_axi_ARQOS;
  assign in_27__m_axi_m_axi_ARREADY = m_axi_in_27_ARREADY;
  assign m_axi_in_27_ARSIZE = in_27__m_axi_m_axi_ARSIZE;
  assign m_axi_in_27_ARVALID = in_27__m_axi_m_axi_ARVALID;
  assign m_axi_in_27_AWADDR = in_27__m_axi_m_axi_AWADDR;
  assign m_axi_in_27_AWBURST = in_27__m_axi_m_axi_AWBURST;
  assign m_axi_in_27_AWCACHE = in_27__m_axi_m_axi_AWCACHE;
  assign m_axi_in_27_AWID = in_27__m_axi_m_axi_AWID;
  assign m_axi_in_27_AWLEN = in_27__m_axi_m_axi_AWLEN;
  assign m_axi_in_27_AWLOCK = in_27__m_axi_m_axi_AWLOCK;
  assign m_axi_in_27_AWPROT = in_27__m_axi_m_axi_AWPROT;
  assign m_axi_in_27_AWQOS = in_27__m_axi_m_axi_AWQOS;
  assign in_27__m_axi_m_axi_AWREADY = m_axi_in_27_AWREADY;
  assign m_axi_in_27_AWSIZE = in_27__m_axi_m_axi_AWSIZE;
  assign m_axi_in_27_AWVALID = in_27__m_axi_m_axi_AWVALID;
  assign in_27__m_axi_m_axi_BID = m_axi_in_27_BID;
  assign m_axi_in_27_BREADY = in_27__m_axi_m_axi_BREADY;
  assign in_27__m_axi_m_axi_BRESP = m_axi_in_27_BRESP;
  assign in_27__m_axi_m_axi_BVALID = m_axi_in_27_BVALID;
  assign in_27__m_axi_m_axi_RDATA = m_axi_in_27_RDATA;
  assign in_27__m_axi_m_axi_RID = m_axi_in_27_RID;
  assign in_27__m_axi_m_axi_RLAST = m_axi_in_27_RLAST;
  assign m_axi_in_27_RREADY = in_27__m_axi_m_axi_RREADY;
  assign in_27__m_axi_m_axi_RRESP = m_axi_in_27_RRESP;
  assign in_27__m_axi_m_axi_RVALID = m_axi_in_27_RVALID;
  assign m_axi_in_27_WDATA = in_27__m_axi_m_axi_WDATA;
  assign m_axi_in_27_WLAST = in_27__m_axi_m_axi_WLAST;
  assign in_27__m_axi_m_axi_WREADY = m_axi_in_27_WREADY;
  assign m_axi_in_27_WSTRB = in_27__m_axi_m_axi_WSTRB;
  assign m_axi_in_27_WVALID = in_27__m_axi_m_axi_WVALID;
  assign in_27__m_axi_read_addr_din = in_27_read_addr__din;
  assign in_27_read_addr__full_n = in_27__m_axi_read_addr_full_n;
  assign in_27__m_axi_read_addr_write = in_27_read_addr__write;
  assign in_27_read_data__dout = in_27__m_axi_read_data_dout;
  assign in_27_read_data__empty_n = in_27__m_axi_read_data_empty_n;
  assign in_27__m_axi_read_data_read = in_27_read_data__read;
  assign in_27__m_axi_rst = ~ ap_rst_n;
  assign in_27__m_axi_write_addr_din = in_27_write_addr__din;
  assign in_27_write_addr__full_n = in_27__m_axi_write_addr_full_n;
  assign in_27__m_axi_write_addr_write = in_27_write_addr__write;
  assign in_27__m_axi_write_data_din = in_27_write_data__din;
  assign in_27_write_data__full_n = in_27__m_axi_write_data_full_n;
  assign in_27__m_axi_write_data_write = in_27_write_data__write;
  assign in_27_write_resp__dout = in_27__m_axi_write_resp_dout;
  assign in_27_write_resp__empty_n = in_27__m_axi_write_resp_empty_n;
  assign in_27__m_axi_write_resp_read = in_27_write_resp__read;
  assign in_28__m_axi_clk = ap_clk;
  assign m_axi_in_28_ARADDR = in_28__m_axi_m_axi_ARADDR;
  assign m_axi_in_28_ARBURST = in_28__m_axi_m_axi_ARBURST;
  assign m_axi_in_28_ARCACHE = in_28__m_axi_m_axi_ARCACHE;
  assign m_axi_in_28_ARID = in_28__m_axi_m_axi_ARID;
  assign m_axi_in_28_ARLEN = in_28__m_axi_m_axi_ARLEN;
  assign m_axi_in_28_ARLOCK = in_28__m_axi_m_axi_ARLOCK;
  assign m_axi_in_28_ARPROT = in_28__m_axi_m_axi_ARPROT;
  assign m_axi_in_28_ARQOS = in_28__m_axi_m_axi_ARQOS;
  assign in_28__m_axi_m_axi_ARREADY = m_axi_in_28_ARREADY;
  assign m_axi_in_28_ARSIZE = in_28__m_axi_m_axi_ARSIZE;
  assign m_axi_in_28_ARVALID = in_28__m_axi_m_axi_ARVALID;
  assign m_axi_in_28_AWADDR = in_28__m_axi_m_axi_AWADDR;
  assign m_axi_in_28_AWBURST = in_28__m_axi_m_axi_AWBURST;
  assign m_axi_in_28_AWCACHE = in_28__m_axi_m_axi_AWCACHE;
  assign m_axi_in_28_AWID = in_28__m_axi_m_axi_AWID;
  assign m_axi_in_28_AWLEN = in_28__m_axi_m_axi_AWLEN;
  assign m_axi_in_28_AWLOCK = in_28__m_axi_m_axi_AWLOCK;
  assign m_axi_in_28_AWPROT = in_28__m_axi_m_axi_AWPROT;
  assign m_axi_in_28_AWQOS = in_28__m_axi_m_axi_AWQOS;
  assign in_28__m_axi_m_axi_AWREADY = m_axi_in_28_AWREADY;
  assign m_axi_in_28_AWSIZE = in_28__m_axi_m_axi_AWSIZE;
  assign m_axi_in_28_AWVALID = in_28__m_axi_m_axi_AWVALID;
  assign in_28__m_axi_m_axi_BID = m_axi_in_28_BID;
  assign m_axi_in_28_BREADY = in_28__m_axi_m_axi_BREADY;
  assign in_28__m_axi_m_axi_BRESP = m_axi_in_28_BRESP;
  assign in_28__m_axi_m_axi_BVALID = m_axi_in_28_BVALID;
  assign in_28__m_axi_m_axi_RDATA = m_axi_in_28_RDATA;
  assign in_28__m_axi_m_axi_RID = m_axi_in_28_RID;
  assign in_28__m_axi_m_axi_RLAST = m_axi_in_28_RLAST;
  assign m_axi_in_28_RREADY = in_28__m_axi_m_axi_RREADY;
  assign in_28__m_axi_m_axi_RRESP = m_axi_in_28_RRESP;
  assign in_28__m_axi_m_axi_RVALID = m_axi_in_28_RVALID;
  assign m_axi_in_28_WDATA = in_28__m_axi_m_axi_WDATA;
  assign m_axi_in_28_WLAST = in_28__m_axi_m_axi_WLAST;
  assign in_28__m_axi_m_axi_WREADY = m_axi_in_28_WREADY;
  assign m_axi_in_28_WSTRB = in_28__m_axi_m_axi_WSTRB;
  assign m_axi_in_28_WVALID = in_28__m_axi_m_axi_WVALID;
  assign in_28__m_axi_read_addr_din = in_28_read_addr__din;
  assign in_28_read_addr__full_n = in_28__m_axi_read_addr_full_n;
  assign in_28__m_axi_read_addr_write = in_28_read_addr__write;
  assign in_28_read_data__dout = in_28__m_axi_read_data_dout;
  assign in_28_read_data__empty_n = in_28__m_axi_read_data_empty_n;
  assign in_28__m_axi_read_data_read = in_28_read_data__read;
  assign in_28__m_axi_rst = ~ ap_rst_n;
  assign in_28__m_axi_write_addr_din = in_28_write_addr__din;
  assign in_28_write_addr__full_n = in_28__m_axi_write_addr_full_n;
  assign in_28__m_axi_write_addr_write = in_28_write_addr__write;
  assign in_28__m_axi_write_data_din = in_28_write_data__din;
  assign in_28_write_data__full_n = in_28__m_axi_write_data_full_n;
  assign in_28__m_axi_write_data_write = in_28_write_data__write;
  assign in_28_write_resp__dout = in_28__m_axi_write_resp_dout;
  assign in_28_write_resp__empty_n = in_28__m_axi_write_resp_empty_n;
  assign in_28__m_axi_write_resp_read = in_28_write_resp__read;
  assign in_29__m_axi_clk = ap_clk;
  assign m_axi_in_29_ARADDR = in_29__m_axi_m_axi_ARADDR;
  assign m_axi_in_29_ARBURST = in_29__m_axi_m_axi_ARBURST;
  assign m_axi_in_29_ARCACHE = in_29__m_axi_m_axi_ARCACHE;
  assign m_axi_in_29_ARID = in_29__m_axi_m_axi_ARID;
  assign m_axi_in_29_ARLEN = in_29__m_axi_m_axi_ARLEN;
  assign m_axi_in_29_ARLOCK = in_29__m_axi_m_axi_ARLOCK;
  assign m_axi_in_29_ARPROT = in_29__m_axi_m_axi_ARPROT;
  assign m_axi_in_29_ARQOS = in_29__m_axi_m_axi_ARQOS;
  assign in_29__m_axi_m_axi_ARREADY = m_axi_in_29_ARREADY;
  assign m_axi_in_29_ARSIZE = in_29__m_axi_m_axi_ARSIZE;
  assign m_axi_in_29_ARVALID = in_29__m_axi_m_axi_ARVALID;
  assign m_axi_in_29_AWADDR = in_29__m_axi_m_axi_AWADDR;
  assign m_axi_in_29_AWBURST = in_29__m_axi_m_axi_AWBURST;
  assign m_axi_in_29_AWCACHE = in_29__m_axi_m_axi_AWCACHE;
  assign m_axi_in_29_AWID = in_29__m_axi_m_axi_AWID;
  assign m_axi_in_29_AWLEN = in_29__m_axi_m_axi_AWLEN;
  assign m_axi_in_29_AWLOCK = in_29__m_axi_m_axi_AWLOCK;
  assign m_axi_in_29_AWPROT = in_29__m_axi_m_axi_AWPROT;
  assign m_axi_in_29_AWQOS = in_29__m_axi_m_axi_AWQOS;
  assign in_29__m_axi_m_axi_AWREADY = m_axi_in_29_AWREADY;
  assign m_axi_in_29_AWSIZE = in_29__m_axi_m_axi_AWSIZE;
  assign m_axi_in_29_AWVALID = in_29__m_axi_m_axi_AWVALID;
  assign in_29__m_axi_m_axi_BID = m_axi_in_29_BID;
  assign m_axi_in_29_BREADY = in_29__m_axi_m_axi_BREADY;
  assign in_29__m_axi_m_axi_BRESP = m_axi_in_29_BRESP;
  assign in_29__m_axi_m_axi_BVALID = m_axi_in_29_BVALID;
  assign in_29__m_axi_m_axi_RDATA = m_axi_in_29_RDATA;
  assign in_29__m_axi_m_axi_RID = m_axi_in_29_RID;
  assign in_29__m_axi_m_axi_RLAST = m_axi_in_29_RLAST;
  assign m_axi_in_29_RREADY = in_29__m_axi_m_axi_RREADY;
  assign in_29__m_axi_m_axi_RRESP = m_axi_in_29_RRESP;
  assign in_29__m_axi_m_axi_RVALID = m_axi_in_29_RVALID;
  assign m_axi_in_29_WDATA = in_29__m_axi_m_axi_WDATA;
  assign m_axi_in_29_WLAST = in_29__m_axi_m_axi_WLAST;
  assign in_29__m_axi_m_axi_WREADY = m_axi_in_29_WREADY;
  assign m_axi_in_29_WSTRB = in_29__m_axi_m_axi_WSTRB;
  assign m_axi_in_29_WVALID = in_29__m_axi_m_axi_WVALID;
  assign in_29__m_axi_read_addr_din = in_29_read_addr__din;
  assign in_29_read_addr__full_n = in_29__m_axi_read_addr_full_n;
  assign in_29__m_axi_read_addr_write = in_29_read_addr__write;
  assign in_29_read_data__dout = in_29__m_axi_read_data_dout;
  assign in_29_read_data__empty_n = in_29__m_axi_read_data_empty_n;
  assign in_29__m_axi_read_data_read = in_29_read_data__read;
  assign in_29__m_axi_rst = ~ ap_rst_n;
  assign in_29__m_axi_write_addr_din = in_29_write_addr__din;
  assign in_29_write_addr__full_n = in_29__m_axi_write_addr_full_n;
  assign in_29__m_axi_write_addr_write = in_29_write_addr__write;
  assign in_29__m_axi_write_data_din = in_29_write_data__din;
  assign in_29_write_data__full_n = in_29__m_axi_write_data_full_n;
  assign in_29__m_axi_write_data_write = in_29_write_data__write;
  assign in_29_write_resp__dout = in_29__m_axi_write_resp_dout;
  assign in_29_write_resp__empty_n = in_29__m_axi_write_resp_empty_n;
  assign in_29__m_axi_write_resp_read = in_29_write_resp__read;
  assign in_3__m_axi_clk = ap_clk;
  assign m_axi_in_3_ARADDR = in_3__m_axi_m_axi_ARADDR;
  assign m_axi_in_3_ARBURST = in_3__m_axi_m_axi_ARBURST;
  assign m_axi_in_3_ARCACHE = in_3__m_axi_m_axi_ARCACHE;
  assign m_axi_in_3_ARID = in_3__m_axi_m_axi_ARID;
  assign m_axi_in_3_ARLEN = in_3__m_axi_m_axi_ARLEN;
  assign m_axi_in_3_ARLOCK = in_3__m_axi_m_axi_ARLOCK;
  assign m_axi_in_3_ARPROT = in_3__m_axi_m_axi_ARPROT;
  assign m_axi_in_3_ARQOS = in_3__m_axi_m_axi_ARQOS;
  assign in_3__m_axi_m_axi_ARREADY = m_axi_in_3_ARREADY;
  assign m_axi_in_3_ARSIZE = in_3__m_axi_m_axi_ARSIZE;
  assign m_axi_in_3_ARVALID = in_3__m_axi_m_axi_ARVALID;
  assign m_axi_in_3_AWADDR = in_3__m_axi_m_axi_AWADDR;
  assign m_axi_in_3_AWBURST = in_3__m_axi_m_axi_AWBURST;
  assign m_axi_in_3_AWCACHE = in_3__m_axi_m_axi_AWCACHE;
  assign m_axi_in_3_AWID = in_3__m_axi_m_axi_AWID;
  assign m_axi_in_3_AWLEN = in_3__m_axi_m_axi_AWLEN;
  assign m_axi_in_3_AWLOCK = in_3__m_axi_m_axi_AWLOCK;
  assign m_axi_in_3_AWPROT = in_3__m_axi_m_axi_AWPROT;
  assign m_axi_in_3_AWQOS = in_3__m_axi_m_axi_AWQOS;
  assign in_3__m_axi_m_axi_AWREADY = m_axi_in_3_AWREADY;
  assign m_axi_in_3_AWSIZE = in_3__m_axi_m_axi_AWSIZE;
  assign m_axi_in_3_AWVALID = in_3__m_axi_m_axi_AWVALID;
  assign in_3__m_axi_m_axi_BID = m_axi_in_3_BID;
  assign m_axi_in_3_BREADY = in_3__m_axi_m_axi_BREADY;
  assign in_3__m_axi_m_axi_BRESP = m_axi_in_3_BRESP;
  assign in_3__m_axi_m_axi_BVALID = m_axi_in_3_BVALID;
  assign in_3__m_axi_m_axi_RDATA = m_axi_in_3_RDATA;
  assign in_3__m_axi_m_axi_RID = m_axi_in_3_RID;
  assign in_3__m_axi_m_axi_RLAST = m_axi_in_3_RLAST;
  assign m_axi_in_3_RREADY = in_3__m_axi_m_axi_RREADY;
  assign in_3__m_axi_m_axi_RRESP = m_axi_in_3_RRESP;
  assign in_3__m_axi_m_axi_RVALID = m_axi_in_3_RVALID;
  assign m_axi_in_3_WDATA = in_3__m_axi_m_axi_WDATA;
  assign m_axi_in_3_WLAST = in_3__m_axi_m_axi_WLAST;
  assign in_3__m_axi_m_axi_WREADY = m_axi_in_3_WREADY;
  assign m_axi_in_3_WSTRB = in_3__m_axi_m_axi_WSTRB;
  assign m_axi_in_3_WVALID = in_3__m_axi_m_axi_WVALID;
  assign in_3__m_axi_read_addr_din = in_3_read_addr__din;
  assign in_3_read_addr__full_n = in_3__m_axi_read_addr_full_n;
  assign in_3__m_axi_read_addr_write = in_3_read_addr__write;
  assign in_3_read_data__dout = in_3__m_axi_read_data_dout;
  assign in_3_read_data__empty_n = in_3__m_axi_read_data_empty_n;
  assign in_3__m_axi_read_data_read = in_3_read_data__read;
  assign in_3__m_axi_rst = ~ ap_rst_n;
  assign in_3__m_axi_write_addr_din = in_3_write_addr__din;
  assign in_3_write_addr__full_n = in_3__m_axi_write_addr_full_n;
  assign in_3__m_axi_write_addr_write = in_3_write_addr__write;
  assign in_3__m_axi_write_data_din = in_3_write_data__din;
  assign in_3_write_data__full_n = in_3__m_axi_write_data_full_n;
  assign in_3__m_axi_write_data_write = in_3_write_data__write;
  assign in_3_write_resp__dout = in_3__m_axi_write_resp_dout;
  assign in_3_write_resp__empty_n = in_3__m_axi_write_resp_empty_n;
  assign in_3__m_axi_write_resp_read = in_3_write_resp__read;
  assign in_30__m_axi_clk = ap_clk;
  assign m_axi_in_30_ARADDR = in_30__m_axi_m_axi_ARADDR;
  assign m_axi_in_30_ARBURST = in_30__m_axi_m_axi_ARBURST;
  assign m_axi_in_30_ARCACHE = in_30__m_axi_m_axi_ARCACHE;
  assign m_axi_in_30_ARID = in_30__m_axi_m_axi_ARID;
  assign m_axi_in_30_ARLEN = in_30__m_axi_m_axi_ARLEN;
  assign m_axi_in_30_ARLOCK = in_30__m_axi_m_axi_ARLOCK;
  assign m_axi_in_30_ARPROT = in_30__m_axi_m_axi_ARPROT;
  assign m_axi_in_30_ARQOS = in_30__m_axi_m_axi_ARQOS;
  assign in_30__m_axi_m_axi_ARREADY = m_axi_in_30_ARREADY;
  assign m_axi_in_30_ARSIZE = in_30__m_axi_m_axi_ARSIZE;
  assign m_axi_in_30_ARVALID = in_30__m_axi_m_axi_ARVALID;
  assign m_axi_in_30_AWADDR = in_30__m_axi_m_axi_AWADDR;
  assign m_axi_in_30_AWBURST = in_30__m_axi_m_axi_AWBURST;
  assign m_axi_in_30_AWCACHE = in_30__m_axi_m_axi_AWCACHE;
  assign m_axi_in_30_AWID = in_30__m_axi_m_axi_AWID;
  assign m_axi_in_30_AWLEN = in_30__m_axi_m_axi_AWLEN;
  assign m_axi_in_30_AWLOCK = in_30__m_axi_m_axi_AWLOCK;
  assign m_axi_in_30_AWPROT = in_30__m_axi_m_axi_AWPROT;
  assign m_axi_in_30_AWQOS = in_30__m_axi_m_axi_AWQOS;
  assign in_30__m_axi_m_axi_AWREADY = m_axi_in_30_AWREADY;
  assign m_axi_in_30_AWSIZE = in_30__m_axi_m_axi_AWSIZE;
  assign m_axi_in_30_AWVALID = in_30__m_axi_m_axi_AWVALID;
  assign in_30__m_axi_m_axi_BID = m_axi_in_30_BID;
  assign m_axi_in_30_BREADY = in_30__m_axi_m_axi_BREADY;
  assign in_30__m_axi_m_axi_BRESP = m_axi_in_30_BRESP;
  assign in_30__m_axi_m_axi_BVALID = m_axi_in_30_BVALID;
  assign in_30__m_axi_m_axi_RDATA = m_axi_in_30_RDATA;
  assign in_30__m_axi_m_axi_RID = m_axi_in_30_RID;
  assign in_30__m_axi_m_axi_RLAST = m_axi_in_30_RLAST;
  assign m_axi_in_30_RREADY = in_30__m_axi_m_axi_RREADY;
  assign in_30__m_axi_m_axi_RRESP = m_axi_in_30_RRESP;
  assign in_30__m_axi_m_axi_RVALID = m_axi_in_30_RVALID;
  assign m_axi_in_30_WDATA = in_30__m_axi_m_axi_WDATA;
  assign m_axi_in_30_WLAST = in_30__m_axi_m_axi_WLAST;
  assign in_30__m_axi_m_axi_WREADY = m_axi_in_30_WREADY;
  assign m_axi_in_30_WSTRB = in_30__m_axi_m_axi_WSTRB;
  assign m_axi_in_30_WVALID = in_30__m_axi_m_axi_WVALID;
  assign in_30__m_axi_read_addr_din = in_30_read_addr__din;
  assign in_30_read_addr__full_n = in_30__m_axi_read_addr_full_n;
  assign in_30__m_axi_read_addr_write = in_30_read_addr__write;
  assign in_30_read_data__dout = in_30__m_axi_read_data_dout;
  assign in_30_read_data__empty_n = in_30__m_axi_read_data_empty_n;
  assign in_30__m_axi_read_data_read = in_30_read_data__read;
  assign in_30__m_axi_rst = ~ ap_rst_n;
  assign in_30__m_axi_write_addr_din = in_30_write_addr__din;
  assign in_30_write_addr__full_n = in_30__m_axi_write_addr_full_n;
  assign in_30__m_axi_write_addr_write = in_30_write_addr__write;
  assign in_30__m_axi_write_data_din = in_30_write_data__din;
  assign in_30_write_data__full_n = in_30__m_axi_write_data_full_n;
  assign in_30__m_axi_write_data_write = in_30_write_data__write;
  assign in_30_write_resp__dout = in_30__m_axi_write_resp_dout;
  assign in_30_write_resp__empty_n = in_30__m_axi_write_resp_empty_n;
  assign in_30__m_axi_write_resp_read = in_30_write_resp__read;
  assign in_31__m_axi_clk = ap_clk;
  assign m_axi_in_31_ARADDR = in_31__m_axi_m_axi_ARADDR;
  assign m_axi_in_31_ARBURST = in_31__m_axi_m_axi_ARBURST;
  assign m_axi_in_31_ARCACHE = in_31__m_axi_m_axi_ARCACHE;
  assign m_axi_in_31_ARID = in_31__m_axi_m_axi_ARID;
  assign m_axi_in_31_ARLEN = in_31__m_axi_m_axi_ARLEN;
  assign m_axi_in_31_ARLOCK = in_31__m_axi_m_axi_ARLOCK;
  assign m_axi_in_31_ARPROT = in_31__m_axi_m_axi_ARPROT;
  assign m_axi_in_31_ARQOS = in_31__m_axi_m_axi_ARQOS;
  assign in_31__m_axi_m_axi_ARREADY = m_axi_in_31_ARREADY;
  assign m_axi_in_31_ARSIZE = in_31__m_axi_m_axi_ARSIZE;
  assign m_axi_in_31_ARVALID = in_31__m_axi_m_axi_ARVALID;
  assign m_axi_in_31_AWADDR = in_31__m_axi_m_axi_AWADDR;
  assign m_axi_in_31_AWBURST = in_31__m_axi_m_axi_AWBURST;
  assign m_axi_in_31_AWCACHE = in_31__m_axi_m_axi_AWCACHE;
  assign m_axi_in_31_AWID = in_31__m_axi_m_axi_AWID;
  assign m_axi_in_31_AWLEN = in_31__m_axi_m_axi_AWLEN;
  assign m_axi_in_31_AWLOCK = in_31__m_axi_m_axi_AWLOCK;
  assign m_axi_in_31_AWPROT = in_31__m_axi_m_axi_AWPROT;
  assign m_axi_in_31_AWQOS = in_31__m_axi_m_axi_AWQOS;
  assign in_31__m_axi_m_axi_AWREADY = m_axi_in_31_AWREADY;
  assign m_axi_in_31_AWSIZE = in_31__m_axi_m_axi_AWSIZE;
  assign m_axi_in_31_AWVALID = in_31__m_axi_m_axi_AWVALID;
  assign in_31__m_axi_m_axi_BID = m_axi_in_31_BID;
  assign m_axi_in_31_BREADY = in_31__m_axi_m_axi_BREADY;
  assign in_31__m_axi_m_axi_BRESP = m_axi_in_31_BRESP;
  assign in_31__m_axi_m_axi_BVALID = m_axi_in_31_BVALID;
  assign in_31__m_axi_m_axi_RDATA = m_axi_in_31_RDATA;
  assign in_31__m_axi_m_axi_RID = m_axi_in_31_RID;
  assign in_31__m_axi_m_axi_RLAST = m_axi_in_31_RLAST;
  assign m_axi_in_31_RREADY = in_31__m_axi_m_axi_RREADY;
  assign in_31__m_axi_m_axi_RRESP = m_axi_in_31_RRESP;
  assign in_31__m_axi_m_axi_RVALID = m_axi_in_31_RVALID;
  assign m_axi_in_31_WDATA = in_31__m_axi_m_axi_WDATA;
  assign m_axi_in_31_WLAST = in_31__m_axi_m_axi_WLAST;
  assign in_31__m_axi_m_axi_WREADY = m_axi_in_31_WREADY;
  assign m_axi_in_31_WSTRB = in_31__m_axi_m_axi_WSTRB;
  assign m_axi_in_31_WVALID = in_31__m_axi_m_axi_WVALID;
  assign in_31__m_axi_read_addr_din = in_31_read_addr__din;
  assign in_31_read_addr__full_n = in_31__m_axi_read_addr_full_n;
  assign in_31__m_axi_read_addr_write = in_31_read_addr__write;
  assign in_31_read_data__dout = in_31__m_axi_read_data_dout;
  assign in_31_read_data__empty_n = in_31__m_axi_read_data_empty_n;
  assign in_31__m_axi_read_data_read = in_31_read_data__read;
  assign in_31__m_axi_rst = ~ ap_rst_n;
  assign in_31__m_axi_write_addr_din = in_31_write_addr__din;
  assign in_31_write_addr__full_n = in_31__m_axi_write_addr_full_n;
  assign in_31__m_axi_write_addr_write = in_31_write_addr__write;
  assign in_31__m_axi_write_data_din = in_31_write_data__din;
  assign in_31_write_data__full_n = in_31__m_axi_write_data_full_n;
  assign in_31__m_axi_write_data_write = in_31_write_data__write;
  assign in_31_write_resp__dout = in_31__m_axi_write_resp_dout;
  assign in_31_write_resp__empty_n = in_31__m_axi_write_resp_empty_n;
  assign in_31__m_axi_write_resp_read = in_31_write_resp__read;
  assign in_32__m_axi_clk = ap_clk;
  assign m_axi_in_32_ARADDR = in_32__m_axi_m_axi_ARADDR;
  assign m_axi_in_32_ARBURST = in_32__m_axi_m_axi_ARBURST;
  assign m_axi_in_32_ARCACHE = in_32__m_axi_m_axi_ARCACHE;
  assign m_axi_in_32_ARID = in_32__m_axi_m_axi_ARID;
  assign m_axi_in_32_ARLEN = in_32__m_axi_m_axi_ARLEN;
  assign m_axi_in_32_ARLOCK = in_32__m_axi_m_axi_ARLOCK;
  assign m_axi_in_32_ARPROT = in_32__m_axi_m_axi_ARPROT;
  assign m_axi_in_32_ARQOS = in_32__m_axi_m_axi_ARQOS;
  assign in_32__m_axi_m_axi_ARREADY = m_axi_in_32_ARREADY;
  assign m_axi_in_32_ARSIZE = in_32__m_axi_m_axi_ARSIZE;
  assign m_axi_in_32_ARVALID = in_32__m_axi_m_axi_ARVALID;
  assign m_axi_in_32_AWADDR = in_32__m_axi_m_axi_AWADDR;
  assign m_axi_in_32_AWBURST = in_32__m_axi_m_axi_AWBURST;
  assign m_axi_in_32_AWCACHE = in_32__m_axi_m_axi_AWCACHE;
  assign m_axi_in_32_AWID = in_32__m_axi_m_axi_AWID;
  assign m_axi_in_32_AWLEN = in_32__m_axi_m_axi_AWLEN;
  assign m_axi_in_32_AWLOCK = in_32__m_axi_m_axi_AWLOCK;
  assign m_axi_in_32_AWPROT = in_32__m_axi_m_axi_AWPROT;
  assign m_axi_in_32_AWQOS = in_32__m_axi_m_axi_AWQOS;
  assign in_32__m_axi_m_axi_AWREADY = m_axi_in_32_AWREADY;
  assign m_axi_in_32_AWSIZE = in_32__m_axi_m_axi_AWSIZE;
  assign m_axi_in_32_AWVALID = in_32__m_axi_m_axi_AWVALID;
  assign in_32__m_axi_m_axi_BID = m_axi_in_32_BID;
  assign m_axi_in_32_BREADY = in_32__m_axi_m_axi_BREADY;
  assign in_32__m_axi_m_axi_BRESP = m_axi_in_32_BRESP;
  assign in_32__m_axi_m_axi_BVALID = m_axi_in_32_BVALID;
  assign in_32__m_axi_m_axi_RDATA = m_axi_in_32_RDATA;
  assign in_32__m_axi_m_axi_RID = m_axi_in_32_RID;
  assign in_32__m_axi_m_axi_RLAST = m_axi_in_32_RLAST;
  assign m_axi_in_32_RREADY = in_32__m_axi_m_axi_RREADY;
  assign in_32__m_axi_m_axi_RRESP = m_axi_in_32_RRESP;
  assign in_32__m_axi_m_axi_RVALID = m_axi_in_32_RVALID;
  assign m_axi_in_32_WDATA = in_32__m_axi_m_axi_WDATA;
  assign m_axi_in_32_WLAST = in_32__m_axi_m_axi_WLAST;
  assign in_32__m_axi_m_axi_WREADY = m_axi_in_32_WREADY;
  assign m_axi_in_32_WSTRB = in_32__m_axi_m_axi_WSTRB;
  assign m_axi_in_32_WVALID = in_32__m_axi_m_axi_WVALID;
  assign in_32__m_axi_read_addr_din = in_32_read_addr__din;
  assign in_32_read_addr__full_n = in_32__m_axi_read_addr_full_n;
  assign in_32__m_axi_read_addr_write = in_32_read_addr__write;
  assign in_32_read_data__dout = in_32__m_axi_read_data_dout;
  assign in_32_read_data__empty_n = in_32__m_axi_read_data_empty_n;
  assign in_32__m_axi_read_data_read = in_32_read_data__read;
  assign in_32__m_axi_rst = ~ ap_rst_n;
  assign in_32__m_axi_write_addr_din = in_32_write_addr__din;
  assign in_32_write_addr__full_n = in_32__m_axi_write_addr_full_n;
  assign in_32__m_axi_write_addr_write = in_32_write_addr__write;
  assign in_32__m_axi_write_data_din = in_32_write_data__din;
  assign in_32_write_data__full_n = in_32__m_axi_write_data_full_n;
  assign in_32__m_axi_write_data_write = in_32_write_data__write;
  assign in_32_write_resp__dout = in_32__m_axi_write_resp_dout;
  assign in_32_write_resp__empty_n = in_32__m_axi_write_resp_empty_n;
  assign in_32__m_axi_write_resp_read = in_32_write_resp__read;
  assign in_33__m_axi_clk = ap_clk;
  assign m_axi_in_33_ARADDR = in_33__m_axi_m_axi_ARADDR;
  assign m_axi_in_33_ARBURST = in_33__m_axi_m_axi_ARBURST;
  assign m_axi_in_33_ARCACHE = in_33__m_axi_m_axi_ARCACHE;
  assign m_axi_in_33_ARID = in_33__m_axi_m_axi_ARID;
  assign m_axi_in_33_ARLEN = in_33__m_axi_m_axi_ARLEN;
  assign m_axi_in_33_ARLOCK = in_33__m_axi_m_axi_ARLOCK;
  assign m_axi_in_33_ARPROT = in_33__m_axi_m_axi_ARPROT;
  assign m_axi_in_33_ARQOS = in_33__m_axi_m_axi_ARQOS;
  assign in_33__m_axi_m_axi_ARREADY = m_axi_in_33_ARREADY;
  assign m_axi_in_33_ARSIZE = in_33__m_axi_m_axi_ARSIZE;
  assign m_axi_in_33_ARVALID = in_33__m_axi_m_axi_ARVALID;
  assign m_axi_in_33_AWADDR = in_33__m_axi_m_axi_AWADDR;
  assign m_axi_in_33_AWBURST = in_33__m_axi_m_axi_AWBURST;
  assign m_axi_in_33_AWCACHE = in_33__m_axi_m_axi_AWCACHE;
  assign m_axi_in_33_AWID = in_33__m_axi_m_axi_AWID;
  assign m_axi_in_33_AWLEN = in_33__m_axi_m_axi_AWLEN;
  assign m_axi_in_33_AWLOCK = in_33__m_axi_m_axi_AWLOCK;
  assign m_axi_in_33_AWPROT = in_33__m_axi_m_axi_AWPROT;
  assign m_axi_in_33_AWQOS = in_33__m_axi_m_axi_AWQOS;
  assign in_33__m_axi_m_axi_AWREADY = m_axi_in_33_AWREADY;
  assign m_axi_in_33_AWSIZE = in_33__m_axi_m_axi_AWSIZE;
  assign m_axi_in_33_AWVALID = in_33__m_axi_m_axi_AWVALID;
  assign in_33__m_axi_m_axi_BID = m_axi_in_33_BID;
  assign m_axi_in_33_BREADY = in_33__m_axi_m_axi_BREADY;
  assign in_33__m_axi_m_axi_BRESP = m_axi_in_33_BRESP;
  assign in_33__m_axi_m_axi_BVALID = m_axi_in_33_BVALID;
  assign in_33__m_axi_m_axi_RDATA = m_axi_in_33_RDATA;
  assign in_33__m_axi_m_axi_RID = m_axi_in_33_RID;
  assign in_33__m_axi_m_axi_RLAST = m_axi_in_33_RLAST;
  assign m_axi_in_33_RREADY = in_33__m_axi_m_axi_RREADY;
  assign in_33__m_axi_m_axi_RRESP = m_axi_in_33_RRESP;
  assign in_33__m_axi_m_axi_RVALID = m_axi_in_33_RVALID;
  assign m_axi_in_33_WDATA = in_33__m_axi_m_axi_WDATA;
  assign m_axi_in_33_WLAST = in_33__m_axi_m_axi_WLAST;
  assign in_33__m_axi_m_axi_WREADY = m_axi_in_33_WREADY;
  assign m_axi_in_33_WSTRB = in_33__m_axi_m_axi_WSTRB;
  assign m_axi_in_33_WVALID = in_33__m_axi_m_axi_WVALID;
  assign in_33__m_axi_read_addr_din = in_33_read_addr__din;
  assign in_33_read_addr__full_n = in_33__m_axi_read_addr_full_n;
  assign in_33__m_axi_read_addr_write = in_33_read_addr__write;
  assign in_33_read_data__dout = in_33__m_axi_read_data_dout;
  assign in_33_read_data__empty_n = in_33__m_axi_read_data_empty_n;
  assign in_33__m_axi_read_data_read = in_33_read_data__read;
  assign in_33__m_axi_rst = ~ ap_rst_n;
  assign in_33__m_axi_write_addr_din = in_33_write_addr__din;
  assign in_33_write_addr__full_n = in_33__m_axi_write_addr_full_n;
  assign in_33__m_axi_write_addr_write = in_33_write_addr__write;
  assign in_33__m_axi_write_data_din = in_33_write_data__din;
  assign in_33_write_data__full_n = in_33__m_axi_write_data_full_n;
  assign in_33__m_axi_write_data_write = in_33_write_data__write;
  assign in_33_write_resp__dout = in_33__m_axi_write_resp_dout;
  assign in_33_write_resp__empty_n = in_33__m_axi_write_resp_empty_n;
  assign in_33__m_axi_write_resp_read = in_33_write_resp__read;
  assign in_34__m_axi_clk = ap_clk;
  assign m_axi_in_34_ARADDR = in_34__m_axi_m_axi_ARADDR;
  assign m_axi_in_34_ARBURST = in_34__m_axi_m_axi_ARBURST;
  assign m_axi_in_34_ARCACHE = in_34__m_axi_m_axi_ARCACHE;
  assign m_axi_in_34_ARID = in_34__m_axi_m_axi_ARID;
  assign m_axi_in_34_ARLEN = in_34__m_axi_m_axi_ARLEN;
  assign m_axi_in_34_ARLOCK = in_34__m_axi_m_axi_ARLOCK;
  assign m_axi_in_34_ARPROT = in_34__m_axi_m_axi_ARPROT;
  assign m_axi_in_34_ARQOS = in_34__m_axi_m_axi_ARQOS;
  assign in_34__m_axi_m_axi_ARREADY = m_axi_in_34_ARREADY;
  assign m_axi_in_34_ARSIZE = in_34__m_axi_m_axi_ARSIZE;
  assign m_axi_in_34_ARVALID = in_34__m_axi_m_axi_ARVALID;
  assign m_axi_in_34_AWADDR = in_34__m_axi_m_axi_AWADDR;
  assign m_axi_in_34_AWBURST = in_34__m_axi_m_axi_AWBURST;
  assign m_axi_in_34_AWCACHE = in_34__m_axi_m_axi_AWCACHE;
  assign m_axi_in_34_AWID = in_34__m_axi_m_axi_AWID;
  assign m_axi_in_34_AWLEN = in_34__m_axi_m_axi_AWLEN;
  assign m_axi_in_34_AWLOCK = in_34__m_axi_m_axi_AWLOCK;
  assign m_axi_in_34_AWPROT = in_34__m_axi_m_axi_AWPROT;
  assign m_axi_in_34_AWQOS = in_34__m_axi_m_axi_AWQOS;
  assign in_34__m_axi_m_axi_AWREADY = m_axi_in_34_AWREADY;
  assign m_axi_in_34_AWSIZE = in_34__m_axi_m_axi_AWSIZE;
  assign m_axi_in_34_AWVALID = in_34__m_axi_m_axi_AWVALID;
  assign in_34__m_axi_m_axi_BID = m_axi_in_34_BID;
  assign m_axi_in_34_BREADY = in_34__m_axi_m_axi_BREADY;
  assign in_34__m_axi_m_axi_BRESP = m_axi_in_34_BRESP;
  assign in_34__m_axi_m_axi_BVALID = m_axi_in_34_BVALID;
  assign in_34__m_axi_m_axi_RDATA = m_axi_in_34_RDATA;
  assign in_34__m_axi_m_axi_RID = m_axi_in_34_RID;
  assign in_34__m_axi_m_axi_RLAST = m_axi_in_34_RLAST;
  assign m_axi_in_34_RREADY = in_34__m_axi_m_axi_RREADY;
  assign in_34__m_axi_m_axi_RRESP = m_axi_in_34_RRESP;
  assign in_34__m_axi_m_axi_RVALID = m_axi_in_34_RVALID;
  assign m_axi_in_34_WDATA = in_34__m_axi_m_axi_WDATA;
  assign m_axi_in_34_WLAST = in_34__m_axi_m_axi_WLAST;
  assign in_34__m_axi_m_axi_WREADY = m_axi_in_34_WREADY;
  assign m_axi_in_34_WSTRB = in_34__m_axi_m_axi_WSTRB;
  assign m_axi_in_34_WVALID = in_34__m_axi_m_axi_WVALID;
  assign in_34__m_axi_read_addr_din = in_34_read_addr__din;
  assign in_34_read_addr__full_n = in_34__m_axi_read_addr_full_n;
  assign in_34__m_axi_read_addr_write = in_34_read_addr__write;
  assign in_34_read_data__dout = in_34__m_axi_read_data_dout;
  assign in_34_read_data__empty_n = in_34__m_axi_read_data_empty_n;
  assign in_34__m_axi_read_data_read = in_34_read_data__read;
  assign in_34__m_axi_rst = ~ ap_rst_n;
  assign in_34__m_axi_write_addr_din = in_34_write_addr__din;
  assign in_34_write_addr__full_n = in_34__m_axi_write_addr_full_n;
  assign in_34__m_axi_write_addr_write = in_34_write_addr__write;
  assign in_34__m_axi_write_data_din = in_34_write_data__din;
  assign in_34_write_data__full_n = in_34__m_axi_write_data_full_n;
  assign in_34__m_axi_write_data_write = in_34_write_data__write;
  assign in_34_write_resp__dout = in_34__m_axi_write_resp_dout;
  assign in_34_write_resp__empty_n = in_34__m_axi_write_resp_empty_n;
  assign in_34__m_axi_write_resp_read = in_34_write_resp__read;
  assign in_35__m_axi_clk = ap_clk;
  assign m_axi_in_35_ARADDR = in_35__m_axi_m_axi_ARADDR;
  assign m_axi_in_35_ARBURST = in_35__m_axi_m_axi_ARBURST;
  assign m_axi_in_35_ARCACHE = in_35__m_axi_m_axi_ARCACHE;
  assign m_axi_in_35_ARID = in_35__m_axi_m_axi_ARID;
  assign m_axi_in_35_ARLEN = in_35__m_axi_m_axi_ARLEN;
  assign m_axi_in_35_ARLOCK = in_35__m_axi_m_axi_ARLOCK;
  assign m_axi_in_35_ARPROT = in_35__m_axi_m_axi_ARPROT;
  assign m_axi_in_35_ARQOS = in_35__m_axi_m_axi_ARQOS;
  assign in_35__m_axi_m_axi_ARREADY = m_axi_in_35_ARREADY;
  assign m_axi_in_35_ARSIZE = in_35__m_axi_m_axi_ARSIZE;
  assign m_axi_in_35_ARVALID = in_35__m_axi_m_axi_ARVALID;
  assign m_axi_in_35_AWADDR = in_35__m_axi_m_axi_AWADDR;
  assign m_axi_in_35_AWBURST = in_35__m_axi_m_axi_AWBURST;
  assign m_axi_in_35_AWCACHE = in_35__m_axi_m_axi_AWCACHE;
  assign m_axi_in_35_AWID = in_35__m_axi_m_axi_AWID;
  assign m_axi_in_35_AWLEN = in_35__m_axi_m_axi_AWLEN;
  assign m_axi_in_35_AWLOCK = in_35__m_axi_m_axi_AWLOCK;
  assign m_axi_in_35_AWPROT = in_35__m_axi_m_axi_AWPROT;
  assign m_axi_in_35_AWQOS = in_35__m_axi_m_axi_AWQOS;
  assign in_35__m_axi_m_axi_AWREADY = m_axi_in_35_AWREADY;
  assign m_axi_in_35_AWSIZE = in_35__m_axi_m_axi_AWSIZE;
  assign m_axi_in_35_AWVALID = in_35__m_axi_m_axi_AWVALID;
  assign in_35__m_axi_m_axi_BID = m_axi_in_35_BID;
  assign m_axi_in_35_BREADY = in_35__m_axi_m_axi_BREADY;
  assign in_35__m_axi_m_axi_BRESP = m_axi_in_35_BRESP;
  assign in_35__m_axi_m_axi_BVALID = m_axi_in_35_BVALID;
  assign in_35__m_axi_m_axi_RDATA = m_axi_in_35_RDATA;
  assign in_35__m_axi_m_axi_RID = m_axi_in_35_RID;
  assign in_35__m_axi_m_axi_RLAST = m_axi_in_35_RLAST;
  assign m_axi_in_35_RREADY = in_35__m_axi_m_axi_RREADY;
  assign in_35__m_axi_m_axi_RRESP = m_axi_in_35_RRESP;
  assign in_35__m_axi_m_axi_RVALID = m_axi_in_35_RVALID;
  assign m_axi_in_35_WDATA = in_35__m_axi_m_axi_WDATA;
  assign m_axi_in_35_WLAST = in_35__m_axi_m_axi_WLAST;
  assign in_35__m_axi_m_axi_WREADY = m_axi_in_35_WREADY;
  assign m_axi_in_35_WSTRB = in_35__m_axi_m_axi_WSTRB;
  assign m_axi_in_35_WVALID = in_35__m_axi_m_axi_WVALID;
  assign in_35__m_axi_read_addr_din = in_35_read_addr__din;
  assign in_35_read_addr__full_n = in_35__m_axi_read_addr_full_n;
  assign in_35__m_axi_read_addr_write = in_35_read_addr__write;
  assign in_35_read_data__dout = in_35__m_axi_read_data_dout;
  assign in_35_read_data__empty_n = in_35__m_axi_read_data_empty_n;
  assign in_35__m_axi_read_data_read = in_35_read_data__read;
  assign in_35__m_axi_rst = ~ ap_rst_n;
  assign in_35__m_axi_write_addr_din = in_35_write_addr__din;
  assign in_35_write_addr__full_n = in_35__m_axi_write_addr_full_n;
  assign in_35__m_axi_write_addr_write = in_35_write_addr__write;
  assign in_35__m_axi_write_data_din = in_35_write_data__din;
  assign in_35_write_data__full_n = in_35__m_axi_write_data_full_n;
  assign in_35__m_axi_write_data_write = in_35_write_data__write;
  assign in_35_write_resp__dout = in_35__m_axi_write_resp_dout;
  assign in_35_write_resp__empty_n = in_35__m_axi_write_resp_empty_n;
  assign in_35__m_axi_write_resp_read = in_35_write_resp__read;
  assign in_36__m_axi_clk = ap_clk;
  assign m_axi_in_36_ARADDR = in_36__m_axi_m_axi_ARADDR;
  assign m_axi_in_36_ARBURST = in_36__m_axi_m_axi_ARBURST;
  assign m_axi_in_36_ARCACHE = in_36__m_axi_m_axi_ARCACHE;
  assign m_axi_in_36_ARID = in_36__m_axi_m_axi_ARID;
  assign m_axi_in_36_ARLEN = in_36__m_axi_m_axi_ARLEN;
  assign m_axi_in_36_ARLOCK = in_36__m_axi_m_axi_ARLOCK;
  assign m_axi_in_36_ARPROT = in_36__m_axi_m_axi_ARPROT;
  assign m_axi_in_36_ARQOS = in_36__m_axi_m_axi_ARQOS;
  assign in_36__m_axi_m_axi_ARREADY = m_axi_in_36_ARREADY;
  assign m_axi_in_36_ARSIZE = in_36__m_axi_m_axi_ARSIZE;
  assign m_axi_in_36_ARVALID = in_36__m_axi_m_axi_ARVALID;
  assign m_axi_in_36_AWADDR = in_36__m_axi_m_axi_AWADDR;
  assign m_axi_in_36_AWBURST = in_36__m_axi_m_axi_AWBURST;
  assign m_axi_in_36_AWCACHE = in_36__m_axi_m_axi_AWCACHE;
  assign m_axi_in_36_AWID = in_36__m_axi_m_axi_AWID;
  assign m_axi_in_36_AWLEN = in_36__m_axi_m_axi_AWLEN;
  assign m_axi_in_36_AWLOCK = in_36__m_axi_m_axi_AWLOCK;
  assign m_axi_in_36_AWPROT = in_36__m_axi_m_axi_AWPROT;
  assign m_axi_in_36_AWQOS = in_36__m_axi_m_axi_AWQOS;
  assign in_36__m_axi_m_axi_AWREADY = m_axi_in_36_AWREADY;
  assign m_axi_in_36_AWSIZE = in_36__m_axi_m_axi_AWSIZE;
  assign m_axi_in_36_AWVALID = in_36__m_axi_m_axi_AWVALID;
  assign in_36__m_axi_m_axi_BID = m_axi_in_36_BID;
  assign m_axi_in_36_BREADY = in_36__m_axi_m_axi_BREADY;
  assign in_36__m_axi_m_axi_BRESP = m_axi_in_36_BRESP;
  assign in_36__m_axi_m_axi_BVALID = m_axi_in_36_BVALID;
  assign in_36__m_axi_m_axi_RDATA = m_axi_in_36_RDATA;
  assign in_36__m_axi_m_axi_RID = m_axi_in_36_RID;
  assign in_36__m_axi_m_axi_RLAST = m_axi_in_36_RLAST;
  assign m_axi_in_36_RREADY = in_36__m_axi_m_axi_RREADY;
  assign in_36__m_axi_m_axi_RRESP = m_axi_in_36_RRESP;
  assign in_36__m_axi_m_axi_RVALID = m_axi_in_36_RVALID;
  assign m_axi_in_36_WDATA = in_36__m_axi_m_axi_WDATA;
  assign m_axi_in_36_WLAST = in_36__m_axi_m_axi_WLAST;
  assign in_36__m_axi_m_axi_WREADY = m_axi_in_36_WREADY;
  assign m_axi_in_36_WSTRB = in_36__m_axi_m_axi_WSTRB;
  assign m_axi_in_36_WVALID = in_36__m_axi_m_axi_WVALID;
  assign in_36__m_axi_read_addr_din = in_36_read_addr__din;
  assign in_36_read_addr__full_n = in_36__m_axi_read_addr_full_n;
  assign in_36__m_axi_read_addr_write = in_36_read_addr__write;
  assign in_36_read_data__dout = in_36__m_axi_read_data_dout;
  assign in_36_read_data__empty_n = in_36__m_axi_read_data_empty_n;
  assign in_36__m_axi_read_data_read = in_36_read_data__read;
  assign in_36__m_axi_rst = ~ ap_rst_n;
  assign in_36__m_axi_write_addr_din = in_36_write_addr__din;
  assign in_36_write_addr__full_n = in_36__m_axi_write_addr_full_n;
  assign in_36__m_axi_write_addr_write = in_36_write_addr__write;
  assign in_36__m_axi_write_data_din = in_36_write_data__din;
  assign in_36_write_data__full_n = in_36__m_axi_write_data_full_n;
  assign in_36__m_axi_write_data_write = in_36_write_data__write;
  assign in_36_write_resp__dout = in_36__m_axi_write_resp_dout;
  assign in_36_write_resp__empty_n = in_36__m_axi_write_resp_empty_n;
  assign in_36__m_axi_write_resp_read = in_36_write_resp__read;
  assign in_37__m_axi_clk = ap_clk;
  assign m_axi_in_37_ARADDR = in_37__m_axi_m_axi_ARADDR;
  assign m_axi_in_37_ARBURST = in_37__m_axi_m_axi_ARBURST;
  assign m_axi_in_37_ARCACHE = in_37__m_axi_m_axi_ARCACHE;
  assign m_axi_in_37_ARID = in_37__m_axi_m_axi_ARID;
  assign m_axi_in_37_ARLEN = in_37__m_axi_m_axi_ARLEN;
  assign m_axi_in_37_ARLOCK = in_37__m_axi_m_axi_ARLOCK;
  assign m_axi_in_37_ARPROT = in_37__m_axi_m_axi_ARPROT;
  assign m_axi_in_37_ARQOS = in_37__m_axi_m_axi_ARQOS;
  assign in_37__m_axi_m_axi_ARREADY = m_axi_in_37_ARREADY;
  assign m_axi_in_37_ARSIZE = in_37__m_axi_m_axi_ARSIZE;
  assign m_axi_in_37_ARVALID = in_37__m_axi_m_axi_ARVALID;
  assign m_axi_in_37_AWADDR = in_37__m_axi_m_axi_AWADDR;
  assign m_axi_in_37_AWBURST = in_37__m_axi_m_axi_AWBURST;
  assign m_axi_in_37_AWCACHE = in_37__m_axi_m_axi_AWCACHE;
  assign m_axi_in_37_AWID = in_37__m_axi_m_axi_AWID;
  assign m_axi_in_37_AWLEN = in_37__m_axi_m_axi_AWLEN;
  assign m_axi_in_37_AWLOCK = in_37__m_axi_m_axi_AWLOCK;
  assign m_axi_in_37_AWPROT = in_37__m_axi_m_axi_AWPROT;
  assign m_axi_in_37_AWQOS = in_37__m_axi_m_axi_AWQOS;
  assign in_37__m_axi_m_axi_AWREADY = m_axi_in_37_AWREADY;
  assign m_axi_in_37_AWSIZE = in_37__m_axi_m_axi_AWSIZE;
  assign m_axi_in_37_AWVALID = in_37__m_axi_m_axi_AWVALID;
  assign in_37__m_axi_m_axi_BID = m_axi_in_37_BID;
  assign m_axi_in_37_BREADY = in_37__m_axi_m_axi_BREADY;
  assign in_37__m_axi_m_axi_BRESP = m_axi_in_37_BRESP;
  assign in_37__m_axi_m_axi_BVALID = m_axi_in_37_BVALID;
  assign in_37__m_axi_m_axi_RDATA = m_axi_in_37_RDATA;
  assign in_37__m_axi_m_axi_RID = m_axi_in_37_RID;
  assign in_37__m_axi_m_axi_RLAST = m_axi_in_37_RLAST;
  assign m_axi_in_37_RREADY = in_37__m_axi_m_axi_RREADY;
  assign in_37__m_axi_m_axi_RRESP = m_axi_in_37_RRESP;
  assign in_37__m_axi_m_axi_RVALID = m_axi_in_37_RVALID;
  assign m_axi_in_37_WDATA = in_37__m_axi_m_axi_WDATA;
  assign m_axi_in_37_WLAST = in_37__m_axi_m_axi_WLAST;
  assign in_37__m_axi_m_axi_WREADY = m_axi_in_37_WREADY;
  assign m_axi_in_37_WSTRB = in_37__m_axi_m_axi_WSTRB;
  assign m_axi_in_37_WVALID = in_37__m_axi_m_axi_WVALID;
  assign in_37__m_axi_read_addr_din = in_37_read_addr__din;
  assign in_37_read_addr__full_n = in_37__m_axi_read_addr_full_n;
  assign in_37__m_axi_read_addr_write = in_37_read_addr__write;
  assign in_37_read_data__dout = in_37__m_axi_read_data_dout;
  assign in_37_read_data__empty_n = in_37__m_axi_read_data_empty_n;
  assign in_37__m_axi_read_data_read = in_37_read_data__read;
  assign in_37__m_axi_rst = ~ ap_rst_n;
  assign in_37__m_axi_write_addr_din = in_37_write_addr__din;
  assign in_37_write_addr__full_n = in_37__m_axi_write_addr_full_n;
  assign in_37__m_axi_write_addr_write = in_37_write_addr__write;
  assign in_37__m_axi_write_data_din = in_37_write_data__din;
  assign in_37_write_data__full_n = in_37__m_axi_write_data_full_n;
  assign in_37__m_axi_write_data_write = in_37_write_data__write;
  assign in_37_write_resp__dout = in_37__m_axi_write_resp_dout;
  assign in_37_write_resp__empty_n = in_37__m_axi_write_resp_empty_n;
  assign in_37__m_axi_write_resp_read = in_37_write_resp__read;
  assign in_38__m_axi_clk = ap_clk;
  assign m_axi_in_38_ARADDR = in_38__m_axi_m_axi_ARADDR;
  assign m_axi_in_38_ARBURST = in_38__m_axi_m_axi_ARBURST;
  assign m_axi_in_38_ARCACHE = in_38__m_axi_m_axi_ARCACHE;
  assign m_axi_in_38_ARID = in_38__m_axi_m_axi_ARID;
  assign m_axi_in_38_ARLEN = in_38__m_axi_m_axi_ARLEN;
  assign m_axi_in_38_ARLOCK = in_38__m_axi_m_axi_ARLOCK;
  assign m_axi_in_38_ARPROT = in_38__m_axi_m_axi_ARPROT;
  assign m_axi_in_38_ARQOS = in_38__m_axi_m_axi_ARQOS;
  assign in_38__m_axi_m_axi_ARREADY = m_axi_in_38_ARREADY;
  assign m_axi_in_38_ARSIZE = in_38__m_axi_m_axi_ARSIZE;
  assign m_axi_in_38_ARVALID = in_38__m_axi_m_axi_ARVALID;
  assign m_axi_in_38_AWADDR = in_38__m_axi_m_axi_AWADDR;
  assign m_axi_in_38_AWBURST = in_38__m_axi_m_axi_AWBURST;
  assign m_axi_in_38_AWCACHE = in_38__m_axi_m_axi_AWCACHE;
  assign m_axi_in_38_AWID = in_38__m_axi_m_axi_AWID;
  assign m_axi_in_38_AWLEN = in_38__m_axi_m_axi_AWLEN;
  assign m_axi_in_38_AWLOCK = in_38__m_axi_m_axi_AWLOCK;
  assign m_axi_in_38_AWPROT = in_38__m_axi_m_axi_AWPROT;
  assign m_axi_in_38_AWQOS = in_38__m_axi_m_axi_AWQOS;
  assign in_38__m_axi_m_axi_AWREADY = m_axi_in_38_AWREADY;
  assign m_axi_in_38_AWSIZE = in_38__m_axi_m_axi_AWSIZE;
  assign m_axi_in_38_AWVALID = in_38__m_axi_m_axi_AWVALID;
  assign in_38__m_axi_m_axi_BID = m_axi_in_38_BID;
  assign m_axi_in_38_BREADY = in_38__m_axi_m_axi_BREADY;
  assign in_38__m_axi_m_axi_BRESP = m_axi_in_38_BRESP;
  assign in_38__m_axi_m_axi_BVALID = m_axi_in_38_BVALID;
  assign in_38__m_axi_m_axi_RDATA = m_axi_in_38_RDATA;
  assign in_38__m_axi_m_axi_RID = m_axi_in_38_RID;
  assign in_38__m_axi_m_axi_RLAST = m_axi_in_38_RLAST;
  assign m_axi_in_38_RREADY = in_38__m_axi_m_axi_RREADY;
  assign in_38__m_axi_m_axi_RRESP = m_axi_in_38_RRESP;
  assign in_38__m_axi_m_axi_RVALID = m_axi_in_38_RVALID;
  assign m_axi_in_38_WDATA = in_38__m_axi_m_axi_WDATA;
  assign m_axi_in_38_WLAST = in_38__m_axi_m_axi_WLAST;
  assign in_38__m_axi_m_axi_WREADY = m_axi_in_38_WREADY;
  assign m_axi_in_38_WSTRB = in_38__m_axi_m_axi_WSTRB;
  assign m_axi_in_38_WVALID = in_38__m_axi_m_axi_WVALID;
  assign in_38__m_axi_read_addr_din = in_38_read_addr__din;
  assign in_38_read_addr__full_n = in_38__m_axi_read_addr_full_n;
  assign in_38__m_axi_read_addr_write = in_38_read_addr__write;
  assign in_38_read_data__dout = in_38__m_axi_read_data_dout;
  assign in_38_read_data__empty_n = in_38__m_axi_read_data_empty_n;
  assign in_38__m_axi_read_data_read = in_38_read_data__read;
  assign in_38__m_axi_rst = ~ ap_rst_n;
  assign in_38__m_axi_write_addr_din = in_38_write_addr__din;
  assign in_38_write_addr__full_n = in_38__m_axi_write_addr_full_n;
  assign in_38__m_axi_write_addr_write = in_38_write_addr__write;
  assign in_38__m_axi_write_data_din = in_38_write_data__din;
  assign in_38_write_data__full_n = in_38__m_axi_write_data_full_n;
  assign in_38__m_axi_write_data_write = in_38_write_data__write;
  assign in_38_write_resp__dout = in_38__m_axi_write_resp_dout;
  assign in_38_write_resp__empty_n = in_38__m_axi_write_resp_empty_n;
  assign in_38__m_axi_write_resp_read = in_38_write_resp__read;
  assign in_39__m_axi_clk = ap_clk;
  assign m_axi_in_39_ARADDR = in_39__m_axi_m_axi_ARADDR;
  assign m_axi_in_39_ARBURST = in_39__m_axi_m_axi_ARBURST;
  assign m_axi_in_39_ARCACHE = in_39__m_axi_m_axi_ARCACHE;
  assign m_axi_in_39_ARID = in_39__m_axi_m_axi_ARID;
  assign m_axi_in_39_ARLEN = in_39__m_axi_m_axi_ARLEN;
  assign m_axi_in_39_ARLOCK = in_39__m_axi_m_axi_ARLOCK;
  assign m_axi_in_39_ARPROT = in_39__m_axi_m_axi_ARPROT;
  assign m_axi_in_39_ARQOS = in_39__m_axi_m_axi_ARQOS;
  assign in_39__m_axi_m_axi_ARREADY = m_axi_in_39_ARREADY;
  assign m_axi_in_39_ARSIZE = in_39__m_axi_m_axi_ARSIZE;
  assign m_axi_in_39_ARVALID = in_39__m_axi_m_axi_ARVALID;
  assign m_axi_in_39_AWADDR = in_39__m_axi_m_axi_AWADDR;
  assign m_axi_in_39_AWBURST = in_39__m_axi_m_axi_AWBURST;
  assign m_axi_in_39_AWCACHE = in_39__m_axi_m_axi_AWCACHE;
  assign m_axi_in_39_AWID = in_39__m_axi_m_axi_AWID;
  assign m_axi_in_39_AWLEN = in_39__m_axi_m_axi_AWLEN;
  assign m_axi_in_39_AWLOCK = in_39__m_axi_m_axi_AWLOCK;
  assign m_axi_in_39_AWPROT = in_39__m_axi_m_axi_AWPROT;
  assign m_axi_in_39_AWQOS = in_39__m_axi_m_axi_AWQOS;
  assign in_39__m_axi_m_axi_AWREADY = m_axi_in_39_AWREADY;
  assign m_axi_in_39_AWSIZE = in_39__m_axi_m_axi_AWSIZE;
  assign m_axi_in_39_AWVALID = in_39__m_axi_m_axi_AWVALID;
  assign in_39__m_axi_m_axi_BID = m_axi_in_39_BID;
  assign m_axi_in_39_BREADY = in_39__m_axi_m_axi_BREADY;
  assign in_39__m_axi_m_axi_BRESP = m_axi_in_39_BRESP;
  assign in_39__m_axi_m_axi_BVALID = m_axi_in_39_BVALID;
  assign in_39__m_axi_m_axi_RDATA = m_axi_in_39_RDATA;
  assign in_39__m_axi_m_axi_RID = m_axi_in_39_RID;
  assign in_39__m_axi_m_axi_RLAST = m_axi_in_39_RLAST;
  assign m_axi_in_39_RREADY = in_39__m_axi_m_axi_RREADY;
  assign in_39__m_axi_m_axi_RRESP = m_axi_in_39_RRESP;
  assign in_39__m_axi_m_axi_RVALID = m_axi_in_39_RVALID;
  assign m_axi_in_39_WDATA = in_39__m_axi_m_axi_WDATA;
  assign m_axi_in_39_WLAST = in_39__m_axi_m_axi_WLAST;
  assign in_39__m_axi_m_axi_WREADY = m_axi_in_39_WREADY;
  assign m_axi_in_39_WSTRB = in_39__m_axi_m_axi_WSTRB;
  assign m_axi_in_39_WVALID = in_39__m_axi_m_axi_WVALID;
  assign in_39__m_axi_read_addr_din = in_39_read_addr__din;
  assign in_39_read_addr__full_n = in_39__m_axi_read_addr_full_n;
  assign in_39__m_axi_read_addr_write = in_39_read_addr__write;
  assign in_39_read_data__dout = in_39__m_axi_read_data_dout;
  assign in_39_read_data__empty_n = in_39__m_axi_read_data_empty_n;
  assign in_39__m_axi_read_data_read = in_39_read_data__read;
  assign in_39__m_axi_rst = ~ ap_rst_n;
  assign in_39__m_axi_write_addr_din = in_39_write_addr__din;
  assign in_39_write_addr__full_n = in_39__m_axi_write_addr_full_n;
  assign in_39__m_axi_write_addr_write = in_39_write_addr__write;
  assign in_39__m_axi_write_data_din = in_39_write_data__din;
  assign in_39_write_data__full_n = in_39__m_axi_write_data_full_n;
  assign in_39__m_axi_write_data_write = in_39_write_data__write;
  assign in_39_write_resp__dout = in_39__m_axi_write_resp_dout;
  assign in_39_write_resp__empty_n = in_39__m_axi_write_resp_empty_n;
  assign in_39__m_axi_write_resp_read = in_39_write_resp__read;
  assign in_4__m_axi_clk = ap_clk;
  assign m_axi_in_4_ARADDR = in_4__m_axi_m_axi_ARADDR;
  assign m_axi_in_4_ARBURST = in_4__m_axi_m_axi_ARBURST;
  assign m_axi_in_4_ARCACHE = in_4__m_axi_m_axi_ARCACHE;
  assign m_axi_in_4_ARID = in_4__m_axi_m_axi_ARID;
  assign m_axi_in_4_ARLEN = in_4__m_axi_m_axi_ARLEN;
  assign m_axi_in_4_ARLOCK = in_4__m_axi_m_axi_ARLOCK;
  assign m_axi_in_4_ARPROT = in_4__m_axi_m_axi_ARPROT;
  assign m_axi_in_4_ARQOS = in_4__m_axi_m_axi_ARQOS;
  assign in_4__m_axi_m_axi_ARREADY = m_axi_in_4_ARREADY;
  assign m_axi_in_4_ARSIZE = in_4__m_axi_m_axi_ARSIZE;
  assign m_axi_in_4_ARVALID = in_4__m_axi_m_axi_ARVALID;
  assign m_axi_in_4_AWADDR = in_4__m_axi_m_axi_AWADDR;
  assign m_axi_in_4_AWBURST = in_4__m_axi_m_axi_AWBURST;
  assign m_axi_in_4_AWCACHE = in_4__m_axi_m_axi_AWCACHE;
  assign m_axi_in_4_AWID = in_4__m_axi_m_axi_AWID;
  assign m_axi_in_4_AWLEN = in_4__m_axi_m_axi_AWLEN;
  assign m_axi_in_4_AWLOCK = in_4__m_axi_m_axi_AWLOCK;
  assign m_axi_in_4_AWPROT = in_4__m_axi_m_axi_AWPROT;
  assign m_axi_in_4_AWQOS = in_4__m_axi_m_axi_AWQOS;
  assign in_4__m_axi_m_axi_AWREADY = m_axi_in_4_AWREADY;
  assign m_axi_in_4_AWSIZE = in_4__m_axi_m_axi_AWSIZE;
  assign m_axi_in_4_AWVALID = in_4__m_axi_m_axi_AWVALID;
  assign in_4__m_axi_m_axi_BID = m_axi_in_4_BID;
  assign m_axi_in_4_BREADY = in_4__m_axi_m_axi_BREADY;
  assign in_4__m_axi_m_axi_BRESP = m_axi_in_4_BRESP;
  assign in_4__m_axi_m_axi_BVALID = m_axi_in_4_BVALID;
  assign in_4__m_axi_m_axi_RDATA = m_axi_in_4_RDATA;
  assign in_4__m_axi_m_axi_RID = m_axi_in_4_RID;
  assign in_4__m_axi_m_axi_RLAST = m_axi_in_4_RLAST;
  assign m_axi_in_4_RREADY = in_4__m_axi_m_axi_RREADY;
  assign in_4__m_axi_m_axi_RRESP = m_axi_in_4_RRESP;
  assign in_4__m_axi_m_axi_RVALID = m_axi_in_4_RVALID;
  assign m_axi_in_4_WDATA = in_4__m_axi_m_axi_WDATA;
  assign m_axi_in_4_WLAST = in_4__m_axi_m_axi_WLAST;
  assign in_4__m_axi_m_axi_WREADY = m_axi_in_4_WREADY;
  assign m_axi_in_4_WSTRB = in_4__m_axi_m_axi_WSTRB;
  assign m_axi_in_4_WVALID = in_4__m_axi_m_axi_WVALID;
  assign in_4__m_axi_read_addr_din = in_4_read_addr__din;
  assign in_4_read_addr__full_n = in_4__m_axi_read_addr_full_n;
  assign in_4__m_axi_read_addr_write = in_4_read_addr__write;
  assign in_4_read_data__dout = in_4__m_axi_read_data_dout;
  assign in_4_read_data__empty_n = in_4__m_axi_read_data_empty_n;
  assign in_4__m_axi_read_data_read = in_4_read_data__read;
  assign in_4__m_axi_rst = ~ ap_rst_n;
  assign in_4__m_axi_write_addr_din = in_4_write_addr__din;
  assign in_4_write_addr__full_n = in_4__m_axi_write_addr_full_n;
  assign in_4__m_axi_write_addr_write = in_4_write_addr__write;
  assign in_4__m_axi_write_data_din = in_4_write_data__din;
  assign in_4_write_data__full_n = in_4__m_axi_write_data_full_n;
  assign in_4__m_axi_write_data_write = in_4_write_data__write;
  assign in_4_write_resp__dout = in_4__m_axi_write_resp_dout;
  assign in_4_write_resp__empty_n = in_4__m_axi_write_resp_empty_n;
  assign in_4__m_axi_write_resp_read = in_4_write_resp__read;
  assign in_40__m_axi_clk = ap_clk;
  assign m_axi_in_40_ARADDR = in_40__m_axi_m_axi_ARADDR;
  assign m_axi_in_40_ARBURST = in_40__m_axi_m_axi_ARBURST;
  assign m_axi_in_40_ARCACHE = in_40__m_axi_m_axi_ARCACHE;
  assign m_axi_in_40_ARID = in_40__m_axi_m_axi_ARID;
  assign m_axi_in_40_ARLEN = in_40__m_axi_m_axi_ARLEN;
  assign m_axi_in_40_ARLOCK = in_40__m_axi_m_axi_ARLOCK;
  assign m_axi_in_40_ARPROT = in_40__m_axi_m_axi_ARPROT;
  assign m_axi_in_40_ARQOS = in_40__m_axi_m_axi_ARQOS;
  assign in_40__m_axi_m_axi_ARREADY = m_axi_in_40_ARREADY;
  assign m_axi_in_40_ARSIZE = in_40__m_axi_m_axi_ARSIZE;
  assign m_axi_in_40_ARVALID = in_40__m_axi_m_axi_ARVALID;
  assign m_axi_in_40_AWADDR = in_40__m_axi_m_axi_AWADDR;
  assign m_axi_in_40_AWBURST = in_40__m_axi_m_axi_AWBURST;
  assign m_axi_in_40_AWCACHE = in_40__m_axi_m_axi_AWCACHE;
  assign m_axi_in_40_AWID = in_40__m_axi_m_axi_AWID;
  assign m_axi_in_40_AWLEN = in_40__m_axi_m_axi_AWLEN;
  assign m_axi_in_40_AWLOCK = in_40__m_axi_m_axi_AWLOCK;
  assign m_axi_in_40_AWPROT = in_40__m_axi_m_axi_AWPROT;
  assign m_axi_in_40_AWQOS = in_40__m_axi_m_axi_AWQOS;
  assign in_40__m_axi_m_axi_AWREADY = m_axi_in_40_AWREADY;
  assign m_axi_in_40_AWSIZE = in_40__m_axi_m_axi_AWSIZE;
  assign m_axi_in_40_AWVALID = in_40__m_axi_m_axi_AWVALID;
  assign in_40__m_axi_m_axi_BID = m_axi_in_40_BID;
  assign m_axi_in_40_BREADY = in_40__m_axi_m_axi_BREADY;
  assign in_40__m_axi_m_axi_BRESP = m_axi_in_40_BRESP;
  assign in_40__m_axi_m_axi_BVALID = m_axi_in_40_BVALID;
  assign in_40__m_axi_m_axi_RDATA = m_axi_in_40_RDATA;
  assign in_40__m_axi_m_axi_RID = m_axi_in_40_RID;
  assign in_40__m_axi_m_axi_RLAST = m_axi_in_40_RLAST;
  assign m_axi_in_40_RREADY = in_40__m_axi_m_axi_RREADY;
  assign in_40__m_axi_m_axi_RRESP = m_axi_in_40_RRESP;
  assign in_40__m_axi_m_axi_RVALID = m_axi_in_40_RVALID;
  assign m_axi_in_40_WDATA = in_40__m_axi_m_axi_WDATA;
  assign m_axi_in_40_WLAST = in_40__m_axi_m_axi_WLAST;
  assign in_40__m_axi_m_axi_WREADY = m_axi_in_40_WREADY;
  assign m_axi_in_40_WSTRB = in_40__m_axi_m_axi_WSTRB;
  assign m_axi_in_40_WVALID = in_40__m_axi_m_axi_WVALID;
  assign in_40__m_axi_read_addr_din = in_40_read_addr__din;
  assign in_40_read_addr__full_n = in_40__m_axi_read_addr_full_n;
  assign in_40__m_axi_read_addr_write = in_40_read_addr__write;
  assign in_40_read_data__dout = in_40__m_axi_read_data_dout;
  assign in_40_read_data__empty_n = in_40__m_axi_read_data_empty_n;
  assign in_40__m_axi_read_data_read = in_40_read_data__read;
  assign in_40__m_axi_rst = ~ ap_rst_n;
  assign in_40__m_axi_write_addr_din = in_40_write_addr__din;
  assign in_40_write_addr__full_n = in_40__m_axi_write_addr_full_n;
  assign in_40__m_axi_write_addr_write = in_40_write_addr__write;
  assign in_40__m_axi_write_data_din = in_40_write_data__din;
  assign in_40_write_data__full_n = in_40__m_axi_write_data_full_n;
  assign in_40__m_axi_write_data_write = in_40_write_data__write;
  assign in_40_write_resp__dout = in_40__m_axi_write_resp_dout;
  assign in_40_write_resp__empty_n = in_40__m_axi_write_resp_empty_n;
  assign in_40__m_axi_write_resp_read = in_40_write_resp__read;
  assign in_41__m_axi_clk = ap_clk;
  assign m_axi_in_41_ARADDR = in_41__m_axi_m_axi_ARADDR;
  assign m_axi_in_41_ARBURST = in_41__m_axi_m_axi_ARBURST;
  assign m_axi_in_41_ARCACHE = in_41__m_axi_m_axi_ARCACHE;
  assign m_axi_in_41_ARID = in_41__m_axi_m_axi_ARID;
  assign m_axi_in_41_ARLEN = in_41__m_axi_m_axi_ARLEN;
  assign m_axi_in_41_ARLOCK = in_41__m_axi_m_axi_ARLOCK;
  assign m_axi_in_41_ARPROT = in_41__m_axi_m_axi_ARPROT;
  assign m_axi_in_41_ARQOS = in_41__m_axi_m_axi_ARQOS;
  assign in_41__m_axi_m_axi_ARREADY = m_axi_in_41_ARREADY;
  assign m_axi_in_41_ARSIZE = in_41__m_axi_m_axi_ARSIZE;
  assign m_axi_in_41_ARVALID = in_41__m_axi_m_axi_ARVALID;
  assign m_axi_in_41_AWADDR = in_41__m_axi_m_axi_AWADDR;
  assign m_axi_in_41_AWBURST = in_41__m_axi_m_axi_AWBURST;
  assign m_axi_in_41_AWCACHE = in_41__m_axi_m_axi_AWCACHE;
  assign m_axi_in_41_AWID = in_41__m_axi_m_axi_AWID;
  assign m_axi_in_41_AWLEN = in_41__m_axi_m_axi_AWLEN;
  assign m_axi_in_41_AWLOCK = in_41__m_axi_m_axi_AWLOCK;
  assign m_axi_in_41_AWPROT = in_41__m_axi_m_axi_AWPROT;
  assign m_axi_in_41_AWQOS = in_41__m_axi_m_axi_AWQOS;
  assign in_41__m_axi_m_axi_AWREADY = m_axi_in_41_AWREADY;
  assign m_axi_in_41_AWSIZE = in_41__m_axi_m_axi_AWSIZE;
  assign m_axi_in_41_AWVALID = in_41__m_axi_m_axi_AWVALID;
  assign in_41__m_axi_m_axi_BID = m_axi_in_41_BID;
  assign m_axi_in_41_BREADY = in_41__m_axi_m_axi_BREADY;
  assign in_41__m_axi_m_axi_BRESP = m_axi_in_41_BRESP;
  assign in_41__m_axi_m_axi_BVALID = m_axi_in_41_BVALID;
  assign in_41__m_axi_m_axi_RDATA = m_axi_in_41_RDATA;
  assign in_41__m_axi_m_axi_RID = m_axi_in_41_RID;
  assign in_41__m_axi_m_axi_RLAST = m_axi_in_41_RLAST;
  assign m_axi_in_41_RREADY = in_41__m_axi_m_axi_RREADY;
  assign in_41__m_axi_m_axi_RRESP = m_axi_in_41_RRESP;
  assign in_41__m_axi_m_axi_RVALID = m_axi_in_41_RVALID;
  assign m_axi_in_41_WDATA = in_41__m_axi_m_axi_WDATA;
  assign m_axi_in_41_WLAST = in_41__m_axi_m_axi_WLAST;
  assign in_41__m_axi_m_axi_WREADY = m_axi_in_41_WREADY;
  assign m_axi_in_41_WSTRB = in_41__m_axi_m_axi_WSTRB;
  assign m_axi_in_41_WVALID = in_41__m_axi_m_axi_WVALID;
  assign in_41__m_axi_read_addr_din = in_41_read_addr__din;
  assign in_41_read_addr__full_n = in_41__m_axi_read_addr_full_n;
  assign in_41__m_axi_read_addr_write = in_41_read_addr__write;
  assign in_41_read_data__dout = in_41__m_axi_read_data_dout;
  assign in_41_read_data__empty_n = in_41__m_axi_read_data_empty_n;
  assign in_41__m_axi_read_data_read = in_41_read_data__read;
  assign in_41__m_axi_rst = ~ ap_rst_n;
  assign in_41__m_axi_write_addr_din = in_41_write_addr__din;
  assign in_41_write_addr__full_n = in_41__m_axi_write_addr_full_n;
  assign in_41__m_axi_write_addr_write = in_41_write_addr__write;
  assign in_41__m_axi_write_data_din = in_41_write_data__din;
  assign in_41_write_data__full_n = in_41__m_axi_write_data_full_n;
  assign in_41__m_axi_write_data_write = in_41_write_data__write;
  assign in_41_write_resp__dout = in_41__m_axi_write_resp_dout;
  assign in_41_write_resp__empty_n = in_41__m_axi_write_resp_empty_n;
  assign in_41__m_axi_write_resp_read = in_41_write_resp__read;
  assign in_42__m_axi_clk = ap_clk;
  assign m_axi_in_42_ARADDR = in_42__m_axi_m_axi_ARADDR;
  assign m_axi_in_42_ARBURST = in_42__m_axi_m_axi_ARBURST;
  assign m_axi_in_42_ARCACHE = in_42__m_axi_m_axi_ARCACHE;
  assign m_axi_in_42_ARID = in_42__m_axi_m_axi_ARID;
  assign m_axi_in_42_ARLEN = in_42__m_axi_m_axi_ARLEN;
  assign m_axi_in_42_ARLOCK = in_42__m_axi_m_axi_ARLOCK;
  assign m_axi_in_42_ARPROT = in_42__m_axi_m_axi_ARPROT;
  assign m_axi_in_42_ARQOS = in_42__m_axi_m_axi_ARQOS;
  assign in_42__m_axi_m_axi_ARREADY = m_axi_in_42_ARREADY;
  assign m_axi_in_42_ARSIZE = in_42__m_axi_m_axi_ARSIZE;
  assign m_axi_in_42_ARVALID = in_42__m_axi_m_axi_ARVALID;
  assign m_axi_in_42_AWADDR = in_42__m_axi_m_axi_AWADDR;
  assign m_axi_in_42_AWBURST = in_42__m_axi_m_axi_AWBURST;
  assign m_axi_in_42_AWCACHE = in_42__m_axi_m_axi_AWCACHE;
  assign m_axi_in_42_AWID = in_42__m_axi_m_axi_AWID;
  assign m_axi_in_42_AWLEN = in_42__m_axi_m_axi_AWLEN;
  assign m_axi_in_42_AWLOCK = in_42__m_axi_m_axi_AWLOCK;
  assign m_axi_in_42_AWPROT = in_42__m_axi_m_axi_AWPROT;
  assign m_axi_in_42_AWQOS = in_42__m_axi_m_axi_AWQOS;
  assign in_42__m_axi_m_axi_AWREADY = m_axi_in_42_AWREADY;
  assign m_axi_in_42_AWSIZE = in_42__m_axi_m_axi_AWSIZE;
  assign m_axi_in_42_AWVALID = in_42__m_axi_m_axi_AWVALID;
  assign in_42__m_axi_m_axi_BID = m_axi_in_42_BID;
  assign m_axi_in_42_BREADY = in_42__m_axi_m_axi_BREADY;
  assign in_42__m_axi_m_axi_BRESP = m_axi_in_42_BRESP;
  assign in_42__m_axi_m_axi_BVALID = m_axi_in_42_BVALID;
  assign in_42__m_axi_m_axi_RDATA = m_axi_in_42_RDATA;
  assign in_42__m_axi_m_axi_RID = m_axi_in_42_RID;
  assign in_42__m_axi_m_axi_RLAST = m_axi_in_42_RLAST;
  assign m_axi_in_42_RREADY = in_42__m_axi_m_axi_RREADY;
  assign in_42__m_axi_m_axi_RRESP = m_axi_in_42_RRESP;
  assign in_42__m_axi_m_axi_RVALID = m_axi_in_42_RVALID;
  assign m_axi_in_42_WDATA = in_42__m_axi_m_axi_WDATA;
  assign m_axi_in_42_WLAST = in_42__m_axi_m_axi_WLAST;
  assign in_42__m_axi_m_axi_WREADY = m_axi_in_42_WREADY;
  assign m_axi_in_42_WSTRB = in_42__m_axi_m_axi_WSTRB;
  assign m_axi_in_42_WVALID = in_42__m_axi_m_axi_WVALID;
  assign in_42__m_axi_read_addr_din = in_42_read_addr__din;
  assign in_42_read_addr__full_n = in_42__m_axi_read_addr_full_n;
  assign in_42__m_axi_read_addr_write = in_42_read_addr__write;
  assign in_42_read_data__dout = in_42__m_axi_read_data_dout;
  assign in_42_read_data__empty_n = in_42__m_axi_read_data_empty_n;
  assign in_42__m_axi_read_data_read = in_42_read_data__read;
  assign in_42__m_axi_rst = ~ ap_rst_n;
  assign in_42__m_axi_write_addr_din = in_42_write_addr__din;
  assign in_42_write_addr__full_n = in_42__m_axi_write_addr_full_n;
  assign in_42__m_axi_write_addr_write = in_42_write_addr__write;
  assign in_42__m_axi_write_data_din = in_42_write_data__din;
  assign in_42_write_data__full_n = in_42__m_axi_write_data_full_n;
  assign in_42__m_axi_write_data_write = in_42_write_data__write;
  assign in_42_write_resp__dout = in_42__m_axi_write_resp_dout;
  assign in_42_write_resp__empty_n = in_42__m_axi_write_resp_empty_n;
  assign in_42__m_axi_write_resp_read = in_42_write_resp__read;
  assign in_43__m_axi_clk = ap_clk;
  assign m_axi_in_43_ARADDR = in_43__m_axi_m_axi_ARADDR;
  assign m_axi_in_43_ARBURST = in_43__m_axi_m_axi_ARBURST;
  assign m_axi_in_43_ARCACHE = in_43__m_axi_m_axi_ARCACHE;
  assign m_axi_in_43_ARID = in_43__m_axi_m_axi_ARID;
  assign m_axi_in_43_ARLEN = in_43__m_axi_m_axi_ARLEN;
  assign m_axi_in_43_ARLOCK = in_43__m_axi_m_axi_ARLOCK;
  assign m_axi_in_43_ARPROT = in_43__m_axi_m_axi_ARPROT;
  assign m_axi_in_43_ARQOS = in_43__m_axi_m_axi_ARQOS;
  assign in_43__m_axi_m_axi_ARREADY = m_axi_in_43_ARREADY;
  assign m_axi_in_43_ARSIZE = in_43__m_axi_m_axi_ARSIZE;
  assign m_axi_in_43_ARVALID = in_43__m_axi_m_axi_ARVALID;
  assign m_axi_in_43_AWADDR = in_43__m_axi_m_axi_AWADDR;
  assign m_axi_in_43_AWBURST = in_43__m_axi_m_axi_AWBURST;
  assign m_axi_in_43_AWCACHE = in_43__m_axi_m_axi_AWCACHE;
  assign m_axi_in_43_AWID = in_43__m_axi_m_axi_AWID;
  assign m_axi_in_43_AWLEN = in_43__m_axi_m_axi_AWLEN;
  assign m_axi_in_43_AWLOCK = in_43__m_axi_m_axi_AWLOCK;
  assign m_axi_in_43_AWPROT = in_43__m_axi_m_axi_AWPROT;
  assign m_axi_in_43_AWQOS = in_43__m_axi_m_axi_AWQOS;
  assign in_43__m_axi_m_axi_AWREADY = m_axi_in_43_AWREADY;
  assign m_axi_in_43_AWSIZE = in_43__m_axi_m_axi_AWSIZE;
  assign m_axi_in_43_AWVALID = in_43__m_axi_m_axi_AWVALID;
  assign in_43__m_axi_m_axi_BID = m_axi_in_43_BID;
  assign m_axi_in_43_BREADY = in_43__m_axi_m_axi_BREADY;
  assign in_43__m_axi_m_axi_BRESP = m_axi_in_43_BRESP;
  assign in_43__m_axi_m_axi_BVALID = m_axi_in_43_BVALID;
  assign in_43__m_axi_m_axi_RDATA = m_axi_in_43_RDATA;
  assign in_43__m_axi_m_axi_RID = m_axi_in_43_RID;
  assign in_43__m_axi_m_axi_RLAST = m_axi_in_43_RLAST;
  assign m_axi_in_43_RREADY = in_43__m_axi_m_axi_RREADY;
  assign in_43__m_axi_m_axi_RRESP = m_axi_in_43_RRESP;
  assign in_43__m_axi_m_axi_RVALID = m_axi_in_43_RVALID;
  assign m_axi_in_43_WDATA = in_43__m_axi_m_axi_WDATA;
  assign m_axi_in_43_WLAST = in_43__m_axi_m_axi_WLAST;
  assign in_43__m_axi_m_axi_WREADY = m_axi_in_43_WREADY;
  assign m_axi_in_43_WSTRB = in_43__m_axi_m_axi_WSTRB;
  assign m_axi_in_43_WVALID = in_43__m_axi_m_axi_WVALID;
  assign in_43__m_axi_read_addr_din = in_43_read_addr__din;
  assign in_43_read_addr__full_n = in_43__m_axi_read_addr_full_n;
  assign in_43__m_axi_read_addr_write = in_43_read_addr__write;
  assign in_43_read_data__dout = in_43__m_axi_read_data_dout;
  assign in_43_read_data__empty_n = in_43__m_axi_read_data_empty_n;
  assign in_43__m_axi_read_data_read = in_43_read_data__read;
  assign in_43__m_axi_rst = ~ ap_rst_n;
  assign in_43__m_axi_write_addr_din = in_43_write_addr__din;
  assign in_43_write_addr__full_n = in_43__m_axi_write_addr_full_n;
  assign in_43__m_axi_write_addr_write = in_43_write_addr__write;
  assign in_43__m_axi_write_data_din = in_43_write_data__din;
  assign in_43_write_data__full_n = in_43__m_axi_write_data_full_n;
  assign in_43__m_axi_write_data_write = in_43_write_data__write;
  assign in_43_write_resp__dout = in_43__m_axi_write_resp_dout;
  assign in_43_write_resp__empty_n = in_43__m_axi_write_resp_empty_n;
  assign in_43__m_axi_write_resp_read = in_43_write_resp__read;
  assign in_44__m_axi_clk = ap_clk;
  assign m_axi_in_44_ARADDR = in_44__m_axi_m_axi_ARADDR;
  assign m_axi_in_44_ARBURST = in_44__m_axi_m_axi_ARBURST;
  assign m_axi_in_44_ARCACHE = in_44__m_axi_m_axi_ARCACHE;
  assign m_axi_in_44_ARID = in_44__m_axi_m_axi_ARID;
  assign m_axi_in_44_ARLEN = in_44__m_axi_m_axi_ARLEN;
  assign m_axi_in_44_ARLOCK = in_44__m_axi_m_axi_ARLOCK;
  assign m_axi_in_44_ARPROT = in_44__m_axi_m_axi_ARPROT;
  assign m_axi_in_44_ARQOS = in_44__m_axi_m_axi_ARQOS;
  assign in_44__m_axi_m_axi_ARREADY = m_axi_in_44_ARREADY;
  assign m_axi_in_44_ARSIZE = in_44__m_axi_m_axi_ARSIZE;
  assign m_axi_in_44_ARVALID = in_44__m_axi_m_axi_ARVALID;
  assign m_axi_in_44_AWADDR = in_44__m_axi_m_axi_AWADDR;
  assign m_axi_in_44_AWBURST = in_44__m_axi_m_axi_AWBURST;
  assign m_axi_in_44_AWCACHE = in_44__m_axi_m_axi_AWCACHE;
  assign m_axi_in_44_AWID = in_44__m_axi_m_axi_AWID;
  assign m_axi_in_44_AWLEN = in_44__m_axi_m_axi_AWLEN;
  assign m_axi_in_44_AWLOCK = in_44__m_axi_m_axi_AWLOCK;
  assign m_axi_in_44_AWPROT = in_44__m_axi_m_axi_AWPROT;
  assign m_axi_in_44_AWQOS = in_44__m_axi_m_axi_AWQOS;
  assign in_44__m_axi_m_axi_AWREADY = m_axi_in_44_AWREADY;
  assign m_axi_in_44_AWSIZE = in_44__m_axi_m_axi_AWSIZE;
  assign m_axi_in_44_AWVALID = in_44__m_axi_m_axi_AWVALID;
  assign in_44__m_axi_m_axi_BID = m_axi_in_44_BID;
  assign m_axi_in_44_BREADY = in_44__m_axi_m_axi_BREADY;
  assign in_44__m_axi_m_axi_BRESP = m_axi_in_44_BRESP;
  assign in_44__m_axi_m_axi_BVALID = m_axi_in_44_BVALID;
  assign in_44__m_axi_m_axi_RDATA = m_axi_in_44_RDATA;
  assign in_44__m_axi_m_axi_RID = m_axi_in_44_RID;
  assign in_44__m_axi_m_axi_RLAST = m_axi_in_44_RLAST;
  assign m_axi_in_44_RREADY = in_44__m_axi_m_axi_RREADY;
  assign in_44__m_axi_m_axi_RRESP = m_axi_in_44_RRESP;
  assign in_44__m_axi_m_axi_RVALID = m_axi_in_44_RVALID;
  assign m_axi_in_44_WDATA = in_44__m_axi_m_axi_WDATA;
  assign m_axi_in_44_WLAST = in_44__m_axi_m_axi_WLAST;
  assign in_44__m_axi_m_axi_WREADY = m_axi_in_44_WREADY;
  assign m_axi_in_44_WSTRB = in_44__m_axi_m_axi_WSTRB;
  assign m_axi_in_44_WVALID = in_44__m_axi_m_axi_WVALID;
  assign in_44__m_axi_read_addr_din = in_44_read_addr__din;
  assign in_44_read_addr__full_n = in_44__m_axi_read_addr_full_n;
  assign in_44__m_axi_read_addr_write = in_44_read_addr__write;
  assign in_44_read_data__dout = in_44__m_axi_read_data_dout;
  assign in_44_read_data__empty_n = in_44__m_axi_read_data_empty_n;
  assign in_44__m_axi_read_data_read = in_44_read_data__read;
  assign in_44__m_axi_rst = ~ ap_rst_n;
  assign in_44__m_axi_write_addr_din = in_44_write_addr__din;
  assign in_44_write_addr__full_n = in_44__m_axi_write_addr_full_n;
  assign in_44__m_axi_write_addr_write = in_44_write_addr__write;
  assign in_44__m_axi_write_data_din = in_44_write_data__din;
  assign in_44_write_data__full_n = in_44__m_axi_write_data_full_n;
  assign in_44__m_axi_write_data_write = in_44_write_data__write;
  assign in_44_write_resp__dout = in_44__m_axi_write_resp_dout;
  assign in_44_write_resp__empty_n = in_44__m_axi_write_resp_empty_n;
  assign in_44__m_axi_write_resp_read = in_44_write_resp__read;
  assign in_45__m_axi_clk = ap_clk;
  assign m_axi_in_45_ARADDR = in_45__m_axi_m_axi_ARADDR;
  assign m_axi_in_45_ARBURST = in_45__m_axi_m_axi_ARBURST;
  assign m_axi_in_45_ARCACHE = in_45__m_axi_m_axi_ARCACHE;
  assign m_axi_in_45_ARID = in_45__m_axi_m_axi_ARID;
  assign m_axi_in_45_ARLEN = in_45__m_axi_m_axi_ARLEN;
  assign m_axi_in_45_ARLOCK = in_45__m_axi_m_axi_ARLOCK;
  assign m_axi_in_45_ARPROT = in_45__m_axi_m_axi_ARPROT;
  assign m_axi_in_45_ARQOS = in_45__m_axi_m_axi_ARQOS;
  assign in_45__m_axi_m_axi_ARREADY = m_axi_in_45_ARREADY;
  assign m_axi_in_45_ARSIZE = in_45__m_axi_m_axi_ARSIZE;
  assign m_axi_in_45_ARVALID = in_45__m_axi_m_axi_ARVALID;
  assign m_axi_in_45_AWADDR = in_45__m_axi_m_axi_AWADDR;
  assign m_axi_in_45_AWBURST = in_45__m_axi_m_axi_AWBURST;
  assign m_axi_in_45_AWCACHE = in_45__m_axi_m_axi_AWCACHE;
  assign m_axi_in_45_AWID = in_45__m_axi_m_axi_AWID;
  assign m_axi_in_45_AWLEN = in_45__m_axi_m_axi_AWLEN;
  assign m_axi_in_45_AWLOCK = in_45__m_axi_m_axi_AWLOCK;
  assign m_axi_in_45_AWPROT = in_45__m_axi_m_axi_AWPROT;
  assign m_axi_in_45_AWQOS = in_45__m_axi_m_axi_AWQOS;
  assign in_45__m_axi_m_axi_AWREADY = m_axi_in_45_AWREADY;
  assign m_axi_in_45_AWSIZE = in_45__m_axi_m_axi_AWSIZE;
  assign m_axi_in_45_AWVALID = in_45__m_axi_m_axi_AWVALID;
  assign in_45__m_axi_m_axi_BID = m_axi_in_45_BID;
  assign m_axi_in_45_BREADY = in_45__m_axi_m_axi_BREADY;
  assign in_45__m_axi_m_axi_BRESP = m_axi_in_45_BRESP;
  assign in_45__m_axi_m_axi_BVALID = m_axi_in_45_BVALID;
  assign in_45__m_axi_m_axi_RDATA = m_axi_in_45_RDATA;
  assign in_45__m_axi_m_axi_RID = m_axi_in_45_RID;
  assign in_45__m_axi_m_axi_RLAST = m_axi_in_45_RLAST;
  assign m_axi_in_45_RREADY = in_45__m_axi_m_axi_RREADY;
  assign in_45__m_axi_m_axi_RRESP = m_axi_in_45_RRESP;
  assign in_45__m_axi_m_axi_RVALID = m_axi_in_45_RVALID;
  assign m_axi_in_45_WDATA = in_45__m_axi_m_axi_WDATA;
  assign m_axi_in_45_WLAST = in_45__m_axi_m_axi_WLAST;
  assign in_45__m_axi_m_axi_WREADY = m_axi_in_45_WREADY;
  assign m_axi_in_45_WSTRB = in_45__m_axi_m_axi_WSTRB;
  assign m_axi_in_45_WVALID = in_45__m_axi_m_axi_WVALID;
  assign in_45__m_axi_read_addr_din = in_45_read_addr__din;
  assign in_45_read_addr__full_n = in_45__m_axi_read_addr_full_n;
  assign in_45__m_axi_read_addr_write = in_45_read_addr__write;
  assign in_45_read_data__dout = in_45__m_axi_read_data_dout;
  assign in_45_read_data__empty_n = in_45__m_axi_read_data_empty_n;
  assign in_45__m_axi_read_data_read = in_45_read_data__read;
  assign in_45__m_axi_rst = ~ ap_rst_n;
  assign in_45__m_axi_write_addr_din = in_45_write_addr__din;
  assign in_45_write_addr__full_n = in_45__m_axi_write_addr_full_n;
  assign in_45__m_axi_write_addr_write = in_45_write_addr__write;
  assign in_45__m_axi_write_data_din = in_45_write_data__din;
  assign in_45_write_data__full_n = in_45__m_axi_write_data_full_n;
  assign in_45__m_axi_write_data_write = in_45_write_data__write;
  assign in_45_write_resp__dout = in_45__m_axi_write_resp_dout;
  assign in_45_write_resp__empty_n = in_45__m_axi_write_resp_empty_n;
  assign in_45__m_axi_write_resp_read = in_45_write_resp__read;
  assign in_46__m_axi_clk = ap_clk;
  assign m_axi_in_46_ARADDR = in_46__m_axi_m_axi_ARADDR;
  assign m_axi_in_46_ARBURST = in_46__m_axi_m_axi_ARBURST;
  assign m_axi_in_46_ARCACHE = in_46__m_axi_m_axi_ARCACHE;
  assign m_axi_in_46_ARID = in_46__m_axi_m_axi_ARID;
  assign m_axi_in_46_ARLEN = in_46__m_axi_m_axi_ARLEN;
  assign m_axi_in_46_ARLOCK = in_46__m_axi_m_axi_ARLOCK;
  assign m_axi_in_46_ARPROT = in_46__m_axi_m_axi_ARPROT;
  assign m_axi_in_46_ARQOS = in_46__m_axi_m_axi_ARQOS;
  assign in_46__m_axi_m_axi_ARREADY = m_axi_in_46_ARREADY;
  assign m_axi_in_46_ARSIZE = in_46__m_axi_m_axi_ARSIZE;
  assign m_axi_in_46_ARVALID = in_46__m_axi_m_axi_ARVALID;
  assign m_axi_in_46_AWADDR = in_46__m_axi_m_axi_AWADDR;
  assign m_axi_in_46_AWBURST = in_46__m_axi_m_axi_AWBURST;
  assign m_axi_in_46_AWCACHE = in_46__m_axi_m_axi_AWCACHE;
  assign m_axi_in_46_AWID = in_46__m_axi_m_axi_AWID;
  assign m_axi_in_46_AWLEN = in_46__m_axi_m_axi_AWLEN;
  assign m_axi_in_46_AWLOCK = in_46__m_axi_m_axi_AWLOCK;
  assign m_axi_in_46_AWPROT = in_46__m_axi_m_axi_AWPROT;
  assign m_axi_in_46_AWQOS = in_46__m_axi_m_axi_AWQOS;
  assign in_46__m_axi_m_axi_AWREADY = m_axi_in_46_AWREADY;
  assign m_axi_in_46_AWSIZE = in_46__m_axi_m_axi_AWSIZE;
  assign m_axi_in_46_AWVALID = in_46__m_axi_m_axi_AWVALID;
  assign in_46__m_axi_m_axi_BID = m_axi_in_46_BID;
  assign m_axi_in_46_BREADY = in_46__m_axi_m_axi_BREADY;
  assign in_46__m_axi_m_axi_BRESP = m_axi_in_46_BRESP;
  assign in_46__m_axi_m_axi_BVALID = m_axi_in_46_BVALID;
  assign in_46__m_axi_m_axi_RDATA = m_axi_in_46_RDATA;
  assign in_46__m_axi_m_axi_RID = m_axi_in_46_RID;
  assign in_46__m_axi_m_axi_RLAST = m_axi_in_46_RLAST;
  assign m_axi_in_46_RREADY = in_46__m_axi_m_axi_RREADY;
  assign in_46__m_axi_m_axi_RRESP = m_axi_in_46_RRESP;
  assign in_46__m_axi_m_axi_RVALID = m_axi_in_46_RVALID;
  assign m_axi_in_46_WDATA = in_46__m_axi_m_axi_WDATA;
  assign m_axi_in_46_WLAST = in_46__m_axi_m_axi_WLAST;
  assign in_46__m_axi_m_axi_WREADY = m_axi_in_46_WREADY;
  assign m_axi_in_46_WSTRB = in_46__m_axi_m_axi_WSTRB;
  assign m_axi_in_46_WVALID = in_46__m_axi_m_axi_WVALID;
  assign in_46__m_axi_read_addr_din = in_46_read_addr__din;
  assign in_46_read_addr__full_n = in_46__m_axi_read_addr_full_n;
  assign in_46__m_axi_read_addr_write = in_46_read_addr__write;
  assign in_46_read_data__dout = in_46__m_axi_read_data_dout;
  assign in_46_read_data__empty_n = in_46__m_axi_read_data_empty_n;
  assign in_46__m_axi_read_data_read = in_46_read_data__read;
  assign in_46__m_axi_rst = ~ ap_rst_n;
  assign in_46__m_axi_write_addr_din = in_46_write_addr__din;
  assign in_46_write_addr__full_n = in_46__m_axi_write_addr_full_n;
  assign in_46__m_axi_write_addr_write = in_46_write_addr__write;
  assign in_46__m_axi_write_data_din = in_46_write_data__din;
  assign in_46_write_data__full_n = in_46__m_axi_write_data_full_n;
  assign in_46__m_axi_write_data_write = in_46_write_data__write;
  assign in_46_write_resp__dout = in_46__m_axi_write_resp_dout;
  assign in_46_write_resp__empty_n = in_46__m_axi_write_resp_empty_n;
  assign in_46__m_axi_write_resp_read = in_46_write_resp__read;
  assign in_47__m_axi_clk = ap_clk;
  assign m_axi_in_47_ARADDR = in_47__m_axi_m_axi_ARADDR;
  assign m_axi_in_47_ARBURST = in_47__m_axi_m_axi_ARBURST;
  assign m_axi_in_47_ARCACHE = in_47__m_axi_m_axi_ARCACHE;
  assign m_axi_in_47_ARID = in_47__m_axi_m_axi_ARID;
  assign m_axi_in_47_ARLEN = in_47__m_axi_m_axi_ARLEN;
  assign m_axi_in_47_ARLOCK = in_47__m_axi_m_axi_ARLOCK;
  assign m_axi_in_47_ARPROT = in_47__m_axi_m_axi_ARPROT;
  assign m_axi_in_47_ARQOS = in_47__m_axi_m_axi_ARQOS;
  assign in_47__m_axi_m_axi_ARREADY = m_axi_in_47_ARREADY;
  assign m_axi_in_47_ARSIZE = in_47__m_axi_m_axi_ARSIZE;
  assign m_axi_in_47_ARVALID = in_47__m_axi_m_axi_ARVALID;
  assign m_axi_in_47_AWADDR = in_47__m_axi_m_axi_AWADDR;
  assign m_axi_in_47_AWBURST = in_47__m_axi_m_axi_AWBURST;
  assign m_axi_in_47_AWCACHE = in_47__m_axi_m_axi_AWCACHE;
  assign m_axi_in_47_AWID = in_47__m_axi_m_axi_AWID;
  assign m_axi_in_47_AWLEN = in_47__m_axi_m_axi_AWLEN;
  assign m_axi_in_47_AWLOCK = in_47__m_axi_m_axi_AWLOCK;
  assign m_axi_in_47_AWPROT = in_47__m_axi_m_axi_AWPROT;
  assign m_axi_in_47_AWQOS = in_47__m_axi_m_axi_AWQOS;
  assign in_47__m_axi_m_axi_AWREADY = m_axi_in_47_AWREADY;
  assign m_axi_in_47_AWSIZE = in_47__m_axi_m_axi_AWSIZE;
  assign m_axi_in_47_AWVALID = in_47__m_axi_m_axi_AWVALID;
  assign in_47__m_axi_m_axi_BID = m_axi_in_47_BID;
  assign m_axi_in_47_BREADY = in_47__m_axi_m_axi_BREADY;
  assign in_47__m_axi_m_axi_BRESP = m_axi_in_47_BRESP;
  assign in_47__m_axi_m_axi_BVALID = m_axi_in_47_BVALID;
  assign in_47__m_axi_m_axi_RDATA = m_axi_in_47_RDATA;
  assign in_47__m_axi_m_axi_RID = m_axi_in_47_RID;
  assign in_47__m_axi_m_axi_RLAST = m_axi_in_47_RLAST;
  assign m_axi_in_47_RREADY = in_47__m_axi_m_axi_RREADY;
  assign in_47__m_axi_m_axi_RRESP = m_axi_in_47_RRESP;
  assign in_47__m_axi_m_axi_RVALID = m_axi_in_47_RVALID;
  assign m_axi_in_47_WDATA = in_47__m_axi_m_axi_WDATA;
  assign m_axi_in_47_WLAST = in_47__m_axi_m_axi_WLAST;
  assign in_47__m_axi_m_axi_WREADY = m_axi_in_47_WREADY;
  assign m_axi_in_47_WSTRB = in_47__m_axi_m_axi_WSTRB;
  assign m_axi_in_47_WVALID = in_47__m_axi_m_axi_WVALID;
  assign in_47__m_axi_read_addr_din = in_47_read_addr__din;
  assign in_47_read_addr__full_n = in_47__m_axi_read_addr_full_n;
  assign in_47__m_axi_read_addr_write = in_47_read_addr__write;
  assign in_47_read_data__dout = in_47__m_axi_read_data_dout;
  assign in_47_read_data__empty_n = in_47__m_axi_read_data_empty_n;
  assign in_47__m_axi_read_data_read = in_47_read_data__read;
  assign in_47__m_axi_rst = ~ ap_rst_n;
  assign in_47__m_axi_write_addr_din = in_47_write_addr__din;
  assign in_47_write_addr__full_n = in_47__m_axi_write_addr_full_n;
  assign in_47__m_axi_write_addr_write = in_47_write_addr__write;
  assign in_47__m_axi_write_data_din = in_47_write_data__din;
  assign in_47_write_data__full_n = in_47__m_axi_write_data_full_n;
  assign in_47__m_axi_write_data_write = in_47_write_data__write;
  assign in_47_write_resp__dout = in_47__m_axi_write_resp_dout;
  assign in_47_write_resp__empty_n = in_47__m_axi_write_resp_empty_n;
  assign in_47__m_axi_write_resp_read = in_47_write_resp__read;
  assign in_48__m_axi_clk = ap_clk;
  assign m_axi_in_48_ARADDR = in_48__m_axi_m_axi_ARADDR;
  assign m_axi_in_48_ARBURST = in_48__m_axi_m_axi_ARBURST;
  assign m_axi_in_48_ARCACHE = in_48__m_axi_m_axi_ARCACHE;
  assign m_axi_in_48_ARID = in_48__m_axi_m_axi_ARID;
  assign m_axi_in_48_ARLEN = in_48__m_axi_m_axi_ARLEN;
  assign m_axi_in_48_ARLOCK = in_48__m_axi_m_axi_ARLOCK;
  assign m_axi_in_48_ARPROT = in_48__m_axi_m_axi_ARPROT;
  assign m_axi_in_48_ARQOS = in_48__m_axi_m_axi_ARQOS;
  assign in_48__m_axi_m_axi_ARREADY = m_axi_in_48_ARREADY;
  assign m_axi_in_48_ARSIZE = in_48__m_axi_m_axi_ARSIZE;
  assign m_axi_in_48_ARVALID = in_48__m_axi_m_axi_ARVALID;
  assign m_axi_in_48_AWADDR = in_48__m_axi_m_axi_AWADDR;
  assign m_axi_in_48_AWBURST = in_48__m_axi_m_axi_AWBURST;
  assign m_axi_in_48_AWCACHE = in_48__m_axi_m_axi_AWCACHE;
  assign m_axi_in_48_AWID = in_48__m_axi_m_axi_AWID;
  assign m_axi_in_48_AWLEN = in_48__m_axi_m_axi_AWLEN;
  assign m_axi_in_48_AWLOCK = in_48__m_axi_m_axi_AWLOCK;
  assign m_axi_in_48_AWPROT = in_48__m_axi_m_axi_AWPROT;
  assign m_axi_in_48_AWQOS = in_48__m_axi_m_axi_AWQOS;
  assign in_48__m_axi_m_axi_AWREADY = m_axi_in_48_AWREADY;
  assign m_axi_in_48_AWSIZE = in_48__m_axi_m_axi_AWSIZE;
  assign m_axi_in_48_AWVALID = in_48__m_axi_m_axi_AWVALID;
  assign in_48__m_axi_m_axi_BID = m_axi_in_48_BID;
  assign m_axi_in_48_BREADY = in_48__m_axi_m_axi_BREADY;
  assign in_48__m_axi_m_axi_BRESP = m_axi_in_48_BRESP;
  assign in_48__m_axi_m_axi_BVALID = m_axi_in_48_BVALID;
  assign in_48__m_axi_m_axi_RDATA = m_axi_in_48_RDATA;
  assign in_48__m_axi_m_axi_RID = m_axi_in_48_RID;
  assign in_48__m_axi_m_axi_RLAST = m_axi_in_48_RLAST;
  assign m_axi_in_48_RREADY = in_48__m_axi_m_axi_RREADY;
  assign in_48__m_axi_m_axi_RRESP = m_axi_in_48_RRESP;
  assign in_48__m_axi_m_axi_RVALID = m_axi_in_48_RVALID;
  assign m_axi_in_48_WDATA = in_48__m_axi_m_axi_WDATA;
  assign m_axi_in_48_WLAST = in_48__m_axi_m_axi_WLAST;
  assign in_48__m_axi_m_axi_WREADY = m_axi_in_48_WREADY;
  assign m_axi_in_48_WSTRB = in_48__m_axi_m_axi_WSTRB;
  assign m_axi_in_48_WVALID = in_48__m_axi_m_axi_WVALID;
  assign in_48__m_axi_read_addr_din = in_48_read_addr__din;
  assign in_48_read_addr__full_n = in_48__m_axi_read_addr_full_n;
  assign in_48__m_axi_read_addr_write = in_48_read_addr__write;
  assign in_48_read_data__dout = in_48__m_axi_read_data_dout;
  assign in_48_read_data__empty_n = in_48__m_axi_read_data_empty_n;
  assign in_48__m_axi_read_data_read = in_48_read_data__read;
  assign in_48__m_axi_rst = ~ ap_rst_n;
  assign in_48__m_axi_write_addr_din = in_48_write_addr__din;
  assign in_48_write_addr__full_n = in_48__m_axi_write_addr_full_n;
  assign in_48__m_axi_write_addr_write = in_48_write_addr__write;
  assign in_48__m_axi_write_data_din = in_48_write_data__din;
  assign in_48_write_data__full_n = in_48__m_axi_write_data_full_n;
  assign in_48__m_axi_write_data_write = in_48_write_data__write;
  assign in_48_write_resp__dout = in_48__m_axi_write_resp_dout;
  assign in_48_write_resp__empty_n = in_48__m_axi_write_resp_empty_n;
  assign in_48__m_axi_write_resp_read = in_48_write_resp__read;
  assign in_49__m_axi_clk = ap_clk;
  assign m_axi_in_49_ARADDR = in_49__m_axi_m_axi_ARADDR;
  assign m_axi_in_49_ARBURST = in_49__m_axi_m_axi_ARBURST;
  assign m_axi_in_49_ARCACHE = in_49__m_axi_m_axi_ARCACHE;
  assign m_axi_in_49_ARID = in_49__m_axi_m_axi_ARID;
  assign m_axi_in_49_ARLEN = in_49__m_axi_m_axi_ARLEN;
  assign m_axi_in_49_ARLOCK = in_49__m_axi_m_axi_ARLOCK;
  assign m_axi_in_49_ARPROT = in_49__m_axi_m_axi_ARPROT;
  assign m_axi_in_49_ARQOS = in_49__m_axi_m_axi_ARQOS;
  assign in_49__m_axi_m_axi_ARREADY = m_axi_in_49_ARREADY;
  assign m_axi_in_49_ARSIZE = in_49__m_axi_m_axi_ARSIZE;
  assign m_axi_in_49_ARVALID = in_49__m_axi_m_axi_ARVALID;
  assign m_axi_in_49_AWADDR = in_49__m_axi_m_axi_AWADDR;
  assign m_axi_in_49_AWBURST = in_49__m_axi_m_axi_AWBURST;
  assign m_axi_in_49_AWCACHE = in_49__m_axi_m_axi_AWCACHE;
  assign m_axi_in_49_AWID = in_49__m_axi_m_axi_AWID;
  assign m_axi_in_49_AWLEN = in_49__m_axi_m_axi_AWLEN;
  assign m_axi_in_49_AWLOCK = in_49__m_axi_m_axi_AWLOCK;
  assign m_axi_in_49_AWPROT = in_49__m_axi_m_axi_AWPROT;
  assign m_axi_in_49_AWQOS = in_49__m_axi_m_axi_AWQOS;
  assign in_49__m_axi_m_axi_AWREADY = m_axi_in_49_AWREADY;
  assign m_axi_in_49_AWSIZE = in_49__m_axi_m_axi_AWSIZE;
  assign m_axi_in_49_AWVALID = in_49__m_axi_m_axi_AWVALID;
  assign in_49__m_axi_m_axi_BID = m_axi_in_49_BID;
  assign m_axi_in_49_BREADY = in_49__m_axi_m_axi_BREADY;
  assign in_49__m_axi_m_axi_BRESP = m_axi_in_49_BRESP;
  assign in_49__m_axi_m_axi_BVALID = m_axi_in_49_BVALID;
  assign in_49__m_axi_m_axi_RDATA = m_axi_in_49_RDATA;
  assign in_49__m_axi_m_axi_RID = m_axi_in_49_RID;
  assign in_49__m_axi_m_axi_RLAST = m_axi_in_49_RLAST;
  assign m_axi_in_49_RREADY = in_49__m_axi_m_axi_RREADY;
  assign in_49__m_axi_m_axi_RRESP = m_axi_in_49_RRESP;
  assign in_49__m_axi_m_axi_RVALID = m_axi_in_49_RVALID;
  assign m_axi_in_49_WDATA = in_49__m_axi_m_axi_WDATA;
  assign m_axi_in_49_WLAST = in_49__m_axi_m_axi_WLAST;
  assign in_49__m_axi_m_axi_WREADY = m_axi_in_49_WREADY;
  assign m_axi_in_49_WSTRB = in_49__m_axi_m_axi_WSTRB;
  assign m_axi_in_49_WVALID = in_49__m_axi_m_axi_WVALID;
  assign in_49__m_axi_read_addr_din = in_49_read_addr__din;
  assign in_49_read_addr__full_n = in_49__m_axi_read_addr_full_n;
  assign in_49__m_axi_read_addr_write = in_49_read_addr__write;
  assign in_49_read_data__dout = in_49__m_axi_read_data_dout;
  assign in_49_read_data__empty_n = in_49__m_axi_read_data_empty_n;
  assign in_49__m_axi_read_data_read = in_49_read_data__read;
  assign in_49__m_axi_rst = ~ ap_rst_n;
  assign in_49__m_axi_write_addr_din = in_49_write_addr__din;
  assign in_49_write_addr__full_n = in_49__m_axi_write_addr_full_n;
  assign in_49__m_axi_write_addr_write = in_49_write_addr__write;
  assign in_49__m_axi_write_data_din = in_49_write_data__din;
  assign in_49_write_data__full_n = in_49__m_axi_write_data_full_n;
  assign in_49__m_axi_write_data_write = in_49_write_data__write;
  assign in_49_write_resp__dout = in_49__m_axi_write_resp_dout;
  assign in_49_write_resp__empty_n = in_49__m_axi_write_resp_empty_n;
  assign in_49__m_axi_write_resp_read = in_49_write_resp__read;
  assign in_5__m_axi_clk = ap_clk;
  assign m_axi_in_5_ARADDR = in_5__m_axi_m_axi_ARADDR;
  assign m_axi_in_5_ARBURST = in_5__m_axi_m_axi_ARBURST;
  assign m_axi_in_5_ARCACHE = in_5__m_axi_m_axi_ARCACHE;
  assign m_axi_in_5_ARID = in_5__m_axi_m_axi_ARID;
  assign m_axi_in_5_ARLEN = in_5__m_axi_m_axi_ARLEN;
  assign m_axi_in_5_ARLOCK = in_5__m_axi_m_axi_ARLOCK;
  assign m_axi_in_5_ARPROT = in_5__m_axi_m_axi_ARPROT;
  assign m_axi_in_5_ARQOS = in_5__m_axi_m_axi_ARQOS;
  assign in_5__m_axi_m_axi_ARREADY = m_axi_in_5_ARREADY;
  assign m_axi_in_5_ARSIZE = in_5__m_axi_m_axi_ARSIZE;
  assign m_axi_in_5_ARVALID = in_5__m_axi_m_axi_ARVALID;
  assign m_axi_in_5_AWADDR = in_5__m_axi_m_axi_AWADDR;
  assign m_axi_in_5_AWBURST = in_5__m_axi_m_axi_AWBURST;
  assign m_axi_in_5_AWCACHE = in_5__m_axi_m_axi_AWCACHE;
  assign m_axi_in_5_AWID = in_5__m_axi_m_axi_AWID;
  assign m_axi_in_5_AWLEN = in_5__m_axi_m_axi_AWLEN;
  assign m_axi_in_5_AWLOCK = in_5__m_axi_m_axi_AWLOCK;
  assign m_axi_in_5_AWPROT = in_5__m_axi_m_axi_AWPROT;
  assign m_axi_in_5_AWQOS = in_5__m_axi_m_axi_AWQOS;
  assign in_5__m_axi_m_axi_AWREADY = m_axi_in_5_AWREADY;
  assign m_axi_in_5_AWSIZE = in_5__m_axi_m_axi_AWSIZE;
  assign m_axi_in_5_AWVALID = in_5__m_axi_m_axi_AWVALID;
  assign in_5__m_axi_m_axi_BID = m_axi_in_5_BID;
  assign m_axi_in_5_BREADY = in_5__m_axi_m_axi_BREADY;
  assign in_5__m_axi_m_axi_BRESP = m_axi_in_5_BRESP;
  assign in_5__m_axi_m_axi_BVALID = m_axi_in_5_BVALID;
  assign in_5__m_axi_m_axi_RDATA = m_axi_in_5_RDATA;
  assign in_5__m_axi_m_axi_RID = m_axi_in_5_RID;
  assign in_5__m_axi_m_axi_RLAST = m_axi_in_5_RLAST;
  assign m_axi_in_5_RREADY = in_5__m_axi_m_axi_RREADY;
  assign in_5__m_axi_m_axi_RRESP = m_axi_in_5_RRESP;
  assign in_5__m_axi_m_axi_RVALID = m_axi_in_5_RVALID;
  assign m_axi_in_5_WDATA = in_5__m_axi_m_axi_WDATA;
  assign m_axi_in_5_WLAST = in_5__m_axi_m_axi_WLAST;
  assign in_5__m_axi_m_axi_WREADY = m_axi_in_5_WREADY;
  assign m_axi_in_5_WSTRB = in_5__m_axi_m_axi_WSTRB;
  assign m_axi_in_5_WVALID = in_5__m_axi_m_axi_WVALID;
  assign in_5__m_axi_read_addr_din = in_5_read_addr__din;
  assign in_5_read_addr__full_n = in_5__m_axi_read_addr_full_n;
  assign in_5__m_axi_read_addr_write = in_5_read_addr__write;
  assign in_5_read_data__dout = in_5__m_axi_read_data_dout;
  assign in_5_read_data__empty_n = in_5__m_axi_read_data_empty_n;
  assign in_5__m_axi_read_data_read = in_5_read_data__read;
  assign in_5__m_axi_rst = ~ ap_rst_n;
  assign in_5__m_axi_write_addr_din = in_5_write_addr__din;
  assign in_5_write_addr__full_n = in_5__m_axi_write_addr_full_n;
  assign in_5__m_axi_write_addr_write = in_5_write_addr__write;
  assign in_5__m_axi_write_data_din = in_5_write_data__din;
  assign in_5_write_data__full_n = in_5__m_axi_write_data_full_n;
  assign in_5__m_axi_write_data_write = in_5_write_data__write;
  assign in_5_write_resp__dout = in_5__m_axi_write_resp_dout;
  assign in_5_write_resp__empty_n = in_5__m_axi_write_resp_empty_n;
  assign in_5__m_axi_write_resp_read = in_5_write_resp__read;
  assign in_50__m_axi_clk = ap_clk;
  assign m_axi_in_50_ARADDR = in_50__m_axi_m_axi_ARADDR;
  assign m_axi_in_50_ARBURST = in_50__m_axi_m_axi_ARBURST;
  assign m_axi_in_50_ARCACHE = in_50__m_axi_m_axi_ARCACHE;
  assign m_axi_in_50_ARID = in_50__m_axi_m_axi_ARID;
  assign m_axi_in_50_ARLEN = in_50__m_axi_m_axi_ARLEN;
  assign m_axi_in_50_ARLOCK = in_50__m_axi_m_axi_ARLOCK;
  assign m_axi_in_50_ARPROT = in_50__m_axi_m_axi_ARPROT;
  assign m_axi_in_50_ARQOS = in_50__m_axi_m_axi_ARQOS;
  assign in_50__m_axi_m_axi_ARREADY = m_axi_in_50_ARREADY;
  assign m_axi_in_50_ARSIZE = in_50__m_axi_m_axi_ARSIZE;
  assign m_axi_in_50_ARVALID = in_50__m_axi_m_axi_ARVALID;
  assign m_axi_in_50_AWADDR = in_50__m_axi_m_axi_AWADDR;
  assign m_axi_in_50_AWBURST = in_50__m_axi_m_axi_AWBURST;
  assign m_axi_in_50_AWCACHE = in_50__m_axi_m_axi_AWCACHE;
  assign m_axi_in_50_AWID = in_50__m_axi_m_axi_AWID;
  assign m_axi_in_50_AWLEN = in_50__m_axi_m_axi_AWLEN;
  assign m_axi_in_50_AWLOCK = in_50__m_axi_m_axi_AWLOCK;
  assign m_axi_in_50_AWPROT = in_50__m_axi_m_axi_AWPROT;
  assign m_axi_in_50_AWQOS = in_50__m_axi_m_axi_AWQOS;
  assign in_50__m_axi_m_axi_AWREADY = m_axi_in_50_AWREADY;
  assign m_axi_in_50_AWSIZE = in_50__m_axi_m_axi_AWSIZE;
  assign m_axi_in_50_AWVALID = in_50__m_axi_m_axi_AWVALID;
  assign in_50__m_axi_m_axi_BID = m_axi_in_50_BID;
  assign m_axi_in_50_BREADY = in_50__m_axi_m_axi_BREADY;
  assign in_50__m_axi_m_axi_BRESP = m_axi_in_50_BRESP;
  assign in_50__m_axi_m_axi_BVALID = m_axi_in_50_BVALID;
  assign in_50__m_axi_m_axi_RDATA = m_axi_in_50_RDATA;
  assign in_50__m_axi_m_axi_RID = m_axi_in_50_RID;
  assign in_50__m_axi_m_axi_RLAST = m_axi_in_50_RLAST;
  assign m_axi_in_50_RREADY = in_50__m_axi_m_axi_RREADY;
  assign in_50__m_axi_m_axi_RRESP = m_axi_in_50_RRESP;
  assign in_50__m_axi_m_axi_RVALID = m_axi_in_50_RVALID;
  assign m_axi_in_50_WDATA = in_50__m_axi_m_axi_WDATA;
  assign m_axi_in_50_WLAST = in_50__m_axi_m_axi_WLAST;
  assign in_50__m_axi_m_axi_WREADY = m_axi_in_50_WREADY;
  assign m_axi_in_50_WSTRB = in_50__m_axi_m_axi_WSTRB;
  assign m_axi_in_50_WVALID = in_50__m_axi_m_axi_WVALID;
  assign in_50__m_axi_read_addr_din = in_50_read_addr__din;
  assign in_50_read_addr__full_n = in_50__m_axi_read_addr_full_n;
  assign in_50__m_axi_read_addr_write = in_50_read_addr__write;
  assign in_50_read_data__dout = in_50__m_axi_read_data_dout;
  assign in_50_read_data__empty_n = in_50__m_axi_read_data_empty_n;
  assign in_50__m_axi_read_data_read = in_50_read_data__read;
  assign in_50__m_axi_rst = ~ ap_rst_n;
  assign in_50__m_axi_write_addr_din = in_50_write_addr__din;
  assign in_50_write_addr__full_n = in_50__m_axi_write_addr_full_n;
  assign in_50__m_axi_write_addr_write = in_50_write_addr__write;
  assign in_50__m_axi_write_data_din = in_50_write_data__din;
  assign in_50_write_data__full_n = in_50__m_axi_write_data_full_n;
  assign in_50__m_axi_write_data_write = in_50_write_data__write;
  assign in_50_write_resp__dout = in_50__m_axi_write_resp_dout;
  assign in_50_write_resp__empty_n = in_50__m_axi_write_resp_empty_n;
  assign in_50__m_axi_write_resp_read = in_50_write_resp__read;
  assign in_51__m_axi_clk = ap_clk;
  assign m_axi_in_51_ARADDR = in_51__m_axi_m_axi_ARADDR;
  assign m_axi_in_51_ARBURST = in_51__m_axi_m_axi_ARBURST;
  assign m_axi_in_51_ARCACHE = in_51__m_axi_m_axi_ARCACHE;
  assign m_axi_in_51_ARID = in_51__m_axi_m_axi_ARID;
  assign m_axi_in_51_ARLEN = in_51__m_axi_m_axi_ARLEN;
  assign m_axi_in_51_ARLOCK = in_51__m_axi_m_axi_ARLOCK;
  assign m_axi_in_51_ARPROT = in_51__m_axi_m_axi_ARPROT;
  assign m_axi_in_51_ARQOS = in_51__m_axi_m_axi_ARQOS;
  assign in_51__m_axi_m_axi_ARREADY = m_axi_in_51_ARREADY;
  assign m_axi_in_51_ARSIZE = in_51__m_axi_m_axi_ARSIZE;
  assign m_axi_in_51_ARVALID = in_51__m_axi_m_axi_ARVALID;
  assign m_axi_in_51_AWADDR = in_51__m_axi_m_axi_AWADDR;
  assign m_axi_in_51_AWBURST = in_51__m_axi_m_axi_AWBURST;
  assign m_axi_in_51_AWCACHE = in_51__m_axi_m_axi_AWCACHE;
  assign m_axi_in_51_AWID = in_51__m_axi_m_axi_AWID;
  assign m_axi_in_51_AWLEN = in_51__m_axi_m_axi_AWLEN;
  assign m_axi_in_51_AWLOCK = in_51__m_axi_m_axi_AWLOCK;
  assign m_axi_in_51_AWPROT = in_51__m_axi_m_axi_AWPROT;
  assign m_axi_in_51_AWQOS = in_51__m_axi_m_axi_AWQOS;
  assign in_51__m_axi_m_axi_AWREADY = m_axi_in_51_AWREADY;
  assign m_axi_in_51_AWSIZE = in_51__m_axi_m_axi_AWSIZE;
  assign m_axi_in_51_AWVALID = in_51__m_axi_m_axi_AWVALID;
  assign in_51__m_axi_m_axi_BID = m_axi_in_51_BID;
  assign m_axi_in_51_BREADY = in_51__m_axi_m_axi_BREADY;
  assign in_51__m_axi_m_axi_BRESP = m_axi_in_51_BRESP;
  assign in_51__m_axi_m_axi_BVALID = m_axi_in_51_BVALID;
  assign in_51__m_axi_m_axi_RDATA = m_axi_in_51_RDATA;
  assign in_51__m_axi_m_axi_RID = m_axi_in_51_RID;
  assign in_51__m_axi_m_axi_RLAST = m_axi_in_51_RLAST;
  assign m_axi_in_51_RREADY = in_51__m_axi_m_axi_RREADY;
  assign in_51__m_axi_m_axi_RRESP = m_axi_in_51_RRESP;
  assign in_51__m_axi_m_axi_RVALID = m_axi_in_51_RVALID;
  assign m_axi_in_51_WDATA = in_51__m_axi_m_axi_WDATA;
  assign m_axi_in_51_WLAST = in_51__m_axi_m_axi_WLAST;
  assign in_51__m_axi_m_axi_WREADY = m_axi_in_51_WREADY;
  assign m_axi_in_51_WSTRB = in_51__m_axi_m_axi_WSTRB;
  assign m_axi_in_51_WVALID = in_51__m_axi_m_axi_WVALID;
  assign in_51__m_axi_read_addr_din = in_51_read_addr__din;
  assign in_51_read_addr__full_n = in_51__m_axi_read_addr_full_n;
  assign in_51__m_axi_read_addr_write = in_51_read_addr__write;
  assign in_51_read_data__dout = in_51__m_axi_read_data_dout;
  assign in_51_read_data__empty_n = in_51__m_axi_read_data_empty_n;
  assign in_51__m_axi_read_data_read = in_51_read_data__read;
  assign in_51__m_axi_rst = ~ ap_rst_n;
  assign in_51__m_axi_write_addr_din = in_51_write_addr__din;
  assign in_51_write_addr__full_n = in_51__m_axi_write_addr_full_n;
  assign in_51__m_axi_write_addr_write = in_51_write_addr__write;
  assign in_51__m_axi_write_data_din = in_51_write_data__din;
  assign in_51_write_data__full_n = in_51__m_axi_write_data_full_n;
  assign in_51__m_axi_write_data_write = in_51_write_data__write;
  assign in_51_write_resp__dout = in_51__m_axi_write_resp_dout;
  assign in_51_write_resp__empty_n = in_51__m_axi_write_resp_empty_n;
  assign in_51__m_axi_write_resp_read = in_51_write_resp__read;
  assign in_52__m_axi_clk = ap_clk;
  assign m_axi_in_52_ARADDR = in_52__m_axi_m_axi_ARADDR;
  assign m_axi_in_52_ARBURST = in_52__m_axi_m_axi_ARBURST;
  assign m_axi_in_52_ARCACHE = in_52__m_axi_m_axi_ARCACHE;
  assign m_axi_in_52_ARID = in_52__m_axi_m_axi_ARID;
  assign m_axi_in_52_ARLEN = in_52__m_axi_m_axi_ARLEN;
  assign m_axi_in_52_ARLOCK = in_52__m_axi_m_axi_ARLOCK;
  assign m_axi_in_52_ARPROT = in_52__m_axi_m_axi_ARPROT;
  assign m_axi_in_52_ARQOS = in_52__m_axi_m_axi_ARQOS;
  assign in_52__m_axi_m_axi_ARREADY = m_axi_in_52_ARREADY;
  assign m_axi_in_52_ARSIZE = in_52__m_axi_m_axi_ARSIZE;
  assign m_axi_in_52_ARVALID = in_52__m_axi_m_axi_ARVALID;
  assign m_axi_in_52_AWADDR = in_52__m_axi_m_axi_AWADDR;
  assign m_axi_in_52_AWBURST = in_52__m_axi_m_axi_AWBURST;
  assign m_axi_in_52_AWCACHE = in_52__m_axi_m_axi_AWCACHE;
  assign m_axi_in_52_AWID = in_52__m_axi_m_axi_AWID;
  assign m_axi_in_52_AWLEN = in_52__m_axi_m_axi_AWLEN;
  assign m_axi_in_52_AWLOCK = in_52__m_axi_m_axi_AWLOCK;
  assign m_axi_in_52_AWPROT = in_52__m_axi_m_axi_AWPROT;
  assign m_axi_in_52_AWQOS = in_52__m_axi_m_axi_AWQOS;
  assign in_52__m_axi_m_axi_AWREADY = m_axi_in_52_AWREADY;
  assign m_axi_in_52_AWSIZE = in_52__m_axi_m_axi_AWSIZE;
  assign m_axi_in_52_AWVALID = in_52__m_axi_m_axi_AWVALID;
  assign in_52__m_axi_m_axi_BID = m_axi_in_52_BID;
  assign m_axi_in_52_BREADY = in_52__m_axi_m_axi_BREADY;
  assign in_52__m_axi_m_axi_BRESP = m_axi_in_52_BRESP;
  assign in_52__m_axi_m_axi_BVALID = m_axi_in_52_BVALID;
  assign in_52__m_axi_m_axi_RDATA = m_axi_in_52_RDATA;
  assign in_52__m_axi_m_axi_RID = m_axi_in_52_RID;
  assign in_52__m_axi_m_axi_RLAST = m_axi_in_52_RLAST;
  assign m_axi_in_52_RREADY = in_52__m_axi_m_axi_RREADY;
  assign in_52__m_axi_m_axi_RRESP = m_axi_in_52_RRESP;
  assign in_52__m_axi_m_axi_RVALID = m_axi_in_52_RVALID;
  assign m_axi_in_52_WDATA = in_52__m_axi_m_axi_WDATA;
  assign m_axi_in_52_WLAST = in_52__m_axi_m_axi_WLAST;
  assign in_52__m_axi_m_axi_WREADY = m_axi_in_52_WREADY;
  assign m_axi_in_52_WSTRB = in_52__m_axi_m_axi_WSTRB;
  assign m_axi_in_52_WVALID = in_52__m_axi_m_axi_WVALID;
  assign in_52__m_axi_read_addr_din = in_52_read_addr__din;
  assign in_52_read_addr__full_n = in_52__m_axi_read_addr_full_n;
  assign in_52__m_axi_read_addr_write = in_52_read_addr__write;
  assign in_52_read_data__dout = in_52__m_axi_read_data_dout;
  assign in_52_read_data__empty_n = in_52__m_axi_read_data_empty_n;
  assign in_52__m_axi_read_data_read = in_52_read_data__read;
  assign in_52__m_axi_rst = ~ ap_rst_n;
  assign in_52__m_axi_write_addr_din = in_52_write_addr__din;
  assign in_52_write_addr__full_n = in_52__m_axi_write_addr_full_n;
  assign in_52__m_axi_write_addr_write = in_52_write_addr__write;
  assign in_52__m_axi_write_data_din = in_52_write_data__din;
  assign in_52_write_data__full_n = in_52__m_axi_write_data_full_n;
  assign in_52__m_axi_write_data_write = in_52_write_data__write;
  assign in_52_write_resp__dout = in_52__m_axi_write_resp_dout;
  assign in_52_write_resp__empty_n = in_52__m_axi_write_resp_empty_n;
  assign in_52__m_axi_write_resp_read = in_52_write_resp__read;
  assign in_53__m_axi_clk = ap_clk;
  assign m_axi_in_53_ARADDR = in_53__m_axi_m_axi_ARADDR;
  assign m_axi_in_53_ARBURST = in_53__m_axi_m_axi_ARBURST;
  assign m_axi_in_53_ARCACHE = in_53__m_axi_m_axi_ARCACHE;
  assign m_axi_in_53_ARID = in_53__m_axi_m_axi_ARID;
  assign m_axi_in_53_ARLEN = in_53__m_axi_m_axi_ARLEN;
  assign m_axi_in_53_ARLOCK = in_53__m_axi_m_axi_ARLOCK;
  assign m_axi_in_53_ARPROT = in_53__m_axi_m_axi_ARPROT;
  assign m_axi_in_53_ARQOS = in_53__m_axi_m_axi_ARQOS;
  assign in_53__m_axi_m_axi_ARREADY = m_axi_in_53_ARREADY;
  assign m_axi_in_53_ARSIZE = in_53__m_axi_m_axi_ARSIZE;
  assign m_axi_in_53_ARVALID = in_53__m_axi_m_axi_ARVALID;
  assign m_axi_in_53_AWADDR = in_53__m_axi_m_axi_AWADDR;
  assign m_axi_in_53_AWBURST = in_53__m_axi_m_axi_AWBURST;
  assign m_axi_in_53_AWCACHE = in_53__m_axi_m_axi_AWCACHE;
  assign m_axi_in_53_AWID = in_53__m_axi_m_axi_AWID;
  assign m_axi_in_53_AWLEN = in_53__m_axi_m_axi_AWLEN;
  assign m_axi_in_53_AWLOCK = in_53__m_axi_m_axi_AWLOCK;
  assign m_axi_in_53_AWPROT = in_53__m_axi_m_axi_AWPROT;
  assign m_axi_in_53_AWQOS = in_53__m_axi_m_axi_AWQOS;
  assign in_53__m_axi_m_axi_AWREADY = m_axi_in_53_AWREADY;
  assign m_axi_in_53_AWSIZE = in_53__m_axi_m_axi_AWSIZE;
  assign m_axi_in_53_AWVALID = in_53__m_axi_m_axi_AWVALID;
  assign in_53__m_axi_m_axi_BID = m_axi_in_53_BID;
  assign m_axi_in_53_BREADY = in_53__m_axi_m_axi_BREADY;
  assign in_53__m_axi_m_axi_BRESP = m_axi_in_53_BRESP;
  assign in_53__m_axi_m_axi_BVALID = m_axi_in_53_BVALID;
  assign in_53__m_axi_m_axi_RDATA = m_axi_in_53_RDATA;
  assign in_53__m_axi_m_axi_RID = m_axi_in_53_RID;
  assign in_53__m_axi_m_axi_RLAST = m_axi_in_53_RLAST;
  assign m_axi_in_53_RREADY = in_53__m_axi_m_axi_RREADY;
  assign in_53__m_axi_m_axi_RRESP = m_axi_in_53_RRESP;
  assign in_53__m_axi_m_axi_RVALID = m_axi_in_53_RVALID;
  assign m_axi_in_53_WDATA = in_53__m_axi_m_axi_WDATA;
  assign m_axi_in_53_WLAST = in_53__m_axi_m_axi_WLAST;
  assign in_53__m_axi_m_axi_WREADY = m_axi_in_53_WREADY;
  assign m_axi_in_53_WSTRB = in_53__m_axi_m_axi_WSTRB;
  assign m_axi_in_53_WVALID = in_53__m_axi_m_axi_WVALID;
  assign in_53__m_axi_read_addr_din = in_53_read_addr__din;
  assign in_53_read_addr__full_n = in_53__m_axi_read_addr_full_n;
  assign in_53__m_axi_read_addr_write = in_53_read_addr__write;
  assign in_53_read_data__dout = in_53__m_axi_read_data_dout;
  assign in_53_read_data__empty_n = in_53__m_axi_read_data_empty_n;
  assign in_53__m_axi_read_data_read = in_53_read_data__read;
  assign in_53__m_axi_rst = ~ ap_rst_n;
  assign in_53__m_axi_write_addr_din = in_53_write_addr__din;
  assign in_53_write_addr__full_n = in_53__m_axi_write_addr_full_n;
  assign in_53__m_axi_write_addr_write = in_53_write_addr__write;
  assign in_53__m_axi_write_data_din = in_53_write_data__din;
  assign in_53_write_data__full_n = in_53__m_axi_write_data_full_n;
  assign in_53__m_axi_write_data_write = in_53_write_data__write;
  assign in_53_write_resp__dout = in_53__m_axi_write_resp_dout;
  assign in_53_write_resp__empty_n = in_53__m_axi_write_resp_empty_n;
  assign in_53__m_axi_write_resp_read = in_53_write_resp__read;
  assign in_6__m_axi_clk = ap_clk;
  assign m_axi_in_6_ARADDR = in_6__m_axi_m_axi_ARADDR;
  assign m_axi_in_6_ARBURST = in_6__m_axi_m_axi_ARBURST;
  assign m_axi_in_6_ARCACHE = in_6__m_axi_m_axi_ARCACHE;
  assign m_axi_in_6_ARID = in_6__m_axi_m_axi_ARID;
  assign m_axi_in_6_ARLEN = in_6__m_axi_m_axi_ARLEN;
  assign m_axi_in_6_ARLOCK = in_6__m_axi_m_axi_ARLOCK;
  assign m_axi_in_6_ARPROT = in_6__m_axi_m_axi_ARPROT;
  assign m_axi_in_6_ARQOS = in_6__m_axi_m_axi_ARQOS;
  assign in_6__m_axi_m_axi_ARREADY = m_axi_in_6_ARREADY;
  assign m_axi_in_6_ARSIZE = in_6__m_axi_m_axi_ARSIZE;
  assign m_axi_in_6_ARVALID = in_6__m_axi_m_axi_ARVALID;
  assign m_axi_in_6_AWADDR = in_6__m_axi_m_axi_AWADDR;
  assign m_axi_in_6_AWBURST = in_6__m_axi_m_axi_AWBURST;
  assign m_axi_in_6_AWCACHE = in_6__m_axi_m_axi_AWCACHE;
  assign m_axi_in_6_AWID = in_6__m_axi_m_axi_AWID;
  assign m_axi_in_6_AWLEN = in_6__m_axi_m_axi_AWLEN;
  assign m_axi_in_6_AWLOCK = in_6__m_axi_m_axi_AWLOCK;
  assign m_axi_in_6_AWPROT = in_6__m_axi_m_axi_AWPROT;
  assign m_axi_in_6_AWQOS = in_6__m_axi_m_axi_AWQOS;
  assign in_6__m_axi_m_axi_AWREADY = m_axi_in_6_AWREADY;
  assign m_axi_in_6_AWSIZE = in_6__m_axi_m_axi_AWSIZE;
  assign m_axi_in_6_AWVALID = in_6__m_axi_m_axi_AWVALID;
  assign in_6__m_axi_m_axi_BID = m_axi_in_6_BID;
  assign m_axi_in_6_BREADY = in_6__m_axi_m_axi_BREADY;
  assign in_6__m_axi_m_axi_BRESP = m_axi_in_6_BRESP;
  assign in_6__m_axi_m_axi_BVALID = m_axi_in_6_BVALID;
  assign in_6__m_axi_m_axi_RDATA = m_axi_in_6_RDATA;
  assign in_6__m_axi_m_axi_RID = m_axi_in_6_RID;
  assign in_6__m_axi_m_axi_RLAST = m_axi_in_6_RLAST;
  assign m_axi_in_6_RREADY = in_6__m_axi_m_axi_RREADY;
  assign in_6__m_axi_m_axi_RRESP = m_axi_in_6_RRESP;
  assign in_6__m_axi_m_axi_RVALID = m_axi_in_6_RVALID;
  assign m_axi_in_6_WDATA = in_6__m_axi_m_axi_WDATA;
  assign m_axi_in_6_WLAST = in_6__m_axi_m_axi_WLAST;
  assign in_6__m_axi_m_axi_WREADY = m_axi_in_6_WREADY;
  assign m_axi_in_6_WSTRB = in_6__m_axi_m_axi_WSTRB;
  assign m_axi_in_6_WVALID = in_6__m_axi_m_axi_WVALID;
  assign in_6__m_axi_read_addr_din = in_6_read_addr__din;
  assign in_6_read_addr__full_n = in_6__m_axi_read_addr_full_n;
  assign in_6__m_axi_read_addr_write = in_6_read_addr__write;
  assign in_6_read_data__dout = in_6__m_axi_read_data_dout;
  assign in_6_read_data__empty_n = in_6__m_axi_read_data_empty_n;
  assign in_6__m_axi_read_data_read = in_6_read_data__read;
  assign in_6__m_axi_rst = ~ ap_rst_n;
  assign in_6__m_axi_write_addr_din = in_6_write_addr__din;
  assign in_6_write_addr__full_n = in_6__m_axi_write_addr_full_n;
  assign in_6__m_axi_write_addr_write = in_6_write_addr__write;
  assign in_6__m_axi_write_data_din = in_6_write_data__din;
  assign in_6_write_data__full_n = in_6__m_axi_write_data_full_n;
  assign in_6__m_axi_write_data_write = in_6_write_data__write;
  assign in_6_write_resp__dout = in_6__m_axi_write_resp_dout;
  assign in_6_write_resp__empty_n = in_6__m_axi_write_resp_empty_n;
  assign in_6__m_axi_write_resp_read = in_6_write_resp__read;
  assign in_7__m_axi_clk = ap_clk;
  assign m_axi_in_7_ARADDR = in_7__m_axi_m_axi_ARADDR;
  assign m_axi_in_7_ARBURST = in_7__m_axi_m_axi_ARBURST;
  assign m_axi_in_7_ARCACHE = in_7__m_axi_m_axi_ARCACHE;
  assign m_axi_in_7_ARID = in_7__m_axi_m_axi_ARID;
  assign m_axi_in_7_ARLEN = in_7__m_axi_m_axi_ARLEN;
  assign m_axi_in_7_ARLOCK = in_7__m_axi_m_axi_ARLOCK;
  assign m_axi_in_7_ARPROT = in_7__m_axi_m_axi_ARPROT;
  assign m_axi_in_7_ARQOS = in_7__m_axi_m_axi_ARQOS;
  assign in_7__m_axi_m_axi_ARREADY = m_axi_in_7_ARREADY;
  assign m_axi_in_7_ARSIZE = in_7__m_axi_m_axi_ARSIZE;
  assign m_axi_in_7_ARVALID = in_7__m_axi_m_axi_ARVALID;
  assign m_axi_in_7_AWADDR = in_7__m_axi_m_axi_AWADDR;
  assign m_axi_in_7_AWBURST = in_7__m_axi_m_axi_AWBURST;
  assign m_axi_in_7_AWCACHE = in_7__m_axi_m_axi_AWCACHE;
  assign m_axi_in_7_AWID = in_7__m_axi_m_axi_AWID;
  assign m_axi_in_7_AWLEN = in_7__m_axi_m_axi_AWLEN;
  assign m_axi_in_7_AWLOCK = in_7__m_axi_m_axi_AWLOCK;
  assign m_axi_in_7_AWPROT = in_7__m_axi_m_axi_AWPROT;
  assign m_axi_in_7_AWQOS = in_7__m_axi_m_axi_AWQOS;
  assign in_7__m_axi_m_axi_AWREADY = m_axi_in_7_AWREADY;
  assign m_axi_in_7_AWSIZE = in_7__m_axi_m_axi_AWSIZE;
  assign m_axi_in_7_AWVALID = in_7__m_axi_m_axi_AWVALID;
  assign in_7__m_axi_m_axi_BID = m_axi_in_7_BID;
  assign m_axi_in_7_BREADY = in_7__m_axi_m_axi_BREADY;
  assign in_7__m_axi_m_axi_BRESP = m_axi_in_7_BRESP;
  assign in_7__m_axi_m_axi_BVALID = m_axi_in_7_BVALID;
  assign in_7__m_axi_m_axi_RDATA = m_axi_in_7_RDATA;
  assign in_7__m_axi_m_axi_RID = m_axi_in_7_RID;
  assign in_7__m_axi_m_axi_RLAST = m_axi_in_7_RLAST;
  assign m_axi_in_7_RREADY = in_7__m_axi_m_axi_RREADY;
  assign in_7__m_axi_m_axi_RRESP = m_axi_in_7_RRESP;
  assign in_7__m_axi_m_axi_RVALID = m_axi_in_7_RVALID;
  assign m_axi_in_7_WDATA = in_7__m_axi_m_axi_WDATA;
  assign m_axi_in_7_WLAST = in_7__m_axi_m_axi_WLAST;
  assign in_7__m_axi_m_axi_WREADY = m_axi_in_7_WREADY;
  assign m_axi_in_7_WSTRB = in_7__m_axi_m_axi_WSTRB;
  assign m_axi_in_7_WVALID = in_7__m_axi_m_axi_WVALID;
  assign in_7__m_axi_read_addr_din = in_7_read_addr__din;
  assign in_7_read_addr__full_n = in_7__m_axi_read_addr_full_n;
  assign in_7__m_axi_read_addr_write = in_7_read_addr__write;
  assign in_7_read_data__dout = in_7__m_axi_read_data_dout;
  assign in_7_read_data__empty_n = in_7__m_axi_read_data_empty_n;
  assign in_7__m_axi_read_data_read = in_7_read_data__read;
  assign in_7__m_axi_rst = ~ ap_rst_n;
  assign in_7__m_axi_write_addr_din = in_7_write_addr__din;
  assign in_7_write_addr__full_n = in_7__m_axi_write_addr_full_n;
  assign in_7__m_axi_write_addr_write = in_7_write_addr__write;
  assign in_7__m_axi_write_data_din = in_7_write_data__din;
  assign in_7_write_data__full_n = in_7__m_axi_write_data_full_n;
  assign in_7__m_axi_write_data_write = in_7_write_data__write;
  assign in_7_write_resp__dout = in_7__m_axi_write_resp_dout;
  assign in_7_write_resp__empty_n = in_7__m_axi_write_resp_empty_n;
  assign in_7__m_axi_write_resp_read = in_7_write_resp__read;
  assign in_8__m_axi_clk = ap_clk;
  assign m_axi_in_8_ARADDR = in_8__m_axi_m_axi_ARADDR;
  assign m_axi_in_8_ARBURST = in_8__m_axi_m_axi_ARBURST;
  assign m_axi_in_8_ARCACHE = in_8__m_axi_m_axi_ARCACHE;
  assign m_axi_in_8_ARID = in_8__m_axi_m_axi_ARID;
  assign m_axi_in_8_ARLEN = in_8__m_axi_m_axi_ARLEN;
  assign m_axi_in_8_ARLOCK = in_8__m_axi_m_axi_ARLOCK;
  assign m_axi_in_8_ARPROT = in_8__m_axi_m_axi_ARPROT;
  assign m_axi_in_8_ARQOS = in_8__m_axi_m_axi_ARQOS;
  assign in_8__m_axi_m_axi_ARREADY = m_axi_in_8_ARREADY;
  assign m_axi_in_8_ARSIZE = in_8__m_axi_m_axi_ARSIZE;
  assign m_axi_in_8_ARVALID = in_8__m_axi_m_axi_ARVALID;
  assign m_axi_in_8_AWADDR = in_8__m_axi_m_axi_AWADDR;
  assign m_axi_in_8_AWBURST = in_8__m_axi_m_axi_AWBURST;
  assign m_axi_in_8_AWCACHE = in_8__m_axi_m_axi_AWCACHE;
  assign m_axi_in_8_AWID = in_8__m_axi_m_axi_AWID;
  assign m_axi_in_8_AWLEN = in_8__m_axi_m_axi_AWLEN;
  assign m_axi_in_8_AWLOCK = in_8__m_axi_m_axi_AWLOCK;
  assign m_axi_in_8_AWPROT = in_8__m_axi_m_axi_AWPROT;
  assign m_axi_in_8_AWQOS = in_8__m_axi_m_axi_AWQOS;
  assign in_8__m_axi_m_axi_AWREADY = m_axi_in_8_AWREADY;
  assign m_axi_in_8_AWSIZE = in_8__m_axi_m_axi_AWSIZE;
  assign m_axi_in_8_AWVALID = in_8__m_axi_m_axi_AWVALID;
  assign in_8__m_axi_m_axi_BID = m_axi_in_8_BID;
  assign m_axi_in_8_BREADY = in_8__m_axi_m_axi_BREADY;
  assign in_8__m_axi_m_axi_BRESP = m_axi_in_8_BRESP;
  assign in_8__m_axi_m_axi_BVALID = m_axi_in_8_BVALID;
  assign in_8__m_axi_m_axi_RDATA = m_axi_in_8_RDATA;
  assign in_8__m_axi_m_axi_RID = m_axi_in_8_RID;
  assign in_8__m_axi_m_axi_RLAST = m_axi_in_8_RLAST;
  assign m_axi_in_8_RREADY = in_8__m_axi_m_axi_RREADY;
  assign in_8__m_axi_m_axi_RRESP = m_axi_in_8_RRESP;
  assign in_8__m_axi_m_axi_RVALID = m_axi_in_8_RVALID;
  assign m_axi_in_8_WDATA = in_8__m_axi_m_axi_WDATA;
  assign m_axi_in_8_WLAST = in_8__m_axi_m_axi_WLAST;
  assign in_8__m_axi_m_axi_WREADY = m_axi_in_8_WREADY;
  assign m_axi_in_8_WSTRB = in_8__m_axi_m_axi_WSTRB;
  assign m_axi_in_8_WVALID = in_8__m_axi_m_axi_WVALID;
  assign in_8__m_axi_read_addr_din = in_8_read_addr__din;
  assign in_8_read_addr__full_n = in_8__m_axi_read_addr_full_n;
  assign in_8__m_axi_read_addr_write = in_8_read_addr__write;
  assign in_8_read_data__dout = in_8__m_axi_read_data_dout;
  assign in_8_read_data__empty_n = in_8__m_axi_read_data_empty_n;
  assign in_8__m_axi_read_data_read = in_8_read_data__read;
  assign in_8__m_axi_rst = ~ ap_rst_n;
  assign in_8__m_axi_write_addr_din = in_8_write_addr__din;
  assign in_8_write_addr__full_n = in_8__m_axi_write_addr_full_n;
  assign in_8__m_axi_write_addr_write = in_8_write_addr__write;
  assign in_8__m_axi_write_data_din = in_8_write_data__din;
  assign in_8_write_data__full_n = in_8__m_axi_write_data_full_n;
  assign in_8__m_axi_write_data_write = in_8_write_data__write;
  assign in_8_write_resp__dout = in_8__m_axi_write_resp_dout;
  assign in_8_write_resp__empty_n = in_8__m_axi_write_resp_empty_n;
  assign in_8__m_axi_write_resp_read = in_8_write_resp__read;
  assign in_9__m_axi_clk = ap_clk;
  assign m_axi_in_9_ARADDR = in_9__m_axi_m_axi_ARADDR;
  assign m_axi_in_9_ARBURST = in_9__m_axi_m_axi_ARBURST;
  assign m_axi_in_9_ARCACHE = in_9__m_axi_m_axi_ARCACHE;
  assign m_axi_in_9_ARID = in_9__m_axi_m_axi_ARID;
  assign m_axi_in_9_ARLEN = in_9__m_axi_m_axi_ARLEN;
  assign m_axi_in_9_ARLOCK = in_9__m_axi_m_axi_ARLOCK;
  assign m_axi_in_9_ARPROT = in_9__m_axi_m_axi_ARPROT;
  assign m_axi_in_9_ARQOS = in_9__m_axi_m_axi_ARQOS;
  assign in_9__m_axi_m_axi_ARREADY = m_axi_in_9_ARREADY;
  assign m_axi_in_9_ARSIZE = in_9__m_axi_m_axi_ARSIZE;
  assign m_axi_in_9_ARVALID = in_9__m_axi_m_axi_ARVALID;
  assign m_axi_in_9_AWADDR = in_9__m_axi_m_axi_AWADDR;
  assign m_axi_in_9_AWBURST = in_9__m_axi_m_axi_AWBURST;
  assign m_axi_in_9_AWCACHE = in_9__m_axi_m_axi_AWCACHE;
  assign m_axi_in_9_AWID = in_9__m_axi_m_axi_AWID;
  assign m_axi_in_9_AWLEN = in_9__m_axi_m_axi_AWLEN;
  assign m_axi_in_9_AWLOCK = in_9__m_axi_m_axi_AWLOCK;
  assign m_axi_in_9_AWPROT = in_9__m_axi_m_axi_AWPROT;
  assign m_axi_in_9_AWQOS = in_9__m_axi_m_axi_AWQOS;
  assign in_9__m_axi_m_axi_AWREADY = m_axi_in_9_AWREADY;
  assign m_axi_in_9_AWSIZE = in_9__m_axi_m_axi_AWSIZE;
  assign m_axi_in_9_AWVALID = in_9__m_axi_m_axi_AWVALID;
  assign in_9__m_axi_m_axi_BID = m_axi_in_9_BID;
  assign m_axi_in_9_BREADY = in_9__m_axi_m_axi_BREADY;
  assign in_9__m_axi_m_axi_BRESP = m_axi_in_9_BRESP;
  assign in_9__m_axi_m_axi_BVALID = m_axi_in_9_BVALID;
  assign in_9__m_axi_m_axi_RDATA = m_axi_in_9_RDATA;
  assign in_9__m_axi_m_axi_RID = m_axi_in_9_RID;
  assign in_9__m_axi_m_axi_RLAST = m_axi_in_9_RLAST;
  assign m_axi_in_9_RREADY = in_9__m_axi_m_axi_RREADY;
  assign in_9__m_axi_m_axi_RRESP = m_axi_in_9_RRESP;
  assign in_9__m_axi_m_axi_RVALID = m_axi_in_9_RVALID;
  assign m_axi_in_9_WDATA = in_9__m_axi_m_axi_WDATA;
  assign m_axi_in_9_WLAST = in_9__m_axi_m_axi_WLAST;
  assign in_9__m_axi_m_axi_WREADY = m_axi_in_9_WREADY;
  assign m_axi_in_9_WSTRB = in_9__m_axi_m_axi_WSTRB;
  assign m_axi_in_9_WVALID = in_9__m_axi_m_axi_WVALID;
  assign in_9__m_axi_read_addr_din = in_9_read_addr__din;
  assign in_9_read_addr__full_n = in_9__m_axi_read_addr_full_n;
  assign in_9__m_axi_read_addr_write = in_9_read_addr__write;
  assign in_9_read_data__dout = in_9__m_axi_read_data_dout;
  assign in_9_read_data__empty_n = in_9__m_axi_read_data_empty_n;
  assign in_9__m_axi_read_data_read = in_9_read_data__read;
  assign in_9__m_axi_rst = ~ ap_rst_n;
  assign in_9__m_axi_write_addr_din = in_9_write_addr__din;
  assign in_9_write_addr__full_n = in_9__m_axi_write_addr_full_n;
  assign in_9__m_axi_write_addr_write = in_9_write_addr__write;
  assign in_9__m_axi_write_data_din = in_9_write_data__din;
  assign in_9_write_data__full_n = in_9__m_axi_write_data_full_n;
  assign in_9__m_axi_write_data_write = in_9_write_data__write;
  assign in_9_write_resp__dout = in_9__m_axi_write_resp_dout;
  assign in_9_write_resp__empty_n = in_9__m_axi_write_resp_empty_n;
  assign in_9__m_axi_write_resp_read = in_9_write_resp__read;
  assign __tapa_fsm_unit_L4_out_dist = L4_out_dist;
  assign __tapa_fsm_unit_L4_out_id = L4_out_id;
  assign __tapa_fsm_unit_ap_clk = ap_clk;
  assign ap_done = __tapa_fsm_unit_ap_done;
  assign ap_idle = __tapa_fsm_unit_ap_idle;
  assign ap_ready = __tapa_fsm_unit_ap_ready;
  assign __tapa_fsm_unit_ap_rst_n = ap_rst_n;
  assign __tapa_fsm_unit_ap_start = ap_start;
  assign __tapa_fsm_unit_in_0 = in_0;
  assign __tapa_fsm_unit_in_1 = in_1;
  assign __tapa_fsm_unit_in_10 = in_10;
  assign __tapa_fsm_unit_in_11 = in_11;
  assign __tapa_fsm_unit_in_12 = in_12;
  assign __tapa_fsm_unit_in_13 = in_13;
  assign __tapa_fsm_unit_in_14 = in_14;
  assign __tapa_fsm_unit_in_15 = in_15;
  assign __tapa_fsm_unit_in_16 = in_16;
  assign __tapa_fsm_unit_in_17 = in_17;
  assign __tapa_fsm_unit_in_18 = in_18;
  assign __tapa_fsm_unit_in_19 = in_19;
  assign __tapa_fsm_unit_in_2 = in_2;
  assign __tapa_fsm_unit_in_20 = in_20;
  assign __tapa_fsm_unit_in_21 = in_21;
  assign __tapa_fsm_unit_in_22 = in_22;
  assign __tapa_fsm_unit_in_23 = in_23;
  assign __tapa_fsm_unit_in_24 = in_24;
  assign __tapa_fsm_unit_in_25 = in_25;
  assign __tapa_fsm_unit_in_26 = in_26;
  assign __tapa_fsm_unit_in_27 = in_27;
  assign __tapa_fsm_unit_in_28 = in_28;
  assign __tapa_fsm_unit_in_29 = in_29;
  assign __tapa_fsm_unit_in_3 = in_3;
  assign __tapa_fsm_unit_in_30 = in_30;
  assign __tapa_fsm_unit_in_31 = in_31;
  assign __tapa_fsm_unit_in_32 = in_32;
  assign __tapa_fsm_unit_in_33 = in_33;
  assign __tapa_fsm_unit_in_34 = in_34;
  assign __tapa_fsm_unit_in_35 = in_35;
  assign __tapa_fsm_unit_in_36 = in_36;
  assign __tapa_fsm_unit_in_37 = in_37;
  assign __tapa_fsm_unit_in_38 = in_38;
  assign __tapa_fsm_unit_in_39 = in_39;
  assign __tapa_fsm_unit_in_4 = in_4;
  assign __tapa_fsm_unit_in_40 = in_40;
  assign __tapa_fsm_unit_in_41 = in_41;
  assign __tapa_fsm_unit_in_42 = in_42;
  assign __tapa_fsm_unit_in_43 = in_43;
  assign __tapa_fsm_unit_in_44 = in_44;
  assign __tapa_fsm_unit_in_45 = in_45;
  assign __tapa_fsm_unit_in_46 = in_46;
  assign __tapa_fsm_unit_in_47 = in_47;
  assign __tapa_fsm_unit_in_48 = in_48;
  assign __tapa_fsm_unit_in_49 = in_49;
  assign __tapa_fsm_unit_in_5 = in_5;
  assign __tapa_fsm_unit_in_50 = in_50;
  assign __tapa_fsm_unit_in_51 = in_51;
  assign __tapa_fsm_unit_in_52 = in_52;
  assign __tapa_fsm_unit_in_53 = in_53;
  assign __tapa_fsm_unit_in_6 = in_6;
  assign __tapa_fsm_unit_in_7 = in_7;
  assign __tapa_fsm_unit_in_8 = in_8;
  assign __tapa_fsm_unit_in_9 = in_9;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_0__ap_done = krnl_globalSort_L1_L2_0__ap_done;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_0__ap_idle = krnl_globalSort_L1_L2_0__ap_idle;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_0__ap_ready = krnl_globalSort_L1_L2_0__ap_ready;
  assign krnl_globalSort_L1_L2_0__ap_start = __tapa_fsm_unit_krnl_globalSort_L1_L2_0__ap_start;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_10__ap_done = krnl_globalSort_L1_L2_10__ap_done;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_10__ap_idle = krnl_globalSort_L1_L2_10__ap_idle;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_10__ap_ready = krnl_globalSort_L1_L2_10__ap_ready;
  assign krnl_globalSort_L1_L2_10__ap_start = __tapa_fsm_unit_krnl_globalSort_L1_L2_10__ap_start;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_11__ap_done = krnl_globalSort_L1_L2_11__ap_done;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_11__ap_idle = krnl_globalSort_L1_L2_11__ap_idle;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_11__ap_ready = krnl_globalSort_L1_L2_11__ap_ready;
  assign krnl_globalSort_L1_L2_11__ap_start = __tapa_fsm_unit_krnl_globalSort_L1_L2_11__ap_start;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_12__ap_done = krnl_globalSort_L1_L2_12__ap_done;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_12__ap_idle = krnl_globalSort_L1_L2_12__ap_idle;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_12__ap_ready = krnl_globalSort_L1_L2_12__ap_ready;
  assign krnl_globalSort_L1_L2_12__ap_start = __tapa_fsm_unit_krnl_globalSort_L1_L2_12__ap_start;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_13__ap_done = krnl_globalSort_L1_L2_13__ap_done;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_13__ap_idle = krnl_globalSort_L1_L2_13__ap_idle;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_13__ap_ready = krnl_globalSort_L1_L2_13__ap_ready;
  assign krnl_globalSort_L1_L2_13__ap_start = __tapa_fsm_unit_krnl_globalSort_L1_L2_13__ap_start;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_14__ap_done = krnl_globalSort_L1_L2_14__ap_done;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_14__ap_idle = krnl_globalSort_L1_L2_14__ap_idle;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_14__ap_ready = krnl_globalSort_L1_L2_14__ap_ready;
  assign krnl_globalSort_L1_L2_14__ap_start = __tapa_fsm_unit_krnl_globalSort_L1_L2_14__ap_start;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_15__ap_done = krnl_globalSort_L1_L2_15__ap_done;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_15__ap_idle = krnl_globalSort_L1_L2_15__ap_idle;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_15__ap_ready = krnl_globalSort_L1_L2_15__ap_ready;
  assign krnl_globalSort_L1_L2_15__ap_start = __tapa_fsm_unit_krnl_globalSort_L1_L2_15__ap_start;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_16__ap_done = krnl_globalSort_L1_L2_16__ap_done;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_16__ap_idle = krnl_globalSort_L1_L2_16__ap_idle;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_16__ap_ready = krnl_globalSort_L1_L2_16__ap_ready;
  assign krnl_globalSort_L1_L2_16__ap_start = __tapa_fsm_unit_krnl_globalSort_L1_L2_16__ap_start;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_17__ap_done = krnl_globalSort_L1_L2_17__ap_done;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_17__ap_idle = krnl_globalSort_L1_L2_17__ap_idle;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_17__ap_ready = krnl_globalSort_L1_L2_17__ap_ready;
  assign krnl_globalSort_L1_L2_17__ap_start = __tapa_fsm_unit_krnl_globalSort_L1_L2_17__ap_start;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_18__ap_done = krnl_globalSort_L1_L2_18__ap_done;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_18__ap_idle = krnl_globalSort_L1_L2_18__ap_idle;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_18__ap_ready = krnl_globalSort_L1_L2_18__ap_ready;
  assign krnl_globalSort_L1_L2_18__ap_start = __tapa_fsm_unit_krnl_globalSort_L1_L2_18__ap_start;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_19__ap_done = krnl_globalSort_L1_L2_19__ap_done;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_19__ap_idle = krnl_globalSort_L1_L2_19__ap_idle;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_19__ap_ready = krnl_globalSort_L1_L2_19__ap_ready;
  assign krnl_globalSort_L1_L2_19__ap_start = __tapa_fsm_unit_krnl_globalSort_L1_L2_19__ap_start;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_1__ap_done = krnl_globalSort_L1_L2_1__ap_done;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_1__ap_idle = krnl_globalSort_L1_L2_1__ap_idle;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_1__ap_ready = krnl_globalSort_L1_L2_1__ap_ready;
  assign krnl_globalSort_L1_L2_1__ap_start = __tapa_fsm_unit_krnl_globalSort_L1_L2_1__ap_start;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_20__ap_done = krnl_globalSort_L1_L2_20__ap_done;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_20__ap_idle = krnl_globalSort_L1_L2_20__ap_idle;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_20__ap_ready = krnl_globalSort_L1_L2_20__ap_ready;
  assign krnl_globalSort_L1_L2_20__ap_start = __tapa_fsm_unit_krnl_globalSort_L1_L2_20__ap_start;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_21__ap_done = krnl_globalSort_L1_L2_21__ap_done;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_21__ap_idle = krnl_globalSort_L1_L2_21__ap_idle;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_21__ap_ready = krnl_globalSort_L1_L2_21__ap_ready;
  assign krnl_globalSort_L1_L2_21__ap_start = __tapa_fsm_unit_krnl_globalSort_L1_L2_21__ap_start;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_22__ap_done = krnl_globalSort_L1_L2_22__ap_done;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_22__ap_idle = krnl_globalSort_L1_L2_22__ap_idle;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_22__ap_ready = krnl_globalSort_L1_L2_22__ap_ready;
  assign krnl_globalSort_L1_L2_22__ap_start = __tapa_fsm_unit_krnl_globalSort_L1_L2_22__ap_start;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_23__ap_done = krnl_globalSort_L1_L2_23__ap_done;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_23__ap_idle = krnl_globalSort_L1_L2_23__ap_idle;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_23__ap_ready = krnl_globalSort_L1_L2_23__ap_ready;
  assign krnl_globalSort_L1_L2_23__ap_start = __tapa_fsm_unit_krnl_globalSort_L1_L2_23__ap_start;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_24__ap_done = krnl_globalSort_L1_L2_24__ap_done;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_24__ap_idle = krnl_globalSort_L1_L2_24__ap_idle;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_24__ap_ready = krnl_globalSort_L1_L2_24__ap_ready;
  assign krnl_globalSort_L1_L2_24__ap_start = __tapa_fsm_unit_krnl_globalSort_L1_L2_24__ap_start;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_25__ap_done = krnl_globalSort_L1_L2_25__ap_done;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_25__ap_idle = krnl_globalSort_L1_L2_25__ap_idle;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_25__ap_ready = krnl_globalSort_L1_L2_25__ap_ready;
  assign krnl_globalSort_L1_L2_25__ap_start = __tapa_fsm_unit_krnl_globalSort_L1_L2_25__ap_start;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_2__ap_done = krnl_globalSort_L1_L2_2__ap_done;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_2__ap_idle = krnl_globalSort_L1_L2_2__ap_idle;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_2__ap_ready = krnl_globalSort_L1_L2_2__ap_ready;
  assign krnl_globalSort_L1_L2_2__ap_start = __tapa_fsm_unit_krnl_globalSort_L1_L2_2__ap_start;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_3__ap_done = krnl_globalSort_L1_L2_3__ap_done;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_3__ap_idle = krnl_globalSort_L1_L2_3__ap_idle;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_3__ap_ready = krnl_globalSort_L1_L2_3__ap_ready;
  assign krnl_globalSort_L1_L2_3__ap_start = __tapa_fsm_unit_krnl_globalSort_L1_L2_3__ap_start;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_4__ap_done = krnl_globalSort_L1_L2_4__ap_done;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_4__ap_idle = krnl_globalSort_L1_L2_4__ap_idle;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_4__ap_ready = krnl_globalSort_L1_L2_4__ap_ready;
  assign krnl_globalSort_L1_L2_4__ap_start = __tapa_fsm_unit_krnl_globalSort_L1_L2_4__ap_start;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_5__ap_done = krnl_globalSort_L1_L2_5__ap_done;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_5__ap_idle = krnl_globalSort_L1_L2_5__ap_idle;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_5__ap_ready = krnl_globalSort_L1_L2_5__ap_ready;
  assign krnl_globalSort_L1_L2_5__ap_start = __tapa_fsm_unit_krnl_globalSort_L1_L2_5__ap_start;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_6__ap_done = krnl_globalSort_L1_L2_6__ap_done;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_6__ap_idle = krnl_globalSort_L1_L2_6__ap_idle;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_6__ap_ready = krnl_globalSort_L1_L2_6__ap_ready;
  assign krnl_globalSort_L1_L2_6__ap_start = __tapa_fsm_unit_krnl_globalSort_L1_L2_6__ap_start;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_7__ap_done = krnl_globalSort_L1_L2_7__ap_done;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_7__ap_idle = krnl_globalSort_L1_L2_7__ap_idle;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_7__ap_ready = krnl_globalSort_L1_L2_7__ap_ready;
  assign krnl_globalSort_L1_L2_7__ap_start = __tapa_fsm_unit_krnl_globalSort_L1_L2_7__ap_start;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_8__ap_done = krnl_globalSort_L1_L2_8__ap_done;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_8__ap_idle = krnl_globalSort_L1_L2_8__ap_idle;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_8__ap_ready = krnl_globalSort_L1_L2_8__ap_ready;
  assign krnl_globalSort_L1_L2_8__ap_start = __tapa_fsm_unit_krnl_globalSort_L1_L2_8__ap_start;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_9__ap_done = krnl_globalSort_L1_L2_9__ap_done;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_9__ap_idle = krnl_globalSort_L1_L2_9__ap_idle;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_9__ap_ready = krnl_globalSort_L1_L2_9__ap_ready;
  assign krnl_globalSort_L1_L2_9__ap_start = __tapa_fsm_unit_krnl_globalSort_L1_L2_9__ap_start;
  assign krnl_globalSort_L3_0___L4_out_dist__q0 = __tapa_fsm_unit_krnl_globalSort_L3_0___L4_out_dist__q0;
  assign krnl_globalSort_L3_0___L4_out_id__q0 = __tapa_fsm_unit_krnl_globalSort_L3_0___L4_out_id__q0;
  assign __tapa_fsm_unit_krnl_globalSort_L3_0__ap_done = krnl_globalSort_L3_0__ap_done;
  assign __tapa_fsm_unit_krnl_globalSort_L3_0__ap_idle = krnl_globalSort_L3_0__ap_idle;
  assign __tapa_fsm_unit_krnl_globalSort_L3_0__ap_ready = krnl_globalSort_L3_0__ap_ready;
  assign krnl_globalSort_L3_0__ap_start = __tapa_fsm_unit_krnl_globalSort_L3_0__ap_start;
  assign krnl_partialKnn_wrapper_0_0___in_0__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_0_0___in_0__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_0_0__ap_done = krnl_partialKnn_wrapper_0_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_0_0__ap_idle = krnl_partialKnn_wrapper_0_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_0_0__ap_ready = krnl_partialKnn_wrapper_0_0__ap_ready;
  assign krnl_partialKnn_wrapper_0_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_0_0__ap_start;
  assign krnl_partialKnn_wrapper_10_0___in_10__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_10_0___in_10__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_10_0__ap_done = krnl_partialKnn_wrapper_10_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_10_0__ap_idle = krnl_partialKnn_wrapper_10_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_10_0__ap_ready = krnl_partialKnn_wrapper_10_0__ap_ready;
  assign krnl_partialKnn_wrapper_10_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_10_0__ap_start;
  assign krnl_partialKnn_wrapper_11_0___in_11__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_11_0___in_11__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_11_0__ap_done = krnl_partialKnn_wrapper_11_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_11_0__ap_idle = krnl_partialKnn_wrapper_11_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_11_0__ap_ready = krnl_partialKnn_wrapper_11_0__ap_ready;
  assign krnl_partialKnn_wrapper_11_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_11_0__ap_start;
  assign krnl_partialKnn_wrapper_12_0___in_12__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_12_0___in_12__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_12_0__ap_done = krnl_partialKnn_wrapper_12_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_12_0__ap_idle = krnl_partialKnn_wrapper_12_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_12_0__ap_ready = krnl_partialKnn_wrapper_12_0__ap_ready;
  assign krnl_partialKnn_wrapper_12_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_12_0__ap_start;
  assign krnl_partialKnn_wrapper_13_0___in_13__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_13_0___in_13__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_13_0__ap_done = krnl_partialKnn_wrapper_13_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_13_0__ap_idle = krnl_partialKnn_wrapper_13_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_13_0__ap_ready = krnl_partialKnn_wrapper_13_0__ap_ready;
  assign krnl_partialKnn_wrapper_13_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_13_0__ap_start;
  assign krnl_partialKnn_wrapper_14_0___in_14__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_14_0___in_14__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_14_0__ap_done = krnl_partialKnn_wrapper_14_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_14_0__ap_idle = krnl_partialKnn_wrapper_14_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_14_0__ap_ready = krnl_partialKnn_wrapper_14_0__ap_ready;
  assign krnl_partialKnn_wrapper_14_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_14_0__ap_start;
  assign krnl_partialKnn_wrapper_15_0___in_15__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_15_0___in_15__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_15_0__ap_done = krnl_partialKnn_wrapper_15_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_15_0__ap_idle = krnl_partialKnn_wrapper_15_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_15_0__ap_ready = krnl_partialKnn_wrapper_15_0__ap_ready;
  assign krnl_partialKnn_wrapper_15_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_15_0__ap_start;
  assign krnl_partialKnn_wrapper_16_0___in_16__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_16_0___in_16__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_16_0__ap_done = krnl_partialKnn_wrapper_16_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_16_0__ap_idle = krnl_partialKnn_wrapper_16_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_16_0__ap_ready = krnl_partialKnn_wrapper_16_0__ap_ready;
  assign krnl_partialKnn_wrapper_16_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_16_0__ap_start;
  assign krnl_partialKnn_wrapper_17_0___in_17__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_17_0___in_17__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_17_0__ap_done = krnl_partialKnn_wrapper_17_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_17_0__ap_idle = krnl_partialKnn_wrapper_17_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_17_0__ap_ready = krnl_partialKnn_wrapper_17_0__ap_ready;
  assign krnl_partialKnn_wrapper_17_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_17_0__ap_start;
  assign krnl_partialKnn_wrapper_18_0___in_18__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_18_0___in_18__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_18_0__ap_done = krnl_partialKnn_wrapper_18_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_18_0__ap_idle = krnl_partialKnn_wrapper_18_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_18_0__ap_ready = krnl_partialKnn_wrapper_18_0__ap_ready;
  assign krnl_partialKnn_wrapper_18_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_18_0__ap_start;
  assign krnl_partialKnn_wrapper_19_0___in_19__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_19_0___in_19__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_19_0__ap_done = krnl_partialKnn_wrapper_19_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_19_0__ap_idle = krnl_partialKnn_wrapper_19_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_19_0__ap_ready = krnl_partialKnn_wrapper_19_0__ap_ready;
  assign krnl_partialKnn_wrapper_19_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_19_0__ap_start;
  assign krnl_partialKnn_wrapper_1_0___in_1__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_1_0___in_1__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_1_0__ap_done = krnl_partialKnn_wrapper_1_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_1_0__ap_idle = krnl_partialKnn_wrapper_1_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_1_0__ap_ready = krnl_partialKnn_wrapper_1_0__ap_ready;
  assign krnl_partialKnn_wrapper_1_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_1_0__ap_start;
  assign krnl_partialKnn_wrapper_20_0___in_20__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_20_0___in_20__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_20_0__ap_done = krnl_partialKnn_wrapper_20_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_20_0__ap_idle = krnl_partialKnn_wrapper_20_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_20_0__ap_ready = krnl_partialKnn_wrapper_20_0__ap_ready;
  assign krnl_partialKnn_wrapper_20_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_20_0__ap_start;
  assign krnl_partialKnn_wrapper_21_0___in_21__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_21_0___in_21__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_21_0__ap_done = krnl_partialKnn_wrapper_21_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_21_0__ap_idle = krnl_partialKnn_wrapper_21_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_21_0__ap_ready = krnl_partialKnn_wrapper_21_0__ap_ready;
  assign krnl_partialKnn_wrapper_21_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_21_0__ap_start;
  assign krnl_partialKnn_wrapper_22_0___in_22__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_22_0___in_22__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_22_0__ap_done = krnl_partialKnn_wrapper_22_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_22_0__ap_idle = krnl_partialKnn_wrapper_22_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_22_0__ap_ready = krnl_partialKnn_wrapper_22_0__ap_ready;
  assign krnl_partialKnn_wrapper_22_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_22_0__ap_start;
  assign krnl_partialKnn_wrapper_23_0___in_23__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_23_0___in_23__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_23_0__ap_done = krnl_partialKnn_wrapper_23_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_23_0__ap_idle = krnl_partialKnn_wrapper_23_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_23_0__ap_ready = krnl_partialKnn_wrapper_23_0__ap_ready;
  assign krnl_partialKnn_wrapper_23_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_23_0__ap_start;
  assign krnl_partialKnn_wrapper_24_0___in_24__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_24_0___in_24__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_24_0__ap_done = krnl_partialKnn_wrapper_24_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_24_0__ap_idle = krnl_partialKnn_wrapper_24_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_24_0__ap_ready = krnl_partialKnn_wrapper_24_0__ap_ready;
  assign krnl_partialKnn_wrapper_24_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_24_0__ap_start;
  assign krnl_partialKnn_wrapper_25_0___in_25__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_25_0___in_25__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_25_0__ap_done = krnl_partialKnn_wrapper_25_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_25_0__ap_idle = krnl_partialKnn_wrapper_25_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_25_0__ap_ready = krnl_partialKnn_wrapper_25_0__ap_ready;
  assign krnl_partialKnn_wrapper_25_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_25_0__ap_start;
  assign krnl_partialKnn_wrapper_26_0___in_26__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_26_0___in_26__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_26_0__ap_done = krnl_partialKnn_wrapper_26_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_26_0__ap_idle = krnl_partialKnn_wrapper_26_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_26_0__ap_ready = krnl_partialKnn_wrapper_26_0__ap_ready;
  assign krnl_partialKnn_wrapper_26_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_26_0__ap_start;
  assign krnl_partialKnn_wrapper_27_0___in_27__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_27_0___in_27__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_27_0__ap_done = krnl_partialKnn_wrapper_27_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_27_0__ap_idle = krnl_partialKnn_wrapper_27_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_27_0__ap_ready = krnl_partialKnn_wrapper_27_0__ap_ready;
  assign krnl_partialKnn_wrapper_27_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_27_0__ap_start;
  assign krnl_partialKnn_wrapper_28_0___in_28__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_28_0___in_28__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_28_0__ap_done = krnl_partialKnn_wrapper_28_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_28_0__ap_idle = krnl_partialKnn_wrapper_28_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_28_0__ap_ready = krnl_partialKnn_wrapper_28_0__ap_ready;
  assign krnl_partialKnn_wrapper_28_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_28_0__ap_start;
  assign krnl_partialKnn_wrapper_29_0___in_29__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_29_0___in_29__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_29_0__ap_done = krnl_partialKnn_wrapper_29_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_29_0__ap_idle = krnl_partialKnn_wrapper_29_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_29_0__ap_ready = krnl_partialKnn_wrapper_29_0__ap_ready;
  assign krnl_partialKnn_wrapper_29_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_29_0__ap_start;
  assign krnl_partialKnn_wrapper_2_0___in_2__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_2_0___in_2__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_2_0__ap_done = krnl_partialKnn_wrapper_2_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_2_0__ap_idle = krnl_partialKnn_wrapper_2_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_2_0__ap_ready = krnl_partialKnn_wrapper_2_0__ap_ready;
  assign krnl_partialKnn_wrapper_2_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_2_0__ap_start;
  assign krnl_partialKnn_wrapper_30_0___in_30__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_30_0___in_30__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_30_0__ap_done = krnl_partialKnn_wrapper_30_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_30_0__ap_idle = krnl_partialKnn_wrapper_30_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_30_0__ap_ready = krnl_partialKnn_wrapper_30_0__ap_ready;
  assign krnl_partialKnn_wrapper_30_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_30_0__ap_start;
  assign krnl_partialKnn_wrapper_31_0___in_31__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_31_0___in_31__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_31_0__ap_done = krnl_partialKnn_wrapper_31_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_31_0__ap_idle = krnl_partialKnn_wrapper_31_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_31_0__ap_ready = krnl_partialKnn_wrapper_31_0__ap_ready;
  assign krnl_partialKnn_wrapper_31_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_31_0__ap_start;
  assign krnl_partialKnn_wrapper_32_0___in_32__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_32_0___in_32__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_32_0__ap_done = krnl_partialKnn_wrapper_32_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_32_0__ap_idle = krnl_partialKnn_wrapper_32_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_32_0__ap_ready = krnl_partialKnn_wrapper_32_0__ap_ready;
  assign krnl_partialKnn_wrapper_32_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_32_0__ap_start;
  assign krnl_partialKnn_wrapper_33_0___in_33__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_33_0___in_33__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_33_0__ap_done = krnl_partialKnn_wrapper_33_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_33_0__ap_idle = krnl_partialKnn_wrapper_33_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_33_0__ap_ready = krnl_partialKnn_wrapper_33_0__ap_ready;
  assign krnl_partialKnn_wrapper_33_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_33_0__ap_start;
  assign krnl_partialKnn_wrapper_34_0___in_34__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_34_0___in_34__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_34_0__ap_done = krnl_partialKnn_wrapper_34_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_34_0__ap_idle = krnl_partialKnn_wrapper_34_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_34_0__ap_ready = krnl_partialKnn_wrapper_34_0__ap_ready;
  assign krnl_partialKnn_wrapper_34_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_34_0__ap_start;
  assign krnl_partialKnn_wrapper_35_0___in_35__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_35_0___in_35__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_35_0__ap_done = krnl_partialKnn_wrapper_35_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_35_0__ap_idle = krnl_partialKnn_wrapper_35_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_35_0__ap_ready = krnl_partialKnn_wrapper_35_0__ap_ready;
  assign krnl_partialKnn_wrapper_35_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_35_0__ap_start;
  assign krnl_partialKnn_wrapper_36_0___in_36__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_36_0___in_36__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_36_0__ap_done = krnl_partialKnn_wrapper_36_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_36_0__ap_idle = krnl_partialKnn_wrapper_36_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_36_0__ap_ready = krnl_partialKnn_wrapper_36_0__ap_ready;
  assign krnl_partialKnn_wrapper_36_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_36_0__ap_start;
  assign krnl_partialKnn_wrapper_37_0___in_37__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_37_0___in_37__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_37_0__ap_done = krnl_partialKnn_wrapper_37_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_37_0__ap_idle = krnl_partialKnn_wrapper_37_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_37_0__ap_ready = krnl_partialKnn_wrapper_37_0__ap_ready;
  assign krnl_partialKnn_wrapper_37_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_37_0__ap_start;
  assign krnl_partialKnn_wrapper_38_0___in_38__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_38_0___in_38__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_38_0__ap_done = krnl_partialKnn_wrapper_38_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_38_0__ap_idle = krnl_partialKnn_wrapper_38_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_38_0__ap_ready = krnl_partialKnn_wrapper_38_0__ap_ready;
  assign krnl_partialKnn_wrapper_38_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_38_0__ap_start;
  assign krnl_partialKnn_wrapper_39_0___in_39__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_39_0___in_39__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_39_0__ap_done = krnl_partialKnn_wrapper_39_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_39_0__ap_idle = krnl_partialKnn_wrapper_39_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_39_0__ap_ready = krnl_partialKnn_wrapper_39_0__ap_ready;
  assign krnl_partialKnn_wrapper_39_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_39_0__ap_start;
  assign krnl_partialKnn_wrapper_3_0___in_3__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_3_0___in_3__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_3_0__ap_done = krnl_partialKnn_wrapper_3_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_3_0__ap_idle = krnl_partialKnn_wrapper_3_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_3_0__ap_ready = krnl_partialKnn_wrapper_3_0__ap_ready;
  assign krnl_partialKnn_wrapper_3_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_3_0__ap_start;
  assign krnl_partialKnn_wrapper_40_0___in_40__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_40_0___in_40__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_40_0__ap_done = krnl_partialKnn_wrapper_40_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_40_0__ap_idle = krnl_partialKnn_wrapper_40_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_40_0__ap_ready = krnl_partialKnn_wrapper_40_0__ap_ready;
  assign krnl_partialKnn_wrapper_40_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_40_0__ap_start;
  assign krnl_partialKnn_wrapper_41_0___in_41__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_41_0___in_41__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_41_0__ap_done = krnl_partialKnn_wrapper_41_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_41_0__ap_idle = krnl_partialKnn_wrapper_41_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_41_0__ap_ready = krnl_partialKnn_wrapper_41_0__ap_ready;
  assign krnl_partialKnn_wrapper_41_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_41_0__ap_start;
  assign krnl_partialKnn_wrapper_42_0___in_42__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_42_0___in_42__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_42_0__ap_done = krnl_partialKnn_wrapper_42_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_42_0__ap_idle = krnl_partialKnn_wrapper_42_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_42_0__ap_ready = krnl_partialKnn_wrapper_42_0__ap_ready;
  assign krnl_partialKnn_wrapper_42_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_42_0__ap_start;
  assign krnl_partialKnn_wrapper_43_0___in_43__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_43_0___in_43__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_43_0__ap_done = krnl_partialKnn_wrapper_43_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_43_0__ap_idle = krnl_partialKnn_wrapper_43_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_43_0__ap_ready = krnl_partialKnn_wrapper_43_0__ap_ready;
  assign krnl_partialKnn_wrapper_43_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_43_0__ap_start;
  assign krnl_partialKnn_wrapper_44_0___in_44__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_44_0___in_44__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_44_0__ap_done = krnl_partialKnn_wrapper_44_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_44_0__ap_idle = krnl_partialKnn_wrapper_44_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_44_0__ap_ready = krnl_partialKnn_wrapper_44_0__ap_ready;
  assign krnl_partialKnn_wrapper_44_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_44_0__ap_start;
  assign krnl_partialKnn_wrapper_45_0___in_45__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_45_0___in_45__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_45_0__ap_done = krnl_partialKnn_wrapper_45_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_45_0__ap_idle = krnl_partialKnn_wrapper_45_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_45_0__ap_ready = krnl_partialKnn_wrapper_45_0__ap_ready;
  assign krnl_partialKnn_wrapper_45_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_45_0__ap_start;
  assign krnl_partialKnn_wrapper_46_0___in_46__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_46_0___in_46__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_46_0__ap_done = krnl_partialKnn_wrapper_46_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_46_0__ap_idle = krnl_partialKnn_wrapper_46_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_46_0__ap_ready = krnl_partialKnn_wrapper_46_0__ap_ready;
  assign krnl_partialKnn_wrapper_46_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_46_0__ap_start;
  assign krnl_partialKnn_wrapper_47_0___in_47__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_47_0___in_47__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_47_0__ap_done = krnl_partialKnn_wrapper_47_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_47_0__ap_idle = krnl_partialKnn_wrapper_47_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_47_0__ap_ready = krnl_partialKnn_wrapper_47_0__ap_ready;
  assign krnl_partialKnn_wrapper_47_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_47_0__ap_start;
  assign krnl_partialKnn_wrapper_48_0___in_48__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_48_0___in_48__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_48_0__ap_done = krnl_partialKnn_wrapper_48_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_48_0__ap_idle = krnl_partialKnn_wrapper_48_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_48_0__ap_ready = krnl_partialKnn_wrapper_48_0__ap_ready;
  assign krnl_partialKnn_wrapper_48_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_48_0__ap_start;
  assign krnl_partialKnn_wrapper_49_0___in_49__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_49_0___in_49__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_49_0__ap_done = krnl_partialKnn_wrapper_49_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_49_0__ap_idle = krnl_partialKnn_wrapper_49_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_49_0__ap_ready = krnl_partialKnn_wrapper_49_0__ap_ready;
  assign krnl_partialKnn_wrapper_49_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_49_0__ap_start;
  assign krnl_partialKnn_wrapper_4_0___in_4__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_4_0___in_4__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_4_0__ap_done = krnl_partialKnn_wrapper_4_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_4_0__ap_idle = krnl_partialKnn_wrapper_4_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_4_0__ap_ready = krnl_partialKnn_wrapper_4_0__ap_ready;
  assign krnl_partialKnn_wrapper_4_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_4_0__ap_start;
  assign krnl_partialKnn_wrapper_50_0___in_50__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_50_0___in_50__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_50_0__ap_done = krnl_partialKnn_wrapper_50_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_50_0__ap_idle = krnl_partialKnn_wrapper_50_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_50_0__ap_ready = krnl_partialKnn_wrapper_50_0__ap_ready;
  assign krnl_partialKnn_wrapper_50_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_50_0__ap_start;
  assign krnl_partialKnn_wrapper_51_0___in_51__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_51_0___in_51__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_51_0__ap_done = krnl_partialKnn_wrapper_51_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_51_0__ap_idle = krnl_partialKnn_wrapper_51_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_51_0__ap_ready = krnl_partialKnn_wrapper_51_0__ap_ready;
  assign krnl_partialKnn_wrapper_51_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_51_0__ap_start;
  assign krnl_partialKnn_wrapper_52_0___in_52__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_52_0___in_52__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_52_0__ap_done = krnl_partialKnn_wrapper_52_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_52_0__ap_idle = krnl_partialKnn_wrapper_52_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_52_0__ap_ready = krnl_partialKnn_wrapper_52_0__ap_ready;
  assign krnl_partialKnn_wrapper_52_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_52_0__ap_start;
  assign krnl_partialKnn_wrapper_53_0___in_53__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_53_0___in_53__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_53_0__ap_done = krnl_partialKnn_wrapper_53_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_53_0__ap_idle = krnl_partialKnn_wrapper_53_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_53_0__ap_ready = krnl_partialKnn_wrapper_53_0__ap_ready;
  assign krnl_partialKnn_wrapper_53_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_53_0__ap_start;
  assign krnl_partialKnn_wrapper_5_0___in_5__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_5_0___in_5__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_5_0__ap_done = krnl_partialKnn_wrapper_5_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_5_0__ap_idle = krnl_partialKnn_wrapper_5_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_5_0__ap_ready = krnl_partialKnn_wrapper_5_0__ap_ready;
  assign krnl_partialKnn_wrapper_5_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_5_0__ap_start;
  assign krnl_partialKnn_wrapper_6_0___in_6__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_6_0___in_6__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_6_0__ap_done = krnl_partialKnn_wrapper_6_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_6_0__ap_idle = krnl_partialKnn_wrapper_6_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_6_0__ap_ready = krnl_partialKnn_wrapper_6_0__ap_ready;
  assign krnl_partialKnn_wrapper_6_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_6_0__ap_start;
  assign krnl_partialKnn_wrapper_7_0___in_7__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_7_0___in_7__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_7_0__ap_done = krnl_partialKnn_wrapper_7_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_7_0__ap_idle = krnl_partialKnn_wrapper_7_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_7_0__ap_ready = krnl_partialKnn_wrapper_7_0__ap_ready;
  assign krnl_partialKnn_wrapper_7_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_7_0__ap_start;
  assign krnl_partialKnn_wrapper_8_0___in_8__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_8_0___in_8__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_8_0__ap_done = krnl_partialKnn_wrapper_8_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_8_0__ap_idle = krnl_partialKnn_wrapper_8_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_8_0__ap_ready = krnl_partialKnn_wrapper_8_0__ap_ready;
  assign krnl_partialKnn_wrapper_8_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_8_0__ap_start;
  assign krnl_partialKnn_wrapper_9_0___in_9__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_9_0___in_9__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_9_0__ap_done = krnl_partialKnn_wrapper_9_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_9_0__ap_idle = krnl_partialKnn_wrapper_9_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_9_0__ap_ready = krnl_partialKnn_wrapper_9_0__ap_ready;
  assign krnl_partialKnn_wrapper_9_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_9_0__ap_start;
endmodule