`timescale 1 ns / 1 ps

module Serpens_fsm
(
  ap_clk,
  ap_rst_n,
  ap_start,
  ap_ready,
  ap_done,
  ap_idle,
  Arbiter_Y_0__ap_start,
  Arbiter_Y_0__ap_ready,
  Arbiter_Y_0__ap_done,
  Arbiter_Y_0__ap_idle,
  Arbiter_Y_1__ap_start,
  Arbiter_Y_1__ap_ready,
  Arbiter_Y_1__ap_done,
  Arbiter_Y_1__ap_idle,
  Arbiter_Y_2__ap_start,
  Arbiter_Y_2__ap_ready,
  Arbiter_Y_2__ap_done,
  Arbiter_Y_2__ap_idle,
  Arbiter_Y_3__ap_start,
  Arbiter_Y_3__ap_ready,
  Arbiter_Y_3__ap_done,
  Arbiter_Y_3__ap_idle,
  Arbiter_Y_4__ap_start,
  Arbiter_Y_4__ap_ready,
  Arbiter_Y_4__ap_done,
  Arbiter_Y_4__ap_idle,
  Arbiter_Y_5__ap_start,
  Arbiter_Y_5__ap_ready,
  Arbiter_Y_5__ap_done,
  Arbiter_Y_5__ap_idle,
  Arbiter_Y_6__ap_start,
  Arbiter_Y_6__ap_ready,
  Arbiter_Y_6__ap_done,
  Arbiter_Y_6__ap_idle,
  Arbiter_Y_7__ap_start,
  Arbiter_Y_7__ap_ready,
  Arbiter_Y_7__ap_done,
  Arbiter_Y_7__ap_idle,
  FloatvAddFloatv_0__ap_start,
  FloatvMultConst_0__ap_start,
  FloatvMultConst_0__ap_ready,
  FloatvMultConst_0__ap_done,
  FloatvMultConst_0__ap_idle,
  FloatvMultConst_1__ap_start,
  FloatvMultConst_1__ap_ready,
  FloatvMultConst_1__ap_done,
  FloatvMultConst_1__ap_idle,
  Merger_Y_0__ap_start,
  PEG_Xvec_0__ap_start,
  PEG_Xvec_0__ap_ready,
  PEG_Xvec_0__ap_done,
  PEG_Xvec_0__ap_idle,
  PEG_Xvec_1__ap_start,
  PEG_Xvec_1__ap_ready,
  PEG_Xvec_1__ap_done,
  PEG_Xvec_1__ap_idle,
  PEG_Xvec_2__ap_start,
  PEG_Xvec_2__ap_ready,
  PEG_Xvec_2__ap_done,
  PEG_Xvec_2__ap_idle,
  PEG_Xvec_3__ap_start,
  PEG_Xvec_3__ap_ready,
  PEG_Xvec_3__ap_done,
  PEG_Xvec_3__ap_idle,
  PEG_Xvec_4__ap_start,
  PEG_Xvec_4__ap_ready,
  PEG_Xvec_4__ap_done,
  PEG_Xvec_4__ap_idle,
  PEG_Xvec_5__ap_start,
  PEG_Xvec_5__ap_ready,
  PEG_Xvec_5__ap_done,
  PEG_Xvec_5__ap_idle,
  PEG_Xvec_6__ap_start,
  PEG_Xvec_6__ap_ready,
  PEG_Xvec_6__ap_done,
  PEG_Xvec_6__ap_idle,
  PEG_Xvec_7__ap_start,
  PEG_Xvec_7__ap_ready,
  PEG_Xvec_7__ap_done,
  PEG_Xvec_7__ap_idle,
  PEG_Xvec_8__ap_start,
  PEG_Xvec_8__ap_ready,
  PEG_Xvec_8__ap_done,
  PEG_Xvec_8__ap_idle,
  PEG_Xvec_9__ap_start,
  PEG_Xvec_9__ap_ready,
  PEG_Xvec_9__ap_done,
  PEG_Xvec_9__ap_idle,
  PEG_Xvec_10__ap_start,
  PEG_Xvec_10__ap_ready,
  PEG_Xvec_10__ap_done,
  PEG_Xvec_10__ap_idle,
  PEG_Xvec_11__ap_start,
  PEG_Xvec_11__ap_ready,
  PEG_Xvec_11__ap_done,
  PEG_Xvec_11__ap_idle,
  PEG_Xvec_12__ap_start,
  PEG_Xvec_12__ap_ready,
  PEG_Xvec_12__ap_done,
  PEG_Xvec_12__ap_idle,
  PEG_Xvec_13__ap_start,
  PEG_Xvec_13__ap_ready,
  PEG_Xvec_13__ap_done,
  PEG_Xvec_13__ap_idle,
  PEG_Xvec_14__ap_start,
  PEG_Xvec_14__ap_ready,
  PEG_Xvec_14__ap_done,
  PEG_Xvec_14__ap_idle,
  PEG_Xvec_15__ap_start,
  PEG_Xvec_15__ap_ready,
  PEG_Xvec_15__ap_done,
  PEG_Xvec_15__ap_idle,
  PEG_Xvec_16__ap_start,
  PEG_Xvec_16__ap_ready,
  PEG_Xvec_16__ap_done,
  PEG_Xvec_16__ap_idle,
  PEG_Xvec_17__ap_start,
  PEG_Xvec_17__ap_ready,
  PEG_Xvec_17__ap_done,
  PEG_Xvec_17__ap_idle,
  PEG_Xvec_18__ap_start,
  PEG_Xvec_18__ap_ready,
  PEG_Xvec_18__ap_done,
  PEG_Xvec_18__ap_idle,
  PEG_Xvec_19__ap_start,
  PEG_Xvec_19__ap_ready,
  PEG_Xvec_19__ap_done,
  PEG_Xvec_19__ap_idle,
  PEG_Xvec_20__ap_start,
  PEG_Xvec_20__ap_ready,
  PEG_Xvec_20__ap_done,
  PEG_Xvec_20__ap_idle,
  PEG_Xvec_21__ap_start,
  PEG_Xvec_21__ap_ready,
  PEG_Xvec_21__ap_done,
  PEG_Xvec_21__ap_idle,
  PEG_Xvec_22__ap_start,
  PEG_Xvec_22__ap_ready,
  PEG_Xvec_22__ap_done,
  PEG_Xvec_22__ap_idle,
  PEG_Xvec_23__ap_start,
  PEG_Xvec_23__ap_ready,
  PEG_Xvec_23__ap_done,
  PEG_Xvec_23__ap_idle,
  PEG_Xvec_24__ap_start,
  PEG_Xvec_24__ap_ready,
  PEG_Xvec_24__ap_done,
  PEG_Xvec_24__ap_idle,
  PEG_Xvec_25__ap_start,
  PEG_Xvec_25__ap_ready,
  PEG_Xvec_25__ap_done,
  PEG_Xvec_25__ap_idle,
  PEG_Xvec_26__ap_start,
  PEG_Xvec_26__ap_ready,
  PEG_Xvec_26__ap_done,
  PEG_Xvec_26__ap_idle,
  PEG_Xvec_27__ap_start,
  PEG_Xvec_27__ap_ready,
  PEG_Xvec_27__ap_done,
  PEG_Xvec_27__ap_idle,
  PEG_Xvec_28__ap_start,
  PEG_Xvec_28__ap_ready,
  PEG_Xvec_28__ap_done,
  PEG_Xvec_28__ap_idle,
  PEG_Xvec_29__ap_start,
  PEG_Xvec_29__ap_ready,
  PEG_Xvec_29__ap_done,
  PEG_Xvec_29__ap_idle,
  PEG_Xvec_30__ap_start,
  PEG_Xvec_30__ap_ready,
  PEG_Xvec_30__ap_done,
  PEG_Xvec_30__ap_idle,
  PEG_Xvec_31__ap_start,
  PEG_Xvec_31__ap_ready,
  PEG_Xvec_31__ap_done,
  PEG_Xvec_31__ap_idle,
  PEG_Xvec_32__ap_start,
  PEG_Xvec_32__ap_ready,
  PEG_Xvec_32__ap_done,
  PEG_Xvec_32__ap_idle,
  PEG_Xvec_33__ap_start,
  PEG_Xvec_33__ap_ready,
  PEG_Xvec_33__ap_done,
  PEG_Xvec_33__ap_idle,
  PEG_Xvec_34__ap_start,
  PEG_Xvec_34__ap_ready,
  PEG_Xvec_34__ap_done,
  PEG_Xvec_34__ap_idle,
  PEG_Xvec_35__ap_start,
  PEG_Xvec_35__ap_ready,
  PEG_Xvec_35__ap_done,
  PEG_Xvec_35__ap_idle,
  PEG_Xvec_36__ap_start,
  PEG_Xvec_36__ap_ready,
  PEG_Xvec_36__ap_done,
  PEG_Xvec_36__ap_idle,
  PEG_Xvec_37__ap_start,
  PEG_Xvec_37__ap_ready,
  PEG_Xvec_37__ap_done,
  PEG_Xvec_37__ap_idle,
  PEG_Xvec_38__ap_start,
  PEG_Xvec_38__ap_ready,
  PEG_Xvec_38__ap_done,
  PEG_Xvec_38__ap_idle,
  PEG_Xvec_39__ap_start,
  PEG_Xvec_39__ap_ready,
  PEG_Xvec_39__ap_done,
  PEG_Xvec_39__ap_idle,
  PEG_Xvec_40__ap_start,
  PEG_Xvec_40__ap_ready,
  PEG_Xvec_40__ap_done,
  PEG_Xvec_40__ap_idle,
  PEG_Xvec_41__ap_start,
  PEG_Xvec_41__ap_ready,
  PEG_Xvec_41__ap_done,
  PEG_Xvec_41__ap_idle,
  PEG_Xvec_42__ap_start,
  PEG_Xvec_42__ap_ready,
  PEG_Xvec_42__ap_done,
  PEG_Xvec_42__ap_idle,
  PEG_Xvec_43__ap_start,
  PEG_Xvec_43__ap_ready,
  PEG_Xvec_43__ap_done,
  PEG_Xvec_43__ap_idle,
  PEG_Xvec_44__ap_start,
  PEG_Xvec_44__ap_ready,
  PEG_Xvec_44__ap_done,
  PEG_Xvec_44__ap_idle,
  PEG_Xvec_45__ap_start,
  PEG_Xvec_45__ap_ready,
  PEG_Xvec_45__ap_done,
  PEG_Xvec_45__ap_idle,
  PEG_Xvec_46__ap_start,
  PEG_Xvec_46__ap_ready,
  PEG_Xvec_46__ap_done,
  PEG_Xvec_46__ap_idle,
  PEG_Xvec_47__ap_start,
  PEG_Xvec_47__ap_ready,
  PEG_Xvec_47__ap_done,
  PEG_Xvec_47__ap_idle,
  PEG_Xvec_48__ap_start,
  PEG_Xvec_48__ap_ready,
  PEG_Xvec_48__ap_done,
  PEG_Xvec_48__ap_idle,
  PEG_Xvec_49__ap_start,
  PEG_Xvec_49__ap_ready,
  PEG_Xvec_49__ap_done,
  PEG_Xvec_49__ap_idle,
  PEG_Xvec_50__ap_start,
  PEG_Xvec_50__ap_ready,
  PEG_Xvec_50__ap_done,
  PEG_Xvec_50__ap_idle,
  PEG_Xvec_51__ap_start,
  PEG_Xvec_51__ap_ready,
  PEG_Xvec_51__ap_done,
  PEG_Xvec_51__ap_idle,
  PEG_Xvec_52__ap_start,
  PEG_Xvec_52__ap_ready,
  PEG_Xvec_52__ap_done,
  PEG_Xvec_52__ap_idle,
  PEG_Xvec_53__ap_start,
  PEG_Xvec_53__ap_ready,
  PEG_Xvec_53__ap_done,
  PEG_Xvec_53__ap_idle,
  PEG_Xvec_54__ap_start,
  PEG_Xvec_54__ap_ready,
  PEG_Xvec_54__ap_done,
  PEG_Xvec_54__ap_idle,
  PEG_Xvec_55__ap_start,
  PEG_Xvec_55__ap_ready,
  PEG_Xvec_55__ap_done,
  PEG_Xvec_55__ap_idle,
  PEG_Yvec_0__ap_start,
  PEG_Yvec_0__ap_ready,
  PEG_Yvec_0__ap_done,
  PEG_Yvec_0__ap_idle,
  PEG_Yvec_1__ap_start,
  PEG_Yvec_1__ap_ready,
  PEG_Yvec_1__ap_done,
  PEG_Yvec_1__ap_idle,
  PEG_Yvec_2__ap_start,
  PEG_Yvec_2__ap_ready,
  PEG_Yvec_2__ap_done,
  PEG_Yvec_2__ap_idle,
  PEG_Yvec_3__ap_start,
  PEG_Yvec_3__ap_ready,
  PEG_Yvec_3__ap_done,
  PEG_Yvec_3__ap_idle,
  PEG_Yvec_4__ap_start,
  PEG_Yvec_4__ap_ready,
  PEG_Yvec_4__ap_done,
  PEG_Yvec_4__ap_idle,
  PEG_Yvec_5__ap_start,
  PEG_Yvec_5__ap_ready,
  PEG_Yvec_5__ap_done,
  PEG_Yvec_5__ap_idle,
  PEG_Yvec_6__ap_start,
  PEG_Yvec_6__ap_ready,
  PEG_Yvec_6__ap_done,
  PEG_Yvec_6__ap_idle,
  PEG_Yvec_7__ap_start,
  PEG_Yvec_7__ap_ready,
  PEG_Yvec_7__ap_done,
  PEG_Yvec_7__ap_idle,
  PEG_Yvec_8__ap_start,
  PEG_Yvec_8__ap_ready,
  PEG_Yvec_8__ap_done,
  PEG_Yvec_8__ap_idle,
  PEG_Yvec_9__ap_start,
  PEG_Yvec_9__ap_ready,
  PEG_Yvec_9__ap_done,
  PEG_Yvec_9__ap_idle,
  PEG_Yvec_10__ap_start,
  PEG_Yvec_10__ap_ready,
  PEG_Yvec_10__ap_done,
  PEG_Yvec_10__ap_idle,
  PEG_Yvec_11__ap_start,
  PEG_Yvec_11__ap_ready,
  PEG_Yvec_11__ap_done,
  PEG_Yvec_11__ap_idle,
  PEG_Yvec_12__ap_start,
  PEG_Yvec_12__ap_ready,
  PEG_Yvec_12__ap_done,
  PEG_Yvec_12__ap_idle,
  PEG_Yvec_13__ap_start,
  PEG_Yvec_13__ap_ready,
  PEG_Yvec_13__ap_done,
  PEG_Yvec_13__ap_idle,
  PEG_Yvec_14__ap_start,
  PEG_Yvec_14__ap_ready,
  PEG_Yvec_14__ap_done,
  PEG_Yvec_14__ap_idle,
  PEG_Yvec_15__ap_start,
  PEG_Yvec_15__ap_ready,
  PEG_Yvec_15__ap_done,
  PEG_Yvec_15__ap_idle,
  PEG_Yvec_16__ap_start,
  PEG_Yvec_16__ap_ready,
  PEG_Yvec_16__ap_done,
  PEG_Yvec_16__ap_idle,
  PEG_Yvec_17__ap_start,
  PEG_Yvec_17__ap_ready,
  PEG_Yvec_17__ap_done,
  PEG_Yvec_17__ap_idle,
  PEG_Yvec_18__ap_start,
  PEG_Yvec_18__ap_ready,
  PEG_Yvec_18__ap_done,
  PEG_Yvec_18__ap_idle,
  PEG_Yvec_19__ap_start,
  PEG_Yvec_19__ap_ready,
  PEG_Yvec_19__ap_done,
  PEG_Yvec_19__ap_idle,
  PEG_Yvec_20__ap_start,
  PEG_Yvec_20__ap_ready,
  PEG_Yvec_20__ap_done,
  PEG_Yvec_20__ap_idle,
  PEG_Yvec_21__ap_start,
  PEG_Yvec_21__ap_ready,
  PEG_Yvec_21__ap_done,
  PEG_Yvec_21__ap_idle,
  PEG_Yvec_22__ap_start,
  PEG_Yvec_22__ap_ready,
  PEG_Yvec_22__ap_done,
  PEG_Yvec_22__ap_idle,
  PEG_Yvec_23__ap_start,
  PEG_Yvec_23__ap_ready,
  PEG_Yvec_23__ap_done,
  PEG_Yvec_23__ap_idle,
  PEG_Yvec_24__ap_start,
  PEG_Yvec_24__ap_ready,
  PEG_Yvec_24__ap_done,
  PEG_Yvec_24__ap_idle,
  PEG_Yvec_25__ap_start,
  PEG_Yvec_25__ap_ready,
  PEG_Yvec_25__ap_done,
  PEG_Yvec_25__ap_idle,
  PEG_Yvec_26__ap_start,
  PEG_Yvec_26__ap_ready,
  PEG_Yvec_26__ap_done,
  PEG_Yvec_26__ap_idle,
  PEG_Yvec_27__ap_start,
  PEG_Yvec_27__ap_ready,
  PEG_Yvec_27__ap_done,
  PEG_Yvec_27__ap_idle,
  PEG_Yvec_28__ap_start,
  PEG_Yvec_28__ap_ready,
  PEG_Yvec_28__ap_done,
  PEG_Yvec_28__ap_idle,
  PEG_Yvec_29__ap_start,
  PEG_Yvec_29__ap_ready,
  PEG_Yvec_29__ap_done,
  PEG_Yvec_29__ap_idle,
  PEG_Yvec_30__ap_start,
  PEG_Yvec_30__ap_ready,
  PEG_Yvec_30__ap_done,
  PEG_Yvec_30__ap_idle,
  PEG_Yvec_31__ap_start,
  PEG_Yvec_31__ap_ready,
  PEG_Yvec_31__ap_done,
  PEG_Yvec_31__ap_idle,
  PEG_Yvec_32__ap_start,
  PEG_Yvec_32__ap_ready,
  PEG_Yvec_32__ap_done,
  PEG_Yvec_32__ap_idle,
  PEG_Yvec_33__ap_start,
  PEG_Yvec_33__ap_ready,
  PEG_Yvec_33__ap_done,
  PEG_Yvec_33__ap_idle,
  PEG_Yvec_34__ap_start,
  PEG_Yvec_34__ap_ready,
  PEG_Yvec_34__ap_done,
  PEG_Yvec_34__ap_idle,
  PEG_Yvec_35__ap_start,
  PEG_Yvec_35__ap_ready,
  PEG_Yvec_35__ap_done,
  PEG_Yvec_35__ap_idle,
  PEG_Yvec_36__ap_start,
  PEG_Yvec_36__ap_ready,
  PEG_Yvec_36__ap_done,
  PEG_Yvec_36__ap_idle,
  PEG_Yvec_37__ap_start,
  PEG_Yvec_37__ap_ready,
  PEG_Yvec_37__ap_done,
  PEG_Yvec_37__ap_idle,
  PEG_Yvec_38__ap_start,
  PEG_Yvec_38__ap_ready,
  PEG_Yvec_38__ap_done,
  PEG_Yvec_38__ap_idle,
  PEG_Yvec_39__ap_start,
  PEG_Yvec_39__ap_ready,
  PEG_Yvec_39__ap_done,
  PEG_Yvec_39__ap_idle,
  PEG_Yvec_40__ap_start,
  PEG_Yvec_40__ap_ready,
  PEG_Yvec_40__ap_done,
  PEG_Yvec_40__ap_idle,
  PEG_Yvec_41__ap_start,
  PEG_Yvec_41__ap_ready,
  PEG_Yvec_41__ap_done,
  PEG_Yvec_41__ap_idle,
  PEG_Yvec_42__ap_start,
  PEG_Yvec_42__ap_ready,
  PEG_Yvec_42__ap_done,
  PEG_Yvec_42__ap_idle,
  PEG_Yvec_43__ap_start,
  PEG_Yvec_43__ap_ready,
  PEG_Yvec_43__ap_done,
  PEG_Yvec_43__ap_idle,
  PEG_Yvec_44__ap_start,
  PEG_Yvec_44__ap_ready,
  PEG_Yvec_44__ap_done,
  PEG_Yvec_44__ap_idle,
  PEG_Yvec_45__ap_start,
  PEG_Yvec_45__ap_ready,
  PEG_Yvec_45__ap_done,
  PEG_Yvec_45__ap_idle,
  PEG_Yvec_46__ap_start,
  PEG_Yvec_46__ap_ready,
  PEG_Yvec_46__ap_done,
  PEG_Yvec_46__ap_idle,
  PEG_Yvec_47__ap_start,
  PEG_Yvec_47__ap_ready,
  PEG_Yvec_47__ap_done,
  PEG_Yvec_47__ap_idle,
  PEG_Yvec_48__ap_start,
  PEG_Yvec_48__ap_ready,
  PEG_Yvec_48__ap_done,
  PEG_Yvec_48__ap_idle,
  PEG_Yvec_49__ap_start,
  PEG_Yvec_49__ap_ready,
  PEG_Yvec_49__ap_done,
  PEG_Yvec_49__ap_idle,
  PEG_Yvec_50__ap_start,
  PEG_Yvec_50__ap_ready,
  PEG_Yvec_50__ap_done,
  PEG_Yvec_50__ap_idle,
  PEG_Yvec_51__ap_start,
  PEG_Yvec_51__ap_ready,
  PEG_Yvec_51__ap_done,
  PEG_Yvec_51__ap_idle,
  PEG_Yvec_52__ap_start,
  PEG_Yvec_52__ap_ready,
  PEG_Yvec_52__ap_done,
  PEG_Yvec_52__ap_idle,
  PEG_Yvec_53__ap_start,
  PEG_Yvec_53__ap_ready,
  PEG_Yvec_53__ap_done,
  PEG_Yvec_53__ap_idle,
  PEG_Yvec_54__ap_start,
  PEG_Yvec_54__ap_ready,
  PEG_Yvec_54__ap_done,
  PEG_Yvec_54__ap_idle,
  PEG_Yvec_55__ap_start,
  PEG_Yvec_55__ap_ready,
  PEG_Yvec_55__ap_done,
  PEG_Yvec_55__ap_idle,
  black_hole_float_v16_0__ap_start,
  black_hole_int_0__ap_start,
  read_A_0__ap_start,
  read_A_0__ap_ready,
  read_A_0__ap_done,
  read_A_0__ap_idle,
  read_A_1__ap_start,
  read_A_1__ap_ready,
  read_A_1__ap_done,
  read_A_1__ap_idle,
  read_A_2__ap_start,
  read_A_2__ap_ready,
  read_A_2__ap_done,
  read_A_2__ap_idle,
  read_A_3__ap_start,
  read_A_3__ap_ready,
  read_A_3__ap_done,
  read_A_3__ap_idle,
  read_A_4__ap_start,
  read_A_4__ap_ready,
  read_A_4__ap_done,
  read_A_4__ap_idle,
  read_A_5__ap_start,
  read_A_5__ap_ready,
  read_A_5__ap_done,
  read_A_5__ap_idle,
  read_A_6__ap_start,
  read_A_6__ap_ready,
  read_A_6__ap_done,
  read_A_6__ap_idle,
  read_A_7__ap_start,
  read_A_7__ap_ready,
  read_A_7__ap_done,
  read_A_7__ap_idle,
  read_A_8__ap_start,
  read_A_8__ap_ready,
  read_A_8__ap_done,
  read_A_8__ap_idle,
  read_A_9__ap_start,
  read_A_9__ap_ready,
  read_A_9__ap_done,
  read_A_9__ap_idle,
  read_A_10__ap_start,
  read_A_10__ap_ready,
  read_A_10__ap_done,
  read_A_10__ap_idle,
  read_A_11__ap_start,
  read_A_11__ap_ready,
  read_A_11__ap_done,
  read_A_11__ap_idle,
  read_A_12__ap_start,
  read_A_12__ap_ready,
  read_A_12__ap_done,
  read_A_12__ap_idle,
  read_A_13__ap_start,
  read_A_13__ap_ready,
  read_A_13__ap_done,
  read_A_13__ap_idle,
  read_A_14__ap_start,
  read_A_14__ap_ready,
  read_A_14__ap_done,
  read_A_14__ap_idle,
  read_A_15__ap_start,
  read_A_15__ap_ready,
  read_A_15__ap_done,
  read_A_15__ap_idle,
  read_A_16__ap_start,
  read_A_16__ap_ready,
  read_A_16__ap_done,
  read_A_16__ap_idle,
  read_A_17__ap_start,
  read_A_17__ap_ready,
  read_A_17__ap_done,
  read_A_17__ap_idle,
  read_A_18__ap_start,
  read_A_18__ap_ready,
  read_A_18__ap_done,
  read_A_18__ap_idle,
  read_A_19__ap_start,
  read_A_19__ap_ready,
  read_A_19__ap_done,
  read_A_19__ap_idle,
  read_A_20__ap_start,
  read_A_20__ap_ready,
  read_A_20__ap_done,
  read_A_20__ap_idle,
  read_A_21__ap_start,
  read_A_21__ap_ready,
  read_A_21__ap_done,
  read_A_21__ap_idle,
  read_A_22__ap_start,
  read_A_22__ap_ready,
  read_A_22__ap_done,
  read_A_22__ap_idle,
  read_A_23__ap_start,
  read_A_23__ap_ready,
  read_A_23__ap_done,
  read_A_23__ap_idle,
  read_A_24__ap_start,
  read_A_24__ap_ready,
  read_A_24__ap_done,
  read_A_24__ap_idle,
  read_A_25__ap_start,
  read_A_25__ap_ready,
  read_A_25__ap_done,
  read_A_25__ap_idle,
  read_A_26__ap_start,
  read_A_26__ap_ready,
  read_A_26__ap_done,
  read_A_26__ap_idle,
  read_A_27__ap_start,
  read_A_27__ap_ready,
  read_A_27__ap_done,
  read_A_27__ap_idle,
  read_A_28__ap_start,
  read_A_28__ap_ready,
  read_A_28__ap_done,
  read_A_28__ap_idle,
  read_A_29__ap_start,
  read_A_29__ap_ready,
  read_A_29__ap_done,
  read_A_29__ap_idle,
  read_A_30__ap_start,
  read_A_30__ap_ready,
  read_A_30__ap_done,
  read_A_30__ap_idle,
  read_A_31__ap_start,
  read_A_31__ap_ready,
  read_A_31__ap_done,
  read_A_31__ap_idle,
  read_A_32__ap_start,
  read_A_32__ap_ready,
  read_A_32__ap_done,
  read_A_32__ap_idle,
  read_A_33__ap_start,
  read_A_33__ap_ready,
  read_A_33__ap_done,
  read_A_33__ap_idle,
  read_A_34__ap_start,
  read_A_34__ap_ready,
  read_A_34__ap_done,
  read_A_34__ap_idle,
  read_A_35__ap_start,
  read_A_35__ap_ready,
  read_A_35__ap_done,
  read_A_35__ap_idle,
  read_A_36__ap_start,
  read_A_36__ap_ready,
  read_A_36__ap_done,
  read_A_36__ap_idle,
  read_A_37__ap_start,
  read_A_37__ap_ready,
  read_A_37__ap_done,
  read_A_37__ap_idle,
  read_A_38__ap_start,
  read_A_38__ap_ready,
  read_A_38__ap_done,
  read_A_38__ap_idle,
  read_A_39__ap_start,
  read_A_39__ap_ready,
  read_A_39__ap_done,
  read_A_39__ap_idle,
  read_A_40__ap_start,
  read_A_40__ap_ready,
  read_A_40__ap_done,
  read_A_40__ap_idle,
  read_A_41__ap_start,
  read_A_41__ap_ready,
  read_A_41__ap_done,
  read_A_41__ap_idle,
  read_A_42__ap_start,
  read_A_42__ap_ready,
  read_A_42__ap_done,
  read_A_42__ap_idle,
  read_A_43__ap_start,
  read_A_43__ap_ready,
  read_A_43__ap_done,
  read_A_43__ap_idle,
  read_A_44__ap_start,
  read_A_44__ap_ready,
  read_A_44__ap_done,
  read_A_44__ap_idle,
  read_A_45__ap_start,
  read_A_45__ap_ready,
  read_A_45__ap_done,
  read_A_45__ap_idle,
  read_A_46__ap_start,
  read_A_46__ap_ready,
  read_A_46__ap_done,
  read_A_46__ap_idle,
  read_A_47__ap_start,
  read_A_47__ap_ready,
  read_A_47__ap_done,
  read_A_47__ap_idle,
  read_A_48__ap_start,
  read_A_48__ap_ready,
  read_A_48__ap_done,
  read_A_48__ap_idle,
  read_A_49__ap_start,
  read_A_49__ap_ready,
  read_A_49__ap_done,
  read_A_49__ap_idle,
  read_A_50__ap_start,
  read_A_50__ap_ready,
  read_A_50__ap_done,
  read_A_50__ap_idle,
  read_A_51__ap_start,
  read_A_51__ap_ready,
  read_A_51__ap_done,
  read_A_51__ap_idle,
  read_A_52__ap_start,
  read_A_52__ap_ready,
  read_A_52__ap_done,
  read_A_52__ap_idle,
  read_A_53__ap_start,
  read_A_53__ap_ready,
  read_A_53__ap_done,
  read_A_53__ap_idle,
  read_A_54__ap_start,
  read_A_54__ap_ready,
  read_A_54__ap_done,
  read_A_54__ap_idle,
  read_A_55__ap_start,
  read_A_55__ap_ready,
  read_A_55__ap_done,
  read_A_55__ap_idle,
  read_X_0__ap_start,
  read_X_0__ap_ready,
  read_X_0__ap_done,
  read_X_0__ap_idle,
  read_Y_0__ap_start,
  read_Y_0__ap_ready,
  read_Y_0__ap_done,
  read_Y_0__ap_idle,
  read_edge_list_ptr_0__ap_start,
  read_edge_list_ptr_0__ap_ready,
  read_edge_list_ptr_0__ap_done,
  read_edge_list_ptr_0__ap_idle,
  write_Y_0__ap_start,
  write_Y_0__ap_ready,
  write_Y_0__ap_done,
  write_Y_0__ap_idle
);
  (* RS_CLK *)input ap_clk;
  (* RS_RST = "ff" *)input ap_rst_n;
  (* RS_AP_CTRL = "Serpens.ap_start" *)input ap_start;
  (* RS_AP_CTRL = "Serpens.ap_ready" *)output ap_ready;
  (* RS_FF = "Serpens__ap_done" *)output ap_done;
  (* RS_FF = "Serpens__ap_idle" *)output ap_idle;
  (* RS_AP_CTRL = "Arbiter_Y_0.ap_start" *)output Arbiter_Y_0__ap_start;
  (* RS_AP_CTRL = "Arbiter_Y_0.ap_ready" *)input Arbiter_Y_0__ap_ready;
  (* RS_FF = "Arbiter_Y_0__ap_done" *)input Arbiter_Y_0__ap_done;
  (* RS_FF = "Arbiter_Y_0__ap_idle" *)input Arbiter_Y_0__ap_idle;
  (* RS_AP_CTRL = "Arbiter_Y_1.ap_start" *)output Arbiter_Y_1__ap_start;
  (* RS_AP_CTRL = "Arbiter_Y_1.ap_ready" *)input Arbiter_Y_1__ap_ready;
  (* RS_FF = "Arbiter_Y_1__ap_done" *)input Arbiter_Y_1__ap_done;
  (* RS_FF = "Arbiter_Y_1__ap_idle" *)input Arbiter_Y_1__ap_idle;
  (* RS_AP_CTRL = "Arbiter_Y_2.ap_start" *)output Arbiter_Y_2__ap_start;
  (* RS_AP_CTRL = "Arbiter_Y_2.ap_ready" *)input Arbiter_Y_2__ap_ready;
  (* RS_FF = "Arbiter_Y_2__ap_done" *)input Arbiter_Y_2__ap_done;
  (* RS_FF = "Arbiter_Y_2__ap_idle" *)input Arbiter_Y_2__ap_idle;
  (* RS_AP_CTRL = "Arbiter_Y_3.ap_start" *)output Arbiter_Y_3__ap_start;
  (* RS_AP_CTRL = "Arbiter_Y_3.ap_ready" *)input Arbiter_Y_3__ap_ready;
  (* RS_FF = "Arbiter_Y_3__ap_done" *)input Arbiter_Y_3__ap_done;
  (* RS_FF = "Arbiter_Y_3__ap_idle" *)input Arbiter_Y_3__ap_idle;
  (* RS_AP_CTRL = "Arbiter_Y_4.ap_start" *)output Arbiter_Y_4__ap_start;
  (* RS_AP_CTRL = "Arbiter_Y_4.ap_ready" *)input Arbiter_Y_4__ap_ready;
  (* RS_FF = "Arbiter_Y_4__ap_done" *)input Arbiter_Y_4__ap_done;
  (* RS_FF = "Arbiter_Y_4__ap_idle" *)input Arbiter_Y_4__ap_idle;
  (* RS_AP_CTRL = "Arbiter_Y_5.ap_start" *)output Arbiter_Y_5__ap_start;
  (* RS_AP_CTRL = "Arbiter_Y_5.ap_ready" *)input Arbiter_Y_5__ap_ready;
  (* RS_FF = "Arbiter_Y_5__ap_done" *)input Arbiter_Y_5__ap_done;
  (* RS_FF = "Arbiter_Y_5__ap_idle" *)input Arbiter_Y_5__ap_idle;
  (* RS_AP_CTRL = "Arbiter_Y_6.ap_start" *)output Arbiter_Y_6__ap_start;
  (* RS_AP_CTRL = "Arbiter_Y_6.ap_ready" *)input Arbiter_Y_6__ap_ready;
  (* RS_FF = "Arbiter_Y_6__ap_done" *)input Arbiter_Y_6__ap_done;
  (* RS_FF = "Arbiter_Y_6__ap_idle" *)input Arbiter_Y_6__ap_idle;
  (* RS_AP_CTRL = "Arbiter_Y_7.ap_start" *)output Arbiter_Y_7__ap_start;
  (* RS_AP_CTRL = "Arbiter_Y_7.ap_ready" *)input Arbiter_Y_7__ap_ready;
  (* RS_FF = "Arbiter_Y_7__ap_done" *)input Arbiter_Y_7__ap_done;
  (* RS_FF = "Arbiter_Y_7__ap_idle" *)input Arbiter_Y_7__ap_idle;
  (* RS_FF = "FloatvAddFloatv_0__ap_start" *)output FloatvAddFloatv_0__ap_start;
  (* RS_AP_CTRL = "FloatvMultConst_0.ap_start" *)output FloatvMultConst_0__ap_start;
  (* RS_AP_CTRL = "FloatvMultConst_0.ap_ready" *)input FloatvMultConst_0__ap_ready;
  (* RS_FF = "FloatvMultConst_0__ap_done" *)input FloatvMultConst_0__ap_done;
  (* RS_FF = "FloatvMultConst_0__ap_idle" *)input FloatvMultConst_0__ap_idle;
  (* RS_AP_CTRL = "FloatvMultConst_1.ap_start" *)output FloatvMultConst_1__ap_start;
  (* RS_AP_CTRL = "FloatvMultConst_1.ap_ready" *)input FloatvMultConst_1__ap_ready;
  (* RS_FF = "FloatvMultConst_1__ap_done" *)input FloatvMultConst_1__ap_done;
  (* RS_FF = "FloatvMultConst_1__ap_idle" *)input FloatvMultConst_1__ap_idle;
  (* RS_FF = "Merger_Y_0__ap_start" *)output Merger_Y_0__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_0.ap_start" *)output PEG_Xvec_0__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_0.ap_ready" *)input PEG_Xvec_0__ap_ready;
  (* RS_FF = "PEG_Xvec_0__ap_done" *)input PEG_Xvec_0__ap_done;
  (* RS_FF = "PEG_Xvec_0__ap_idle" *)input PEG_Xvec_0__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_1.ap_start" *)output PEG_Xvec_1__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_1.ap_ready" *)input PEG_Xvec_1__ap_ready;
  (* RS_FF = "PEG_Xvec_1__ap_done" *)input PEG_Xvec_1__ap_done;
  (* RS_FF = "PEG_Xvec_1__ap_idle" *)input PEG_Xvec_1__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_2.ap_start" *)output PEG_Xvec_2__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_2.ap_ready" *)input PEG_Xvec_2__ap_ready;
  (* RS_FF = "PEG_Xvec_2__ap_done" *)input PEG_Xvec_2__ap_done;
  (* RS_FF = "PEG_Xvec_2__ap_idle" *)input PEG_Xvec_2__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_3.ap_start" *)output PEG_Xvec_3__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_3.ap_ready" *)input PEG_Xvec_3__ap_ready;
  (* RS_FF = "PEG_Xvec_3__ap_done" *)input PEG_Xvec_3__ap_done;
  (* RS_FF = "PEG_Xvec_3__ap_idle" *)input PEG_Xvec_3__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_4.ap_start" *)output PEG_Xvec_4__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_4.ap_ready" *)input PEG_Xvec_4__ap_ready;
  (* RS_FF = "PEG_Xvec_4__ap_done" *)input PEG_Xvec_4__ap_done;
  (* RS_FF = "PEG_Xvec_4__ap_idle" *)input PEG_Xvec_4__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_5.ap_start" *)output PEG_Xvec_5__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_5.ap_ready" *)input PEG_Xvec_5__ap_ready;
  (* RS_FF = "PEG_Xvec_5__ap_done" *)input PEG_Xvec_5__ap_done;
  (* RS_FF = "PEG_Xvec_5__ap_idle" *)input PEG_Xvec_5__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_6.ap_start" *)output PEG_Xvec_6__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_6.ap_ready" *)input PEG_Xvec_6__ap_ready;
  (* RS_FF = "PEG_Xvec_6__ap_done" *)input PEG_Xvec_6__ap_done;
  (* RS_FF = "PEG_Xvec_6__ap_idle" *)input PEG_Xvec_6__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_7.ap_start" *)output PEG_Xvec_7__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_7.ap_ready" *)input PEG_Xvec_7__ap_ready;
  (* RS_FF = "PEG_Xvec_7__ap_done" *)input PEG_Xvec_7__ap_done;
  (* RS_FF = "PEG_Xvec_7__ap_idle" *)input PEG_Xvec_7__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_8.ap_start" *)output PEG_Xvec_8__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_8.ap_ready" *)input PEG_Xvec_8__ap_ready;
  (* RS_FF = "PEG_Xvec_8__ap_done" *)input PEG_Xvec_8__ap_done;
  (* RS_FF = "PEG_Xvec_8__ap_idle" *)input PEG_Xvec_8__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_9.ap_start" *)output PEG_Xvec_9__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_9.ap_ready" *)input PEG_Xvec_9__ap_ready;
  (* RS_FF = "PEG_Xvec_9__ap_done" *)input PEG_Xvec_9__ap_done;
  (* RS_FF = "PEG_Xvec_9__ap_idle" *)input PEG_Xvec_9__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_10.ap_start" *)output PEG_Xvec_10__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_10.ap_ready" *)input PEG_Xvec_10__ap_ready;
  (* RS_FF = "PEG_Xvec_10__ap_done" *)input PEG_Xvec_10__ap_done;
  (* RS_FF = "PEG_Xvec_10__ap_idle" *)input PEG_Xvec_10__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_11.ap_start" *)output PEG_Xvec_11__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_11.ap_ready" *)input PEG_Xvec_11__ap_ready;
  (* RS_FF = "PEG_Xvec_11__ap_done" *)input PEG_Xvec_11__ap_done;
  (* RS_FF = "PEG_Xvec_11__ap_idle" *)input PEG_Xvec_11__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_12.ap_start" *)output PEG_Xvec_12__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_12.ap_ready" *)input PEG_Xvec_12__ap_ready;
  (* RS_FF = "PEG_Xvec_12__ap_done" *)input PEG_Xvec_12__ap_done;
  (* RS_FF = "PEG_Xvec_12__ap_idle" *)input PEG_Xvec_12__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_13.ap_start" *)output PEG_Xvec_13__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_13.ap_ready" *)input PEG_Xvec_13__ap_ready;
  (* RS_FF = "PEG_Xvec_13__ap_done" *)input PEG_Xvec_13__ap_done;
  (* RS_FF = "PEG_Xvec_13__ap_idle" *)input PEG_Xvec_13__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_14.ap_start" *)output PEG_Xvec_14__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_14.ap_ready" *)input PEG_Xvec_14__ap_ready;
  (* RS_FF = "PEG_Xvec_14__ap_done" *)input PEG_Xvec_14__ap_done;
  (* RS_FF = "PEG_Xvec_14__ap_idle" *)input PEG_Xvec_14__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_15.ap_start" *)output PEG_Xvec_15__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_15.ap_ready" *)input PEG_Xvec_15__ap_ready;
  (* RS_FF = "PEG_Xvec_15__ap_done" *)input PEG_Xvec_15__ap_done;
  (* RS_FF = "PEG_Xvec_15__ap_idle" *)input PEG_Xvec_15__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_16.ap_start" *)output PEG_Xvec_16__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_16.ap_ready" *)input PEG_Xvec_16__ap_ready;
  (* RS_FF = "PEG_Xvec_16__ap_done" *)input PEG_Xvec_16__ap_done;
  (* RS_FF = "PEG_Xvec_16__ap_idle" *)input PEG_Xvec_16__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_17.ap_start" *)output PEG_Xvec_17__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_17.ap_ready" *)input PEG_Xvec_17__ap_ready;
  (* RS_FF = "PEG_Xvec_17__ap_done" *)input PEG_Xvec_17__ap_done;
  (* RS_FF = "PEG_Xvec_17__ap_idle" *)input PEG_Xvec_17__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_18.ap_start" *)output PEG_Xvec_18__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_18.ap_ready" *)input PEG_Xvec_18__ap_ready;
  (* RS_FF = "PEG_Xvec_18__ap_done" *)input PEG_Xvec_18__ap_done;
  (* RS_FF = "PEG_Xvec_18__ap_idle" *)input PEG_Xvec_18__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_19.ap_start" *)output PEG_Xvec_19__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_19.ap_ready" *)input PEG_Xvec_19__ap_ready;
  (* RS_FF = "PEG_Xvec_19__ap_done" *)input PEG_Xvec_19__ap_done;
  (* RS_FF = "PEG_Xvec_19__ap_idle" *)input PEG_Xvec_19__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_20.ap_start" *)output PEG_Xvec_20__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_20.ap_ready" *)input PEG_Xvec_20__ap_ready;
  (* RS_FF = "PEG_Xvec_20__ap_done" *)input PEG_Xvec_20__ap_done;
  (* RS_FF = "PEG_Xvec_20__ap_idle" *)input PEG_Xvec_20__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_21.ap_start" *)output PEG_Xvec_21__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_21.ap_ready" *)input PEG_Xvec_21__ap_ready;
  (* RS_FF = "PEG_Xvec_21__ap_done" *)input PEG_Xvec_21__ap_done;
  (* RS_FF = "PEG_Xvec_21__ap_idle" *)input PEG_Xvec_21__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_22.ap_start" *)output PEG_Xvec_22__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_22.ap_ready" *)input PEG_Xvec_22__ap_ready;
  (* RS_FF = "PEG_Xvec_22__ap_done" *)input PEG_Xvec_22__ap_done;
  (* RS_FF = "PEG_Xvec_22__ap_idle" *)input PEG_Xvec_22__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_23.ap_start" *)output PEG_Xvec_23__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_23.ap_ready" *)input PEG_Xvec_23__ap_ready;
  (* RS_FF = "PEG_Xvec_23__ap_done" *)input PEG_Xvec_23__ap_done;
  (* RS_FF = "PEG_Xvec_23__ap_idle" *)input PEG_Xvec_23__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_24.ap_start" *)output PEG_Xvec_24__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_24.ap_ready" *)input PEG_Xvec_24__ap_ready;
  (* RS_FF = "PEG_Xvec_24__ap_done" *)input PEG_Xvec_24__ap_done;
  (* RS_FF = "PEG_Xvec_24__ap_idle" *)input PEG_Xvec_24__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_25.ap_start" *)output PEG_Xvec_25__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_25.ap_ready" *)input PEG_Xvec_25__ap_ready;
  (* RS_FF = "PEG_Xvec_25__ap_done" *)input PEG_Xvec_25__ap_done;
  (* RS_FF = "PEG_Xvec_25__ap_idle" *)input PEG_Xvec_25__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_26.ap_start" *)output PEG_Xvec_26__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_26.ap_ready" *)input PEG_Xvec_26__ap_ready;
  (* RS_FF = "PEG_Xvec_26__ap_done" *)input PEG_Xvec_26__ap_done;
  (* RS_FF = "PEG_Xvec_26__ap_idle" *)input PEG_Xvec_26__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_27.ap_start" *)output PEG_Xvec_27__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_27.ap_ready" *)input PEG_Xvec_27__ap_ready;
  (* RS_FF = "PEG_Xvec_27__ap_done" *)input PEG_Xvec_27__ap_done;
  (* RS_FF = "PEG_Xvec_27__ap_idle" *)input PEG_Xvec_27__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_28.ap_start" *)output PEG_Xvec_28__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_28.ap_ready" *)input PEG_Xvec_28__ap_ready;
  (* RS_FF = "PEG_Xvec_28__ap_done" *)input PEG_Xvec_28__ap_done;
  (* RS_FF = "PEG_Xvec_28__ap_idle" *)input PEG_Xvec_28__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_29.ap_start" *)output PEG_Xvec_29__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_29.ap_ready" *)input PEG_Xvec_29__ap_ready;
  (* RS_FF = "PEG_Xvec_29__ap_done" *)input PEG_Xvec_29__ap_done;
  (* RS_FF = "PEG_Xvec_29__ap_idle" *)input PEG_Xvec_29__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_30.ap_start" *)output PEG_Xvec_30__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_30.ap_ready" *)input PEG_Xvec_30__ap_ready;
  (* RS_FF = "PEG_Xvec_30__ap_done" *)input PEG_Xvec_30__ap_done;
  (* RS_FF = "PEG_Xvec_30__ap_idle" *)input PEG_Xvec_30__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_31.ap_start" *)output PEG_Xvec_31__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_31.ap_ready" *)input PEG_Xvec_31__ap_ready;
  (* RS_FF = "PEG_Xvec_31__ap_done" *)input PEG_Xvec_31__ap_done;
  (* RS_FF = "PEG_Xvec_31__ap_idle" *)input PEG_Xvec_31__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_32.ap_start" *)output PEG_Xvec_32__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_32.ap_ready" *)input PEG_Xvec_32__ap_ready;
  (* RS_FF = "PEG_Xvec_32__ap_done" *)input PEG_Xvec_32__ap_done;
  (* RS_FF = "PEG_Xvec_32__ap_idle" *)input PEG_Xvec_32__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_33.ap_start" *)output PEG_Xvec_33__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_33.ap_ready" *)input PEG_Xvec_33__ap_ready;
  (* RS_FF = "PEG_Xvec_33__ap_done" *)input PEG_Xvec_33__ap_done;
  (* RS_FF = "PEG_Xvec_33__ap_idle" *)input PEG_Xvec_33__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_34.ap_start" *)output PEG_Xvec_34__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_34.ap_ready" *)input PEG_Xvec_34__ap_ready;
  (* RS_FF = "PEG_Xvec_34__ap_done" *)input PEG_Xvec_34__ap_done;
  (* RS_FF = "PEG_Xvec_34__ap_idle" *)input PEG_Xvec_34__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_35.ap_start" *)output PEG_Xvec_35__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_35.ap_ready" *)input PEG_Xvec_35__ap_ready;
  (* RS_FF = "PEG_Xvec_35__ap_done" *)input PEG_Xvec_35__ap_done;
  (* RS_FF = "PEG_Xvec_35__ap_idle" *)input PEG_Xvec_35__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_36.ap_start" *)output PEG_Xvec_36__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_36.ap_ready" *)input PEG_Xvec_36__ap_ready;
  (* RS_FF = "PEG_Xvec_36__ap_done" *)input PEG_Xvec_36__ap_done;
  (* RS_FF = "PEG_Xvec_36__ap_idle" *)input PEG_Xvec_36__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_37.ap_start" *)output PEG_Xvec_37__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_37.ap_ready" *)input PEG_Xvec_37__ap_ready;
  (* RS_FF = "PEG_Xvec_37__ap_done" *)input PEG_Xvec_37__ap_done;
  (* RS_FF = "PEG_Xvec_37__ap_idle" *)input PEG_Xvec_37__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_38.ap_start" *)output PEG_Xvec_38__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_38.ap_ready" *)input PEG_Xvec_38__ap_ready;
  (* RS_FF = "PEG_Xvec_38__ap_done" *)input PEG_Xvec_38__ap_done;
  (* RS_FF = "PEG_Xvec_38__ap_idle" *)input PEG_Xvec_38__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_39.ap_start" *)output PEG_Xvec_39__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_39.ap_ready" *)input PEG_Xvec_39__ap_ready;
  (* RS_FF = "PEG_Xvec_39__ap_done" *)input PEG_Xvec_39__ap_done;
  (* RS_FF = "PEG_Xvec_39__ap_idle" *)input PEG_Xvec_39__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_40.ap_start" *)output PEG_Xvec_40__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_40.ap_ready" *)input PEG_Xvec_40__ap_ready;
  (* RS_FF = "PEG_Xvec_40__ap_done" *)input PEG_Xvec_40__ap_done;
  (* RS_FF = "PEG_Xvec_40__ap_idle" *)input PEG_Xvec_40__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_41.ap_start" *)output PEG_Xvec_41__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_41.ap_ready" *)input PEG_Xvec_41__ap_ready;
  (* RS_FF = "PEG_Xvec_41__ap_done" *)input PEG_Xvec_41__ap_done;
  (* RS_FF = "PEG_Xvec_41__ap_idle" *)input PEG_Xvec_41__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_42.ap_start" *)output PEG_Xvec_42__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_42.ap_ready" *)input PEG_Xvec_42__ap_ready;
  (* RS_FF = "PEG_Xvec_42__ap_done" *)input PEG_Xvec_42__ap_done;
  (* RS_FF = "PEG_Xvec_42__ap_idle" *)input PEG_Xvec_42__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_43.ap_start" *)output PEG_Xvec_43__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_43.ap_ready" *)input PEG_Xvec_43__ap_ready;
  (* RS_FF = "PEG_Xvec_43__ap_done" *)input PEG_Xvec_43__ap_done;
  (* RS_FF = "PEG_Xvec_43__ap_idle" *)input PEG_Xvec_43__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_44.ap_start" *)output PEG_Xvec_44__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_44.ap_ready" *)input PEG_Xvec_44__ap_ready;
  (* RS_FF = "PEG_Xvec_44__ap_done" *)input PEG_Xvec_44__ap_done;
  (* RS_FF = "PEG_Xvec_44__ap_idle" *)input PEG_Xvec_44__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_45.ap_start" *)output PEG_Xvec_45__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_45.ap_ready" *)input PEG_Xvec_45__ap_ready;
  (* RS_FF = "PEG_Xvec_45__ap_done" *)input PEG_Xvec_45__ap_done;
  (* RS_FF = "PEG_Xvec_45__ap_idle" *)input PEG_Xvec_45__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_46.ap_start" *)output PEG_Xvec_46__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_46.ap_ready" *)input PEG_Xvec_46__ap_ready;
  (* RS_FF = "PEG_Xvec_46__ap_done" *)input PEG_Xvec_46__ap_done;
  (* RS_FF = "PEG_Xvec_46__ap_idle" *)input PEG_Xvec_46__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_47.ap_start" *)output PEG_Xvec_47__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_47.ap_ready" *)input PEG_Xvec_47__ap_ready;
  (* RS_FF = "PEG_Xvec_47__ap_done" *)input PEG_Xvec_47__ap_done;
  (* RS_FF = "PEG_Xvec_47__ap_idle" *)input PEG_Xvec_47__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_48.ap_start" *)output PEG_Xvec_48__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_48.ap_ready" *)input PEG_Xvec_48__ap_ready;
  (* RS_FF = "PEG_Xvec_48__ap_done" *)input PEG_Xvec_48__ap_done;
  (* RS_FF = "PEG_Xvec_48__ap_idle" *)input PEG_Xvec_48__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_49.ap_start" *)output PEG_Xvec_49__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_49.ap_ready" *)input PEG_Xvec_49__ap_ready;
  (* RS_FF = "PEG_Xvec_49__ap_done" *)input PEG_Xvec_49__ap_done;
  (* RS_FF = "PEG_Xvec_49__ap_idle" *)input PEG_Xvec_49__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_50.ap_start" *)output PEG_Xvec_50__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_50.ap_ready" *)input PEG_Xvec_50__ap_ready;
  (* RS_FF = "PEG_Xvec_50__ap_done" *)input PEG_Xvec_50__ap_done;
  (* RS_FF = "PEG_Xvec_50__ap_idle" *)input PEG_Xvec_50__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_51.ap_start" *)output PEG_Xvec_51__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_51.ap_ready" *)input PEG_Xvec_51__ap_ready;
  (* RS_FF = "PEG_Xvec_51__ap_done" *)input PEG_Xvec_51__ap_done;
  (* RS_FF = "PEG_Xvec_51__ap_idle" *)input PEG_Xvec_51__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_52.ap_start" *)output PEG_Xvec_52__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_52.ap_ready" *)input PEG_Xvec_52__ap_ready;
  (* RS_FF = "PEG_Xvec_52__ap_done" *)input PEG_Xvec_52__ap_done;
  (* RS_FF = "PEG_Xvec_52__ap_idle" *)input PEG_Xvec_52__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_53.ap_start" *)output PEG_Xvec_53__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_53.ap_ready" *)input PEG_Xvec_53__ap_ready;
  (* RS_FF = "PEG_Xvec_53__ap_done" *)input PEG_Xvec_53__ap_done;
  (* RS_FF = "PEG_Xvec_53__ap_idle" *)input PEG_Xvec_53__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_54.ap_start" *)output PEG_Xvec_54__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_54.ap_ready" *)input PEG_Xvec_54__ap_ready;
  (* RS_FF = "PEG_Xvec_54__ap_done" *)input PEG_Xvec_54__ap_done;
  (* RS_FF = "PEG_Xvec_54__ap_idle" *)input PEG_Xvec_54__ap_idle;
  (* RS_AP_CTRL = "PEG_Xvec_55.ap_start" *)output PEG_Xvec_55__ap_start;
  (* RS_AP_CTRL = "PEG_Xvec_55.ap_ready" *)input PEG_Xvec_55__ap_ready;
  (* RS_FF = "PEG_Xvec_55__ap_done" *)input PEG_Xvec_55__ap_done;
  (* RS_FF = "PEG_Xvec_55__ap_idle" *)input PEG_Xvec_55__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_0.ap_start" *)output PEG_Yvec_0__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_0.ap_ready" *)input PEG_Yvec_0__ap_ready;
  (* RS_FF = "PEG_Yvec_0__ap_done" *)input PEG_Yvec_0__ap_done;
  (* RS_FF = "PEG_Yvec_0__ap_idle" *)input PEG_Yvec_0__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_1.ap_start" *)output PEG_Yvec_1__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_1.ap_ready" *)input PEG_Yvec_1__ap_ready;
  (* RS_FF = "PEG_Yvec_1__ap_done" *)input PEG_Yvec_1__ap_done;
  (* RS_FF = "PEG_Yvec_1__ap_idle" *)input PEG_Yvec_1__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_2.ap_start" *)output PEG_Yvec_2__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_2.ap_ready" *)input PEG_Yvec_2__ap_ready;
  (* RS_FF = "PEG_Yvec_2__ap_done" *)input PEG_Yvec_2__ap_done;
  (* RS_FF = "PEG_Yvec_2__ap_idle" *)input PEG_Yvec_2__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_3.ap_start" *)output PEG_Yvec_3__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_3.ap_ready" *)input PEG_Yvec_3__ap_ready;
  (* RS_FF = "PEG_Yvec_3__ap_done" *)input PEG_Yvec_3__ap_done;
  (* RS_FF = "PEG_Yvec_3__ap_idle" *)input PEG_Yvec_3__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_4.ap_start" *)output PEG_Yvec_4__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_4.ap_ready" *)input PEG_Yvec_4__ap_ready;
  (* RS_FF = "PEG_Yvec_4__ap_done" *)input PEG_Yvec_4__ap_done;
  (* RS_FF = "PEG_Yvec_4__ap_idle" *)input PEG_Yvec_4__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_5.ap_start" *)output PEG_Yvec_5__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_5.ap_ready" *)input PEG_Yvec_5__ap_ready;
  (* RS_FF = "PEG_Yvec_5__ap_done" *)input PEG_Yvec_5__ap_done;
  (* RS_FF = "PEG_Yvec_5__ap_idle" *)input PEG_Yvec_5__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_6.ap_start" *)output PEG_Yvec_6__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_6.ap_ready" *)input PEG_Yvec_6__ap_ready;
  (* RS_FF = "PEG_Yvec_6__ap_done" *)input PEG_Yvec_6__ap_done;
  (* RS_FF = "PEG_Yvec_6__ap_idle" *)input PEG_Yvec_6__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_7.ap_start" *)output PEG_Yvec_7__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_7.ap_ready" *)input PEG_Yvec_7__ap_ready;
  (* RS_FF = "PEG_Yvec_7__ap_done" *)input PEG_Yvec_7__ap_done;
  (* RS_FF = "PEG_Yvec_7__ap_idle" *)input PEG_Yvec_7__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_8.ap_start" *)output PEG_Yvec_8__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_8.ap_ready" *)input PEG_Yvec_8__ap_ready;
  (* RS_FF = "PEG_Yvec_8__ap_done" *)input PEG_Yvec_8__ap_done;
  (* RS_FF = "PEG_Yvec_8__ap_idle" *)input PEG_Yvec_8__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_9.ap_start" *)output PEG_Yvec_9__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_9.ap_ready" *)input PEG_Yvec_9__ap_ready;
  (* RS_FF = "PEG_Yvec_9__ap_done" *)input PEG_Yvec_9__ap_done;
  (* RS_FF = "PEG_Yvec_9__ap_idle" *)input PEG_Yvec_9__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_10.ap_start" *)output PEG_Yvec_10__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_10.ap_ready" *)input PEG_Yvec_10__ap_ready;
  (* RS_FF = "PEG_Yvec_10__ap_done" *)input PEG_Yvec_10__ap_done;
  (* RS_FF = "PEG_Yvec_10__ap_idle" *)input PEG_Yvec_10__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_11.ap_start" *)output PEG_Yvec_11__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_11.ap_ready" *)input PEG_Yvec_11__ap_ready;
  (* RS_FF = "PEG_Yvec_11__ap_done" *)input PEG_Yvec_11__ap_done;
  (* RS_FF = "PEG_Yvec_11__ap_idle" *)input PEG_Yvec_11__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_12.ap_start" *)output PEG_Yvec_12__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_12.ap_ready" *)input PEG_Yvec_12__ap_ready;
  (* RS_FF = "PEG_Yvec_12__ap_done" *)input PEG_Yvec_12__ap_done;
  (* RS_FF = "PEG_Yvec_12__ap_idle" *)input PEG_Yvec_12__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_13.ap_start" *)output PEG_Yvec_13__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_13.ap_ready" *)input PEG_Yvec_13__ap_ready;
  (* RS_FF = "PEG_Yvec_13__ap_done" *)input PEG_Yvec_13__ap_done;
  (* RS_FF = "PEG_Yvec_13__ap_idle" *)input PEG_Yvec_13__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_14.ap_start" *)output PEG_Yvec_14__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_14.ap_ready" *)input PEG_Yvec_14__ap_ready;
  (* RS_FF = "PEG_Yvec_14__ap_done" *)input PEG_Yvec_14__ap_done;
  (* RS_FF = "PEG_Yvec_14__ap_idle" *)input PEG_Yvec_14__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_15.ap_start" *)output PEG_Yvec_15__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_15.ap_ready" *)input PEG_Yvec_15__ap_ready;
  (* RS_FF = "PEG_Yvec_15__ap_done" *)input PEG_Yvec_15__ap_done;
  (* RS_FF = "PEG_Yvec_15__ap_idle" *)input PEG_Yvec_15__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_16.ap_start" *)output PEG_Yvec_16__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_16.ap_ready" *)input PEG_Yvec_16__ap_ready;
  (* RS_FF = "PEG_Yvec_16__ap_done" *)input PEG_Yvec_16__ap_done;
  (* RS_FF = "PEG_Yvec_16__ap_idle" *)input PEG_Yvec_16__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_17.ap_start" *)output PEG_Yvec_17__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_17.ap_ready" *)input PEG_Yvec_17__ap_ready;
  (* RS_FF = "PEG_Yvec_17__ap_done" *)input PEG_Yvec_17__ap_done;
  (* RS_FF = "PEG_Yvec_17__ap_idle" *)input PEG_Yvec_17__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_18.ap_start" *)output PEG_Yvec_18__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_18.ap_ready" *)input PEG_Yvec_18__ap_ready;
  (* RS_FF = "PEG_Yvec_18__ap_done" *)input PEG_Yvec_18__ap_done;
  (* RS_FF = "PEG_Yvec_18__ap_idle" *)input PEG_Yvec_18__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_19.ap_start" *)output PEG_Yvec_19__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_19.ap_ready" *)input PEG_Yvec_19__ap_ready;
  (* RS_FF = "PEG_Yvec_19__ap_done" *)input PEG_Yvec_19__ap_done;
  (* RS_FF = "PEG_Yvec_19__ap_idle" *)input PEG_Yvec_19__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_20.ap_start" *)output PEG_Yvec_20__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_20.ap_ready" *)input PEG_Yvec_20__ap_ready;
  (* RS_FF = "PEG_Yvec_20__ap_done" *)input PEG_Yvec_20__ap_done;
  (* RS_FF = "PEG_Yvec_20__ap_idle" *)input PEG_Yvec_20__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_21.ap_start" *)output PEG_Yvec_21__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_21.ap_ready" *)input PEG_Yvec_21__ap_ready;
  (* RS_FF = "PEG_Yvec_21__ap_done" *)input PEG_Yvec_21__ap_done;
  (* RS_FF = "PEG_Yvec_21__ap_idle" *)input PEG_Yvec_21__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_22.ap_start" *)output PEG_Yvec_22__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_22.ap_ready" *)input PEG_Yvec_22__ap_ready;
  (* RS_FF = "PEG_Yvec_22__ap_done" *)input PEG_Yvec_22__ap_done;
  (* RS_FF = "PEG_Yvec_22__ap_idle" *)input PEG_Yvec_22__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_23.ap_start" *)output PEG_Yvec_23__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_23.ap_ready" *)input PEG_Yvec_23__ap_ready;
  (* RS_FF = "PEG_Yvec_23__ap_done" *)input PEG_Yvec_23__ap_done;
  (* RS_FF = "PEG_Yvec_23__ap_idle" *)input PEG_Yvec_23__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_24.ap_start" *)output PEG_Yvec_24__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_24.ap_ready" *)input PEG_Yvec_24__ap_ready;
  (* RS_FF = "PEG_Yvec_24__ap_done" *)input PEG_Yvec_24__ap_done;
  (* RS_FF = "PEG_Yvec_24__ap_idle" *)input PEG_Yvec_24__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_25.ap_start" *)output PEG_Yvec_25__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_25.ap_ready" *)input PEG_Yvec_25__ap_ready;
  (* RS_FF = "PEG_Yvec_25__ap_done" *)input PEG_Yvec_25__ap_done;
  (* RS_FF = "PEG_Yvec_25__ap_idle" *)input PEG_Yvec_25__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_26.ap_start" *)output PEG_Yvec_26__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_26.ap_ready" *)input PEG_Yvec_26__ap_ready;
  (* RS_FF = "PEG_Yvec_26__ap_done" *)input PEG_Yvec_26__ap_done;
  (* RS_FF = "PEG_Yvec_26__ap_idle" *)input PEG_Yvec_26__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_27.ap_start" *)output PEG_Yvec_27__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_27.ap_ready" *)input PEG_Yvec_27__ap_ready;
  (* RS_FF = "PEG_Yvec_27__ap_done" *)input PEG_Yvec_27__ap_done;
  (* RS_FF = "PEG_Yvec_27__ap_idle" *)input PEG_Yvec_27__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_28.ap_start" *)output PEG_Yvec_28__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_28.ap_ready" *)input PEG_Yvec_28__ap_ready;
  (* RS_FF = "PEG_Yvec_28__ap_done" *)input PEG_Yvec_28__ap_done;
  (* RS_FF = "PEG_Yvec_28__ap_idle" *)input PEG_Yvec_28__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_29.ap_start" *)output PEG_Yvec_29__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_29.ap_ready" *)input PEG_Yvec_29__ap_ready;
  (* RS_FF = "PEG_Yvec_29__ap_done" *)input PEG_Yvec_29__ap_done;
  (* RS_FF = "PEG_Yvec_29__ap_idle" *)input PEG_Yvec_29__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_30.ap_start" *)output PEG_Yvec_30__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_30.ap_ready" *)input PEG_Yvec_30__ap_ready;
  (* RS_FF = "PEG_Yvec_30__ap_done" *)input PEG_Yvec_30__ap_done;
  (* RS_FF = "PEG_Yvec_30__ap_idle" *)input PEG_Yvec_30__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_31.ap_start" *)output PEG_Yvec_31__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_31.ap_ready" *)input PEG_Yvec_31__ap_ready;
  (* RS_FF = "PEG_Yvec_31__ap_done" *)input PEG_Yvec_31__ap_done;
  (* RS_FF = "PEG_Yvec_31__ap_idle" *)input PEG_Yvec_31__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_32.ap_start" *)output PEG_Yvec_32__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_32.ap_ready" *)input PEG_Yvec_32__ap_ready;
  (* RS_FF = "PEG_Yvec_32__ap_done" *)input PEG_Yvec_32__ap_done;
  (* RS_FF = "PEG_Yvec_32__ap_idle" *)input PEG_Yvec_32__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_33.ap_start" *)output PEG_Yvec_33__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_33.ap_ready" *)input PEG_Yvec_33__ap_ready;
  (* RS_FF = "PEG_Yvec_33__ap_done" *)input PEG_Yvec_33__ap_done;
  (* RS_FF = "PEG_Yvec_33__ap_idle" *)input PEG_Yvec_33__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_34.ap_start" *)output PEG_Yvec_34__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_34.ap_ready" *)input PEG_Yvec_34__ap_ready;
  (* RS_FF = "PEG_Yvec_34__ap_done" *)input PEG_Yvec_34__ap_done;
  (* RS_FF = "PEG_Yvec_34__ap_idle" *)input PEG_Yvec_34__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_35.ap_start" *)output PEG_Yvec_35__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_35.ap_ready" *)input PEG_Yvec_35__ap_ready;
  (* RS_FF = "PEG_Yvec_35__ap_done" *)input PEG_Yvec_35__ap_done;
  (* RS_FF = "PEG_Yvec_35__ap_idle" *)input PEG_Yvec_35__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_36.ap_start" *)output PEG_Yvec_36__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_36.ap_ready" *)input PEG_Yvec_36__ap_ready;
  (* RS_FF = "PEG_Yvec_36__ap_done" *)input PEG_Yvec_36__ap_done;
  (* RS_FF = "PEG_Yvec_36__ap_idle" *)input PEG_Yvec_36__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_37.ap_start" *)output PEG_Yvec_37__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_37.ap_ready" *)input PEG_Yvec_37__ap_ready;
  (* RS_FF = "PEG_Yvec_37__ap_done" *)input PEG_Yvec_37__ap_done;
  (* RS_FF = "PEG_Yvec_37__ap_idle" *)input PEG_Yvec_37__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_38.ap_start" *)output PEG_Yvec_38__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_38.ap_ready" *)input PEG_Yvec_38__ap_ready;
  (* RS_FF = "PEG_Yvec_38__ap_done" *)input PEG_Yvec_38__ap_done;
  (* RS_FF = "PEG_Yvec_38__ap_idle" *)input PEG_Yvec_38__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_39.ap_start" *)output PEG_Yvec_39__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_39.ap_ready" *)input PEG_Yvec_39__ap_ready;
  (* RS_FF = "PEG_Yvec_39__ap_done" *)input PEG_Yvec_39__ap_done;
  (* RS_FF = "PEG_Yvec_39__ap_idle" *)input PEG_Yvec_39__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_40.ap_start" *)output PEG_Yvec_40__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_40.ap_ready" *)input PEG_Yvec_40__ap_ready;
  (* RS_FF = "PEG_Yvec_40__ap_done" *)input PEG_Yvec_40__ap_done;
  (* RS_FF = "PEG_Yvec_40__ap_idle" *)input PEG_Yvec_40__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_41.ap_start" *)output PEG_Yvec_41__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_41.ap_ready" *)input PEG_Yvec_41__ap_ready;
  (* RS_FF = "PEG_Yvec_41__ap_done" *)input PEG_Yvec_41__ap_done;
  (* RS_FF = "PEG_Yvec_41__ap_idle" *)input PEG_Yvec_41__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_42.ap_start" *)output PEG_Yvec_42__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_42.ap_ready" *)input PEG_Yvec_42__ap_ready;
  (* RS_FF = "PEG_Yvec_42__ap_done" *)input PEG_Yvec_42__ap_done;
  (* RS_FF = "PEG_Yvec_42__ap_idle" *)input PEG_Yvec_42__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_43.ap_start" *)output PEG_Yvec_43__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_43.ap_ready" *)input PEG_Yvec_43__ap_ready;
  (* RS_FF = "PEG_Yvec_43__ap_done" *)input PEG_Yvec_43__ap_done;
  (* RS_FF = "PEG_Yvec_43__ap_idle" *)input PEG_Yvec_43__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_44.ap_start" *)output PEG_Yvec_44__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_44.ap_ready" *)input PEG_Yvec_44__ap_ready;
  (* RS_FF = "PEG_Yvec_44__ap_done" *)input PEG_Yvec_44__ap_done;
  (* RS_FF = "PEG_Yvec_44__ap_idle" *)input PEG_Yvec_44__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_45.ap_start" *)output PEG_Yvec_45__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_45.ap_ready" *)input PEG_Yvec_45__ap_ready;
  (* RS_FF = "PEG_Yvec_45__ap_done" *)input PEG_Yvec_45__ap_done;
  (* RS_FF = "PEG_Yvec_45__ap_idle" *)input PEG_Yvec_45__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_46.ap_start" *)output PEG_Yvec_46__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_46.ap_ready" *)input PEG_Yvec_46__ap_ready;
  (* RS_FF = "PEG_Yvec_46__ap_done" *)input PEG_Yvec_46__ap_done;
  (* RS_FF = "PEG_Yvec_46__ap_idle" *)input PEG_Yvec_46__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_47.ap_start" *)output PEG_Yvec_47__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_47.ap_ready" *)input PEG_Yvec_47__ap_ready;
  (* RS_FF = "PEG_Yvec_47__ap_done" *)input PEG_Yvec_47__ap_done;
  (* RS_FF = "PEG_Yvec_47__ap_idle" *)input PEG_Yvec_47__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_48.ap_start" *)output PEG_Yvec_48__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_48.ap_ready" *)input PEG_Yvec_48__ap_ready;
  (* RS_FF = "PEG_Yvec_48__ap_done" *)input PEG_Yvec_48__ap_done;
  (* RS_FF = "PEG_Yvec_48__ap_idle" *)input PEG_Yvec_48__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_49.ap_start" *)output PEG_Yvec_49__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_49.ap_ready" *)input PEG_Yvec_49__ap_ready;
  (* RS_FF = "PEG_Yvec_49__ap_done" *)input PEG_Yvec_49__ap_done;
  (* RS_FF = "PEG_Yvec_49__ap_idle" *)input PEG_Yvec_49__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_50.ap_start" *)output PEG_Yvec_50__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_50.ap_ready" *)input PEG_Yvec_50__ap_ready;
  (* RS_FF = "PEG_Yvec_50__ap_done" *)input PEG_Yvec_50__ap_done;
  (* RS_FF = "PEG_Yvec_50__ap_idle" *)input PEG_Yvec_50__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_51.ap_start" *)output PEG_Yvec_51__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_51.ap_ready" *)input PEG_Yvec_51__ap_ready;
  (* RS_FF = "PEG_Yvec_51__ap_done" *)input PEG_Yvec_51__ap_done;
  (* RS_FF = "PEG_Yvec_51__ap_idle" *)input PEG_Yvec_51__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_52.ap_start" *)output PEG_Yvec_52__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_52.ap_ready" *)input PEG_Yvec_52__ap_ready;
  (* RS_FF = "PEG_Yvec_52__ap_done" *)input PEG_Yvec_52__ap_done;
  (* RS_FF = "PEG_Yvec_52__ap_idle" *)input PEG_Yvec_52__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_53.ap_start" *)output PEG_Yvec_53__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_53.ap_ready" *)input PEG_Yvec_53__ap_ready;
  (* RS_FF = "PEG_Yvec_53__ap_done" *)input PEG_Yvec_53__ap_done;
  (* RS_FF = "PEG_Yvec_53__ap_idle" *)input PEG_Yvec_53__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_54.ap_start" *)output PEG_Yvec_54__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_54.ap_ready" *)input PEG_Yvec_54__ap_ready;
  (* RS_FF = "PEG_Yvec_54__ap_done" *)input PEG_Yvec_54__ap_done;
  (* RS_FF = "PEG_Yvec_54__ap_idle" *)input PEG_Yvec_54__ap_idle;
  (* RS_AP_CTRL = "PEG_Yvec_55.ap_start" *)output PEG_Yvec_55__ap_start;
  (* RS_AP_CTRL = "PEG_Yvec_55.ap_ready" *)input PEG_Yvec_55__ap_ready;
  (* RS_FF = "PEG_Yvec_55__ap_done" *)input PEG_Yvec_55__ap_done;
  (* RS_FF = "PEG_Yvec_55__ap_idle" *)input PEG_Yvec_55__ap_idle;
  (* RS_FF = "black_hole_float_v16_0__ap_start" *)output black_hole_float_v16_0__ap_start;
  (* RS_FF = "black_hole_int_0__ap_start" *)output black_hole_int_0__ap_start;
  (* RS_AP_CTRL = "read_A_0.ap_start" *)output read_A_0__ap_start;
  (* RS_AP_CTRL = "read_A_0.ap_ready" *)input read_A_0__ap_ready;
  (* RS_FF = "read_A_0__ap_done" *)input read_A_0__ap_done;
  (* RS_FF = "read_A_0__ap_idle" *)input read_A_0__ap_idle;
  (* RS_AP_CTRL = "read_A_1.ap_start" *)output read_A_1__ap_start;
  (* RS_AP_CTRL = "read_A_1.ap_ready" *)input read_A_1__ap_ready;
  (* RS_FF = "read_A_1__ap_done" *)input read_A_1__ap_done;
  (* RS_FF = "read_A_1__ap_idle" *)input read_A_1__ap_idle;
  (* RS_AP_CTRL = "read_A_2.ap_start" *)output read_A_2__ap_start;
  (* RS_AP_CTRL = "read_A_2.ap_ready" *)input read_A_2__ap_ready;
  (* RS_FF = "read_A_2__ap_done" *)input read_A_2__ap_done;
  (* RS_FF = "read_A_2__ap_idle" *)input read_A_2__ap_idle;
  (* RS_AP_CTRL = "read_A_3.ap_start" *)output read_A_3__ap_start;
  (* RS_AP_CTRL = "read_A_3.ap_ready" *)input read_A_3__ap_ready;
  (* RS_FF = "read_A_3__ap_done" *)input read_A_3__ap_done;
  (* RS_FF = "read_A_3__ap_idle" *)input read_A_3__ap_idle;
  (* RS_AP_CTRL = "read_A_4.ap_start" *)output read_A_4__ap_start;
  (* RS_AP_CTRL = "read_A_4.ap_ready" *)input read_A_4__ap_ready;
  (* RS_FF = "read_A_4__ap_done" *)input read_A_4__ap_done;
  (* RS_FF = "read_A_4__ap_idle" *)input read_A_4__ap_idle;
  (* RS_AP_CTRL = "read_A_5.ap_start" *)output read_A_5__ap_start;
  (* RS_AP_CTRL = "read_A_5.ap_ready" *)input read_A_5__ap_ready;
  (* RS_FF = "read_A_5__ap_done" *)input read_A_5__ap_done;
  (* RS_FF = "read_A_5__ap_idle" *)input read_A_5__ap_idle;
  (* RS_AP_CTRL = "read_A_6.ap_start" *)output read_A_6__ap_start;
  (* RS_AP_CTRL = "read_A_6.ap_ready" *)input read_A_6__ap_ready;
  (* RS_FF = "read_A_6__ap_done" *)input read_A_6__ap_done;
  (* RS_FF = "read_A_6__ap_idle" *)input read_A_6__ap_idle;
  (* RS_AP_CTRL = "read_A_7.ap_start" *)output read_A_7__ap_start;
  (* RS_AP_CTRL = "read_A_7.ap_ready" *)input read_A_7__ap_ready;
  (* RS_FF = "read_A_7__ap_done" *)input read_A_7__ap_done;
  (* RS_FF = "read_A_7__ap_idle" *)input read_A_7__ap_idle;
  (* RS_AP_CTRL = "read_A_8.ap_start" *)output read_A_8__ap_start;
  (* RS_AP_CTRL = "read_A_8.ap_ready" *)input read_A_8__ap_ready;
  (* RS_FF = "read_A_8__ap_done" *)input read_A_8__ap_done;
  (* RS_FF = "read_A_8__ap_idle" *)input read_A_8__ap_idle;
  (* RS_AP_CTRL = "read_A_9.ap_start" *)output read_A_9__ap_start;
  (* RS_AP_CTRL = "read_A_9.ap_ready" *)input read_A_9__ap_ready;
  (* RS_FF = "read_A_9__ap_done" *)input read_A_9__ap_done;
  (* RS_FF = "read_A_9__ap_idle" *)input read_A_9__ap_idle;
  (* RS_AP_CTRL = "read_A_10.ap_start" *)output read_A_10__ap_start;
  (* RS_AP_CTRL = "read_A_10.ap_ready" *)input read_A_10__ap_ready;
  (* RS_FF = "read_A_10__ap_done" *)input read_A_10__ap_done;
  (* RS_FF = "read_A_10__ap_idle" *)input read_A_10__ap_idle;
  (* RS_AP_CTRL = "read_A_11.ap_start" *)output read_A_11__ap_start;
  (* RS_AP_CTRL = "read_A_11.ap_ready" *)input read_A_11__ap_ready;
  (* RS_FF = "read_A_11__ap_done" *)input read_A_11__ap_done;
  (* RS_FF = "read_A_11__ap_idle" *)input read_A_11__ap_idle;
  (* RS_AP_CTRL = "read_A_12.ap_start" *)output read_A_12__ap_start;
  (* RS_AP_CTRL = "read_A_12.ap_ready" *)input read_A_12__ap_ready;
  (* RS_FF = "read_A_12__ap_done" *)input read_A_12__ap_done;
  (* RS_FF = "read_A_12__ap_idle" *)input read_A_12__ap_idle;
  (* RS_AP_CTRL = "read_A_13.ap_start" *)output read_A_13__ap_start;
  (* RS_AP_CTRL = "read_A_13.ap_ready" *)input read_A_13__ap_ready;
  (* RS_FF = "read_A_13__ap_done" *)input read_A_13__ap_done;
  (* RS_FF = "read_A_13__ap_idle" *)input read_A_13__ap_idle;
  (* RS_AP_CTRL = "read_A_14.ap_start" *)output read_A_14__ap_start;
  (* RS_AP_CTRL = "read_A_14.ap_ready" *)input read_A_14__ap_ready;
  (* RS_FF = "read_A_14__ap_done" *)input read_A_14__ap_done;
  (* RS_FF = "read_A_14__ap_idle" *)input read_A_14__ap_idle;
  (* RS_AP_CTRL = "read_A_15.ap_start" *)output read_A_15__ap_start;
  (* RS_AP_CTRL = "read_A_15.ap_ready" *)input read_A_15__ap_ready;
  (* RS_FF = "read_A_15__ap_done" *)input read_A_15__ap_done;
  (* RS_FF = "read_A_15__ap_idle" *)input read_A_15__ap_idle;
  (* RS_AP_CTRL = "read_A_16.ap_start" *)output read_A_16__ap_start;
  (* RS_AP_CTRL = "read_A_16.ap_ready" *)input read_A_16__ap_ready;
  (* RS_FF = "read_A_16__ap_done" *)input read_A_16__ap_done;
  (* RS_FF = "read_A_16__ap_idle" *)input read_A_16__ap_idle;
  (* RS_AP_CTRL = "read_A_17.ap_start" *)output read_A_17__ap_start;
  (* RS_AP_CTRL = "read_A_17.ap_ready" *)input read_A_17__ap_ready;
  (* RS_FF = "read_A_17__ap_done" *)input read_A_17__ap_done;
  (* RS_FF = "read_A_17__ap_idle" *)input read_A_17__ap_idle;
  (* RS_AP_CTRL = "read_A_18.ap_start" *)output read_A_18__ap_start;
  (* RS_AP_CTRL = "read_A_18.ap_ready" *)input read_A_18__ap_ready;
  (* RS_FF = "read_A_18__ap_done" *)input read_A_18__ap_done;
  (* RS_FF = "read_A_18__ap_idle" *)input read_A_18__ap_idle;
  (* RS_AP_CTRL = "read_A_19.ap_start" *)output read_A_19__ap_start;
  (* RS_AP_CTRL = "read_A_19.ap_ready" *)input read_A_19__ap_ready;
  (* RS_FF = "read_A_19__ap_done" *)input read_A_19__ap_done;
  (* RS_FF = "read_A_19__ap_idle" *)input read_A_19__ap_idle;
  (* RS_AP_CTRL = "read_A_20.ap_start" *)output read_A_20__ap_start;
  (* RS_AP_CTRL = "read_A_20.ap_ready" *)input read_A_20__ap_ready;
  (* RS_FF = "read_A_20__ap_done" *)input read_A_20__ap_done;
  (* RS_FF = "read_A_20__ap_idle" *)input read_A_20__ap_idle;
  (* RS_AP_CTRL = "read_A_21.ap_start" *)output read_A_21__ap_start;
  (* RS_AP_CTRL = "read_A_21.ap_ready" *)input read_A_21__ap_ready;
  (* RS_FF = "read_A_21__ap_done" *)input read_A_21__ap_done;
  (* RS_FF = "read_A_21__ap_idle" *)input read_A_21__ap_idle;
  (* RS_AP_CTRL = "read_A_22.ap_start" *)output read_A_22__ap_start;
  (* RS_AP_CTRL = "read_A_22.ap_ready" *)input read_A_22__ap_ready;
  (* RS_FF = "read_A_22__ap_done" *)input read_A_22__ap_done;
  (* RS_FF = "read_A_22__ap_idle" *)input read_A_22__ap_idle;
  (* RS_AP_CTRL = "read_A_23.ap_start" *)output read_A_23__ap_start;
  (* RS_AP_CTRL = "read_A_23.ap_ready" *)input read_A_23__ap_ready;
  (* RS_FF = "read_A_23__ap_done" *)input read_A_23__ap_done;
  (* RS_FF = "read_A_23__ap_idle" *)input read_A_23__ap_idle;
  (* RS_AP_CTRL = "read_A_24.ap_start" *)output read_A_24__ap_start;
  (* RS_AP_CTRL = "read_A_24.ap_ready" *)input read_A_24__ap_ready;
  (* RS_FF = "read_A_24__ap_done" *)input read_A_24__ap_done;
  (* RS_FF = "read_A_24__ap_idle" *)input read_A_24__ap_idle;
  (* RS_AP_CTRL = "read_A_25.ap_start" *)output read_A_25__ap_start;
  (* RS_AP_CTRL = "read_A_25.ap_ready" *)input read_A_25__ap_ready;
  (* RS_FF = "read_A_25__ap_done" *)input read_A_25__ap_done;
  (* RS_FF = "read_A_25__ap_idle" *)input read_A_25__ap_idle;
  (* RS_AP_CTRL = "read_A_26.ap_start" *)output read_A_26__ap_start;
  (* RS_AP_CTRL = "read_A_26.ap_ready" *)input read_A_26__ap_ready;
  (* RS_FF = "read_A_26__ap_done" *)input read_A_26__ap_done;
  (* RS_FF = "read_A_26__ap_idle" *)input read_A_26__ap_idle;
  (* RS_AP_CTRL = "read_A_27.ap_start" *)output read_A_27__ap_start;
  (* RS_AP_CTRL = "read_A_27.ap_ready" *)input read_A_27__ap_ready;
  (* RS_FF = "read_A_27__ap_done" *)input read_A_27__ap_done;
  (* RS_FF = "read_A_27__ap_idle" *)input read_A_27__ap_idle;
  (* RS_AP_CTRL = "read_A_28.ap_start" *)output read_A_28__ap_start;
  (* RS_AP_CTRL = "read_A_28.ap_ready" *)input read_A_28__ap_ready;
  (* RS_FF = "read_A_28__ap_done" *)input read_A_28__ap_done;
  (* RS_FF = "read_A_28__ap_idle" *)input read_A_28__ap_idle;
  (* RS_AP_CTRL = "read_A_29.ap_start" *)output read_A_29__ap_start;
  (* RS_AP_CTRL = "read_A_29.ap_ready" *)input read_A_29__ap_ready;
  (* RS_FF = "read_A_29__ap_done" *)input read_A_29__ap_done;
  (* RS_FF = "read_A_29__ap_idle" *)input read_A_29__ap_idle;
  (* RS_AP_CTRL = "read_A_30.ap_start" *)output read_A_30__ap_start;
  (* RS_AP_CTRL = "read_A_30.ap_ready" *)input read_A_30__ap_ready;
  (* RS_FF = "read_A_30__ap_done" *)input read_A_30__ap_done;
  (* RS_FF = "read_A_30__ap_idle" *)input read_A_30__ap_idle;
  (* RS_AP_CTRL = "read_A_31.ap_start" *)output read_A_31__ap_start;
  (* RS_AP_CTRL = "read_A_31.ap_ready" *)input read_A_31__ap_ready;
  (* RS_FF = "read_A_31__ap_done" *)input read_A_31__ap_done;
  (* RS_FF = "read_A_31__ap_idle" *)input read_A_31__ap_idle;
  (* RS_AP_CTRL = "read_A_32.ap_start" *)output read_A_32__ap_start;
  (* RS_AP_CTRL = "read_A_32.ap_ready" *)input read_A_32__ap_ready;
  (* RS_FF = "read_A_32__ap_done" *)input read_A_32__ap_done;
  (* RS_FF = "read_A_32__ap_idle" *)input read_A_32__ap_idle;
  (* RS_AP_CTRL = "read_A_33.ap_start" *)output read_A_33__ap_start;
  (* RS_AP_CTRL = "read_A_33.ap_ready" *)input read_A_33__ap_ready;
  (* RS_FF = "read_A_33__ap_done" *)input read_A_33__ap_done;
  (* RS_FF = "read_A_33__ap_idle" *)input read_A_33__ap_idle;
  (* RS_AP_CTRL = "read_A_34.ap_start" *)output read_A_34__ap_start;
  (* RS_AP_CTRL = "read_A_34.ap_ready" *)input read_A_34__ap_ready;
  (* RS_FF = "read_A_34__ap_done" *)input read_A_34__ap_done;
  (* RS_FF = "read_A_34__ap_idle" *)input read_A_34__ap_idle;
  (* RS_AP_CTRL = "read_A_35.ap_start" *)output read_A_35__ap_start;
  (* RS_AP_CTRL = "read_A_35.ap_ready" *)input read_A_35__ap_ready;
  (* RS_FF = "read_A_35__ap_done" *)input read_A_35__ap_done;
  (* RS_FF = "read_A_35__ap_idle" *)input read_A_35__ap_idle;
  (* RS_AP_CTRL = "read_A_36.ap_start" *)output read_A_36__ap_start;
  (* RS_AP_CTRL = "read_A_36.ap_ready" *)input read_A_36__ap_ready;
  (* RS_FF = "read_A_36__ap_done" *)input read_A_36__ap_done;
  (* RS_FF = "read_A_36__ap_idle" *)input read_A_36__ap_idle;
  (* RS_AP_CTRL = "read_A_37.ap_start" *)output read_A_37__ap_start;
  (* RS_AP_CTRL = "read_A_37.ap_ready" *)input read_A_37__ap_ready;
  (* RS_FF = "read_A_37__ap_done" *)input read_A_37__ap_done;
  (* RS_FF = "read_A_37__ap_idle" *)input read_A_37__ap_idle;
  (* RS_AP_CTRL = "read_A_38.ap_start" *)output read_A_38__ap_start;
  (* RS_AP_CTRL = "read_A_38.ap_ready" *)input read_A_38__ap_ready;
  (* RS_FF = "read_A_38__ap_done" *)input read_A_38__ap_done;
  (* RS_FF = "read_A_38__ap_idle" *)input read_A_38__ap_idle;
  (* RS_AP_CTRL = "read_A_39.ap_start" *)output read_A_39__ap_start;
  (* RS_AP_CTRL = "read_A_39.ap_ready" *)input read_A_39__ap_ready;
  (* RS_FF = "read_A_39__ap_done" *)input read_A_39__ap_done;
  (* RS_FF = "read_A_39__ap_idle" *)input read_A_39__ap_idle;
  (* RS_AP_CTRL = "read_A_40.ap_start" *)output read_A_40__ap_start;
  (* RS_AP_CTRL = "read_A_40.ap_ready" *)input read_A_40__ap_ready;
  (* RS_FF = "read_A_40__ap_done" *)input read_A_40__ap_done;
  (* RS_FF = "read_A_40__ap_idle" *)input read_A_40__ap_idle;
  (* RS_AP_CTRL = "read_A_41.ap_start" *)output read_A_41__ap_start;
  (* RS_AP_CTRL = "read_A_41.ap_ready" *)input read_A_41__ap_ready;
  (* RS_FF = "read_A_41__ap_done" *)input read_A_41__ap_done;
  (* RS_FF = "read_A_41__ap_idle" *)input read_A_41__ap_idle;
  (* RS_AP_CTRL = "read_A_42.ap_start" *)output read_A_42__ap_start;
  (* RS_AP_CTRL = "read_A_42.ap_ready" *)input read_A_42__ap_ready;
  (* RS_FF = "read_A_42__ap_done" *)input read_A_42__ap_done;
  (* RS_FF = "read_A_42__ap_idle" *)input read_A_42__ap_idle;
  (* RS_AP_CTRL = "read_A_43.ap_start" *)output read_A_43__ap_start;
  (* RS_AP_CTRL = "read_A_43.ap_ready" *)input read_A_43__ap_ready;
  (* RS_FF = "read_A_43__ap_done" *)input read_A_43__ap_done;
  (* RS_FF = "read_A_43__ap_idle" *)input read_A_43__ap_idle;
  (* RS_AP_CTRL = "read_A_44.ap_start" *)output read_A_44__ap_start;
  (* RS_AP_CTRL = "read_A_44.ap_ready" *)input read_A_44__ap_ready;
  (* RS_FF = "read_A_44__ap_done" *)input read_A_44__ap_done;
  (* RS_FF = "read_A_44__ap_idle" *)input read_A_44__ap_idle;
  (* RS_AP_CTRL = "read_A_45.ap_start" *)output read_A_45__ap_start;
  (* RS_AP_CTRL = "read_A_45.ap_ready" *)input read_A_45__ap_ready;
  (* RS_FF = "read_A_45__ap_done" *)input read_A_45__ap_done;
  (* RS_FF = "read_A_45__ap_idle" *)input read_A_45__ap_idle;
  (* RS_AP_CTRL = "read_A_46.ap_start" *)output read_A_46__ap_start;
  (* RS_AP_CTRL = "read_A_46.ap_ready" *)input read_A_46__ap_ready;
  (* RS_FF = "read_A_46__ap_done" *)input read_A_46__ap_done;
  (* RS_FF = "read_A_46__ap_idle" *)input read_A_46__ap_idle;
  (* RS_AP_CTRL = "read_A_47.ap_start" *)output read_A_47__ap_start;
  (* RS_AP_CTRL = "read_A_47.ap_ready" *)input read_A_47__ap_ready;
  (* RS_FF = "read_A_47__ap_done" *)input read_A_47__ap_done;
  (* RS_FF = "read_A_47__ap_idle" *)input read_A_47__ap_idle;
  (* RS_AP_CTRL = "read_A_48.ap_start" *)output read_A_48__ap_start;
  (* RS_AP_CTRL = "read_A_48.ap_ready" *)input read_A_48__ap_ready;
  (* RS_FF = "read_A_48__ap_done" *)input read_A_48__ap_done;
  (* RS_FF = "read_A_48__ap_idle" *)input read_A_48__ap_idle;
  (* RS_AP_CTRL = "read_A_49.ap_start" *)output read_A_49__ap_start;
  (* RS_AP_CTRL = "read_A_49.ap_ready" *)input read_A_49__ap_ready;
  (* RS_FF = "read_A_49__ap_done" *)input read_A_49__ap_done;
  (* RS_FF = "read_A_49__ap_idle" *)input read_A_49__ap_idle;
  (* RS_AP_CTRL = "read_A_50.ap_start" *)output read_A_50__ap_start;
  (* RS_AP_CTRL = "read_A_50.ap_ready" *)input read_A_50__ap_ready;
  (* RS_FF = "read_A_50__ap_done" *)input read_A_50__ap_done;
  (* RS_FF = "read_A_50__ap_idle" *)input read_A_50__ap_idle;
  (* RS_AP_CTRL = "read_A_51.ap_start" *)output read_A_51__ap_start;
  (* RS_AP_CTRL = "read_A_51.ap_ready" *)input read_A_51__ap_ready;
  (* RS_FF = "read_A_51__ap_done" *)input read_A_51__ap_done;
  (* RS_FF = "read_A_51__ap_idle" *)input read_A_51__ap_idle;
  (* RS_AP_CTRL = "read_A_52.ap_start" *)output read_A_52__ap_start;
  (* RS_AP_CTRL = "read_A_52.ap_ready" *)input read_A_52__ap_ready;
  (* RS_FF = "read_A_52__ap_done" *)input read_A_52__ap_done;
  (* RS_FF = "read_A_52__ap_idle" *)input read_A_52__ap_idle;
  (* RS_AP_CTRL = "read_A_53.ap_start" *)output read_A_53__ap_start;
  (* RS_AP_CTRL = "read_A_53.ap_ready" *)input read_A_53__ap_ready;
  (* RS_FF = "read_A_53__ap_done" *)input read_A_53__ap_done;
  (* RS_FF = "read_A_53__ap_idle" *)input read_A_53__ap_idle;
  (* RS_AP_CTRL = "read_A_54.ap_start" *)output read_A_54__ap_start;
  (* RS_AP_CTRL = "read_A_54.ap_ready" *)input read_A_54__ap_ready;
  (* RS_FF = "read_A_54__ap_done" *)input read_A_54__ap_done;
  (* RS_FF = "read_A_54__ap_idle" *)input read_A_54__ap_idle;
  (* RS_AP_CTRL = "read_A_55.ap_start" *)output read_A_55__ap_start;
  (* RS_AP_CTRL = "read_A_55.ap_ready" *)input read_A_55__ap_ready;
  (* RS_FF = "read_A_55__ap_done" *)input read_A_55__ap_done;
  (* RS_FF = "read_A_55__ap_idle" *)input read_A_55__ap_idle;
  (* RS_AP_CTRL = "read_X_0.ap_start" *)output read_X_0__ap_start;
  (* RS_AP_CTRL = "read_X_0.ap_ready" *)input read_X_0__ap_ready;
  (* RS_FF = "read_X_0__ap_done" *)input read_X_0__ap_done;
  (* RS_FF = "read_X_0__ap_idle" *)input read_X_0__ap_idle;
  (* RS_AP_CTRL = "read_Y_0.ap_start" *)output read_Y_0__ap_start;
  (* RS_AP_CTRL = "read_Y_0.ap_ready" *)input read_Y_0__ap_ready;
  (* RS_FF = "read_Y_0__ap_done" *)input read_Y_0__ap_done;
  (* RS_FF = "read_Y_0__ap_idle" *)input read_Y_0__ap_idle;
  (* RS_AP_CTRL = "read_edge_list_ptr_0.ap_start" *)output read_edge_list_ptr_0__ap_start;
  (* RS_AP_CTRL = "read_edge_list_ptr_0.ap_ready" *)input read_edge_list_ptr_0__ap_ready;
  (* RS_FF = "read_edge_list_ptr_0__ap_done" *)input read_edge_list_ptr_0__ap_done;
  (* RS_FF = "read_edge_list_ptr_0__ap_idle" *)input read_edge_list_ptr_0__ap_idle;
  (* RS_AP_CTRL = "write_Y_0.ap_start" *)output write_Y_0__ap_start;
  (* RS_AP_CTRL = "write_Y_0.ap_ready" *)input write_Y_0__ap_ready;
  (* RS_FF = "write_Y_0__ap_done" *)input write_Y_0__ap_done;
  (* RS_FF = "write_Y_0__ap_idle" *)input write_Y_0__ap_idle;
  wire Arbiter_Y_0__ap_start_global__q0;
  wire Arbiter_Y_0__is_done__q0;
  wire Arbiter_Y_0__ap_done_global__q0;
  wire Arbiter_Y_0__ap_start;
  wire Arbiter_Y_0__ap_ready;
  wire Arbiter_Y_0__ap_done;
  wire Arbiter_Y_0__ap_idle;
  reg [1:0] Arbiter_Y_0__state;
  wire Arbiter_Y_1__ap_start_global__q0;
  wire Arbiter_Y_1__is_done__q0;
  wire Arbiter_Y_1__ap_done_global__q0;
  wire Arbiter_Y_1__ap_start;
  wire Arbiter_Y_1__ap_ready;
  wire Arbiter_Y_1__ap_done;
  wire Arbiter_Y_1__ap_idle;
  reg [1:0] Arbiter_Y_1__state;
  wire Arbiter_Y_2__ap_start_global__q0;
  wire Arbiter_Y_2__is_done__q0;
  wire Arbiter_Y_2__ap_done_global__q0;
  wire Arbiter_Y_2__ap_start;
  wire Arbiter_Y_2__ap_ready;
  wire Arbiter_Y_2__ap_done;
  wire Arbiter_Y_2__ap_idle;
  reg [1:0] Arbiter_Y_2__state;
  wire Arbiter_Y_3__ap_start_global__q0;
  wire Arbiter_Y_3__is_done__q0;
  wire Arbiter_Y_3__ap_done_global__q0;
  wire Arbiter_Y_3__ap_start;
  wire Arbiter_Y_3__ap_ready;
  wire Arbiter_Y_3__ap_done;
  wire Arbiter_Y_3__ap_idle;
  reg [1:0] Arbiter_Y_3__state;
  wire Arbiter_Y_4__ap_start_global__q0;
  wire Arbiter_Y_4__is_done__q0;
  wire Arbiter_Y_4__ap_done_global__q0;
  wire Arbiter_Y_4__ap_start;
  wire Arbiter_Y_4__ap_ready;
  wire Arbiter_Y_4__ap_done;
  wire Arbiter_Y_4__ap_idle;
  reg [1:0] Arbiter_Y_4__state;
  wire Arbiter_Y_5__ap_start_global__q0;
  wire Arbiter_Y_5__is_done__q0;
  wire Arbiter_Y_5__ap_done_global__q0;
  wire Arbiter_Y_5__ap_start;
  wire Arbiter_Y_5__ap_ready;
  wire Arbiter_Y_5__ap_done;
  wire Arbiter_Y_5__ap_idle;
  reg [1:0] Arbiter_Y_5__state;
  wire Arbiter_Y_6__ap_start_global__q0;
  wire Arbiter_Y_6__is_done__q0;
  wire Arbiter_Y_6__ap_done_global__q0;
  wire Arbiter_Y_6__ap_start;
  wire Arbiter_Y_6__ap_ready;
  wire Arbiter_Y_6__ap_done;
  wire Arbiter_Y_6__ap_idle;
  reg [1:0] Arbiter_Y_6__state;
  wire Arbiter_Y_7__ap_start_global__q0;
  wire Arbiter_Y_7__is_done__q0;
  wire Arbiter_Y_7__ap_done_global__q0;
  wire Arbiter_Y_7__ap_start;
  wire Arbiter_Y_7__ap_ready;
  wire Arbiter_Y_7__ap_done;
  wire Arbiter_Y_7__ap_idle;
  reg [1:0] Arbiter_Y_7__state;
  wire FloatvAddFloatv_0__ap_start_global__q0;
  reg FloatvAddFloatv_0__ap_start;
  wire FloatvMultConst_0__ap_start_global__q0;
  wire FloatvMultConst_0__is_done__q0;
  wire FloatvMultConst_0__ap_done_global__q0;
  wire FloatvMultConst_0__ap_start;
  wire FloatvMultConst_0__ap_ready;
  wire FloatvMultConst_0__ap_done;
  wire FloatvMultConst_0__ap_idle;
  reg [1:0] FloatvMultConst_0__state;
  wire FloatvMultConst_1__ap_start_global__q0;
  wire FloatvMultConst_1__is_done__q0;
  wire FloatvMultConst_1__ap_done_global__q0;
  wire FloatvMultConst_1__ap_start;
  wire FloatvMultConst_1__ap_ready;
  wire FloatvMultConst_1__ap_done;
  wire FloatvMultConst_1__ap_idle;
  reg [1:0] FloatvMultConst_1__state;
  wire Merger_Y_0__ap_start_global__q0;
  reg Merger_Y_0__ap_start;
  wire PEG_Xvec_0__ap_start_global__q0;
  wire PEG_Xvec_0__is_done__q0;
  wire PEG_Xvec_0__ap_done_global__q0;
  wire PEG_Xvec_0__ap_start;
  wire PEG_Xvec_0__ap_ready;
  wire PEG_Xvec_0__ap_done;
  wire PEG_Xvec_0__ap_idle;
  reg [1:0] PEG_Xvec_0__state;
  wire PEG_Xvec_1__ap_start_global__q0;
  wire PEG_Xvec_1__is_done__q0;
  wire PEG_Xvec_1__ap_done_global__q0;
  wire PEG_Xvec_1__ap_start;
  wire PEG_Xvec_1__ap_ready;
  wire PEG_Xvec_1__ap_done;
  wire PEG_Xvec_1__ap_idle;
  reg [1:0] PEG_Xvec_1__state;
  wire PEG_Xvec_2__ap_start_global__q0;
  wire PEG_Xvec_2__is_done__q0;
  wire PEG_Xvec_2__ap_done_global__q0;
  wire PEG_Xvec_2__ap_start;
  wire PEG_Xvec_2__ap_ready;
  wire PEG_Xvec_2__ap_done;
  wire PEG_Xvec_2__ap_idle;
  reg [1:0] PEG_Xvec_2__state;
  wire PEG_Xvec_3__ap_start_global__q0;
  wire PEG_Xvec_3__is_done__q0;
  wire PEG_Xvec_3__ap_done_global__q0;
  wire PEG_Xvec_3__ap_start;
  wire PEG_Xvec_3__ap_ready;
  wire PEG_Xvec_3__ap_done;
  wire PEG_Xvec_3__ap_idle;
  reg [1:0] PEG_Xvec_3__state;
  wire PEG_Xvec_4__ap_start_global__q0;
  wire PEG_Xvec_4__is_done__q0;
  wire PEG_Xvec_4__ap_done_global__q0;
  wire PEG_Xvec_4__ap_start;
  wire PEG_Xvec_4__ap_ready;
  wire PEG_Xvec_4__ap_done;
  wire PEG_Xvec_4__ap_idle;
  reg [1:0] PEG_Xvec_4__state;
  wire PEG_Xvec_5__ap_start_global__q0;
  wire PEG_Xvec_5__is_done__q0;
  wire PEG_Xvec_5__ap_done_global__q0;
  wire PEG_Xvec_5__ap_start;
  wire PEG_Xvec_5__ap_ready;
  wire PEG_Xvec_5__ap_done;
  wire PEG_Xvec_5__ap_idle;
  reg [1:0] PEG_Xvec_5__state;
  wire PEG_Xvec_6__ap_start_global__q0;
  wire PEG_Xvec_6__is_done__q0;
  wire PEG_Xvec_6__ap_done_global__q0;
  wire PEG_Xvec_6__ap_start;
  wire PEG_Xvec_6__ap_ready;
  wire PEG_Xvec_6__ap_done;
  wire PEG_Xvec_6__ap_idle;
  reg [1:0] PEG_Xvec_6__state;
  wire PEG_Xvec_7__ap_start_global__q0;
  wire PEG_Xvec_7__is_done__q0;
  wire PEG_Xvec_7__ap_done_global__q0;
  wire PEG_Xvec_7__ap_start;
  wire PEG_Xvec_7__ap_ready;
  wire PEG_Xvec_7__ap_done;
  wire PEG_Xvec_7__ap_idle;
  reg [1:0] PEG_Xvec_7__state;
  wire PEG_Xvec_8__ap_start_global__q0;
  wire PEG_Xvec_8__is_done__q0;
  wire PEG_Xvec_8__ap_done_global__q0;
  wire PEG_Xvec_8__ap_start;
  wire PEG_Xvec_8__ap_ready;
  wire PEG_Xvec_8__ap_done;
  wire PEG_Xvec_8__ap_idle;
  reg [1:0] PEG_Xvec_8__state;
  wire PEG_Xvec_9__ap_start_global__q0;
  wire PEG_Xvec_9__is_done__q0;
  wire PEG_Xvec_9__ap_done_global__q0;
  wire PEG_Xvec_9__ap_start;
  wire PEG_Xvec_9__ap_ready;
  wire PEG_Xvec_9__ap_done;
  wire PEG_Xvec_9__ap_idle;
  reg [1:0] PEG_Xvec_9__state;
  wire PEG_Xvec_10__ap_start_global__q0;
  wire PEG_Xvec_10__is_done__q0;
  wire PEG_Xvec_10__ap_done_global__q0;
  wire PEG_Xvec_10__ap_start;
  wire PEG_Xvec_10__ap_ready;
  wire PEG_Xvec_10__ap_done;
  wire PEG_Xvec_10__ap_idle;
  reg [1:0] PEG_Xvec_10__state;
  wire PEG_Xvec_11__ap_start_global__q0;
  wire PEG_Xvec_11__is_done__q0;
  wire PEG_Xvec_11__ap_done_global__q0;
  wire PEG_Xvec_11__ap_start;
  wire PEG_Xvec_11__ap_ready;
  wire PEG_Xvec_11__ap_done;
  wire PEG_Xvec_11__ap_idle;
  reg [1:0] PEG_Xvec_11__state;
  wire PEG_Xvec_12__ap_start_global__q0;
  wire PEG_Xvec_12__is_done__q0;
  wire PEG_Xvec_12__ap_done_global__q0;
  wire PEG_Xvec_12__ap_start;
  wire PEG_Xvec_12__ap_ready;
  wire PEG_Xvec_12__ap_done;
  wire PEG_Xvec_12__ap_idle;
  reg [1:0] PEG_Xvec_12__state;
  wire PEG_Xvec_13__ap_start_global__q0;
  wire PEG_Xvec_13__is_done__q0;
  wire PEG_Xvec_13__ap_done_global__q0;
  wire PEG_Xvec_13__ap_start;
  wire PEG_Xvec_13__ap_ready;
  wire PEG_Xvec_13__ap_done;
  wire PEG_Xvec_13__ap_idle;
  reg [1:0] PEG_Xvec_13__state;
  wire PEG_Xvec_14__ap_start_global__q0;
  wire PEG_Xvec_14__is_done__q0;
  wire PEG_Xvec_14__ap_done_global__q0;
  wire PEG_Xvec_14__ap_start;
  wire PEG_Xvec_14__ap_ready;
  wire PEG_Xvec_14__ap_done;
  wire PEG_Xvec_14__ap_idle;
  reg [1:0] PEG_Xvec_14__state;
  wire PEG_Xvec_15__ap_start_global__q0;
  wire PEG_Xvec_15__is_done__q0;
  wire PEG_Xvec_15__ap_done_global__q0;
  wire PEG_Xvec_15__ap_start;
  wire PEG_Xvec_15__ap_ready;
  wire PEG_Xvec_15__ap_done;
  wire PEG_Xvec_15__ap_idle;
  reg [1:0] PEG_Xvec_15__state;
  wire PEG_Xvec_16__ap_start_global__q0;
  wire PEG_Xvec_16__is_done__q0;
  wire PEG_Xvec_16__ap_done_global__q0;
  wire PEG_Xvec_16__ap_start;
  wire PEG_Xvec_16__ap_ready;
  wire PEG_Xvec_16__ap_done;
  wire PEG_Xvec_16__ap_idle;
  reg [1:0] PEG_Xvec_16__state;
  wire PEG_Xvec_17__ap_start_global__q0;
  wire PEG_Xvec_17__is_done__q0;
  wire PEG_Xvec_17__ap_done_global__q0;
  wire PEG_Xvec_17__ap_start;
  wire PEG_Xvec_17__ap_ready;
  wire PEG_Xvec_17__ap_done;
  wire PEG_Xvec_17__ap_idle;
  reg [1:0] PEG_Xvec_17__state;
  wire PEG_Xvec_18__ap_start_global__q0;
  wire PEG_Xvec_18__is_done__q0;
  wire PEG_Xvec_18__ap_done_global__q0;
  wire PEG_Xvec_18__ap_start;
  wire PEG_Xvec_18__ap_ready;
  wire PEG_Xvec_18__ap_done;
  wire PEG_Xvec_18__ap_idle;
  reg [1:0] PEG_Xvec_18__state;
  wire PEG_Xvec_19__ap_start_global__q0;
  wire PEG_Xvec_19__is_done__q0;
  wire PEG_Xvec_19__ap_done_global__q0;
  wire PEG_Xvec_19__ap_start;
  wire PEG_Xvec_19__ap_ready;
  wire PEG_Xvec_19__ap_done;
  wire PEG_Xvec_19__ap_idle;
  reg [1:0] PEG_Xvec_19__state;
  wire PEG_Xvec_20__ap_start_global__q0;
  wire PEG_Xvec_20__is_done__q0;
  wire PEG_Xvec_20__ap_done_global__q0;
  wire PEG_Xvec_20__ap_start;
  wire PEG_Xvec_20__ap_ready;
  wire PEG_Xvec_20__ap_done;
  wire PEG_Xvec_20__ap_idle;
  reg [1:0] PEG_Xvec_20__state;
  wire PEG_Xvec_21__ap_start_global__q0;
  wire PEG_Xvec_21__is_done__q0;
  wire PEG_Xvec_21__ap_done_global__q0;
  wire PEG_Xvec_21__ap_start;
  wire PEG_Xvec_21__ap_ready;
  wire PEG_Xvec_21__ap_done;
  wire PEG_Xvec_21__ap_idle;
  reg [1:0] PEG_Xvec_21__state;
  wire PEG_Xvec_22__ap_start_global__q0;
  wire PEG_Xvec_22__is_done__q0;
  wire PEG_Xvec_22__ap_done_global__q0;
  wire PEG_Xvec_22__ap_start;
  wire PEG_Xvec_22__ap_ready;
  wire PEG_Xvec_22__ap_done;
  wire PEG_Xvec_22__ap_idle;
  reg [1:0] PEG_Xvec_22__state;
  wire PEG_Xvec_23__ap_start_global__q0;
  wire PEG_Xvec_23__is_done__q0;
  wire PEG_Xvec_23__ap_done_global__q0;
  wire PEG_Xvec_23__ap_start;
  wire PEG_Xvec_23__ap_ready;
  wire PEG_Xvec_23__ap_done;
  wire PEG_Xvec_23__ap_idle;
  reg [1:0] PEG_Xvec_23__state;
  wire PEG_Xvec_24__ap_start_global__q0;
  wire PEG_Xvec_24__is_done__q0;
  wire PEG_Xvec_24__ap_done_global__q0;
  wire PEG_Xvec_24__ap_start;
  wire PEG_Xvec_24__ap_ready;
  wire PEG_Xvec_24__ap_done;
  wire PEG_Xvec_24__ap_idle;
  reg [1:0] PEG_Xvec_24__state;
  wire PEG_Xvec_25__ap_start_global__q0;
  wire PEG_Xvec_25__is_done__q0;
  wire PEG_Xvec_25__ap_done_global__q0;
  wire PEG_Xvec_25__ap_start;
  wire PEG_Xvec_25__ap_ready;
  wire PEG_Xvec_25__ap_done;
  wire PEG_Xvec_25__ap_idle;
  reg [1:0] PEG_Xvec_25__state;
  wire PEG_Xvec_26__ap_start_global__q0;
  wire PEG_Xvec_26__is_done__q0;
  wire PEG_Xvec_26__ap_done_global__q0;
  wire PEG_Xvec_26__ap_start;
  wire PEG_Xvec_26__ap_ready;
  wire PEG_Xvec_26__ap_done;
  wire PEG_Xvec_26__ap_idle;
  reg [1:0] PEG_Xvec_26__state;
  wire PEG_Xvec_27__ap_start_global__q0;
  wire PEG_Xvec_27__is_done__q0;
  wire PEG_Xvec_27__ap_done_global__q0;
  wire PEG_Xvec_27__ap_start;
  wire PEG_Xvec_27__ap_ready;
  wire PEG_Xvec_27__ap_done;
  wire PEG_Xvec_27__ap_idle;
  reg [1:0] PEG_Xvec_27__state;
  wire PEG_Xvec_28__ap_start_global__q0;
  wire PEG_Xvec_28__is_done__q0;
  wire PEG_Xvec_28__ap_done_global__q0;
  wire PEG_Xvec_28__ap_start;
  wire PEG_Xvec_28__ap_ready;
  wire PEG_Xvec_28__ap_done;
  wire PEG_Xvec_28__ap_idle;
  reg [1:0] PEG_Xvec_28__state;
  wire PEG_Xvec_29__ap_start_global__q0;
  wire PEG_Xvec_29__is_done__q0;
  wire PEG_Xvec_29__ap_done_global__q0;
  wire PEG_Xvec_29__ap_start;
  wire PEG_Xvec_29__ap_ready;
  wire PEG_Xvec_29__ap_done;
  wire PEG_Xvec_29__ap_idle;
  reg [1:0] PEG_Xvec_29__state;
  wire PEG_Xvec_30__ap_start_global__q0;
  wire PEG_Xvec_30__is_done__q0;
  wire PEG_Xvec_30__ap_done_global__q0;
  wire PEG_Xvec_30__ap_start;
  wire PEG_Xvec_30__ap_ready;
  wire PEG_Xvec_30__ap_done;
  wire PEG_Xvec_30__ap_idle;
  reg [1:0] PEG_Xvec_30__state;
  wire PEG_Xvec_31__ap_start_global__q0;
  wire PEG_Xvec_31__is_done__q0;
  wire PEG_Xvec_31__ap_done_global__q0;
  wire PEG_Xvec_31__ap_start;
  wire PEG_Xvec_31__ap_ready;
  wire PEG_Xvec_31__ap_done;
  wire PEG_Xvec_31__ap_idle;
  reg [1:0] PEG_Xvec_31__state;
  wire PEG_Xvec_32__ap_start_global__q0;
  wire PEG_Xvec_32__is_done__q0;
  wire PEG_Xvec_32__ap_done_global__q0;
  wire PEG_Xvec_32__ap_start;
  wire PEG_Xvec_32__ap_ready;
  wire PEG_Xvec_32__ap_done;
  wire PEG_Xvec_32__ap_idle;
  reg [1:0] PEG_Xvec_32__state;
  wire PEG_Xvec_33__ap_start_global__q0;
  wire PEG_Xvec_33__is_done__q0;
  wire PEG_Xvec_33__ap_done_global__q0;
  wire PEG_Xvec_33__ap_start;
  wire PEG_Xvec_33__ap_ready;
  wire PEG_Xvec_33__ap_done;
  wire PEG_Xvec_33__ap_idle;
  reg [1:0] PEG_Xvec_33__state;
  wire PEG_Xvec_34__ap_start_global__q0;
  wire PEG_Xvec_34__is_done__q0;
  wire PEG_Xvec_34__ap_done_global__q0;
  wire PEG_Xvec_34__ap_start;
  wire PEG_Xvec_34__ap_ready;
  wire PEG_Xvec_34__ap_done;
  wire PEG_Xvec_34__ap_idle;
  reg [1:0] PEG_Xvec_34__state;
  wire PEG_Xvec_35__ap_start_global__q0;
  wire PEG_Xvec_35__is_done__q0;
  wire PEG_Xvec_35__ap_done_global__q0;
  wire PEG_Xvec_35__ap_start;
  wire PEG_Xvec_35__ap_ready;
  wire PEG_Xvec_35__ap_done;
  wire PEG_Xvec_35__ap_idle;
  reg [1:0] PEG_Xvec_35__state;
  wire PEG_Xvec_36__ap_start_global__q0;
  wire PEG_Xvec_36__is_done__q0;
  wire PEG_Xvec_36__ap_done_global__q0;
  wire PEG_Xvec_36__ap_start;
  wire PEG_Xvec_36__ap_ready;
  wire PEG_Xvec_36__ap_done;
  wire PEG_Xvec_36__ap_idle;
  reg [1:0] PEG_Xvec_36__state;
  wire PEG_Xvec_37__ap_start_global__q0;
  wire PEG_Xvec_37__is_done__q0;
  wire PEG_Xvec_37__ap_done_global__q0;
  wire PEG_Xvec_37__ap_start;
  wire PEG_Xvec_37__ap_ready;
  wire PEG_Xvec_37__ap_done;
  wire PEG_Xvec_37__ap_idle;
  reg [1:0] PEG_Xvec_37__state;
  wire PEG_Xvec_38__ap_start_global__q0;
  wire PEG_Xvec_38__is_done__q0;
  wire PEG_Xvec_38__ap_done_global__q0;
  wire PEG_Xvec_38__ap_start;
  wire PEG_Xvec_38__ap_ready;
  wire PEG_Xvec_38__ap_done;
  wire PEG_Xvec_38__ap_idle;
  reg [1:0] PEG_Xvec_38__state;
  wire PEG_Xvec_39__ap_start_global__q0;
  wire PEG_Xvec_39__is_done__q0;
  wire PEG_Xvec_39__ap_done_global__q0;
  wire PEG_Xvec_39__ap_start;
  wire PEG_Xvec_39__ap_ready;
  wire PEG_Xvec_39__ap_done;
  wire PEG_Xvec_39__ap_idle;
  reg [1:0] PEG_Xvec_39__state;
  wire PEG_Xvec_40__ap_start_global__q0;
  wire PEG_Xvec_40__is_done__q0;
  wire PEG_Xvec_40__ap_done_global__q0;
  wire PEG_Xvec_40__ap_start;
  wire PEG_Xvec_40__ap_ready;
  wire PEG_Xvec_40__ap_done;
  wire PEG_Xvec_40__ap_idle;
  reg [1:0] PEG_Xvec_40__state;
  wire PEG_Xvec_41__ap_start_global__q0;
  wire PEG_Xvec_41__is_done__q0;
  wire PEG_Xvec_41__ap_done_global__q0;
  wire PEG_Xvec_41__ap_start;
  wire PEG_Xvec_41__ap_ready;
  wire PEG_Xvec_41__ap_done;
  wire PEG_Xvec_41__ap_idle;
  reg [1:0] PEG_Xvec_41__state;
  wire PEG_Xvec_42__ap_start_global__q0;
  wire PEG_Xvec_42__is_done__q0;
  wire PEG_Xvec_42__ap_done_global__q0;
  wire PEG_Xvec_42__ap_start;
  wire PEG_Xvec_42__ap_ready;
  wire PEG_Xvec_42__ap_done;
  wire PEG_Xvec_42__ap_idle;
  reg [1:0] PEG_Xvec_42__state;
  wire PEG_Xvec_43__ap_start_global__q0;
  wire PEG_Xvec_43__is_done__q0;
  wire PEG_Xvec_43__ap_done_global__q0;
  wire PEG_Xvec_43__ap_start;
  wire PEG_Xvec_43__ap_ready;
  wire PEG_Xvec_43__ap_done;
  wire PEG_Xvec_43__ap_idle;
  reg [1:0] PEG_Xvec_43__state;
  wire PEG_Xvec_44__ap_start_global__q0;
  wire PEG_Xvec_44__is_done__q0;
  wire PEG_Xvec_44__ap_done_global__q0;
  wire PEG_Xvec_44__ap_start;
  wire PEG_Xvec_44__ap_ready;
  wire PEG_Xvec_44__ap_done;
  wire PEG_Xvec_44__ap_idle;
  reg [1:0] PEG_Xvec_44__state;
  wire PEG_Xvec_45__ap_start_global__q0;
  wire PEG_Xvec_45__is_done__q0;
  wire PEG_Xvec_45__ap_done_global__q0;
  wire PEG_Xvec_45__ap_start;
  wire PEG_Xvec_45__ap_ready;
  wire PEG_Xvec_45__ap_done;
  wire PEG_Xvec_45__ap_idle;
  reg [1:0] PEG_Xvec_45__state;
  wire PEG_Xvec_46__ap_start_global__q0;
  wire PEG_Xvec_46__is_done__q0;
  wire PEG_Xvec_46__ap_done_global__q0;
  wire PEG_Xvec_46__ap_start;
  wire PEG_Xvec_46__ap_ready;
  wire PEG_Xvec_46__ap_done;
  wire PEG_Xvec_46__ap_idle;
  reg [1:0] PEG_Xvec_46__state;
  wire PEG_Xvec_47__ap_start_global__q0;
  wire PEG_Xvec_47__is_done__q0;
  wire PEG_Xvec_47__ap_done_global__q0;
  wire PEG_Xvec_47__ap_start;
  wire PEG_Xvec_47__ap_ready;
  wire PEG_Xvec_47__ap_done;
  wire PEG_Xvec_47__ap_idle;
  reg [1:0] PEG_Xvec_47__state;
  wire PEG_Xvec_48__ap_start_global__q0;
  wire PEG_Xvec_48__is_done__q0;
  wire PEG_Xvec_48__ap_done_global__q0;
  wire PEG_Xvec_48__ap_start;
  wire PEG_Xvec_48__ap_ready;
  wire PEG_Xvec_48__ap_done;
  wire PEG_Xvec_48__ap_idle;
  reg [1:0] PEG_Xvec_48__state;
  wire PEG_Xvec_49__ap_start_global__q0;
  wire PEG_Xvec_49__is_done__q0;
  wire PEG_Xvec_49__ap_done_global__q0;
  wire PEG_Xvec_49__ap_start;
  wire PEG_Xvec_49__ap_ready;
  wire PEG_Xvec_49__ap_done;
  wire PEG_Xvec_49__ap_idle;
  reg [1:0] PEG_Xvec_49__state;
  wire PEG_Xvec_50__ap_start_global__q0;
  wire PEG_Xvec_50__is_done__q0;
  wire PEG_Xvec_50__ap_done_global__q0;
  wire PEG_Xvec_50__ap_start;
  wire PEG_Xvec_50__ap_ready;
  wire PEG_Xvec_50__ap_done;
  wire PEG_Xvec_50__ap_idle;
  reg [1:0] PEG_Xvec_50__state;
  wire PEG_Xvec_51__ap_start_global__q0;
  wire PEG_Xvec_51__is_done__q0;
  wire PEG_Xvec_51__ap_done_global__q0;
  wire PEG_Xvec_51__ap_start;
  wire PEG_Xvec_51__ap_ready;
  wire PEG_Xvec_51__ap_done;
  wire PEG_Xvec_51__ap_idle;
  reg [1:0] PEG_Xvec_51__state;
  wire PEG_Xvec_52__ap_start_global__q0;
  wire PEG_Xvec_52__is_done__q0;
  wire PEG_Xvec_52__ap_done_global__q0;
  wire PEG_Xvec_52__ap_start;
  wire PEG_Xvec_52__ap_ready;
  wire PEG_Xvec_52__ap_done;
  wire PEG_Xvec_52__ap_idle;
  reg [1:0] PEG_Xvec_52__state;
  wire PEG_Xvec_53__ap_start_global__q0;
  wire PEG_Xvec_53__is_done__q0;
  wire PEG_Xvec_53__ap_done_global__q0;
  wire PEG_Xvec_53__ap_start;
  wire PEG_Xvec_53__ap_ready;
  wire PEG_Xvec_53__ap_done;
  wire PEG_Xvec_53__ap_idle;
  reg [1:0] PEG_Xvec_53__state;
  wire PEG_Xvec_54__ap_start_global__q0;
  wire PEG_Xvec_54__is_done__q0;
  wire PEG_Xvec_54__ap_done_global__q0;
  wire PEG_Xvec_54__ap_start;
  wire PEG_Xvec_54__ap_ready;
  wire PEG_Xvec_54__ap_done;
  wire PEG_Xvec_54__ap_idle;
  reg [1:0] PEG_Xvec_54__state;
  wire PEG_Xvec_55__ap_start_global__q0;
  wire PEG_Xvec_55__is_done__q0;
  wire PEG_Xvec_55__ap_done_global__q0;
  wire PEG_Xvec_55__ap_start;
  wire PEG_Xvec_55__ap_ready;
  wire PEG_Xvec_55__ap_done;
  wire PEG_Xvec_55__ap_idle;
  reg [1:0] PEG_Xvec_55__state;
  wire PEG_Yvec_0__ap_start_global__q0;
  wire PEG_Yvec_0__is_done__q0;
  wire PEG_Yvec_0__ap_done_global__q0;
  wire PEG_Yvec_0__ap_start;
  wire PEG_Yvec_0__ap_ready;
  wire PEG_Yvec_0__ap_done;
  wire PEG_Yvec_0__ap_idle;
  reg [1:0] PEG_Yvec_0__state;
  wire PEG_Yvec_1__ap_start_global__q0;
  wire PEG_Yvec_1__is_done__q0;
  wire PEG_Yvec_1__ap_done_global__q0;
  wire PEG_Yvec_1__ap_start;
  wire PEG_Yvec_1__ap_ready;
  wire PEG_Yvec_1__ap_done;
  wire PEG_Yvec_1__ap_idle;
  reg [1:0] PEG_Yvec_1__state;
  wire PEG_Yvec_2__ap_start_global__q0;
  wire PEG_Yvec_2__is_done__q0;
  wire PEG_Yvec_2__ap_done_global__q0;
  wire PEG_Yvec_2__ap_start;
  wire PEG_Yvec_2__ap_ready;
  wire PEG_Yvec_2__ap_done;
  wire PEG_Yvec_2__ap_idle;
  reg [1:0] PEG_Yvec_2__state;
  wire PEG_Yvec_3__ap_start_global__q0;
  wire PEG_Yvec_3__is_done__q0;
  wire PEG_Yvec_3__ap_done_global__q0;
  wire PEG_Yvec_3__ap_start;
  wire PEG_Yvec_3__ap_ready;
  wire PEG_Yvec_3__ap_done;
  wire PEG_Yvec_3__ap_idle;
  reg [1:0] PEG_Yvec_3__state;
  wire PEG_Yvec_4__ap_start_global__q0;
  wire PEG_Yvec_4__is_done__q0;
  wire PEG_Yvec_4__ap_done_global__q0;
  wire PEG_Yvec_4__ap_start;
  wire PEG_Yvec_4__ap_ready;
  wire PEG_Yvec_4__ap_done;
  wire PEG_Yvec_4__ap_idle;
  reg [1:0] PEG_Yvec_4__state;
  wire PEG_Yvec_5__ap_start_global__q0;
  wire PEG_Yvec_5__is_done__q0;
  wire PEG_Yvec_5__ap_done_global__q0;
  wire PEG_Yvec_5__ap_start;
  wire PEG_Yvec_5__ap_ready;
  wire PEG_Yvec_5__ap_done;
  wire PEG_Yvec_5__ap_idle;
  reg [1:0] PEG_Yvec_5__state;
  wire PEG_Yvec_6__ap_start_global__q0;
  wire PEG_Yvec_6__is_done__q0;
  wire PEG_Yvec_6__ap_done_global__q0;
  wire PEG_Yvec_6__ap_start;
  wire PEG_Yvec_6__ap_ready;
  wire PEG_Yvec_6__ap_done;
  wire PEG_Yvec_6__ap_idle;
  reg [1:0] PEG_Yvec_6__state;
  wire PEG_Yvec_7__ap_start_global__q0;
  wire PEG_Yvec_7__is_done__q0;
  wire PEG_Yvec_7__ap_done_global__q0;
  wire PEG_Yvec_7__ap_start;
  wire PEG_Yvec_7__ap_ready;
  wire PEG_Yvec_7__ap_done;
  wire PEG_Yvec_7__ap_idle;
  reg [1:0] PEG_Yvec_7__state;
  wire PEG_Yvec_8__ap_start_global__q0;
  wire PEG_Yvec_8__is_done__q0;
  wire PEG_Yvec_8__ap_done_global__q0;
  wire PEG_Yvec_8__ap_start;
  wire PEG_Yvec_8__ap_ready;
  wire PEG_Yvec_8__ap_done;
  wire PEG_Yvec_8__ap_idle;
  reg [1:0] PEG_Yvec_8__state;
  wire PEG_Yvec_9__ap_start_global__q0;
  wire PEG_Yvec_9__is_done__q0;
  wire PEG_Yvec_9__ap_done_global__q0;
  wire PEG_Yvec_9__ap_start;
  wire PEG_Yvec_9__ap_ready;
  wire PEG_Yvec_9__ap_done;
  wire PEG_Yvec_9__ap_idle;
  reg [1:0] PEG_Yvec_9__state;
  wire PEG_Yvec_10__ap_start_global__q0;
  wire PEG_Yvec_10__is_done__q0;
  wire PEG_Yvec_10__ap_done_global__q0;
  wire PEG_Yvec_10__ap_start;
  wire PEG_Yvec_10__ap_ready;
  wire PEG_Yvec_10__ap_done;
  wire PEG_Yvec_10__ap_idle;
  reg [1:0] PEG_Yvec_10__state;
  wire PEG_Yvec_11__ap_start_global__q0;
  wire PEG_Yvec_11__is_done__q0;
  wire PEG_Yvec_11__ap_done_global__q0;
  wire PEG_Yvec_11__ap_start;
  wire PEG_Yvec_11__ap_ready;
  wire PEG_Yvec_11__ap_done;
  wire PEG_Yvec_11__ap_idle;
  reg [1:0] PEG_Yvec_11__state;
  wire PEG_Yvec_12__ap_start_global__q0;
  wire PEG_Yvec_12__is_done__q0;
  wire PEG_Yvec_12__ap_done_global__q0;
  wire PEG_Yvec_12__ap_start;
  wire PEG_Yvec_12__ap_ready;
  wire PEG_Yvec_12__ap_done;
  wire PEG_Yvec_12__ap_idle;
  reg [1:0] PEG_Yvec_12__state;
  wire PEG_Yvec_13__ap_start_global__q0;
  wire PEG_Yvec_13__is_done__q0;
  wire PEG_Yvec_13__ap_done_global__q0;
  wire PEG_Yvec_13__ap_start;
  wire PEG_Yvec_13__ap_ready;
  wire PEG_Yvec_13__ap_done;
  wire PEG_Yvec_13__ap_idle;
  reg [1:0] PEG_Yvec_13__state;
  wire PEG_Yvec_14__ap_start_global__q0;
  wire PEG_Yvec_14__is_done__q0;
  wire PEG_Yvec_14__ap_done_global__q0;
  wire PEG_Yvec_14__ap_start;
  wire PEG_Yvec_14__ap_ready;
  wire PEG_Yvec_14__ap_done;
  wire PEG_Yvec_14__ap_idle;
  reg [1:0] PEG_Yvec_14__state;
  wire PEG_Yvec_15__ap_start_global__q0;
  wire PEG_Yvec_15__is_done__q0;
  wire PEG_Yvec_15__ap_done_global__q0;
  wire PEG_Yvec_15__ap_start;
  wire PEG_Yvec_15__ap_ready;
  wire PEG_Yvec_15__ap_done;
  wire PEG_Yvec_15__ap_idle;
  reg [1:0] PEG_Yvec_15__state;
  wire PEG_Yvec_16__ap_start_global__q0;
  wire PEG_Yvec_16__is_done__q0;
  wire PEG_Yvec_16__ap_done_global__q0;
  wire PEG_Yvec_16__ap_start;
  wire PEG_Yvec_16__ap_ready;
  wire PEG_Yvec_16__ap_done;
  wire PEG_Yvec_16__ap_idle;
  reg [1:0] PEG_Yvec_16__state;
  wire PEG_Yvec_17__ap_start_global__q0;
  wire PEG_Yvec_17__is_done__q0;
  wire PEG_Yvec_17__ap_done_global__q0;
  wire PEG_Yvec_17__ap_start;
  wire PEG_Yvec_17__ap_ready;
  wire PEG_Yvec_17__ap_done;
  wire PEG_Yvec_17__ap_idle;
  reg [1:0] PEG_Yvec_17__state;
  wire PEG_Yvec_18__ap_start_global__q0;
  wire PEG_Yvec_18__is_done__q0;
  wire PEG_Yvec_18__ap_done_global__q0;
  wire PEG_Yvec_18__ap_start;
  wire PEG_Yvec_18__ap_ready;
  wire PEG_Yvec_18__ap_done;
  wire PEG_Yvec_18__ap_idle;
  reg [1:0] PEG_Yvec_18__state;
  wire PEG_Yvec_19__ap_start_global__q0;
  wire PEG_Yvec_19__is_done__q0;
  wire PEG_Yvec_19__ap_done_global__q0;
  wire PEG_Yvec_19__ap_start;
  wire PEG_Yvec_19__ap_ready;
  wire PEG_Yvec_19__ap_done;
  wire PEG_Yvec_19__ap_idle;
  reg [1:0] PEG_Yvec_19__state;
  wire PEG_Yvec_20__ap_start_global__q0;
  wire PEG_Yvec_20__is_done__q0;
  wire PEG_Yvec_20__ap_done_global__q0;
  wire PEG_Yvec_20__ap_start;
  wire PEG_Yvec_20__ap_ready;
  wire PEG_Yvec_20__ap_done;
  wire PEG_Yvec_20__ap_idle;
  reg [1:0] PEG_Yvec_20__state;
  wire PEG_Yvec_21__ap_start_global__q0;
  wire PEG_Yvec_21__is_done__q0;
  wire PEG_Yvec_21__ap_done_global__q0;
  wire PEG_Yvec_21__ap_start;
  wire PEG_Yvec_21__ap_ready;
  wire PEG_Yvec_21__ap_done;
  wire PEG_Yvec_21__ap_idle;
  reg [1:0] PEG_Yvec_21__state;
  wire PEG_Yvec_22__ap_start_global__q0;
  wire PEG_Yvec_22__is_done__q0;
  wire PEG_Yvec_22__ap_done_global__q0;
  wire PEG_Yvec_22__ap_start;
  wire PEG_Yvec_22__ap_ready;
  wire PEG_Yvec_22__ap_done;
  wire PEG_Yvec_22__ap_idle;
  reg [1:0] PEG_Yvec_22__state;
  wire PEG_Yvec_23__ap_start_global__q0;
  wire PEG_Yvec_23__is_done__q0;
  wire PEG_Yvec_23__ap_done_global__q0;
  wire PEG_Yvec_23__ap_start;
  wire PEG_Yvec_23__ap_ready;
  wire PEG_Yvec_23__ap_done;
  wire PEG_Yvec_23__ap_idle;
  reg [1:0] PEG_Yvec_23__state;
  wire PEG_Yvec_24__ap_start_global__q0;
  wire PEG_Yvec_24__is_done__q0;
  wire PEG_Yvec_24__ap_done_global__q0;
  wire PEG_Yvec_24__ap_start;
  wire PEG_Yvec_24__ap_ready;
  wire PEG_Yvec_24__ap_done;
  wire PEG_Yvec_24__ap_idle;
  reg [1:0] PEG_Yvec_24__state;
  wire PEG_Yvec_25__ap_start_global__q0;
  wire PEG_Yvec_25__is_done__q0;
  wire PEG_Yvec_25__ap_done_global__q0;
  wire PEG_Yvec_25__ap_start;
  wire PEG_Yvec_25__ap_ready;
  wire PEG_Yvec_25__ap_done;
  wire PEG_Yvec_25__ap_idle;
  reg [1:0] PEG_Yvec_25__state;
  wire PEG_Yvec_26__ap_start_global__q0;
  wire PEG_Yvec_26__is_done__q0;
  wire PEG_Yvec_26__ap_done_global__q0;
  wire PEG_Yvec_26__ap_start;
  wire PEG_Yvec_26__ap_ready;
  wire PEG_Yvec_26__ap_done;
  wire PEG_Yvec_26__ap_idle;
  reg [1:0] PEG_Yvec_26__state;
  wire PEG_Yvec_27__ap_start_global__q0;
  wire PEG_Yvec_27__is_done__q0;
  wire PEG_Yvec_27__ap_done_global__q0;
  wire PEG_Yvec_27__ap_start;
  wire PEG_Yvec_27__ap_ready;
  wire PEG_Yvec_27__ap_done;
  wire PEG_Yvec_27__ap_idle;
  reg [1:0] PEG_Yvec_27__state;
  wire PEG_Yvec_28__ap_start_global__q0;
  wire PEG_Yvec_28__is_done__q0;
  wire PEG_Yvec_28__ap_done_global__q0;
  wire PEG_Yvec_28__ap_start;
  wire PEG_Yvec_28__ap_ready;
  wire PEG_Yvec_28__ap_done;
  wire PEG_Yvec_28__ap_idle;
  reg [1:0] PEG_Yvec_28__state;
  wire PEG_Yvec_29__ap_start_global__q0;
  wire PEG_Yvec_29__is_done__q0;
  wire PEG_Yvec_29__ap_done_global__q0;
  wire PEG_Yvec_29__ap_start;
  wire PEG_Yvec_29__ap_ready;
  wire PEG_Yvec_29__ap_done;
  wire PEG_Yvec_29__ap_idle;
  reg [1:0] PEG_Yvec_29__state;
  wire PEG_Yvec_30__ap_start_global__q0;
  wire PEG_Yvec_30__is_done__q0;
  wire PEG_Yvec_30__ap_done_global__q0;
  wire PEG_Yvec_30__ap_start;
  wire PEG_Yvec_30__ap_ready;
  wire PEG_Yvec_30__ap_done;
  wire PEG_Yvec_30__ap_idle;
  reg [1:0] PEG_Yvec_30__state;
  wire PEG_Yvec_31__ap_start_global__q0;
  wire PEG_Yvec_31__is_done__q0;
  wire PEG_Yvec_31__ap_done_global__q0;
  wire PEG_Yvec_31__ap_start;
  wire PEG_Yvec_31__ap_ready;
  wire PEG_Yvec_31__ap_done;
  wire PEG_Yvec_31__ap_idle;
  reg [1:0] PEG_Yvec_31__state;
  wire PEG_Yvec_32__ap_start_global__q0;
  wire PEG_Yvec_32__is_done__q0;
  wire PEG_Yvec_32__ap_done_global__q0;
  wire PEG_Yvec_32__ap_start;
  wire PEG_Yvec_32__ap_ready;
  wire PEG_Yvec_32__ap_done;
  wire PEG_Yvec_32__ap_idle;
  reg [1:0] PEG_Yvec_32__state;
  wire PEG_Yvec_33__ap_start_global__q0;
  wire PEG_Yvec_33__is_done__q0;
  wire PEG_Yvec_33__ap_done_global__q0;
  wire PEG_Yvec_33__ap_start;
  wire PEG_Yvec_33__ap_ready;
  wire PEG_Yvec_33__ap_done;
  wire PEG_Yvec_33__ap_idle;
  reg [1:0] PEG_Yvec_33__state;
  wire PEG_Yvec_34__ap_start_global__q0;
  wire PEG_Yvec_34__is_done__q0;
  wire PEG_Yvec_34__ap_done_global__q0;
  wire PEG_Yvec_34__ap_start;
  wire PEG_Yvec_34__ap_ready;
  wire PEG_Yvec_34__ap_done;
  wire PEG_Yvec_34__ap_idle;
  reg [1:0] PEG_Yvec_34__state;
  wire PEG_Yvec_35__ap_start_global__q0;
  wire PEG_Yvec_35__is_done__q0;
  wire PEG_Yvec_35__ap_done_global__q0;
  wire PEG_Yvec_35__ap_start;
  wire PEG_Yvec_35__ap_ready;
  wire PEG_Yvec_35__ap_done;
  wire PEG_Yvec_35__ap_idle;
  reg [1:0] PEG_Yvec_35__state;
  wire PEG_Yvec_36__ap_start_global__q0;
  wire PEG_Yvec_36__is_done__q0;
  wire PEG_Yvec_36__ap_done_global__q0;
  wire PEG_Yvec_36__ap_start;
  wire PEG_Yvec_36__ap_ready;
  wire PEG_Yvec_36__ap_done;
  wire PEG_Yvec_36__ap_idle;
  reg [1:0] PEG_Yvec_36__state;
  wire PEG_Yvec_37__ap_start_global__q0;
  wire PEG_Yvec_37__is_done__q0;
  wire PEG_Yvec_37__ap_done_global__q0;
  wire PEG_Yvec_37__ap_start;
  wire PEG_Yvec_37__ap_ready;
  wire PEG_Yvec_37__ap_done;
  wire PEG_Yvec_37__ap_idle;
  reg [1:0] PEG_Yvec_37__state;
  wire PEG_Yvec_38__ap_start_global__q0;
  wire PEG_Yvec_38__is_done__q0;
  wire PEG_Yvec_38__ap_done_global__q0;
  wire PEG_Yvec_38__ap_start;
  wire PEG_Yvec_38__ap_ready;
  wire PEG_Yvec_38__ap_done;
  wire PEG_Yvec_38__ap_idle;
  reg [1:0] PEG_Yvec_38__state;
  wire PEG_Yvec_39__ap_start_global__q0;
  wire PEG_Yvec_39__is_done__q0;
  wire PEG_Yvec_39__ap_done_global__q0;
  wire PEG_Yvec_39__ap_start;
  wire PEG_Yvec_39__ap_ready;
  wire PEG_Yvec_39__ap_done;
  wire PEG_Yvec_39__ap_idle;
  reg [1:0] PEG_Yvec_39__state;
  wire PEG_Yvec_40__ap_start_global__q0;
  wire PEG_Yvec_40__is_done__q0;
  wire PEG_Yvec_40__ap_done_global__q0;
  wire PEG_Yvec_40__ap_start;
  wire PEG_Yvec_40__ap_ready;
  wire PEG_Yvec_40__ap_done;
  wire PEG_Yvec_40__ap_idle;
  reg [1:0] PEG_Yvec_40__state;
  wire PEG_Yvec_41__ap_start_global__q0;
  wire PEG_Yvec_41__is_done__q0;
  wire PEG_Yvec_41__ap_done_global__q0;
  wire PEG_Yvec_41__ap_start;
  wire PEG_Yvec_41__ap_ready;
  wire PEG_Yvec_41__ap_done;
  wire PEG_Yvec_41__ap_idle;
  reg [1:0] PEG_Yvec_41__state;
  wire PEG_Yvec_42__ap_start_global__q0;
  wire PEG_Yvec_42__is_done__q0;
  wire PEG_Yvec_42__ap_done_global__q0;
  wire PEG_Yvec_42__ap_start;
  wire PEG_Yvec_42__ap_ready;
  wire PEG_Yvec_42__ap_done;
  wire PEG_Yvec_42__ap_idle;
  reg [1:0] PEG_Yvec_42__state;
  wire PEG_Yvec_43__ap_start_global__q0;
  wire PEG_Yvec_43__is_done__q0;
  wire PEG_Yvec_43__ap_done_global__q0;
  wire PEG_Yvec_43__ap_start;
  wire PEG_Yvec_43__ap_ready;
  wire PEG_Yvec_43__ap_done;
  wire PEG_Yvec_43__ap_idle;
  reg [1:0] PEG_Yvec_43__state;
  wire PEG_Yvec_44__ap_start_global__q0;
  wire PEG_Yvec_44__is_done__q0;
  wire PEG_Yvec_44__ap_done_global__q0;
  wire PEG_Yvec_44__ap_start;
  wire PEG_Yvec_44__ap_ready;
  wire PEG_Yvec_44__ap_done;
  wire PEG_Yvec_44__ap_idle;
  reg [1:0] PEG_Yvec_44__state;
  wire PEG_Yvec_45__ap_start_global__q0;
  wire PEG_Yvec_45__is_done__q0;
  wire PEG_Yvec_45__ap_done_global__q0;
  wire PEG_Yvec_45__ap_start;
  wire PEG_Yvec_45__ap_ready;
  wire PEG_Yvec_45__ap_done;
  wire PEG_Yvec_45__ap_idle;
  reg [1:0] PEG_Yvec_45__state;
  wire PEG_Yvec_46__ap_start_global__q0;
  wire PEG_Yvec_46__is_done__q0;
  wire PEG_Yvec_46__ap_done_global__q0;
  wire PEG_Yvec_46__ap_start;
  wire PEG_Yvec_46__ap_ready;
  wire PEG_Yvec_46__ap_done;
  wire PEG_Yvec_46__ap_idle;
  reg [1:0] PEG_Yvec_46__state;
  wire PEG_Yvec_47__ap_start_global__q0;
  wire PEG_Yvec_47__is_done__q0;
  wire PEG_Yvec_47__ap_done_global__q0;
  wire PEG_Yvec_47__ap_start;
  wire PEG_Yvec_47__ap_ready;
  wire PEG_Yvec_47__ap_done;
  wire PEG_Yvec_47__ap_idle;
  reg [1:0] PEG_Yvec_47__state;
  wire PEG_Yvec_48__ap_start_global__q0;
  wire PEG_Yvec_48__is_done__q0;
  wire PEG_Yvec_48__ap_done_global__q0;
  wire PEG_Yvec_48__ap_start;
  wire PEG_Yvec_48__ap_ready;
  wire PEG_Yvec_48__ap_done;
  wire PEG_Yvec_48__ap_idle;
  reg [1:0] PEG_Yvec_48__state;
  wire PEG_Yvec_49__ap_start_global__q0;
  wire PEG_Yvec_49__is_done__q0;
  wire PEG_Yvec_49__ap_done_global__q0;
  wire PEG_Yvec_49__ap_start;
  wire PEG_Yvec_49__ap_ready;
  wire PEG_Yvec_49__ap_done;
  wire PEG_Yvec_49__ap_idle;
  reg [1:0] PEG_Yvec_49__state;
  wire PEG_Yvec_50__ap_start_global__q0;
  wire PEG_Yvec_50__is_done__q0;
  wire PEG_Yvec_50__ap_done_global__q0;
  wire PEG_Yvec_50__ap_start;
  wire PEG_Yvec_50__ap_ready;
  wire PEG_Yvec_50__ap_done;
  wire PEG_Yvec_50__ap_idle;
  reg [1:0] PEG_Yvec_50__state;
  wire PEG_Yvec_51__ap_start_global__q0;
  wire PEG_Yvec_51__is_done__q0;
  wire PEG_Yvec_51__ap_done_global__q0;
  wire PEG_Yvec_51__ap_start;
  wire PEG_Yvec_51__ap_ready;
  wire PEG_Yvec_51__ap_done;
  wire PEG_Yvec_51__ap_idle;
  reg [1:0] PEG_Yvec_51__state;
  wire PEG_Yvec_52__ap_start_global__q0;
  wire PEG_Yvec_52__is_done__q0;
  wire PEG_Yvec_52__ap_done_global__q0;
  wire PEG_Yvec_52__ap_start;
  wire PEG_Yvec_52__ap_ready;
  wire PEG_Yvec_52__ap_done;
  wire PEG_Yvec_52__ap_idle;
  reg [1:0] PEG_Yvec_52__state;
  wire PEG_Yvec_53__ap_start_global__q0;
  wire PEG_Yvec_53__is_done__q0;
  wire PEG_Yvec_53__ap_done_global__q0;
  wire PEG_Yvec_53__ap_start;
  wire PEG_Yvec_53__ap_ready;
  wire PEG_Yvec_53__ap_done;
  wire PEG_Yvec_53__ap_idle;
  reg [1:0] PEG_Yvec_53__state;
  wire PEG_Yvec_54__ap_start_global__q0;
  wire PEG_Yvec_54__is_done__q0;
  wire PEG_Yvec_54__ap_done_global__q0;
  wire PEG_Yvec_54__ap_start;
  wire PEG_Yvec_54__ap_ready;
  wire PEG_Yvec_54__ap_done;
  wire PEG_Yvec_54__ap_idle;
  reg [1:0] PEG_Yvec_54__state;
  wire PEG_Yvec_55__ap_start_global__q0;
  wire PEG_Yvec_55__is_done__q0;
  wire PEG_Yvec_55__ap_done_global__q0;
  wire PEG_Yvec_55__ap_start;
  wire PEG_Yvec_55__ap_ready;
  wire PEG_Yvec_55__ap_done;
  wire PEG_Yvec_55__ap_idle;
  reg [1:0] PEG_Yvec_55__state;
  wire black_hole_float_v16_0__ap_start_global__q0;
  reg black_hole_float_v16_0__ap_start;
  wire black_hole_int_0__ap_start_global__q0;
  reg black_hole_int_0__ap_start;
  wire read_A_0__ap_start_global__q0;
  wire read_A_0__is_done__q0;
  wire read_A_0__ap_done_global__q0;
  wire read_A_0__ap_start;
  wire read_A_0__ap_ready;
  wire read_A_0__ap_done;
  wire read_A_0__ap_idle;
  reg [1:0] read_A_0__state;
  wire read_A_1__ap_start_global__q0;
  wire read_A_1__is_done__q0;
  wire read_A_1__ap_done_global__q0;
  wire read_A_1__ap_start;
  wire read_A_1__ap_ready;
  wire read_A_1__ap_done;
  wire read_A_1__ap_idle;
  reg [1:0] read_A_1__state;
  wire read_A_2__ap_start_global__q0;
  wire read_A_2__is_done__q0;
  wire read_A_2__ap_done_global__q0;
  wire read_A_2__ap_start;
  wire read_A_2__ap_ready;
  wire read_A_2__ap_done;
  wire read_A_2__ap_idle;
  reg [1:0] read_A_2__state;
  wire read_A_3__ap_start_global__q0;
  wire read_A_3__is_done__q0;
  wire read_A_3__ap_done_global__q0;
  wire read_A_3__ap_start;
  wire read_A_3__ap_ready;
  wire read_A_3__ap_done;
  wire read_A_3__ap_idle;
  reg [1:0] read_A_3__state;
  wire read_A_4__ap_start_global__q0;
  wire read_A_4__is_done__q0;
  wire read_A_4__ap_done_global__q0;
  wire read_A_4__ap_start;
  wire read_A_4__ap_ready;
  wire read_A_4__ap_done;
  wire read_A_4__ap_idle;
  reg [1:0] read_A_4__state;
  wire read_A_5__ap_start_global__q0;
  wire read_A_5__is_done__q0;
  wire read_A_5__ap_done_global__q0;
  wire read_A_5__ap_start;
  wire read_A_5__ap_ready;
  wire read_A_5__ap_done;
  wire read_A_5__ap_idle;
  reg [1:0] read_A_5__state;
  wire read_A_6__ap_start_global__q0;
  wire read_A_6__is_done__q0;
  wire read_A_6__ap_done_global__q0;
  wire read_A_6__ap_start;
  wire read_A_6__ap_ready;
  wire read_A_6__ap_done;
  wire read_A_6__ap_idle;
  reg [1:0] read_A_6__state;
  wire read_A_7__ap_start_global__q0;
  wire read_A_7__is_done__q0;
  wire read_A_7__ap_done_global__q0;
  wire read_A_7__ap_start;
  wire read_A_7__ap_ready;
  wire read_A_7__ap_done;
  wire read_A_7__ap_idle;
  reg [1:0] read_A_7__state;
  wire read_A_8__ap_start_global__q0;
  wire read_A_8__is_done__q0;
  wire read_A_8__ap_done_global__q0;
  wire read_A_8__ap_start;
  wire read_A_8__ap_ready;
  wire read_A_8__ap_done;
  wire read_A_8__ap_idle;
  reg [1:0] read_A_8__state;
  wire read_A_9__ap_start_global__q0;
  wire read_A_9__is_done__q0;
  wire read_A_9__ap_done_global__q0;
  wire read_A_9__ap_start;
  wire read_A_9__ap_ready;
  wire read_A_9__ap_done;
  wire read_A_9__ap_idle;
  reg [1:0] read_A_9__state;
  wire read_A_10__ap_start_global__q0;
  wire read_A_10__is_done__q0;
  wire read_A_10__ap_done_global__q0;
  wire read_A_10__ap_start;
  wire read_A_10__ap_ready;
  wire read_A_10__ap_done;
  wire read_A_10__ap_idle;
  reg [1:0] read_A_10__state;
  wire read_A_11__ap_start_global__q0;
  wire read_A_11__is_done__q0;
  wire read_A_11__ap_done_global__q0;
  wire read_A_11__ap_start;
  wire read_A_11__ap_ready;
  wire read_A_11__ap_done;
  wire read_A_11__ap_idle;
  reg [1:0] read_A_11__state;
  wire read_A_12__ap_start_global__q0;
  wire read_A_12__is_done__q0;
  wire read_A_12__ap_done_global__q0;
  wire read_A_12__ap_start;
  wire read_A_12__ap_ready;
  wire read_A_12__ap_done;
  wire read_A_12__ap_idle;
  reg [1:0] read_A_12__state;
  wire read_A_13__ap_start_global__q0;
  wire read_A_13__is_done__q0;
  wire read_A_13__ap_done_global__q0;
  wire read_A_13__ap_start;
  wire read_A_13__ap_ready;
  wire read_A_13__ap_done;
  wire read_A_13__ap_idle;
  reg [1:0] read_A_13__state;
  wire read_A_14__ap_start_global__q0;
  wire read_A_14__is_done__q0;
  wire read_A_14__ap_done_global__q0;
  wire read_A_14__ap_start;
  wire read_A_14__ap_ready;
  wire read_A_14__ap_done;
  wire read_A_14__ap_idle;
  reg [1:0] read_A_14__state;
  wire read_A_15__ap_start_global__q0;
  wire read_A_15__is_done__q0;
  wire read_A_15__ap_done_global__q0;
  wire read_A_15__ap_start;
  wire read_A_15__ap_ready;
  wire read_A_15__ap_done;
  wire read_A_15__ap_idle;
  reg [1:0] read_A_15__state;
  wire read_A_16__ap_start_global__q0;
  wire read_A_16__is_done__q0;
  wire read_A_16__ap_done_global__q0;
  wire read_A_16__ap_start;
  wire read_A_16__ap_ready;
  wire read_A_16__ap_done;
  wire read_A_16__ap_idle;
  reg [1:0] read_A_16__state;
  wire read_A_17__ap_start_global__q0;
  wire read_A_17__is_done__q0;
  wire read_A_17__ap_done_global__q0;
  wire read_A_17__ap_start;
  wire read_A_17__ap_ready;
  wire read_A_17__ap_done;
  wire read_A_17__ap_idle;
  reg [1:0] read_A_17__state;
  wire read_A_18__ap_start_global__q0;
  wire read_A_18__is_done__q0;
  wire read_A_18__ap_done_global__q0;
  wire read_A_18__ap_start;
  wire read_A_18__ap_ready;
  wire read_A_18__ap_done;
  wire read_A_18__ap_idle;
  reg [1:0] read_A_18__state;
  wire read_A_19__ap_start_global__q0;
  wire read_A_19__is_done__q0;
  wire read_A_19__ap_done_global__q0;
  wire read_A_19__ap_start;
  wire read_A_19__ap_ready;
  wire read_A_19__ap_done;
  wire read_A_19__ap_idle;
  reg [1:0] read_A_19__state;
  wire read_A_20__ap_start_global__q0;
  wire read_A_20__is_done__q0;
  wire read_A_20__ap_done_global__q0;
  wire read_A_20__ap_start;
  wire read_A_20__ap_ready;
  wire read_A_20__ap_done;
  wire read_A_20__ap_idle;
  reg [1:0] read_A_20__state;
  wire read_A_21__ap_start_global__q0;
  wire read_A_21__is_done__q0;
  wire read_A_21__ap_done_global__q0;
  wire read_A_21__ap_start;
  wire read_A_21__ap_ready;
  wire read_A_21__ap_done;
  wire read_A_21__ap_idle;
  reg [1:0] read_A_21__state;
  wire read_A_22__ap_start_global__q0;
  wire read_A_22__is_done__q0;
  wire read_A_22__ap_done_global__q0;
  wire read_A_22__ap_start;
  wire read_A_22__ap_ready;
  wire read_A_22__ap_done;
  wire read_A_22__ap_idle;
  reg [1:0] read_A_22__state;
  wire read_A_23__ap_start_global__q0;
  wire read_A_23__is_done__q0;
  wire read_A_23__ap_done_global__q0;
  wire read_A_23__ap_start;
  wire read_A_23__ap_ready;
  wire read_A_23__ap_done;
  wire read_A_23__ap_idle;
  reg [1:0] read_A_23__state;
  wire read_A_24__ap_start_global__q0;
  wire read_A_24__is_done__q0;
  wire read_A_24__ap_done_global__q0;
  wire read_A_24__ap_start;
  wire read_A_24__ap_ready;
  wire read_A_24__ap_done;
  wire read_A_24__ap_idle;
  reg [1:0] read_A_24__state;
  wire read_A_25__ap_start_global__q0;
  wire read_A_25__is_done__q0;
  wire read_A_25__ap_done_global__q0;
  wire read_A_25__ap_start;
  wire read_A_25__ap_ready;
  wire read_A_25__ap_done;
  wire read_A_25__ap_idle;
  reg [1:0] read_A_25__state;
  wire read_A_26__ap_start_global__q0;
  wire read_A_26__is_done__q0;
  wire read_A_26__ap_done_global__q0;
  wire read_A_26__ap_start;
  wire read_A_26__ap_ready;
  wire read_A_26__ap_done;
  wire read_A_26__ap_idle;
  reg [1:0] read_A_26__state;
  wire read_A_27__ap_start_global__q0;
  wire read_A_27__is_done__q0;
  wire read_A_27__ap_done_global__q0;
  wire read_A_27__ap_start;
  wire read_A_27__ap_ready;
  wire read_A_27__ap_done;
  wire read_A_27__ap_idle;
  reg [1:0] read_A_27__state;
  wire read_A_28__ap_start_global__q0;
  wire read_A_28__is_done__q0;
  wire read_A_28__ap_done_global__q0;
  wire read_A_28__ap_start;
  wire read_A_28__ap_ready;
  wire read_A_28__ap_done;
  wire read_A_28__ap_idle;
  reg [1:0] read_A_28__state;
  wire read_A_29__ap_start_global__q0;
  wire read_A_29__is_done__q0;
  wire read_A_29__ap_done_global__q0;
  wire read_A_29__ap_start;
  wire read_A_29__ap_ready;
  wire read_A_29__ap_done;
  wire read_A_29__ap_idle;
  reg [1:0] read_A_29__state;
  wire read_A_30__ap_start_global__q0;
  wire read_A_30__is_done__q0;
  wire read_A_30__ap_done_global__q0;
  wire read_A_30__ap_start;
  wire read_A_30__ap_ready;
  wire read_A_30__ap_done;
  wire read_A_30__ap_idle;
  reg [1:0] read_A_30__state;
  wire read_A_31__ap_start_global__q0;
  wire read_A_31__is_done__q0;
  wire read_A_31__ap_done_global__q0;
  wire read_A_31__ap_start;
  wire read_A_31__ap_ready;
  wire read_A_31__ap_done;
  wire read_A_31__ap_idle;
  reg [1:0] read_A_31__state;
  wire read_A_32__ap_start_global__q0;
  wire read_A_32__is_done__q0;
  wire read_A_32__ap_done_global__q0;
  wire read_A_32__ap_start;
  wire read_A_32__ap_ready;
  wire read_A_32__ap_done;
  wire read_A_32__ap_idle;
  reg [1:0] read_A_32__state;
  wire read_A_33__ap_start_global__q0;
  wire read_A_33__is_done__q0;
  wire read_A_33__ap_done_global__q0;
  wire read_A_33__ap_start;
  wire read_A_33__ap_ready;
  wire read_A_33__ap_done;
  wire read_A_33__ap_idle;
  reg [1:0] read_A_33__state;
  wire read_A_34__ap_start_global__q0;
  wire read_A_34__is_done__q0;
  wire read_A_34__ap_done_global__q0;
  wire read_A_34__ap_start;
  wire read_A_34__ap_ready;
  wire read_A_34__ap_done;
  wire read_A_34__ap_idle;
  reg [1:0] read_A_34__state;
  wire read_A_35__ap_start_global__q0;
  wire read_A_35__is_done__q0;
  wire read_A_35__ap_done_global__q0;
  wire read_A_35__ap_start;
  wire read_A_35__ap_ready;
  wire read_A_35__ap_done;
  wire read_A_35__ap_idle;
  reg [1:0] read_A_35__state;
  wire read_A_36__ap_start_global__q0;
  wire read_A_36__is_done__q0;
  wire read_A_36__ap_done_global__q0;
  wire read_A_36__ap_start;
  wire read_A_36__ap_ready;
  wire read_A_36__ap_done;
  wire read_A_36__ap_idle;
  reg [1:0] read_A_36__state;
  wire read_A_37__ap_start_global__q0;
  wire read_A_37__is_done__q0;
  wire read_A_37__ap_done_global__q0;
  wire read_A_37__ap_start;
  wire read_A_37__ap_ready;
  wire read_A_37__ap_done;
  wire read_A_37__ap_idle;
  reg [1:0] read_A_37__state;
  wire read_A_38__ap_start_global__q0;
  wire read_A_38__is_done__q0;
  wire read_A_38__ap_done_global__q0;
  wire read_A_38__ap_start;
  wire read_A_38__ap_ready;
  wire read_A_38__ap_done;
  wire read_A_38__ap_idle;
  reg [1:0] read_A_38__state;
  wire read_A_39__ap_start_global__q0;
  wire read_A_39__is_done__q0;
  wire read_A_39__ap_done_global__q0;
  wire read_A_39__ap_start;
  wire read_A_39__ap_ready;
  wire read_A_39__ap_done;
  wire read_A_39__ap_idle;
  reg [1:0] read_A_39__state;
  wire read_A_40__ap_start_global__q0;
  wire read_A_40__is_done__q0;
  wire read_A_40__ap_done_global__q0;
  wire read_A_40__ap_start;
  wire read_A_40__ap_ready;
  wire read_A_40__ap_done;
  wire read_A_40__ap_idle;
  reg [1:0] read_A_40__state;
  wire read_A_41__ap_start_global__q0;
  wire read_A_41__is_done__q0;
  wire read_A_41__ap_done_global__q0;
  wire read_A_41__ap_start;
  wire read_A_41__ap_ready;
  wire read_A_41__ap_done;
  wire read_A_41__ap_idle;
  reg [1:0] read_A_41__state;
  wire read_A_42__ap_start_global__q0;
  wire read_A_42__is_done__q0;
  wire read_A_42__ap_done_global__q0;
  wire read_A_42__ap_start;
  wire read_A_42__ap_ready;
  wire read_A_42__ap_done;
  wire read_A_42__ap_idle;
  reg [1:0] read_A_42__state;
  wire read_A_43__ap_start_global__q0;
  wire read_A_43__is_done__q0;
  wire read_A_43__ap_done_global__q0;
  wire read_A_43__ap_start;
  wire read_A_43__ap_ready;
  wire read_A_43__ap_done;
  wire read_A_43__ap_idle;
  reg [1:0] read_A_43__state;
  wire read_A_44__ap_start_global__q0;
  wire read_A_44__is_done__q0;
  wire read_A_44__ap_done_global__q0;
  wire read_A_44__ap_start;
  wire read_A_44__ap_ready;
  wire read_A_44__ap_done;
  wire read_A_44__ap_idle;
  reg [1:0] read_A_44__state;
  wire read_A_45__ap_start_global__q0;
  wire read_A_45__is_done__q0;
  wire read_A_45__ap_done_global__q0;
  wire read_A_45__ap_start;
  wire read_A_45__ap_ready;
  wire read_A_45__ap_done;
  wire read_A_45__ap_idle;
  reg [1:0] read_A_45__state;
  wire read_A_46__ap_start_global__q0;
  wire read_A_46__is_done__q0;
  wire read_A_46__ap_done_global__q0;
  wire read_A_46__ap_start;
  wire read_A_46__ap_ready;
  wire read_A_46__ap_done;
  wire read_A_46__ap_idle;
  reg [1:0] read_A_46__state;
  wire read_A_47__ap_start_global__q0;
  wire read_A_47__is_done__q0;
  wire read_A_47__ap_done_global__q0;
  wire read_A_47__ap_start;
  wire read_A_47__ap_ready;
  wire read_A_47__ap_done;
  wire read_A_47__ap_idle;
  reg [1:0] read_A_47__state;
  wire read_A_48__ap_start_global__q0;
  wire read_A_48__is_done__q0;
  wire read_A_48__ap_done_global__q0;
  wire read_A_48__ap_start;
  wire read_A_48__ap_ready;
  wire read_A_48__ap_done;
  wire read_A_48__ap_idle;
  reg [1:0] read_A_48__state;
  wire read_A_49__ap_start_global__q0;
  wire read_A_49__is_done__q0;
  wire read_A_49__ap_done_global__q0;
  wire read_A_49__ap_start;
  wire read_A_49__ap_ready;
  wire read_A_49__ap_done;
  wire read_A_49__ap_idle;
  reg [1:0] read_A_49__state;
  wire read_A_50__ap_start_global__q0;
  wire read_A_50__is_done__q0;
  wire read_A_50__ap_done_global__q0;
  wire read_A_50__ap_start;
  wire read_A_50__ap_ready;
  wire read_A_50__ap_done;
  wire read_A_50__ap_idle;
  reg [1:0] read_A_50__state;
  wire read_A_51__ap_start_global__q0;
  wire read_A_51__is_done__q0;
  wire read_A_51__ap_done_global__q0;
  wire read_A_51__ap_start;
  wire read_A_51__ap_ready;
  wire read_A_51__ap_done;
  wire read_A_51__ap_idle;
  reg [1:0] read_A_51__state;
  wire read_A_52__ap_start_global__q0;
  wire read_A_52__is_done__q0;
  wire read_A_52__ap_done_global__q0;
  wire read_A_52__ap_start;
  wire read_A_52__ap_ready;
  wire read_A_52__ap_done;
  wire read_A_52__ap_idle;
  reg [1:0] read_A_52__state;
  wire read_A_53__ap_start_global__q0;
  wire read_A_53__is_done__q0;
  wire read_A_53__ap_done_global__q0;
  wire read_A_53__ap_start;
  wire read_A_53__ap_ready;
  wire read_A_53__ap_done;
  wire read_A_53__ap_idle;
  reg [1:0] read_A_53__state;
  wire read_A_54__ap_start_global__q0;
  wire read_A_54__is_done__q0;
  wire read_A_54__ap_done_global__q0;
  wire read_A_54__ap_start;
  wire read_A_54__ap_ready;
  wire read_A_54__ap_done;
  wire read_A_54__ap_idle;
  reg [1:0] read_A_54__state;
  wire read_A_55__ap_start_global__q0;
  wire read_A_55__is_done__q0;
  wire read_A_55__ap_done_global__q0;
  wire read_A_55__ap_start;
  wire read_A_55__ap_ready;
  wire read_A_55__ap_done;
  wire read_A_55__ap_idle;
  reg [1:0] read_A_55__state;
  wire read_X_0__ap_start_global__q0;
  wire read_X_0__is_done__q0;
  wire read_X_0__ap_done_global__q0;
  wire read_X_0__ap_start;
  wire read_X_0__ap_ready;
  wire read_X_0__ap_done;
  wire read_X_0__ap_idle;
  reg [1:0] read_X_0__state;
  wire read_Y_0__ap_start_global__q0;
  wire read_Y_0__is_done__q0;
  wire read_Y_0__ap_done_global__q0;
  wire read_Y_0__ap_start;
  wire read_Y_0__ap_ready;
  wire read_Y_0__ap_done;
  wire read_Y_0__ap_idle;
  reg [1:0] read_Y_0__state;
  wire read_edge_list_ptr_0__ap_start_global__q0;
  wire read_edge_list_ptr_0__is_done__q0;
  wire read_edge_list_ptr_0__ap_done_global__q0;
  wire read_edge_list_ptr_0__ap_start;
  wire read_edge_list_ptr_0__ap_ready;
  wire read_edge_list_ptr_0__ap_done;
  wire read_edge_list_ptr_0__ap_idle;
  reg [1:0] read_edge_list_ptr_0__state;
  wire write_Y_0__ap_start_global__q0;
  wire write_Y_0__is_done__q0;
  wire write_Y_0__ap_done_global__q0;
  wire write_Y_0__ap_start;
  wire write_Y_0__ap_ready;
  wire write_Y_0__ap_done;
  wire write_Y_0__ap_idle;
  reg [1:0] write_Y_0__state;
  reg [1:0] tapa_state;
  reg [0:0] countdown;
  wire ap_start__q0;
  wire ap_done__q0;
  assign Arbiter_Y_0__ap_start_global__q0 = ap_start__q0;
  assign Arbiter_Y_0__is_done__q0 = (Arbiter_Y_0__state == 2'b10);
  assign Arbiter_Y_0__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Arbiter_Y_0__state <= 2'b00;
    end else begin
      if(Arbiter_Y_0__state == 2'b00) begin
        if(Arbiter_Y_0__ap_start_global__q0) begin
          Arbiter_Y_0__state <= 2'b01;
        end 
      end 
      if(Arbiter_Y_0__state == 2'b01) begin
        if(Arbiter_Y_0__ap_ready) begin
          if(Arbiter_Y_0__ap_done) begin
            Arbiter_Y_0__state <= 2'b10;
          end else begin
            Arbiter_Y_0__state <= 2'b11;
          end
        end 
      end 
      if(Arbiter_Y_0__state == 2'b11) begin
        if(Arbiter_Y_0__ap_done) begin
          Arbiter_Y_0__state <= 2'b10;
        end 
      end 
      if(Arbiter_Y_0__state == 2'b10) begin
        if(Arbiter_Y_0__ap_done_global__q0) begin
          Arbiter_Y_0__state <= 2'b00;
        end 
      end 
    end
  end
  assign Arbiter_Y_0__ap_start = (Arbiter_Y_0__state == 2'b01);
  assign Arbiter_Y_1__ap_start_global__q0 = ap_start__q0;
  assign Arbiter_Y_1__is_done__q0 = (Arbiter_Y_1__state == 2'b10);
  assign Arbiter_Y_1__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Arbiter_Y_1__state <= 2'b00;
    end else begin
      if(Arbiter_Y_1__state == 2'b00) begin
        if(Arbiter_Y_1__ap_start_global__q0) begin
          Arbiter_Y_1__state <= 2'b01;
        end 
      end 
      if(Arbiter_Y_1__state == 2'b01) begin
        if(Arbiter_Y_1__ap_ready) begin
          if(Arbiter_Y_1__ap_done) begin
            Arbiter_Y_1__state <= 2'b10;
          end else begin
            Arbiter_Y_1__state <= 2'b11;
          end
        end 
      end 
      if(Arbiter_Y_1__state == 2'b11) begin
        if(Arbiter_Y_1__ap_done) begin
          Arbiter_Y_1__state <= 2'b10;
        end 
      end 
      if(Arbiter_Y_1__state == 2'b10) begin
        if(Arbiter_Y_1__ap_done_global__q0) begin
          Arbiter_Y_1__state <= 2'b00;
        end 
      end 
    end
  end
  assign Arbiter_Y_1__ap_start = (Arbiter_Y_1__state == 2'b01);
  assign Arbiter_Y_2__ap_start_global__q0 = ap_start__q0;
  assign Arbiter_Y_2__is_done__q0 = (Arbiter_Y_2__state == 2'b10);
  assign Arbiter_Y_2__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Arbiter_Y_2__state <= 2'b00;
    end else begin
      if(Arbiter_Y_2__state == 2'b00) begin
        if(Arbiter_Y_2__ap_start_global__q0) begin
          Arbiter_Y_2__state <= 2'b01;
        end 
      end 
      if(Arbiter_Y_2__state == 2'b01) begin
        if(Arbiter_Y_2__ap_ready) begin
          if(Arbiter_Y_2__ap_done) begin
            Arbiter_Y_2__state <= 2'b10;
          end else begin
            Arbiter_Y_2__state <= 2'b11;
          end
        end 
      end 
      if(Arbiter_Y_2__state == 2'b11) begin
        if(Arbiter_Y_2__ap_done) begin
          Arbiter_Y_2__state <= 2'b10;
        end 
      end 
      if(Arbiter_Y_2__state == 2'b10) begin
        if(Arbiter_Y_2__ap_done_global__q0) begin
          Arbiter_Y_2__state <= 2'b00;
        end 
      end 
    end
  end
  assign Arbiter_Y_2__ap_start = (Arbiter_Y_2__state == 2'b01);
  assign Arbiter_Y_3__ap_start_global__q0 = ap_start__q0;
  assign Arbiter_Y_3__is_done__q0 = (Arbiter_Y_3__state == 2'b10);
  assign Arbiter_Y_3__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Arbiter_Y_3__state <= 2'b00;
    end else begin
      if(Arbiter_Y_3__state == 2'b00) begin
        if(Arbiter_Y_3__ap_start_global__q0) begin
          Arbiter_Y_3__state <= 2'b01;
        end 
      end 
      if(Arbiter_Y_3__state == 2'b01) begin
        if(Arbiter_Y_3__ap_ready) begin
          if(Arbiter_Y_3__ap_done) begin
            Arbiter_Y_3__state <= 2'b10;
          end else begin
            Arbiter_Y_3__state <= 2'b11;
          end
        end 
      end 
      if(Arbiter_Y_3__state == 2'b11) begin
        if(Arbiter_Y_3__ap_done) begin
          Arbiter_Y_3__state <= 2'b10;
        end 
      end 
      if(Arbiter_Y_3__state == 2'b10) begin
        if(Arbiter_Y_3__ap_done_global__q0) begin
          Arbiter_Y_3__state <= 2'b00;
        end 
      end 
    end
  end
  assign Arbiter_Y_3__ap_start = (Arbiter_Y_3__state == 2'b01);
  assign Arbiter_Y_4__ap_start_global__q0 = ap_start__q0;
  assign Arbiter_Y_4__is_done__q0 = (Arbiter_Y_4__state == 2'b10);
  assign Arbiter_Y_4__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Arbiter_Y_4__state <= 2'b00;
    end else begin
      if(Arbiter_Y_4__state == 2'b00) begin
        if(Arbiter_Y_4__ap_start_global__q0) begin
          Arbiter_Y_4__state <= 2'b01;
        end 
      end 
      if(Arbiter_Y_4__state == 2'b01) begin
        if(Arbiter_Y_4__ap_ready) begin
          if(Arbiter_Y_4__ap_done) begin
            Arbiter_Y_4__state <= 2'b10;
          end else begin
            Arbiter_Y_4__state <= 2'b11;
          end
        end 
      end 
      if(Arbiter_Y_4__state == 2'b11) begin
        if(Arbiter_Y_4__ap_done) begin
          Arbiter_Y_4__state <= 2'b10;
        end 
      end 
      if(Arbiter_Y_4__state == 2'b10) begin
        if(Arbiter_Y_4__ap_done_global__q0) begin
          Arbiter_Y_4__state <= 2'b00;
        end 
      end 
    end
  end
  assign Arbiter_Y_4__ap_start = (Arbiter_Y_4__state == 2'b01);
  assign Arbiter_Y_5__ap_start_global__q0 = ap_start__q0;
  assign Arbiter_Y_5__is_done__q0 = (Arbiter_Y_5__state == 2'b10);
  assign Arbiter_Y_5__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Arbiter_Y_5__state <= 2'b00;
    end else begin
      if(Arbiter_Y_5__state == 2'b00) begin
        if(Arbiter_Y_5__ap_start_global__q0) begin
          Arbiter_Y_5__state <= 2'b01;
        end 
      end 
      if(Arbiter_Y_5__state == 2'b01) begin
        if(Arbiter_Y_5__ap_ready) begin
          if(Arbiter_Y_5__ap_done) begin
            Arbiter_Y_5__state <= 2'b10;
          end else begin
            Arbiter_Y_5__state <= 2'b11;
          end
        end 
      end 
      if(Arbiter_Y_5__state == 2'b11) begin
        if(Arbiter_Y_5__ap_done) begin
          Arbiter_Y_5__state <= 2'b10;
        end 
      end 
      if(Arbiter_Y_5__state == 2'b10) begin
        if(Arbiter_Y_5__ap_done_global__q0) begin
          Arbiter_Y_5__state <= 2'b00;
        end 
      end 
    end
  end
  assign Arbiter_Y_5__ap_start = (Arbiter_Y_5__state == 2'b01);
  assign Arbiter_Y_6__ap_start_global__q0 = ap_start__q0;
  assign Arbiter_Y_6__is_done__q0 = (Arbiter_Y_6__state == 2'b10);
  assign Arbiter_Y_6__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Arbiter_Y_6__state <= 2'b00;
    end else begin
      if(Arbiter_Y_6__state == 2'b00) begin
        if(Arbiter_Y_6__ap_start_global__q0) begin
          Arbiter_Y_6__state <= 2'b01;
        end 
      end 
      if(Arbiter_Y_6__state == 2'b01) begin
        if(Arbiter_Y_6__ap_ready) begin
          if(Arbiter_Y_6__ap_done) begin
            Arbiter_Y_6__state <= 2'b10;
          end else begin
            Arbiter_Y_6__state <= 2'b11;
          end
        end 
      end 
      if(Arbiter_Y_6__state == 2'b11) begin
        if(Arbiter_Y_6__ap_done) begin
          Arbiter_Y_6__state <= 2'b10;
        end 
      end 
      if(Arbiter_Y_6__state == 2'b10) begin
        if(Arbiter_Y_6__ap_done_global__q0) begin
          Arbiter_Y_6__state <= 2'b00;
        end 
      end 
    end
  end
  assign Arbiter_Y_6__ap_start = (Arbiter_Y_6__state == 2'b01);
  assign Arbiter_Y_7__ap_start_global__q0 = ap_start__q0;
  assign Arbiter_Y_7__is_done__q0 = (Arbiter_Y_7__state == 2'b10);
  assign Arbiter_Y_7__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Arbiter_Y_7__state <= 2'b00;
    end else begin
      if(Arbiter_Y_7__state == 2'b00) begin
        if(Arbiter_Y_7__ap_start_global__q0) begin
          Arbiter_Y_7__state <= 2'b01;
        end 
      end 
      if(Arbiter_Y_7__state == 2'b01) begin
        if(Arbiter_Y_7__ap_ready) begin
          if(Arbiter_Y_7__ap_done) begin
            Arbiter_Y_7__state <= 2'b10;
          end else begin
            Arbiter_Y_7__state <= 2'b11;
          end
        end 
      end 
      if(Arbiter_Y_7__state == 2'b11) begin
        if(Arbiter_Y_7__ap_done) begin
          Arbiter_Y_7__state <= 2'b10;
        end 
      end 
      if(Arbiter_Y_7__state == 2'b10) begin
        if(Arbiter_Y_7__ap_done_global__q0) begin
          Arbiter_Y_7__state <= 2'b00;
        end 
      end 
    end
  end
  assign Arbiter_Y_7__ap_start = (Arbiter_Y_7__state == 2'b01);
  assign FloatvAddFloatv_0__ap_start_global__q0 = ap_start__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      FloatvAddFloatv_0__ap_start <= 1'b0;
    end else if(FloatvAddFloatv_0__ap_start_global__q0) begin
      FloatvAddFloatv_0__ap_start <= 1'b1;
    end 
  end
  assign FloatvMultConst_0__ap_start_global__q0 = ap_start__q0;
  assign FloatvMultConst_0__is_done__q0 = (FloatvMultConst_0__state == 2'b10);
  assign FloatvMultConst_0__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      FloatvMultConst_0__state <= 2'b00;
    end else begin
      if(FloatvMultConst_0__state == 2'b00) begin
        if(FloatvMultConst_0__ap_start_global__q0) begin
          FloatvMultConst_0__state <= 2'b01;
        end 
      end 
      if(FloatvMultConst_0__state == 2'b01) begin
        if(FloatvMultConst_0__ap_ready) begin
          if(FloatvMultConst_0__ap_done) begin
            FloatvMultConst_0__state <= 2'b10;
          end else begin
            FloatvMultConst_0__state <= 2'b11;
          end
        end 
      end 
      if(FloatvMultConst_0__state == 2'b11) begin
        if(FloatvMultConst_0__ap_done) begin
          FloatvMultConst_0__state <= 2'b10;
        end 
      end 
      if(FloatvMultConst_0__state == 2'b10) begin
        if(FloatvMultConst_0__ap_done_global__q0) begin
          FloatvMultConst_0__state <= 2'b00;
        end 
      end 
    end
  end
  assign FloatvMultConst_0__ap_start = (FloatvMultConst_0__state == 2'b01);
  assign FloatvMultConst_1__ap_start_global__q0 = ap_start__q0;
  assign FloatvMultConst_1__is_done__q0 = (FloatvMultConst_1__state == 2'b10);
  assign FloatvMultConst_1__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      FloatvMultConst_1__state <= 2'b00;
    end else begin
      if(FloatvMultConst_1__state == 2'b00) begin
        if(FloatvMultConst_1__ap_start_global__q0) begin
          FloatvMultConst_1__state <= 2'b01;
        end 
      end 
      if(FloatvMultConst_1__state == 2'b01) begin
        if(FloatvMultConst_1__ap_ready) begin
          if(FloatvMultConst_1__ap_done) begin
            FloatvMultConst_1__state <= 2'b10;
          end else begin
            FloatvMultConst_1__state <= 2'b11;
          end
        end 
      end 
      if(FloatvMultConst_1__state == 2'b11) begin
        if(FloatvMultConst_1__ap_done) begin
          FloatvMultConst_1__state <= 2'b10;
        end 
      end 
      if(FloatvMultConst_1__state == 2'b10) begin
        if(FloatvMultConst_1__ap_done_global__q0) begin
          FloatvMultConst_1__state <= 2'b00;
        end 
      end 
    end
  end
  assign FloatvMultConst_1__ap_start = (FloatvMultConst_1__state == 2'b01);
  assign Merger_Y_0__ap_start_global__q0 = ap_start__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Merger_Y_0__ap_start <= 1'b0;
    end else if(Merger_Y_0__ap_start_global__q0) begin
      Merger_Y_0__ap_start <= 1'b1;
    end 
  end
  assign PEG_Xvec_0__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_0__is_done__q0 = (PEG_Xvec_0__state == 2'b10);
  assign PEG_Xvec_0__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_0__state <= 2'b00;
    end else begin
      if(PEG_Xvec_0__state == 2'b00) begin
        if(PEG_Xvec_0__ap_start_global__q0) begin
          PEG_Xvec_0__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_0__state == 2'b01) begin
        if(PEG_Xvec_0__ap_ready) begin
          if(PEG_Xvec_0__ap_done) begin
            PEG_Xvec_0__state <= 2'b10;
          end else begin
            PEG_Xvec_0__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_0__state == 2'b11) begin
        if(PEG_Xvec_0__ap_done) begin
          PEG_Xvec_0__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_0__state == 2'b10) begin
        if(PEG_Xvec_0__ap_done_global__q0) begin
          PEG_Xvec_0__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_0__ap_start = (PEG_Xvec_0__state == 2'b01);
  assign PEG_Xvec_1__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_1__is_done__q0 = (PEG_Xvec_1__state == 2'b10);
  assign PEG_Xvec_1__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_1__state <= 2'b00;
    end else begin
      if(PEG_Xvec_1__state == 2'b00) begin
        if(PEG_Xvec_1__ap_start_global__q0) begin
          PEG_Xvec_1__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_1__state == 2'b01) begin
        if(PEG_Xvec_1__ap_ready) begin
          if(PEG_Xvec_1__ap_done) begin
            PEG_Xvec_1__state <= 2'b10;
          end else begin
            PEG_Xvec_1__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_1__state == 2'b11) begin
        if(PEG_Xvec_1__ap_done) begin
          PEG_Xvec_1__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_1__state == 2'b10) begin
        if(PEG_Xvec_1__ap_done_global__q0) begin
          PEG_Xvec_1__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_1__ap_start = (PEG_Xvec_1__state == 2'b01);
  assign PEG_Xvec_2__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_2__is_done__q0 = (PEG_Xvec_2__state == 2'b10);
  assign PEG_Xvec_2__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_2__state <= 2'b00;
    end else begin
      if(PEG_Xvec_2__state == 2'b00) begin
        if(PEG_Xvec_2__ap_start_global__q0) begin
          PEG_Xvec_2__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_2__state == 2'b01) begin
        if(PEG_Xvec_2__ap_ready) begin
          if(PEG_Xvec_2__ap_done) begin
            PEG_Xvec_2__state <= 2'b10;
          end else begin
            PEG_Xvec_2__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_2__state == 2'b11) begin
        if(PEG_Xvec_2__ap_done) begin
          PEG_Xvec_2__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_2__state == 2'b10) begin
        if(PEG_Xvec_2__ap_done_global__q0) begin
          PEG_Xvec_2__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_2__ap_start = (PEG_Xvec_2__state == 2'b01);
  assign PEG_Xvec_3__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_3__is_done__q0 = (PEG_Xvec_3__state == 2'b10);
  assign PEG_Xvec_3__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_3__state <= 2'b00;
    end else begin
      if(PEG_Xvec_3__state == 2'b00) begin
        if(PEG_Xvec_3__ap_start_global__q0) begin
          PEG_Xvec_3__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_3__state == 2'b01) begin
        if(PEG_Xvec_3__ap_ready) begin
          if(PEG_Xvec_3__ap_done) begin
            PEG_Xvec_3__state <= 2'b10;
          end else begin
            PEG_Xvec_3__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_3__state == 2'b11) begin
        if(PEG_Xvec_3__ap_done) begin
          PEG_Xvec_3__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_3__state == 2'b10) begin
        if(PEG_Xvec_3__ap_done_global__q0) begin
          PEG_Xvec_3__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_3__ap_start = (PEG_Xvec_3__state == 2'b01);
  assign PEG_Xvec_4__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_4__is_done__q0 = (PEG_Xvec_4__state == 2'b10);
  assign PEG_Xvec_4__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_4__state <= 2'b00;
    end else begin
      if(PEG_Xvec_4__state == 2'b00) begin
        if(PEG_Xvec_4__ap_start_global__q0) begin
          PEG_Xvec_4__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_4__state == 2'b01) begin
        if(PEG_Xvec_4__ap_ready) begin
          if(PEG_Xvec_4__ap_done) begin
            PEG_Xvec_4__state <= 2'b10;
          end else begin
            PEG_Xvec_4__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_4__state == 2'b11) begin
        if(PEG_Xvec_4__ap_done) begin
          PEG_Xvec_4__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_4__state == 2'b10) begin
        if(PEG_Xvec_4__ap_done_global__q0) begin
          PEG_Xvec_4__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_4__ap_start = (PEG_Xvec_4__state == 2'b01);
  assign PEG_Xvec_5__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_5__is_done__q0 = (PEG_Xvec_5__state == 2'b10);
  assign PEG_Xvec_5__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_5__state <= 2'b00;
    end else begin
      if(PEG_Xvec_5__state == 2'b00) begin
        if(PEG_Xvec_5__ap_start_global__q0) begin
          PEG_Xvec_5__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_5__state == 2'b01) begin
        if(PEG_Xvec_5__ap_ready) begin
          if(PEG_Xvec_5__ap_done) begin
            PEG_Xvec_5__state <= 2'b10;
          end else begin
            PEG_Xvec_5__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_5__state == 2'b11) begin
        if(PEG_Xvec_5__ap_done) begin
          PEG_Xvec_5__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_5__state == 2'b10) begin
        if(PEG_Xvec_5__ap_done_global__q0) begin
          PEG_Xvec_5__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_5__ap_start = (PEG_Xvec_5__state == 2'b01);
  assign PEG_Xvec_6__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_6__is_done__q0 = (PEG_Xvec_6__state == 2'b10);
  assign PEG_Xvec_6__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_6__state <= 2'b00;
    end else begin
      if(PEG_Xvec_6__state == 2'b00) begin
        if(PEG_Xvec_6__ap_start_global__q0) begin
          PEG_Xvec_6__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_6__state == 2'b01) begin
        if(PEG_Xvec_6__ap_ready) begin
          if(PEG_Xvec_6__ap_done) begin
            PEG_Xvec_6__state <= 2'b10;
          end else begin
            PEG_Xvec_6__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_6__state == 2'b11) begin
        if(PEG_Xvec_6__ap_done) begin
          PEG_Xvec_6__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_6__state == 2'b10) begin
        if(PEG_Xvec_6__ap_done_global__q0) begin
          PEG_Xvec_6__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_6__ap_start = (PEG_Xvec_6__state == 2'b01);
  assign PEG_Xvec_7__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_7__is_done__q0 = (PEG_Xvec_7__state == 2'b10);
  assign PEG_Xvec_7__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_7__state <= 2'b00;
    end else begin
      if(PEG_Xvec_7__state == 2'b00) begin
        if(PEG_Xvec_7__ap_start_global__q0) begin
          PEG_Xvec_7__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_7__state == 2'b01) begin
        if(PEG_Xvec_7__ap_ready) begin
          if(PEG_Xvec_7__ap_done) begin
            PEG_Xvec_7__state <= 2'b10;
          end else begin
            PEG_Xvec_7__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_7__state == 2'b11) begin
        if(PEG_Xvec_7__ap_done) begin
          PEG_Xvec_7__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_7__state == 2'b10) begin
        if(PEG_Xvec_7__ap_done_global__q0) begin
          PEG_Xvec_7__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_7__ap_start = (PEG_Xvec_7__state == 2'b01);
  assign PEG_Xvec_8__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_8__is_done__q0 = (PEG_Xvec_8__state == 2'b10);
  assign PEG_Xvec_8__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_8__state <= 2'b00;
    end else begin
      if(PEG_Xvec_8__state == 2'b00) begin
        if(PEG_Xvec_8__ap_start_global__q0) begin
          PEG_Xvec_8__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_8__state == 2'b01) begin
        if(PEG_Xvec_8__ap_ready) begin
          if(PEG_Xvec_8__ap_done) begin
            PEG_Xvec_8__state <= 2'b10;
          end else begin
            PEG_Xvec_8__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_8__state == 2'b11) begin
        if(PEG_Xvec_8__ap_done) begin
          PEG_Xvec_8__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_8__state == 2'b10) begin
        if(PEG_Xvec_8__ap_done_global__q0) begin
          PEG_Xvec_8__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_8__ap_start = (PEG_Xvec_8__state == 2'b01);
  assign PEG_Xvec_9__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_9__is_done__q0 = (PEG_Xvec_9__state == 2'b10);
  assign PEG_Xvec_9__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_9__state <= 2'b00;
    end else begin
      if(PEG_Xvec_9__state == 2'b00) begin
        if(PEG_Xvec_9__ap_start_global__q0) begin
          PEG_Xvec_9__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_9__state == 2'b01) begin
        if(PEG_Xvec_9__ap_ready) begin
          if(PEG_Xvec_9__ap_done) begin
            PEG_Xvec_9__state <= 2'b10;
          end else begin
            PEG_Xvec_9__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_9__state == 2'b11) begin
        if(PEG_Xvec_9__ap_done) begin
          PEG_Xvec_9__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_9__state == 2'b10) begin
        if(PEG_Xvec_9__ap_done_global__q0) begin
          PEG_Xvec_9__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_9__ap_start = (PEG_Xvec_9__state == 2'b01);
  assign PEG_Xvec_10__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_10__is_done__q0 = (PEG_Xvec_10__state == 2'b10);
  assign PEG_Xvec_10__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_10__state <= 2'b00;
    end else begin
      if(PEG_Xvec_10__state == 2'b00) begin
        if(PEG_Xvec_10__ap_start_global__q0) begin
          PEG_Xvec_10__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_10__state == 2'b01) begin
        if(PEG_Xvec_10__ap_ready) begin
          if(PEG_Xvec_10__ap_done) begin
            PEG_Xvec_10__state <= 2'b10;
          end else begin
            PEG_Xvec_10__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_10__state == 2'b11) begin
        if(PEG_Xvec_10__ap_done) begin
          PEG_Xvec_10__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_10__state == 2'b10) begin
        if(PEG_Xvec_10__ap_done_global__q0) begin
          PEG_Xvec_10__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_10__ap_start = (PEG_Xvec_10__state == 2'b01);
  assign PEG_Xvec_11__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_11__is_done__q0 = (PEG_Xvec_11__state == 2'b10);
  assign PEG_Xvec_11__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_11__state <= 2'b00;
    end else begin
      if(PEG_Xvec_11__state == 2'b00) begin
        if(PEG_Xvec_11__ap_start_global__q0) begin
          PEG_Xvec_11__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_11__state == 2'b01) begin
        if(PEG_Xvec_11__ap_ready) begin
          if(PEG_Xvec_11__ap_done) begin
            PEG_Xvec_11__state <= 2'b10;
          end else begin
            PEG_Xvec_11__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_11__state == 2'b11) begin
        if(PEG_Xvec_11__ap_done) begin
          PEG_Xvec_11__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_11__state == 2'b10) begin
        if(PEG_Xvec_11__ap_done_global__q0) begin
          PEG_Xvec_11__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_11__ap_start = (PEG_Xvec_11__state == 2'b01);
  assign PEG_Xvec_12__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_12__is_done__q0 = (PEG_Xvec_12__state == 2'b10);
  assign PEG_Xvec_12__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_12__state <= 2'b00;
    end else begin
      if(PEG_Xvec_12__state == 2'b00) begin
        if(PEG_Xvec_12__ap_start_global__q0) begin
          PEG_Xvec_12__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_12__state == 2'b01) begin
        if(PEG_Xvec_12__ap_ready) begin
          if(PEG_Xvec_12__ap_done) begin
            PEG_Xvec_12__state <= 2'b10;
          end else begin
            PEG_Xvec_12__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_12__state == 2'b11) begin
        if(PEG_Xvec_12__ap_done) begin
          PEG_Xvec_12__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_12__state == 2'b10) begin
        if(PEG_Xvec_12__ap_done_global__q0) begin
          PEG_Xvec_12__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_12__ap_start = (PEG_Xvec_12__state == 2'b01);
  assign PEG_Xvec_13__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_13__is_done__q0 = (PEG_Xvec_13__state == 2'b10);
  assign PEG_Xvec_13__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_13__state <= 2'b00;
    end else begin
      if(PEG_Xvec_13__state == 2'b00) begin
        if(PEG_Xvec_13__ap_start_global__q0) begin
          PEG_Xvec_13__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_13__state == 2'b01) begin
        if(PEG_Xvec_13__ap_ready) begin
          if(PEG_Xvec_13__ap_done) begin
            PEG_Xvec_13__state <= 2'b10;
          end else begin
            PEG_Xvec_13__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_13__state == 2'b11) begin
        if(PEG_Xvec_13__ap_done) begin
          PEG_Xvec_13__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_13__state == 2'b10) begin
        if(PEG_Xvec_13__ap_done_global__q0) begin
          PEG_Xvec_13__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_13__ap_start = (PEG_Xvec_13__state == 2'b01);
  assign PEG_Xvec_14__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_14__is_done__q0 = (PEG_Xvec_14__state == 2'b10);
  assign PEG_Xvec_14__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_14__state <= 2'b00;
    end else begin
      if(PEG_Xvec_14__state == 2'b00) begin
        if(PEG_Xvec_14__ap_start_global__q0) begin
          PEG_Xvec_14__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_14__state == 2'b01) begin
        if(PEG_Xvec_14__ap_ready) begin
          if(PEG_Xvec_14__ap_done) begin
            PEG_Xvec_14__state <= 2'b10;
          end else begin
            PEG_Xvec_14__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_14__state == 2'b11) begin
        if(PEG_Xvec_14__ap_done) begin
          PEG_Xvec_14__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_14__state == 2'b10) begin
        if(PEG_Xvec_14__ap_done_global__q0) begin
          PEG_Xvec_14__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_14__ap_start = (PEG_Xvec_14__state == 2'b01);
  assign PEG_Xvec_15__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_15__is_done__q0 = (PEG_Xvec_15__state == 2'b10);
  assign PEG_Xvec_15__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_15__state <= 2'b00;
    end else begin
      if(PEG_Xvec_15__state == 2'b00) begin
        if(PEG_Xvec_15__ap_start_global__q0) begin
          PEG_Xvec_15__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_15__state == 2'b01) begin
        if(PEG_Xvec_15__ap_ready) begin
          if(PEG_Xvec_15__ap_done) begin
            PEG_Xvec_15__state <= 2'b10;
          end else begin
            PEG_Xvec_15__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_15__state == 2'b11) begin
        if(PEG_Xvec_15__ap_done) begin
          PEG_Xvec_15__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_15__state == 2'b10) begin
        if(PEG_Xvec_15__ap_done_global__q0) begin
          PEG_Xvec_15__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_15__ap_start = (PEG_Xvec_15__state == 2'b01);
  assign PEG_Xvec_16__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_16__is_done__q0 = (PEG_Xvec_16__state == 2'b10);
  assign PEG_Xvec_16__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_16__state <= 2'b00;
    end else begin
      if(PEG_Xvec_16__state == 2'b00) begin
        if(PEG_Xvec_16__ap_start_global__q0) begin
          PEG_Xvec_16__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_16__state == 2'b01) begin
        if(PEG_Xvec_16__ap_ready) begin
          if(PEG_Xvec_16__ap_done) begin
            PEG_Xvec_16__state <= 2'b10;
          end else begin
            PEG_Xvec_16__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_16__state == 2'b11) begin
        if(PEG_Xvec_16__ap_done) begin
          PEG_Xvec_16__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_16__state == 2'b10) begin
        if(PEG_Xvec_16__ap_done_global__q0) begin
          PEG_Xvec_16__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_16__ap_start = (PEG_Xvec_16__state == 2'b01);
  assign PEG_Xvec_17__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_17__is_done__q0 = (PEG_Xvec_17__state == 2'b10);
  assign PEG_Xvec_17__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_17__state <= 2'b00;
    end else begin
      if(PEG_Xvec_17__state == 2'b00) begin
        if(PEG_Xvec_17__ap_start_global__q0) begin
          PEG_Xvec_17__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_17__state == 2'b01) begin
        if(PEG_Xvec_17__ap_ready) begin
          if(PEG_Xvec_17__ap_done) begin
            PEG_Xvec_17__state <= 2'b10;
          end else begin
            PEG_Xvec_17__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_17__state == 2'b11) begin
        if(PEG_Xvec_17__ap_done) begin
          PEG_Xvec_17__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_17__state == 2'b10) begin
        if(PEG_Xvec_17__ap_done_global__q0) begin
          PEG_Xvec_17__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_17__ap_start = (PEG_Xvec_17__state == 2'b01);
  assign PEG_Xvec_18__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_18__is_done__q0 = (PEG_Xvec_18__state == 2'b10);
  assign PEG_Xvec_18__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_18__state <= 2'b00;
    end else begin
      if(PEG_Xvec_18__state == 2'b00) begin
        if(PEG_Xvec_18__ap_start_global__q0) begin
          PEG_Xvec_18__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_18__state == 2'b01) begin
        if(PEG_Xvec_18__ap_ready) begin
          if(PEG_Xvec_18__ap_done) begin
            PEG_Xvec_18__state <= 2'b10;
          end else begin
            PEG_Xvec_18__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_18__state == 2'b11) begin
        if(PEG_Xvec_18__ap_done) begin
          PEG_Xvec_18__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_18__state == 2'b10) begin
        if(PEG_Xvec_18__ap_done_global__q0) begin
          PEG_Xvec_18__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_18__ap_start = (PEG_Xvec_18__state == 2'b01);
  assign PEG_Xvec_19__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_19__is_done__q0 = (PEG_Xvec_19__state == 2'b10);
  assign PEG_Xvec_19__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_19__state <= 2'b00;
    end else begin
      if(PEG_Xvec_19__state == 2'b00) begin
        if(PEG_Xvec_19__ap_start_global__q0) begin
          PEG_Xvec_19__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_19__state == 2'b01) begin
        if(PEG_Xvec_19__ap_ready) begin
          if(PEG_Xvec_19__ap_done) begin
            PEG_Xvec_19__state <= 2'b10;
          end else begin
            PEG_Xvec_19__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_19__state == 2'b11) begin
        if(PEG_Xvec_19__ap_done) begin
          PEG_Xvec_19__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_19__state == 2'b10) begin
        if(PEG_Xvec_19__ap_done_global__q0) begin
          PEG_Xvec_19__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_19__ap_start = (PEG_Xvec_19__state == 2'b01);
  assign PEG_Xvec_20__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_20__is_done__q0 = (PEG_Xvec_20__state == 2'b10);
  assign PEG_Xvec_20__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_20__state <= 2'b00;
    end else begin
      if(PEG_Xvec_20__state == 2'b00) begin
        if(PEG_Xvec_20__ap_start_global__q0) begin
          PEG_Xvec_20__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_20__state == 2'b01) begin
        if(PEG_Xvec_20__ap_ready) begin
          if(PEG_Xvec_20__ap_done) begin
            PEG_Xvec_20__state <= 2'b10;
          end else begin
            PEG_Xvec_20__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_20__state == 2'b11) begin
        if(PEG_Xvec_20__ap_done) begin
          PEG_Xvec_20__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_20__state == 2'b10) begin
        if(PEG_Xvec_20__ap_done_global__q0) begin
          PEG_Xvec_20__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_20__ap_start = (PEG_Xvec_20__state == 2'b01);
  assign PEG_Xvec_21__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_21__is_done__q0 = (PEG_Xvec_21__state == 2'b10);
  assign PEG_Xvec_21__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_21__state <= 2'b00;
    end else begin
      if(PEG_Xvec_21__state == 2'b00) begin
        if(PEG_Xvec_21__ap_start_global__q0) begin
          PEG_Xvec_21__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_21__state == 2'b01) begin
        if(PEG_Xvec_21__ap_ready) begin
          if(PEG_Xvec_21__ap_done) begin
            PEG_Xvec_21__state <= 2'b10;
          end else begin
            PEG_Xvec_21__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_21__state == 2'b11) begin
        if(PEG_Xvec_21__ap_done) begin
          PEG_Xvec_21__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_21__state == 2'b10) begin
        if(PEG_Xvec_21__ap_done_global__q0) begin
          PEG_Xvec_21__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_21__ap_start = (PEG_Xvec_21__state == 2'b01);
  assign PEG_Xvec_22__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_22__is_done__q0 = (PEG_Xvec_22__state == 2'b10);
  assign PEG_Xvec_22__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_22__state <= 2'b00;
    end else begin
      if(PEG_Xvec_22__state == 2'b00) begin
        if(PEG_Xvec_22__ap_start_global__q0) begin
          PEG_Xvec_22__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_22__state == 2'b01) begin
        if(PEG_Xvec_22__ap_ready) begin
          if(PEG_Xvec_22__ap_done) begin
            PEG_Xvec_22__state <= 2'b10;
          end else begin
            PEG_Xvec_22__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_22__state == 2'b11) begin
        if(PEG_Xvec_22__ap_done) begin
          PEG_Xvec_22__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_22__state == 2'b10) begin
        if(PEG_Xvec_22__ap_done_global__q0) begin
          PEG_Xvec_22__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_22__ap_start = (PEG_Xvec_22__state == 2'b01);
  assign PEG_Xvec_23__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_23__is_done__q0 = (PEG_Xvec_23__state == 2'b10);
  assign PEG_Xvec_23__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_23__state <= 2'b00;
    end else begin
      if(PEG_Xvec_23__state == 2'b00) begin
        if(PEG_Xvec_23__ap_start_global__q0) begin
          PEG_Xvec_23__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_23__state == 2'b01) begin
        if(PEG_Xvec_23__ap_ready) begin
          if(PEG_Xvec_23__ap_done) begin
            PEG_Xvec_23__state <= 2'b10;
          end else begin
            PEG_Xvec_23__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_23__state == 2'b11) begin
        if(PEG_Xvec_23__ap_done) begin
          PEG_Xvec_23__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_23__state == 2'b10) begin
        if(PEG_Xvec_23__ap_done_global__q0) begin
          PEG_Xvec_23__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_23__ap_start = (PEG_Xvec_23__state == 2'b01);
  assign PEG_Xvec_24__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_24__is_done__q0 = (PEG_Xvec_24__state == 2'b10);
  assign PEG_Xvec_24__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_24__state <= 2'b00;
    end else begin
      if(PEG_Xvec_24__state == 2'b00) begin
        if(PEG_Xvec_24__ap_start_global__q0) begin
          PEG_Xvec_24__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_24__state == 2'b01) begin
        if(PEG_Xvec_24__ap_ready) begin
          if(PEG_Xvec_24__ap_done) begin
            PEG_Xvec_24__state <= 2'b10;
          end else begin
            PEG_Xvec_24__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_24__state == 2'b11) begin
        if(PEG_Xvec_24__ap_done) begin
          PEG_Xvec_24__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_24__state == 2'b10) begin
        if(PEG_Xvec_24__ap_done_global__q0) begin
          PEG_Xvec_24__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_24__ap_start = (PEG_Xvec_24__state == 2'b01);
  assign PEG_Xvec_25__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_25__is_done__q0 = (PEG_Xvec_25__state == 2'b10);
  assign PEG_Xvec_25__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_25__state <= 2'b00;
    end else begin
      if(PEG_Xvec_25__state == 2'b00) begin
        if(PEG_Xvec_25__ap_start_global__q0) begin
          PEG_Xvec_25__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_25__state == 2'b01) begin
        if(PEG_Xvec_25__ap_ready) begin
          if(PEG_Xvec_25__ap_done) begin
            PEG_Xvec_25__state <= 2'b10;
          end else begin
            PEG_Xvec_25__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_25__state == 2'b11) begin
        if(PEG_Xvec_25__ap_done) begin
          PEG_Xvec_25__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_25__state == 2'b10) begin
        if(PEG_Xvec_25__ap_done_global__q0) begin
          PEG_Xvec_25__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_25__ap_start = (PEG_Xvec_25__state == 2'b01);
  assign PEG_Xvec_26__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_26__is_done__q0 = (PEG_Xvec_26__state == 2'b10);
  assign PEG_Xvec_26__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_26__state <= 2'b00;
    end else begin
      if(PEG_Xvec_26__state == 2'b00) begin
        if(PEG_Xvec_26__ap_start_global__q0) begin
          PEG_Xvec_26__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_26__state == 2'b01) begin
        if(PEG_Xvec_26__ap_ready) begin
          if(PEG_Xvec_26__ap_done) begin
            PEG_Xvec_26__state <= 2'b10;
          end else begin
            PEG_Xvec_26__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_26__state == 2'b11) begin
        if(PEG_Xvec_26__ap_done) begin
          PEG_Xvec_26__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_26__state == 2'b10) begin
        if(PEG_Xvec_26__ap_done_global__q0) begin
          PEG_Xvec_26__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_26__ap_start = (PEG_Xvec_26__state == 2'b01);
  assign PEG_Xvec_27__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_27__is_done__q0 = (PEG_Xvec_27__state == 2'b10);
  assign PEG_Xvec_27__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_27__state <= 2'b00;
    end else begin
      if(PEG_Xvec_27__state == 2'b00) begin
        if(PEG_Xvec_27__ap_start_global__q0) begin
          PEG_Xvec_27__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_27__state == 2'b01) begin
        if(PEG_Xvec_27__ap_ready) begin
          if(PEG_Xvec_27__ap_done) begin
            PEG_Xvec_27__state <= 2'b10;
          end else begin
            PEG_Xvec_27__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_27__state == 2'b11) begin
        if(PEG_Xvec_27__ap_done) begin
          PEG_Xvec_27__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_27__state == 2'b10) begin
        if(PEG_Xvec_27__ap_done_global__q0) begin
          PEG_Xvec_27__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_27__ap_start = (PEG_Xvec_27__state == 2'b01);
  assign PEG_Xvec_28__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_28__is_done__q0 = (PEG_Xvec_28__state == 2'b10);
  assign PEG_Xvec_28__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_28__state <= 2'b00;
    end else begin
      if(PEG_Xvec_28__state == 2'b00) begin
        if(PEG_Xvec_28__ap_start_global__q0) begin
          PEG_Xvec_28__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_28__state == 2'b01) begin
        if(PEG_Xvec_28__ap_ready) begin
          if(PEG_Xvec_28__ap_done) begin
            PEG_Xvec_28__state <= 2'b10;
          end else begin
            PEG_Xvec_28__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_28__state == 2'b11) begin
        if(PEG_Xvec_28__ap_done) begin
          PEG_Xvec_28__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_28__state == 2'b10) begin
        if(PEG_Xvec_28__ap_done_global__q0) begin
          PEG_Xvec_28__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_28__ap_start = (PEG_Xvec_28__state == 2'b01);
  assign PEG_Xvec_29__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_29__is_done__q0 = (PEG_Xvec_29__state == 2'b10);
  assign PEG_Xvec_29__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_29__state <= 2'b00;
    end else begin
      if(PEG_Xvec_29__state == 2'b00) begin
        if(PEG_Xvec_29__ap_start_global__q0) begin
          PEG_Xvec_29__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_29__state == 2'b01) begin
        if(PEG_Xvec_29__ap_ready) begin
          if(PEG_Xvec_29__ap_done) begin
            PEG_Xvec_29__state <= 2'b10;
          end else begin
            PEG_Xvec_29__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_29__state == 2'b11) begin
        if(PEG_Xvec_29__ap_done) begin
          PEG_Xvec_29__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_29__state == 2'b10) begin
        if(PEG_Xvec_29__ap_done_global__q0) begin
          PEG_Xvec_29__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_29__ap_start = (PEG_Xvec_29__state == 2'b01);
  assign PEG_Xvec_30__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_30__is_done__q0 = (PEG_Xvec_30__state == 2'b10);
  assign PEG_Xvec_30__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_30__state <= 2'b00;
    end else begin
      if(PEG_Xvec_30__state == 2'b00) begin
        if(PEG_Xvec_30__ap_start_global__q0) begin
          PEG_Xvec_30__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_30__state == 2'b01) begin
        if(PEG_Xvec_30__ap_ready) begin
          if(PEG_Xvec_30__ap_done) begin
            PEG_Xvec_30__state <= 2'b10;
          end else begin
            PEG_Xvec_30__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_30__state == 2'b11) begin
        if(PEG_Xvec_30__ap_done) begin
          PEG_Xvec_30__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_30__state == 2'b10) begin
        if(PEG_Xvec_30__ap_done_global__q0) begin
          PEG_Xvec_30__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_30__ap_start = (PEG_Xvec_30__state == 2'b01);
  assign PEG_Xvec_31__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_31__is_done__q0 = (PEG_Xvec_31__state == 2'b10);
  assign PEG_Xvec_31__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_31__state <= 2'b00;
    end else begin
      if(PEG_Xvec_31__state == 2'b00) begin
        if(PEG_Xvec_31__ap_start_global__q0) begin
          PEG_Xvec_31__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_31__state == 2'b01) begin
        if(PEG_Xvec_31__ap_ready) begin
          if(PEG_Xvec_31__ap_done) begin
            PEG_Xvec_31__state <= 2'b10;
          end else begin
            PEG_Xvec_31__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_31__state == 2'b11) begin
        if(PEG_Xvec_31__ap_done) begin
          PEG_Xvec_31__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_31__state == 2'b10) begin
        if(PEG_Xvec_31__ap_done_global__q0) begin
          PEG_Xvec_31__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_31__ap_start = (PEG_Xvec_31__state == 2'b01);
  assign PEG_Xvec_32__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_32__is_done__q0 = (PEG_Xvec_32__state == 2'b10);
  assign PEG_Xvec_32__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_32__state <= 2'b00;
    end else begin
      if(PEG_Xvec_32__state == 2'b00) begin
        if(PEG_Xvec_32__ap_start_global__q0) begin
          PEG_Xvec_32__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_32__state == 2'b01) begin
        if(PEG_Xvec_32__ap_ready) begin
          if(PEG_Xvec_32__ap_done) begin
            PEG_Xvec_32__state <= 2'b10;
          end else begin
            PEG_Xvec_32__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_32__state == 2'b11) begin
        if(PEG_Xvec_32__ap_done) begin
          PEG_Xvec_32__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_32__state == 2'b10) begin
        if(PEG_Xvec_32__ap_done_global__q0) begin
          PEG_Xvec_32__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_32__ap_start = (PEG_Xvec_32__state == 2'b01);
  assign PEG_Xvec_33__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_33__is_done__q0 = (PEG_Xvec_33__state == 2'b10);
  assign PEG_Xvec_33__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_33__state <= 2'b00;
    end else begin
      if(PEG_Xvec_33__state == 2'b00) begin
        if(PEG_Xvec_33__ap_start_global__q0) begin
          PEG_Xvec_33__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_33__state == 2'b01) begin
        if(PEG_Xvec_33__ap_ready) begin
          if(PEG_Xvec_33__ap_done) begin
            PEG_Xvec_33__state <= 2'b10;
          end else begin
            PEG_Xvec_33__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_33__state == 2'b11) begin
        if(PEG_Xvec_33__ap_done) begin
          PEG_Xvec_33__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_33__state == 2'b10) begin
        if(PEG_Xvec_33__ap_done_global__q0) begin
          PEG_Xvec_33__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_33__ap_start = (PEG_Xvec_33__state == 2'b01);
  assign PEG_Xvec_34__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_34__is_done__q0 = (PEG_Xvec_34__state == 2'b10);
  assign PEG_Xvec_34__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_34__state <= 2'b00;
    end else begin
      if(PEG_Xvec_34__state == 2'b00) begin
        if(PEG_Xvec_34__ap_start_global__q0) begin
          PEG_Xvec_34__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_34__state == 2'b01) begin
        if(PEG_Xvec_34__ap_ready) begin
          if(PEG_Xvec_34__ap_done) begin
            PEG_Xvec_34__state <= 2'b10;
          end else begin
            PEG_Xvec_34__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_34__state == 2'b11) begin
        if(PEG_Xvec_34__ap_done) begin
          PEG_Xvec_34__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_34__state == 2'b10) begin
        if(PEG_Xvec_34__ap_done_global__q0) begin
          PEG_Xvec_34__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_34__ap_start = (PEG_Xvec_34__state == 2'b01);
  assign PEG_Xvec_35__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_35__is_done__q0 = (PEG_Xvec_35__state == 2'b10);
  assign PEG_Xvec_35__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_35__state <= 2'b00;
    end else begin
      if(PEG_Xvec_35__state == 2'b00) begin
        if(PEG_Xvec_35__ap_start_global__q0) begin
          PEG_Xvec_35__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_35__state == 2'b01) begin
        if(PEG_Xvec_35__ap_ready) begin
          if(PEG_Xvec_35__ap_done) begin
            PEG_Xvec_35__state <= 2'b10;
          end else begin
            PEG_Xvec_35__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_35__state == 2'b11) begin
        if(PEG_Xvec_35__ap_done) begin
          PEG_Xvec_35__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_35__state == 2'b10) begin
        if(PEG_Xvec_35__ap_done_global__q0) begin
          PEG_Xvec_35__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_35__ap_start = (PEG_Xvec_35__state == 2'b01);
  assign PEG_Xvec_36__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_36__is_done__q0 = (PEG_Xvec_36__state == 2'b10);
  assign PEG_Xvec_36__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_36__state <= 2'b00;
    end else begin
      if(PEG_Xvec_36__state == 2'b00) begin
        if(PEG_Xvec_36__ap_start_global__q0) begin
          PEG_Xvec_36__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_36__state == 2'b01) begin
        if(PEG_Xvec_36__ap_ready) begin
          if(PEG_Xvec_36__ap_done) begin
            PEG_Xvec_36__state <= 2'b10;
          end else begin
            PEG_Xvec_36__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_36__state == 2'b11) begin
        if(PEG_Xvec_36__ap_done) begin
          PEG_Xvec_36__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_36__state == 2'b10) begin
        if(PEG_Xvec_36__ap_done_global__q0) begin
          PEG_Xvec_36__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_36__ap_start = (PEG_Xvec_36__state == 2'b01);
  assign PEG_Xvec_37__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_37__is_done__q0 = (PEG_Xvec_37__state == 2'b10);
  assign PEG_Xvec_37__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_37__state <= 2'b00;
    end else begin
      if(PEG_Xvec_37__state == 2'b00) begin
        if(PEG_Xvec_37__ap_start_global__q0) begin
          PEG_Xvec_37__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_37__state == 2'b01) begin
        if(PEG_Xvec_37__ap_ready) begin
          if(PEG_Xvec_37__ap_done) begin
            PEG_Xvec_37__state <= 2'b10;
          end else begin
            PEG_Xvec_37__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_37__state == 2'b11) begin
        if(PEG_Xvec_37__ap_done) begin
          PEG_Xvec_37__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_37__state == 2'b10) begin
        if(PEG_Xvec_37__ap_done_global__q0) begin
          PEG_Xvec_37__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_37__ap_start = (PEG_Xvec_37__state == 2'b01);
  assign PEG_Xvec_38__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_38__is_done__q0 = (PEG_Xvec_38__state == 2'b10);
  assign PEG_Xvec_38__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_38__state <= 2'b00;
    end else begin
      if(PEG_Xvec_38__state == 2'b00) begin
        if(PEG_Xvec_38__ap_start_global__q0) begin
          PEG_Xvec_38__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_38__state == 2'b01) begin
        if(PEG_Xvec_38__ap_ready) begin
          if(PEG_Xvec_38__ap_done) begin
            PEG_Xvec_38__state <= 2'b10;
          end else begin
            PEG_Xvec_38__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_38__state == 2'b11) begin
        if(PEG_Xvec_38__ap_done) begin
          PEG_Xvec_38__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_38__state == 2'b10) begin
        if(PEG_Xvec_38__ap_done_global__q0) begin
          PEG_Xvec_38__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_38__ap_start = (PEG_Xvec_38__state == 2'b01);
  assign PEG_Xvec_39__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_39__is_done__q0 = (PEG_Xvec_39__state == 2'b10);
  assign PEG_Xvec_39__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_39__state <= 2'b00;
    end else begin
      if(PEG_Xvec_39__state == 2'b00) begin
        if(PEG_Xvec_39__ap_start_global__q0) begin
          PEG_Xvec_39__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_39__state == 2'b01) begin
        if(PEG_Xvec_39__ap_ready) begin
          if(PEG_Xvec_39__ap_done) begin
            PEG_Xvec_39__state <= 2'b10;
          end else begin
            PEG_Xvec_39__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_39__state == 2'b11) begin
        if(PEG_Xvec_39__ap_done) begin
          PEG_Xvec_39__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_39__state == 2'b10) begin
        if(PEG_Xvec_39__ap_done_global__q0) begin
          PEG_Xvec_39__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_39__ap_start = (PEG_Xvec_39__state == 2'b01);
  assign PEG_Xvec_40__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_40__is_done__q0 = (PEG_Xvec_40__state == 2'b10);
  assign PEG_Xvec_40__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_40__state <= 2'b00;
    end else begin
      if(PEG_Xvec_40__state == 2'b00) begin
        if(PEG_Xvec_40__ap_start_global__q0) begin
          PEG_Xvec_40__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_40__state == 2'b01) begin
        if(PEG_Xvec_40__ap_ready) begin
          if(PEG_Xvec_40__ap_done) begin
            PEG_Xvec_40__state <= 2'b10;
          end else begin
            PEG_Xvec_40__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_40__state == 2'b11) begin
        if(PEG_Xvec_40__ap_done) begin
          PEG_Xvec_40__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_40__state == 2'b10) begin
        if(PEG_Xvec_40__ap_done_global__q0) begin
          PEG_Xvec_40__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_40__ap_start = (PEG_Xvec_40__state == 2'b01);
  assign PEG_Xvec_41__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_41__is_done__q0 = (PEG_Xvec_41__state == 2'b10);
  assign PEG_Xvec_41__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_41__state <= 2'b00;
    end else begin
      if(PEG_Xvec_41__state == 2'b00) begin
        if(PEG_Xvec_41__ap_start_global__q0) begin
          PEG_Xvec_41__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_41__state == 2'b01) begin
        if(PEG_Xvec_41__ap_ready) begin
          if(PEG_Xvec_41__ap_done) begin
            PEG_Xvec_41__state <= 2'b10;
          end else begin
            PEG_Xvec_41__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_41__state == 2'b11) begin
        if(PEG_Xvec_41__ap_done) begin
          PEG_Xvec_41__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_41__state == 2'b10) begin
        if(PEG_Xvec_41__ap_done_global__q0) begin
          PEG_Xvec_41__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_41__ap_start = (PEG_Xvec_41__state == 2'b01);
  assign PEG_Xvec_42__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_42__is_done__q0 = (PEG_Xvec_42__state == 2'b10);
  assign PEG_Xvec_42__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_42__state <= 2'b00;
    end else begin
      if(PEG_Xvec_42__state == 2'b00) begin
        if(PEG_Xvec_42__ap_start_global__q0) begin
          PEG_Xvec_42__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_42__state == 2'b01) begin
        if(PEG_Xvec_42__ap_ready) begin
          if(PEG_Xvec_42__ap_done) begin
            PEG_Xvec_42__state <= 2'b10;
          end else begin
            PEG_Xvec_42__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_42__state == 2'b11) begin
        if(PEG_Xvec_42__ap_done) begin
          PEG_Xvec_42__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_42__state == 2'b10) begin
        if(PEG_Xvec_42__ap_done_global__q0) begin
          PEG_Xvec_42__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_42__ap_start = (PEG_Xvec_42__state == 2'b01);
  assign PEG_Xvec_43__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_43__is_done__q0 = (PEG_Xvec_43__state == 2'b10);
  assign PEG_Xvec_43__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_43__state <= 2'b00;
    end else begin
      if(PEG_Xvec_43__state == 2'b00) begin
        if(PEG_Xvec_43__ap_start_global__q0) begin
          PEG_Xvec_43__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_43__state == 2'b01) begin
        if(PEG_Xvec_43__ap_ready) begin
          if(PEG_Xvec_43__ap_done) begin
            PEG_Xvec_43__state <= 2'b10;
          end else begin
            PEG_Xvec_43__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_43__state == 2'b11) begin
        if(PEG_Xvec_43__ap_done) begin
          PEG_Xvec_43__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_43__state == 2'b10) begin
        if(PEG_Xvec_43__ap_done_global__q0) begin
          PEG_Xvec_43__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_43__ap_start = (PEG_Xvec_43__state == 2'b01);
  assign PEG_Xvec_44__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_44__is_done__q0 = (PEG_Xvec_44__state == 2'b10);
  assign PEG_Xvec_44__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_44__state <= 2'b00;
    end else begin
      if(PEG_Xvec_44__state == 2'b00) begin
        if(PEG_Xvec_44__ap_start_global__q0) begin
          PEG_Xvec_44__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_44__state == 2'b01) begin
        if(PEG_Xvec_44__ap_ready) begin
          if(PEG_Xvec_44__ap_done) begin
            PEG_Xvec_44__state <= 2'b10;
          end else begin
            PEG_Xvec_44__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_44__state == 2'b11) begin
        if(PEG_Xvec_44__ap_done) begin
          PEG_Xvec_44__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_44__state == 2'b10) begin
        if(PEG_Xvec_44__ap_done_global__q0) begin
          PEG_Xvec_44__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_44__ap_start = (PEG_Xvec_44__state == 2'b01);
  assign PEG_Xvec_45__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_45__is_done__q0 = (PEG_Xvec_45__state == 2'b10);
  assign PEG_Xvec_45__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_45__state <= 2'b00;
    end else begin
      if(PEG_Xvec_45__state == 2'b00) begin
        if(PEG_Xvec_45__ap_start_global__q0) begin
          PEG_Xvec_45__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_45__state == 2'b01) begin
        if(PEG_Xvec_45__ap_ready) begin
          if(PEG_Xvec_45__ap_done) begin
            PEG_Xvec_45__state <= 2'b10;
          end else begin
            PEG_Xvec_45__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_45__state == 2'b11) begin
        if(PEG_Xvec_45__ap_done) begin
          PEG_Xvec_45__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_45__state == 2'b10) begin
        if(PEG_Xvec_45__ap_done_global__q0) begin
          PEG_Xvec_45__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_45__ap_start = (PEG_Xvec_45__state == 2'b01);
  assign PEG_Xvec_46__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_46__is_done__q0 = (PEG_Xvec_46__state == 2'b10);
  assign PEG_Xvec_46__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_46__state <= 2'b00;
    end else begin
      if(PEG_Xvec_46__state == 2'b00) begin
        if(PEG_Xvec_46__ap_start_global__q0) begin
          PEG_Xvec_46__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_46__state == 2'b01) begin
        if(PEG_Xvec_46__ap_ready) begin
          if(PEG_Xvec_46__ap_done) begin
            PEG_Xvec_46__state <= 2'b10;
          end else begin
            PEG_Xvec_46__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_46__state == 2'b11) begin
        if(PEG_Xvec_46__ap_done) begin
          PEG_Xvec_46__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_46__state == 2'b10) begin
        if(PEG_Xvec_46__ap_done_global__q0) begin
          PEG_Xvec_46__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_46__ap_start = (PEG_Xvec_46__state == 2'b01);
  assign PEG_Xvec_47__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_47__is_done__q0 = (PEG_Xvec_47__state == 2'b10);
  assign PEG_Xvec_47__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_47__state <= 2'b00;
    end else begin
      if(PEG_Xvec_47__state == 2'b00) begin
        if(PEG_Xvec_47__ap_start_global__q0) begin
          PEG_Xvec_47__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_47__state == 2'b01) begin
        if(PEG_Xvec_47__ap_ready) begin
          if(PEG_Xvec_47__ap_done) begin
            PEG_Xvec_47__state <= 2'b10;
          end else begin
            PEG_Xvec_47__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_47__state == 2'b11) begin
        if(PEG_Xvec_47__ap_done) begin
          PEG_Xvec_47__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_47__state == 2'b10) begin
        if(PEG_Xvec_47__ap_done_global__q0) begin
          PEG_Xvec_47__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_47__ap_start = (PEG_Xvec_47__state == 2'b01);
  assign PEG_Xvec_48__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_48__is_done__q0 = (PEG_Xvec_48__state == 2'b10);
  assign PEG_Xvec_48__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_48__state <= 2'b00;
    end else begin
      if(PEG_Xvec_48__state == 2'b00) begin
        if(PEG_Xvec_48__ap_start_global__q0) begin
          PEG_Xvec_48__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_48__state == 2'b01) begin
        if(PEG_Xvec_48__ap_ready) begin
          if(PEG_Xvec_48__ap_done) begin
            PEG_Xvec_48__state <= 2'b10;
          end else begin
            PEG_Xvec_48__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_48__state == 2'b11) begin
        if(PEG_Xvec_48__ap_done) begin
          PEG_Xvec_48__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_48__state == 2'b10) begin
        if(PEG_Xvec_48__ap_done_global__q0) begin
          PEG_Xvec_48__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_48__ap_start = (PEG_Xvec_48__state == 2'b01);
  assign PEG_Xvec_49__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_49__is_done__q0 = (PEG_Xvec_49__state == 2'b10);
  assign PEG_Xvec_49__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_49__state <= 2'b00;
    end else begin
      if(PEG_Xvec_49__state == 2'b00) begin
        if(PEG_Xvec_49__ap_start_global__q0) begin
          PEG_Xvec_49__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_49__state == 2'b01) begin
        if(PEG_Xvec_49__ap_ready) begin
          if(PEG_Xvec_49__ap_done) begin
            PEG_Xvec_49__state <= 2'b10;
          end else begin
            PEG_Xvec_49__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_49__state == 2'b11) begin
        if(PEG_Xvec_49__ap_done) begin
          PEG_Xvec_49__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_49__state == 2'b10) begin
        if(PEG_Xvec_49__ap_done_global__q0) begin
          PEG_Xvec_49__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_49__ap_start = (PEG_Xvec_49__state == 2'b01);
  assign PEG_Xvec_50__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_50__is_done__q0 = (PEG_Xvec_50__state == 2'b10);
  assign PEG_Xvec_50__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_50__state <= 2'b00;
    end else begin
      if(PEG_Xvec_50__state == 2'b00) begin
        if(PEG_Xvec_50__ap_start_global__q0) begin
          PEG_Xvec_50__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_50__state == 2'b01) begin
        if(PEG_Xvec_50__ap_ready) begin
          if(PEG_Xvec_50__ap_done) begin
            PEG_Xvec_50__state <= 2'b10;
          end else begin
            PEG_Xvec_50__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_50__state == 2'b11) begin
        if(PEG_Xvec_50__ap_done) begin
          PEG_Xvec_50__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_50__state == 2'b10) begin
        if(PEG_Xvec_50__ap_done_global__q0) begin
          PEG_Xvec_50__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_50__ap_start = (PEG_Xvec_50__state == 2'b01);
  assign PEG_Xvec_51__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_51__is_done__q0 = (PEG_Xvec_51__state == 2'b10);
  assign PEG_Xvec_51__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_51__state <= 2'b00;
    end else begin
      if(PEG_Xvec_51__state == 2'b00) begin
        if(PEG_Xvec_51__ap_start_global__q0) begin
          PEG_Xvec_51__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_51__state == 2'b01) begin
        if(PEG_Xvec_51__ap_ready) begin
          if(PEG_Xvec_51__ap_done) begin
            PEG_Xvec_51__state <= 2'b10;
          end else begin
            PEG_Xvec_51__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_51__state == 2'b11) begin
        if(PEG_Xvec_51__ap_done) begin
          PEG_Xvec_51__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_51__state == 2'b10) begin
        if(PEG_Xvec_51__ap_done_global__q0) begin
          PEG_Xvec_51__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_51__ap_start = (PEG_Xvec_51__state == 2'b01);
  assign PEG_Xvec_52__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_52__is_done__q0 = (PEG_Xvec_52__state == 2'b10);
  assign PEG_Xvec_52__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_52__state <= 2'b00;
    end else begin
      if(PEG_Xvec_52__state == 2'b00) begin
        if(PEG_Xvec_52__ap_start_global__q0) begin
          PEG_Xvec_52__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_52__state == 2'b01) begin
        if(PEG_Xvec_52__ap_ready) begin
          if(PEG_Xvec_52__ap_done) begin
            PEG_Xvec_52__state <= 2'b10;
          end else begin
            PEG_Xvec_52__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_52__state == 2'b11) begin
        if(PEG_Xvec_52__ap_done) begin
          PEG_Xvec_52__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_52__state == 2'b10) begin
        if(PEG_Xvec_52__ap_done_global__q0) begin
          PEG_Xvec_52__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_52__ap_start = (PEG_Xvec_52__state == 2'b01);
  assign PEG_Xvec_53__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_53__is_done__q0 = (PEG_Xvec_53__state == 2'b10);
  assign PEG_Xvec_53__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_53__state <= 2'b00;
    end else begin
      if(PEG_Xvec_53__state == 2'b00) begin
        if(PEG_Xvec_53__ap_start_global__q0) begin
          PEG_Xvec_53__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_53__state == 2'b01) begin
        if(PEG_Xvec_53__ap_ready) begin
          if(PEG_Xvec_53__ap_done) begin
            PEG_Xvec_53__state <= 2'b10;
          end else begin
            PEG_Xvec_53__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_53__state == 2'b11) begin
        if(PEG_Xvec_53__ap_done) begin
          PEG_Xvec_53__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_53__state == 2'b10) begin
        if(PEG_Xvec_53__ap_done_global__q0) begin
          PEG_Xvec_53__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_53__ap_start = (PEG_Xvec_53__state == 2'b01);
  assign PEG_Xvec_54__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_54__is_done__q0 = (PEG_Xvec_54__state == 2'b10);
  assign PEG_Xvec_54__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_54__state <= 2'b00;
    end else begin
      if(PEG_Xvec_54__state == 2'b00) begin
        if(PEG_Xvec_54__ap_start_global__q0) begin
          PEG_Xvec_54__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_54__state == 2'b01) begin
        if(PEG_Xvec_54__ap_ready) begin
          if(PEG_Xvec_54__ap_done) begin
            PEG_Xvec_54__state <= 2'b10;
          end else begin
            PEG_Xvec_54__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_54__state == 2'b11) begin
        if(PEG_Xvec_54__ap_done) begin
          PEG_Xvec_54__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_54__state == 2'b10) begin
        if(PEG_Xvec_54__ap_done_global__q0) begin
          PEG_Xvec_54__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_54__ap_start = (PEG_Xvec_54__state == 2'b01);
  assign PEG_Xvec_55__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_55__is_done__q0 = (PEG_Xvec_55__state == 2'b10);
  assign PEG_Xvec_55__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_55__state <= 2'b00;
    end else begin
      if(PEG_Xvec_55__state == 2'b00) begin
        if(PEG_Xvec_55__ap_start_global__q0) begin
          PEG_Xvec_55__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_55__state == 2'b01) begin
        if(PEG_Xvec_55__ap_ready) begin
          if(PEG_Xvec_55__ap_done) begin
            PEG_Xvec_55__state <= 2'b10;
          end else begin
            PEG_Xvec_55__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_55__state == 2'b11) begin
        if(PEG_Xvec_55__ap_done) begin
          PEG_Xvec_55__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_55__state == 2'b10) begin
        if(PEG_Xvec_55__ap_done_global__q0) begin
          PEG_Xvec_55__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Xvec_55__ap_start = (PEG_Xvec_55__state == 2'b01);
  assign PEG_Yvec_0__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_0__is_done__q0 = (PEG_Yvec_0__state == 2'b10);
  assign PEG_Yvec_0__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_0__state <= 2'b00;
    end else begin
      if(PEG_Yvec_0__state == 2'b00) begin
        if(PEG_Yvec_0__ap_start_global__q0) begin
          PEG_Yvec_0__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_0__state == 2'b01) begin
        if(PEG_Yvec_0__ap_ready) begin
          if(PEG_Yvec_0__ap_done) begin
            PEG_Yvec_0__state <= 2'b10;
          end else begin
            PEG_Yvec_0__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_0__state == 2'b11) begin
        if(PEG_Yvec_0__ap_done) begin
          PEG_Yvec_0__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_0__state == 2'b10) begin
        if(PEG_Yvec_0__ap_done_global__q0) begin
          PEG_Yvec_0__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_0__ap_start = (PEG_Yvec_0__state == 2'b01);
  assign PEG_Yvec_1__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_1__is_done__q0 = (PEG_Yvec_1__state == 2'b10);
  assign PEG_Yvec_1__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_1__state <= 2'b00;
    end else begin
      if(PEG_Yvec_1__state == 2'b00) begin
        if(PEG_Yvec_1__ap_start_global__q0) begin
          PEG_Yvec_1__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_1__state == 2'b01) begin
        if(PEG_Yvec_1__ap_ready) begin
          if(PEG_Yvec_1__ap_done) begin
            PEG_Yvec_1__state <= 2'b10;
          end else begin
            PEG_Yvec_1__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_1__state == 2'b11) begin
        if(PEG_Yvec_1__ap_done) begin
          PEG_Yvec_1__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_1__state == 2'b10) begin
        if(PEG_Yvec_1__ap_done_global__q0) begin
          PEG_Yvec_1__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_1__ap_start = (PEG_Yvec_1__state == 2'b01);
  assign PEG_Yvec_2__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_2__is_done__q0 = (PEG_Yvec_2__state == 2'b10);
  assign PEG_Yvec_2__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_2__state <= 2'b00;
    end else begin
      if(PEG_Yvec_2__state == 2'b00) begin
        if(PEG_Yvec_2__ap_start_global__q0) begin
          PEG_Yvec_2__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_2__state == 2'b01) begin
        if(PEG_Yvec_2__ap_ready) begin
          if(PEG_Yvec_2__ap_done) begin
            PEG_Yvec_2__state <= 2'b10;
          end else begin
            PEG_Yvec_2__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_2__state == 2'b11) begin
        if(PEG_Yvec_2__ap_done) begin
          PEG_Yvec_2__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_2__state == 2'b10) begin
        if(PEG_Yvec_2__ap_done_global__q0) begin
          PEG_Yvec_2__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_2__ap_start = (PEG_Yvec_2__state == 2'b01);
  assign PEG_Yvec_3__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_3__is_done__q0 = (PEG_Yvec_3__state == 2'b10);
  assign PEG_Yvec_3__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_3__state <= 2'b00;
    end else begin
      if(PEG_Yvec_3__state == 2'b00) begin
        if(PEG_Yvec_3__ap_start_global__q0) begin
          PEG_Yvec_3__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_3__state == 2'b01) begin
        if(PEG_Yvec_3__ap_ready) begin
          if(PEG_Yvec_3__ap_done) begin
            PEG_Yvec_3__state <= 2'b10;
          end else begin
            PEG_Yvec_3__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_3__state == 2'b11) begin
        if(PEG_Yvec_3__ap_done) begin
          PEG_Yvec_3__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_3__state == 2'b10) begin
        if(PEG_Yvec_3__ap_done_global__q0) begin
          PEG_Yvec_3__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_3__ap_start = (PEG_Yvec_3__state == 2'b01);
  assign PEG_Yvec_4__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_4__is_done__q0 = (PEG_Yvec_4__state == 2'b10);
  assign PEG_Yvec_4__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_4__state <= 2'b00;
    end else begin
      if(PEG_Yvec_4__state == 2'b00) begin
        if(PEG_Yvec_4__ap_start_global__q0) begin
          PEG_Yvec_4__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_4__state == 2'b01) begin
        if(PEG_Yvec_4__ap_ready) begin
          if(PEG_Yvec_4__ap_done) begin
            PEG_Yvec_4__state <= 2'b10;
          end else begin
            PEG_Yvec_4__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_4__state == 2'b11) begin
        if(PEG_Yvec_4__ap_done) begin
          PEG_Yvec_4__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_4__state == 2'b10) begin
        if(PEG_Yvec_4__ap_done_global__q0) begin
          PEG_Yvec_4__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_4__ap_start = (PEG_Yvec_4__state == 2'b01);
  assign PEG_Yvec_5__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_5__is_done__q0 = (PEG_Yvec_5__state == 2'b10);
  assign PEG_Yvec_5__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_5__state <= 2'b00;
    end else begin
      if(PEG_Yvec_5__state == 2'b00) begin
        if(PEG_Yvec_5__ap_start_global__q0) begin
          PEG_Yvec_5__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_5__state == 2'b01) begin
        if(PEG_Yvec_5__ap_ready) begin
          if(PEG_Yvec_5__ap_done) begin
            PEG_Yvec_5__state <= 2'b10;
          end else begin
            PEG_Yvec_5__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_5__state == 2'b11) begin
        if(PEG_Yvec_5__ap_done) begin
          PEG_Yvec_5__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_5__state == 2'b10) begin
        if(PEG_Yvec_5__ap_done_global__q0) begin
          PEG_Yvec_5__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_5__ap_start = (PEG_Yvec_5__state == 2'b01);
  assign PEG_Yvec_6__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_6__is_done__q0 = (PEG_Yvec_6__state == 2'b10);
  assign PEG_Yvec_6__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_6__state <= 2'b00;
    end else begin
      if(PEG_Yvec_6__state == 2'b00) begin
        if(PEG_Yvec_6__ap_start_global__q0) begin
          PEG_Yvec_6__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_6__state == 2'b01) begin
        if(PEG_Yvec_6__ap_ready) begin
          if(PEG_Yvec_6__ap_done) begin
            PEG_Yvec_6__state <= 2'b10;
          end else begin
            PEG_Yvec_6__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_6__state == 2'b11) begin
        if(PEG_Yvec_6__ap_done) begin
          PEG_Yvec_6__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_6__state == 2'b10) begin
        if(PEG_Yvec_6__ap_done_global__q0) begin
          PEG_Yvec_6__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_6__ap_start = (PEG_Yvec_6__state == 2'b01);
  assign PEG_Yvec_7__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_7__is_done__q0 = (PEG_Yvec_7__state == 2'b10);
  assign PEG_Yvec_7__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_7__state <= 2'b00;
    end else begin
      if(PEG_Yvec_7__state == 2'b00) begin
        if(PEG_Yvec_7__ap_start_global__q0) begin
          PEG_Yvec_7__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_7__state == 2'b01) begin
        if(PEG_Yvec_7__ap_ready) begin
          if(PEG_Yvec_7__ap_done) begin
            PEG_Yvec_7__state <= 2'b10;
          end else begin
            PEG_Yvec_7__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_7__state == 2'b11) begin
        if(PEG_Yvec_7__ap_done) begin
          PEG_Yvec_7__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_7__state == 2'b10) begin
        if(PEG_Yvec_7__ap_done_global__q0) begin
          PEG_Yvec_7__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_7__ap_start = (PEG_Yvec_7__state == 2'b01);
  assign PEG_Yvec_8__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_8__is_done__q0 = (PEG_Yvec_8__state == 2'b10);
  assign PEG_Yvec_8__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_8__state <= 2'b00;
    end else begin
      if(PEG_Yvec_8__state == 2'b00) begin
        if(PEG_Yvec_8__ap_start_global__q0) begin
          PEG_Yvec_8__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_8__state == 2'b01) begin
        if(PEG_Yvec_8__ap_ready) begin
          if(PEG_Yvec_8__ap_done) begin
            PEG_Yvec_8__state <= 2'b10;
          end else begin
            PEG_Yvec_8__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_8__state == 2'b11) begin
        if(PEG_Yvec_8__ap_done) begin
          PEG_Yvec_8__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_8__state == 2'b10) begin
        if(PEG_Yvec_8__ap_done_global__q0) begin
          PEG_Yvec_8__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_8__ap_start = (PEG_Yvec_8__state == 2'b01);
  assign PEG_Yvec_9__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_9__is_done__q0 = (PEG_Yvec_9__state == 2'b10);
  assign PEG_Yvec_9__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_9__state <= 2'b00;
    end else begin
      if(PEG_Yvec_9__state == 2'b00) begin
        if(PEG_Yvec_9__ap_start_global__q0) begin
          PEG_Yvec_9__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_9__state == 2'b01) begin
        if(PEG_Yvec_9__ap_ready) begin
          if(PEG_Yvec_9__ap_done) begin
            PEG_Yvec_9__state <= 2'b10;
          end else begin
            PEG_Yvec_9__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_9__state == 2'b11) begin
        if(PEG_Yvec_9__ap_done) begin
          PEG_Yvec_9__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_9__state == 2'b10) begin
        if(PEG_Yvec_9__ap_done_global__q0) begin
          PEG_Yvec_9__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_9__ap_start = (PEG_Yvec_9__state == 2'b01);
  assign PEG_Yvec_10__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_10__is_done__q0 = (PEG_Yvec_10__state == 2'b10);
  assign PEG_Yvec_10__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_10__state <= 2'b00;
    end else begin
      if(PEG_Yvec_10__state == 2'b00) begin
        if(PEG_Yvec_10__ap_start_global__q0) begin
          PEG_Yvec_10__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_10__state == 2'b01) begin
        if(PEG_Yvec_10__ap_ready) begin
          if(PEG_Yvec_10__ap_done) begin
            PEG_Yvec_10__state <= 2'b10;
          end else begin
            PEG_Yvec_10__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_10__state == 2'b11) begin
        if(PEG_Yvec_10__ap_done) begin
          PEG_Yvec_10__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_10__state == 2'b10) begin
        if(PEG_Yvec_10__ap_done_global__q0) begin
          PEG_Yvec_10__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_10__ap_start = (PEG_Yvec_10__state == 2'b01);
  assign PEG_Yvec_11__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_11__is_done__q0 = (PEG_Yvec_11__state == 2'b10);
  assign PEG_Yvec_11__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_11__state <= 2'b00;
    end else begin
      if(PEG_Yvec_11__state == 2'b00) begin
        if(PEG_Yvec_11__ap_start_global__q0) begin
          PEG_Yvec_11__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_11__state == 2'b01) begin
        if(PEG_Yvec_11__ap_ready) begin
          if(PEG_Yvec_11__ap_done) begin
            PEG_Yvec_11__state <= 2'b10;
          end else begin
            PEG_Yvec_11__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_11__state == 2'b11) begin
        if(PEG_Yvec_11__ap_done) begin
          PEG_Yvec_11__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_11__state == 2'b10) begin
        if(PEG_Yvec_11__ap_done_global__q0) begin
          PEG_Yvec_11__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_11__ap_start = (PEG_Yvec_11__state == 2'b01);
  assign PEG_Yvec_12__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_12__is_done__q0 = (PEG_Yvec_12__state == 2'b10);
  assign PEG_Yvec_12__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_12__state <= 2'b00;
    end else begin
      if(PEG_Yvec_12__state == 2'b00) begin
        if(PEG_Yvec_12__ap_start_global__q0) begin
          PEG_Yvec_12__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_12__state == 2'b01) begin
        if(PEG_Yvec_12__ap_ready) begin
          if(PEG_Yvec_12__ap_done) begin
            PEG_Yvec_12__state <= 2'b10;
          end else begin
            PEG_Yvec_12__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_12__state == 2'b11) begin
        if(PEG_Yvec_12__ap_done) begin
          PEG_Yvec_12__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_12__state == 2'b10) begin
        if(PEG_Yvec_12__ap_done_global__q0) begin
          PEG_Yvec_12__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_12__ap_start = (PEG_Yvec_12__state == 2'b01);
  assign PEG_Yvec_13__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_13__is_done__q0 = (PEG_Yvec_13__state == 2'b10);
  assign PEG_Yvec_13__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_13__state <= 2'b00;
    end else begin
      if(PEG_Yvec_13__state == 2'b00) begin
        if(PEG_Yvec_13__ap_start_global__q0) begin
          PEG_Yvec_13__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_13__state == 2'b01) begin
        if(PEG_Yvec_13__ap_ready) begin
          if(PEG_Yvec_13__ap_done) begin
            PEG_Yvec_13__state <= 2'b10;
          end else begin
            PEG_Yvec_13__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_13__state == 2'b11) begin
        if(PEG_Yvec_13__ap_done) begin
          PEG_Yvec_13__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_13__state == 2'b10) begin
        if(PEG_Yvec_13__ap_done_global__q0) begin
          PEG_Yvec_13__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_13__ap_start = (PEG_Yvec_13__state == 2'b01);
  assign PEG_Yvec_14__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_14__is_done__q0 = (PEG_Yvec_14__state == 2'b10);
  assign PEG_Yvec_14__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_14__state <= 2'b00;
    end else begin
      if(PEG_Yvec_14__state == 2'b00) begin
        if(PEG_Yvec_14__ap_start_global__q0) begin
          PEG_Yvec_14__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_14__state == 2'b01) begin
        if(PEG_Yvec_14__ap_ready) begin
          if(PEG_Yvec_14__ap_done) begin
            PEG_Yvec_14__state <= 2'b10;
          end else begin
            PEG_Yvec_14__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_14__state == 2'b11) begin
        if(PEG_Yvec_14__ap_done) begin
          PEG_Yvec_14__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_14__state == 2'b10) begin
        if(PEG_Yvec_14__ap_done_global__q0) begin
          PEG_Yvec_14__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_14__ap_start = (PEG_Yvec_14__state == 2'b01);
  assign PEG_Yvec_15__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_15__is_done__q0 = (PEG_Yvec_15__state == 2'b10);
  assign PEG_Yvec_15__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_15__state <= 2'b00;
    end else begin
      if(PEG_Yvec_15__state == 2'b00) begin
        if(PEG_Yvec_15__ap_start_global__q0) begin
          PEG_Yvec_15__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_15__state == 2'b01) begin
        if(PEG_Yvec_15__ap_ready) begin
          if(PEG_Yvec_15__ap_done) begin
            PEG_Yvec_15__state <= 2'b10;
          end else begin
            PEG_Yvec_15__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_15__state == 2'b11) begin
        if(PEG_Yvec_15__ap_done) begin
          PEG_Yvec_15__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_15__state == 2'b10) begin
        if(PEG_Yvec_15__ap_done_global__q0) begin
          PEG_Yvec_15__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_15__ap_start = (PEG_Yvec_15__state == 2'b01);
  assign PEG_Yvec_16__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_16__is_done__q0 = (PEG_Yvec_16__state == 2'b10);
  assign PEG_Yvec_16__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_16__state <= 2'b00;
    end else begin
      if(PEG_Yvec_16__state == 2'b00) begin
        if(PEG_Yvec_16__ap_start_global__q0) begin
          PEG_Yvec_16__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_16__state == 2'b01) begin
        if(PEG_Yvec_16__ap_ready) begin
          if(PEG_Yvec_16__ap_done) begin
            PEG_Yvec_16__state <= 2'b10;
          end else begin
            PEG_Yvec_16__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_16__state == 2'b11) begin
        if(PEG_Yvec_16__ap_done) begin
          PEG_Yvec_16__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_16__state == 2'b10) begin
        if(PEG_Yvec_16__ap_done_global__q0) begin
          PEG_Yvec_16__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_16__ap_start = (PEG_Yvec_16__state == 2'b01);
  assign PEG_Yvec_17__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_17__is_done__q0 = (PEG_Yvec_17__state == 2'b10);
  assign PEG_Yvec_17__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_17__state <= 2'b00;
    end else begin
      if(PEG_Yvec_17__state == 2'b00) begin
        if(PEG_Yvec_17__ap_start_global__q0) begin
          PEG_Yvec_17__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_17__state == 2'b01) begin
        if(PEG_Yvec_17__ap_ready) begin
          if(PEG_Yvec_17__ap_done) begin
            PEG_Yvec_17__state <= 2'b10;
          end else begin
            PEG_Yvec_17__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_17__state == 2'b11) begin
        if(PEG_Yvec_17__ap_done) begin
          PEG_Yvec_17__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_17__state == 2'b10) begin
        if(PEG_Yvec_17__ap_done_global__q0) begin
          PEG_Yvec_17__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_17__ap_start = (PEG_Yvec_17__state == 2'b01);
  assign PEG_Yvec_18__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_18__is_done__q0 = (PEG_Yvec_18__state == 2'b10);
  assign PEG_Yvec_18__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_18__state <= 2'b00;
    end else begin
      if(PEG_Yvec_18__state == 2'b00) begin
        if(PEG_Yvec_18__ap_start_global__q0) begin
          PEG_Yvec_18__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_18__state == 2'b01) begin
        if(PEG_Yvec_18__ap_ready) begin
          if(PEG_Yvec_18__ap_done) begin
            PEG_Yvec_18__state <= 2'b10;
          end else begin
            PEG_Yvec_18__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_18__state == 2'b11) begin
        if(PEG_Yvec_18__ap_done) begin
          PEG_Yvec_18__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_18__state == 2'b10) begin
        if(PEG_Yvec_18__ap_done_global__q0) begin
          PEG_Yvec_18__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_18__ap_start = (PEG_Yvec_18__state == 2'b01);
  assign PEG_Yvec_19__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_19__is_done__q0 = (PEG_Yvec_19__state == 2'b10);
  assign PEG_Yvec_19__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_19__state <= 2'b00;
    end else begin
      if(PEG_Yvec_19__state == 2'b00) begin
        if(PEG_Yvec_19__ap_start_global__q0) begin
          PEG_Yvec_19__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_19__state == 2'b01) begin
        if(PEG_Yvec_19__ap_ready) begin
          if(PEG_Yvec_19__ap_done) begin
            PEG_Yvec_19__state <= 2'b10;
          end else begin
            PEG_Yvec_19__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_19__state == 2'b11) begin
        if(PEG_Yvec_19__ap_done) begin
          PEG_Yvec_19__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_19__state == 2'b10) begin
        if(PEG_Yvec_19__ap_done_global__q0) begin
          PEG_Yvec_19__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_19__ap_start = (PEG_Yvec_19__state == 2'b01);
  assign PEG_Yvec_20__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_20__is_done__q0 = (PEG_Yvec_20__state == 2'b10);
  assign PEG_Yvec_20__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_20__state <= 2'b00;
    end else begin
      if(PEG_Yvec_20__state == 2'b00) begin
        if(PEG_Yvec_20__ap_start_global__q0) begin
          PEG_Yvec_20__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_20__state == 2'b01) begin
        if(PEG_Yvec_20__ap_ready) begin
          if(PEG_Yvec_20__ap_done) begin
            PEG_Yvec_20__state <= 2'b10;
          end else begin
            PEG_Yvec_20__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_20__state == 2'b11) begin
        if(PEG_Yvec_20__ap_done) begin
          PEG_Yvec_20__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_20__state == 2'b10) begin
        if(PEG_Yvec_20__ap_done_global__q0) begin
          PEG_Yvec_20__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_20__ap_start = (PEG_Yvec_20__state == 2'b01);
  assign PEG_Yvec_21__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_21__is_done__q0 = (PEG_Yvec_21__state == 2'b10);
  assign PEG_Yvec_21__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_21__state <= 2'b00;
    end else begin
      if(PEG_Yvec_21__state == 2'b00) begin
        if(PEG_Yvec_21__ap_start_global__q0) begin
          PEG_Yvec_21__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_21__state == 2'b01) begin
        if(PEG_Yvec_21__ap_ready) begin
          if(PEG_Yvec_21__ap_done) begin
            PEG_Yvec_21__state <= 2'b10;
          end else begin
            PEG_Yvec_21__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_21__state == 2'b11) begin
        if(PEG_Yvec_21__ap_done) begin
          PEG_Yvec_21__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_21__state == 2'b10) begin
        if(PEG_Yvec_21__ap_done_global__q0) begin
          PEG_Yvec_21__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_21__ap_start = (PEG_Yvec_21__state == 2'b01);
  assign PEG_Yvec_22__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_22__is_done__q0 = (PEG_Yvec_22__state == 2'b10);
  assign PEG_Yvec_22__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_22__state <= 2'b00;
    end else begin
      if(PEG_Yvec_22__state == 2'b00) begin
        if(PEG_Yvec_22__ap_start_global__q0) begin
          PEG_Yvec_22__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_22__state == 2'b01) begin
        if(PEG_Yvec_22__ap_ready) begin
          if(PEG_Yvec_22__ap_done) begin
            PEG_Yvec_22__state <= 2'b10;
          end else begin
            PEG_Yvec_22__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_22__state == 2'b11) begin
        if(PEG_Yvec_22__ap_done) begin
          PEG_Yvec_22__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_22__state == 2'b10) begin
        if(PEG_Yvec_22__ap_done_global__q0) begin
          PEG_Yvec_22__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_22__ap_start = (PEG_Yvec_22__state == 2'b01);
  assign PEG_Yvec_23__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_23__is_done__q0 = (PEG_Yvec_23__state == 2'b10);
  assign PEG_Yvec_23__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_23__state <= 2'b00;
    end else begin
      if(PEG_Yvec_23__state == 2'b00) begin
        if(PEG_Yvec_23__ap_start_global__q0) begin
          PEG_Yvec_23__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_23__state == 2'b01) begin
        if(PEG_Yvec_23__ap_ready) begin
          if(PEG_Yvec_23__ap_done) begin
            PEG_Yvec_23__state <= 2'b10;
          end else begin
            PEG_Yvec_23__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_23__state == 2'b11) begin
        if(PEG_Yvec_23__ap_done) begin
          PEG_Yvec_23__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_23__state == 2'b10) begin
        if(PEG_Yvec_23__ap_done_global__q0) begin
          PEG_Yvec_23__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_23__ap_start = (PEG_Yvec_23__state == 2'b01);
  assign PEG_Yvec_24__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_24__is_done__q0 = (PEG_Yvec_24__state == 2'b10);
  assign PEG_Yvec_24__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_24__state <= 2'b00;
    end else begin
      if(PEG_Yvec_24__state == 2'b00) begin
        if(PEG_Yvec_24__ap_start_global__q0) begin
          PEG_Yvec_24__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_24__state == 2'b01) begin
        if(PEG_Yvec_24__ap_ready) begin
          if(PEG_Yvec_24__ap_done) begin
            PEG_Yvec_24__state <= 2'b10;
          end else begin
            PEG_Yvec_24__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_24__state == 2'b11) begin
        if(PEG_Yvec_24__ap_done) begin
          PEG_Yvec_24__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_24__state == 2'b10) begin
        if(PEG_Yvec_24__ap_done_global__q0) begin
          PEG_Yvec_24__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_24__ap_start = (PEG_Yvec_24__state == 2'b01);
  assign PEG_Yvec_25__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_25__is_done__q0 = (PEG_Yvec_25__state == 2'b10);
  assign PEG_Yvec_25__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_25__state <= 2'b00;
    end else begin
      if(PEG_Yvec_25__state == 2'b00) begin
        if(PEG_Yvec_25__ap_start_global__q0) begin
          PEG_Yvec_25__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_25__state == 2'b01) begin
        if(PEG_Yvec_25__ap_ready) begin
          if(PEG_Yvec_25__ap_done) begin
            PEG_Yvec_25__state <= 2'b10;
          end else begin
            PEG_Yvec_25__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_25__state == 2'b11) begin
        if(PEG_Yvec_25__ap_done) begin
          PEG_Yvec_25__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_25__state == 2'b10) begin
        if(PEG_Yvec_25__ap_done_global__q0) begin
          PEG_Yvec_25__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_25__ap_start = (PEG_Yvec_25__state == 2'b01);
  assign PEG_Yvec_26__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_26__is_done__q0 = (PEG_Yvec_26__state == 2'b10);
  assign PEG_Yvec_26__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_26__state <= 2'b00;
    end else begin
      if(PEG_Yvec_26__state == 2'b00) begin
        if(PEG_Yvec_26__ap_start_global__q0) begin
          PEG_Yvec_26__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_26__state == 2'b01) begin
        if(PEG_Yvec_26__ap_ready) begin
          if(PEG_Yvec_26__ap_done) begin
            PEG_Yvec_26__state <= 2'b10;
          end else begin
            PEG_Yvec_26__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_26__state == 2'b11) begin
        if(PEG_Yvec_26__ap_done) begin
          PEG_Yvec_26__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_26__state == 2'b10) begin
        if(PEG_Yvec_26__ap_done_global__q0) begin
          PEG_Yvec_26__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_26__ap_start = (PEG_Yvec_26__state == 2'b01);
  assign PEG_Yvec_27__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_27__is_done__q0 = (PEG_Yvec_27__state == 2'b10);
  assign PEG_Yvec_27__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_27__state <= 2'b00;
    end else begin
      if(PEG_Yvec_27__state == 2'b00) begin
        if(PEG_Yvec_27__ap_start_global__q0) begin
          PEG_Yvec_27__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_27__state == 2'b01) begin
        if(PEG_Yvec_27__ap_ready) begin
          if(PEG_Yvec_27__ap_done) begin
            PEG_Yvec_27__state <= 2'b10;
          end else begin
            PEG_Yvec_27__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_27__state == 2'b11) begin
        if(PEG_Yvec_27__ap_done) begin
          PEG_Yvec_27__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_27__state == 2'b10) begin
        if(PEG_Yvec_27__ap_done_global__q0) begin
          PEG_Yvec_27__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_27__ap_start = (PEG_Yvec_27__state == 2'b01);
  assign PEG_Yvec_28__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_28__is_done__q0 = (PEG_Yvec_28__state == 2'b10);
  assign PEG_Yvec_28__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_28__state <= 2'b00;
    end else begin
      if(PEG_Yvec_28__state == 2'b00) begin
        if(PEG_Yvec_28__ap_start_global__q0) begin
          PEG_Yvec_28__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_28__state == 2'b01) begin
        if(PEG_Yvec_28__ap_ready) begin
          if(PEG_Yvec_28__ap_done) begin
            PEG_Yvec_28__state <= 2'b10;
          end else begin
            PEG_Yvec_28__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_28__state == 2'b11) begin
        if(PEG_Yvec_28__ap_done) begin
          PEG_Yvec_28__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_28__state == 2'b10) begin
        if(PEG_Yvec_28__ap_done_global__q0) begin
          PEG_Yvec_28__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_28__ap_start = (PEG_Yvec_28__state == 2'b01);
  assign PEG_Yvec_29__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_29__is_done__q0 = (PEG_Yvec_29__state == 2'b10);
  assign PEG_Yvec_29__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_29__state <= 2'b00;
    end else begin
      if(PEG_Yvec_29__state == 2'b00) begin
        if(PEG_Yvec_29__ap_start_global__q0) begin
          PEG_Yvec_29__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_29__state == 2'b01) begin
        if(PEG_Yvec_29__ap_ready) begin
          if(PEG_Yvec_29__ap_done) begin
            PEG_Yvec_29__state <= 2'b10;
          end else begin
            PEG_Yvec_29__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_29__state == 2'b11) begin
        if(PEG_Yvec_29__ap_done) begin
          PEG_Yvec_29__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_29__state == 2'b10) begin
        if(PEG_Yvec_29__ap_done_global__q0) begin
          PEG_Yvec_29__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_29__ap_start = (PEG_Yvec_29__state == 2'b01);
  assign PEG_Yvec_30__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_30__is_done__q0 = (PEG_Yvec_30__state == 2'b10);
  assign PEG_Yvec_30__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_30__state <= 2'b00;
    end else begin
      if(PEG_Yvec_30__state == 2'b00) begin
        if(PEG_Yvec_30__ap_start_global__q0) begin
          PEG_Yvec_30__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_30__state == 2'b01) begin
        if(PEG_Yvec_30__ap_ready) begin
          if(PEG_Yvec_30__ap_done) begin
            PEG_Yvec_30__state <= 2'b10;
          end else begin
            PEG_Yvec_30__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_30__state == 2'b11) begin
        if(PEG_Yvec_30__ap_done) begin
          PEG_Yvec_30__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_30__state == 2'b10) begin
        if(PEG_Yvec_30__ap_done_global__q0) begin
          PEG_Yvec_30__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_30__ap_start = (PEG_Yvec_30__state == 2'b01);
  assign PEG_Yvec_31__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_31__is_done__q0 = (PEG_Yvec_31__state == 2'b10);
  assign PEG_Yvec_31__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_31__state <= 2'b00;
    end else begin
      if(PEG_Yvec_31__state == 2'b00) begin
        if(PEG_Yvec_31__ap_start_global__q0) begin
          PEG_Yvec_31__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_31__state == 2'b01) begin
        if(PEG_Yvec_31__ap_ready) begin
          if(PEG_Yvec_31__ap_done) begin
            PEG_Yvec_31__state <= 2'b10;
          end else begin
            PEG_Yvec_31__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_31__state == 2'b11) begin
        if(PEG_Yvec_31__ap_done) begin
          PEG_Yvec_31__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_31__state == 2'b10) begin
        if(PEG_Yvec_31__ap_done_global__q0) begin
          PEG_Yvec_31__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_31__ap_start = (PEG_Yvec_31__state == 2'b01);
  assign PEG_Yvec_32__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_32__is_done__q0 = (PEG_Yvec_32__state == 2'b10);
  assign PEG_Yvec_32__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_32__state <= 2'b00;
    end else begin
      if(PEG_Yvec_32__state == 2'b00) begin
        if(PEG_Yvec_32__ap_start_global__q0) begin
          PEG_Yvec_32__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_32__state == 2'b01) begin
        if(PEG_Yvec_32__ap_ready) begin
          if(PEG_Yvec_32__ap_done) begin
            PEG_Yvec_32__state <= 2'b10;
          end else begin
            PEG_Yvec_32__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_32__state == 2'b11) begin
        if(PEG_Yvec_32__ap_done) begin
          PEG_Yvec_32__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_32__state == 2'b10) begin
        if(PEG_Yvec_32__ap_done_global__q0) begin
          PEG_Yvec_32__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_32__ap_start = (PEG_Yvec_32__state == 2'b01);
  assign PEG_Yvec_33__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_33__is_done__q0 = (PEG_Yvec_33__state == 2'b10);
  assign PEG_Yvec_33__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_33__state <= 2'b00;
    end else begin
      if(PEG_Yvec_33__state == 2'b00) begin
        if(PEG_Yvec_33__ap_start_global__q0) begin
          PEG_Yvec_33__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_33__state == 2'b01) begin
        if(PEG_Yvec_33__ap_ready) begin
          if(PEG_Yvec_33__ap_done) begin
            PEG_Yvec_33__state <= 2'b10;
          end else begin
            PEG_Yvec_33__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_33__state == 2'b11) begin
        if(PEG_Yvec_33__ap_done) begin
          PEG_Yvec_33__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_33__state == 2'b10) begin
        if(PEG_Yvec_33__ap_done_global__q0) begin
          PEG_Yvec_33__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_33__ap_start = (PEG_Yvec_33__state == 2'b01);
  assign PEG_Yvec_34__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_34__is_done__q0 = (PEG_Yvec_34__state == 2'b10);
  assign PEG_Yvec_34__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_34__state <= 2'b00;
    end else begin
      if(PEG_Yvec_34__state == 2'b00) begin
        if(PEG_Yvec_34__ap_start_global__q0) begin
          PEG_Yvec_34__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_34__state == 2'b01) begin
        if(PEG_Yvec_34__ap_ready) begin
          if(PEG_Yvec_34__ap_done) begin
            PEG_Yvec_34__state <= 2'b10;
          end else begin
            PEG_Yvec_34__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_34__state == 2'b11) begin
        if(PEG_Yvec_34__ap_done) begin
          PEG_Yvec_34__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_34__state == 2'b10) begin
        if(PEG_Yvec_34__ap_done_global__q0) begin
          PEG_Yvec_34__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_34__ap_start = (PEG_Yvec_34__state == 2'b01);
  assign PEG_Yvec_35__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_35__is_done__q0 = (PEG_Yvec_35__state == 2'b10);
  assign PEG_Yvec_35__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_35__state <= 2'b00;
    end else begin
      if(PEG_Yvec_35__state == 2'b00) begin
        if(PEG_Yvec_35__ap_start_global__q0) begin
          PEG_Yvec_35__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_35__state == 2'b01) begin
        if(PEG_Yvec_35__ap_ready) begin
          if(PEG_Yvec_35__ap_done) begin
            PEG_Yvec_35__state <= 2'b10;
          end else begin
            PEG_Yvec_35__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_35__state == 2'b11) begin
        if(PEG_Yvec_35__ap_done) begin
          PEG_Yvec_35__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_35__state == 2'b10) begin
        if(PEG_Yvec_35__ap_done_global__q0) begin
          PEG_Yvec_35__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_35__ap_start = (PEG_Yvec_35__state == 2'b01);
  assign PEG_Yvec_36__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_36__is_done__q0 = (PEG_Yvec_36__state == 2'b10);
  assign PEG_Yvec_36__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_36__state <= 2'b00;
    end else begin
      if(PEG_Yvec_36__state == 2'b00) begin
        if(PEG_Yvec_36__ap_start_global__q0) begin
          PEG_Yvec_36__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_36__state == 2'b01) begin
        if(PEG_Yvec_36__ap_ready) begin
          if(PEG_Yvec_36__ap_done) begin
            PEG_Yvec_36__state <= 2'b10;
          end else begin
            PEG_Yvec_36__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_36__state == 2'b11) begin
        if(PEG_Yvec_36__ap_done) begin
          PEG_Yvec_36__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_36__state == 2'b10) begin
        if(PEG_Yvec_36__ap_done_global__q0) begin
          PEG_Yvec_36__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_36__ap_start = (PEG_Yvec_36__state == 2'b01);
  assign PEG_Yvec_37__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_37__is_done__q0 = (PEG_Yvec_37__state == 2'b10);
  assign PEG_Yvec_37__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_37__state <= 2'b00;
    end else begin
      if(PEG_Yvec_37__state == 2'b00) begin
        if(PEG_Yvec_37__ap_start_global__q0) begin
          PEG_Yvec_37__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_37__state == 2'b01) begin
        if(PEG_Yvec_37__ap_ready) begin
          if(PEG_Yvec_37__ap_done) begin
            PEG_Yvec_37__state <= 2'b10;
          end else begin
            PEG_Yvec_37__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_37__state == 2'b11) begin
        if(PEG_Yvec_37__ap_done) begin
          PEG_Yvec_37__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_37__state == 2'b10) begin
        if(PEG_Yvec_37__ap_done_global__q0) begin
          PEG_Yvec_37__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_37__ap_start = (PEG_Yvec_37__state == 2'b01);
  assign PEG_Yvec_38__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_38__is_done__q0 = (PEG_Yvec_38__state == 2'b10);
  assign PEG_Yvec_38__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_38__state <= 2'b00;
    end else begin
      if(PEG_Yvec_38__state == 2'b00) begin
        if(PEG_Yvec_38__ap_start_global__q0) begin
          PEG_Yvec_38__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_38__state == 2'b01) begin
        if(PEG_Yvec_38__ap_ready) begin
          if(PEG_Yvec_38__ap_done) begin
            PEG_Yvec_38__state <= 2'b10;
          end else begin
            PEG_Yvec_38__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_38__state == 2'b11) begin
        if(PEG_Yvec_38__ap_done) begin
          PEG_Yvec_38__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_38__state == 2'b10) begin
        if(PEG_Yvec_38__ap_done_global__q0) begin
          PEG_Yvec_38__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_38__ap_start = (PEG_Yvec_38__state == 2'b01);
  assign PEG_Yvec_39__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_39__is_done__q0 = (PEG_Yvec_39__state == 2'b10);
  assign PEG_Yvec_39__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_39__state <= 2'b00;
    end else begin
      if(PEG_Yvec_39__state == 2'b00) begin
        if(PEG_Yvec_39__ap_start_global__q0) begin
          PEG_Yvec_39__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_39__state == 2'b01) begin
        if(PEG_Yvec_39__ap_ready) begin
          if(PEG_Yvec_39__ap_done) begin
            PEG_Yvec_39__state <= 2'b10;
          end else begin
            PEG_Yvec_39__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_39__state == 2'b11) begin
        if(PEG_Yvec_39__ap_done) begin
          PEG_Yvec_39__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_39__state == 2'b10) begin
        if(PEG_Yvec_39__ap_done_global__q0) begin
          PEG_Yvec_39__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_39__ap_start = (PEG_Yvec_39__state == 2'b01);
  assign PEG_Yvec_40__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_40__is_done__q0 = (PEG_Yvec_40__state == 2'b10);
  assign PEG_Yvec_40__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_40__state <= 2'b00;
    end else begin
      if(PEG_Yvec_40__state == 2'b00) begin
        if(PEG_Yvec_40__ap_start_global__q0) begin
          PEG_Yvec_40__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_40__state == 2'b01) begin
        if(PEG_Yvec_40__ap_ready) begin
          if(PEG_Yvec_40__ap_done) begin
            PEG_Yvec_40__state <= 2'b10;
          end else begin
            PEG_Yvec_40__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_40__state == 2'b11) begin
        if(PEG_Yvec_40__ap_done) begin
          PEG_Yvec_40__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_40__state == 2'b10) begin
        if(PEG_Yvec_40__ap_done_global__q0) begin
          PEG_Yvec_40__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_40__ap_start = (PEG_Yvec_40__state == 2'b01);
  assign PEG_Yvec_41__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_41__is_done__q0 = (PEG_Yvec_41__state == 2'b10);
  assign PEG_Yvec_41__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_41__state <= 2'b00;
    end else begin
      if(PEG_Yvec_41__state == 2'b00) begin
        if(PEG_Yvec_41__ap_start_global__q0) begin
          PEG_Yvec_41__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_41__state == 2'b01) begin
        if(PEG_Yvec_41__ap_ready) begin
          if(PEG_Yvec_41__ap_done) begin
            PEG_Yvec_41__state <= 2'b10;
          end else begin
            PEG_Yvec_41__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_41__state == 2'b11) begin
        if(PEG_Yvec_41__ap_done) begin
          PEG_Yvec_41__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_41__state == 2'b10) begin
        if(PEG_Yvec_41__ap_done_global__q0) begin
          PEG_Yvec_41__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_41__ap_start = (PEG_Yvec_41__state == 2'b01);
  assign PEG_Yvec_42__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_42__is_done__q0 = (PEG_Yvec_42__state == 2'b10);
  assign PEG_Yvec_42__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_42__state <= 2'b00;
    end else begin
      if(PEG_Yvec_42__state == 2'b00) begin
        if(PEG_Yvec_42__ap_start_global__q0) begin
          PEG_Yvec_42__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_42__state == 2'b01) begin
        if(PEG_Yvec_42__ap_ready) begin
          if(PEG_Yvec_42__ap_done) begin
            PEG_Yvec_42__state <= 2'b10;
          end else begin
            PEG_Yvec_42__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_42__state == 2'b11) begin
        if(PEG_Yvec_42__ap_done) begin
          PEG_Yvec_42__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_42__state == 2'b10) begin
        if(PEG_Yvec_42__ap_done_global__q0) begin
          PEG_Yvec_42__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_42__ap_start = (PEG_Yvec_42__state == 2'b01);
  assign PEG_Yvec_43__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_43__is_done__q0 = (PEG_Yvec_43__state == 2'b10);
  assign PEG_Yvec_43__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_43__state <= 2'b00;
    end else begin
      if(PEG_Yvec_43__state == 2'b00) begin
        if(PEG_Yvec_43__ap_start_global__q0) begin
          PEG_Yvec_43__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_43__state == 2'b01) begin
        if(PEG_Yvec_43__ap_ready) begin
          if(PEG_Yvec_43__ap_done) begin
            PEG_Yvec_43__state <= 2'b10;
          end else begin
            PEG_Yvec_43__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_43__state == 2'b11) begin
        if(PEG_Yvec_43__ap_done) begin
          PEG_Yvec_43__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_43__state == 2'b10) begin
        if(PEG_Yvec_43__ap_done_global__q0) begin
          PEG_Yvec_43__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_43__ap_start = (PEG_Yvec_43__state == 2'b01);
  assign PEG_Yvec_44__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_44__is_done__q0 = (PEG_Yvec_44__state == 2'b10);
  assign PEG_Yvec_44__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_44__state <= 2'b00;
    end else begin
      if(PEG_Yvec_44__state == 2'b00) begin
        if(PEG_Yvec_44__ap_start_global__q0) begin
          PEG_Yvec_44__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_44__state == 2'b01) begin
        if(PEG_Yvec_44__ap_ready) begin
          if(PEG_Yvec_44__ap_done) begin
            PEG_Yvec_44__state <= 2'b10;
          end else begin
            PEG_Yvec_44__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_44__state == 2'b11) begin
        if(PEG_Yvec_44__ap_done) begin
          PEG_Yvec_44__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_44__state == 2'b10) begin
        if(PEG_Yvec_44__ap_done_global__q0) begin
          PEG_Yvec_44__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_44__ap_start = (PEG_Yvec_44__state == 2'b01);
  assign PEG_Yvec_45__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_45__is_done__q0 = (PEG_Yvec_45__state == 2'b10);
  assign PEG_Yvec_45__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_45__state <= 2'b00;
    end else begin
      if(PEG_Yvec_45__state == 2'b00) begin
        if(PEG_Yvec_45__ap_start_global__q0) begin
          PEG_Yvec_45__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_45__state == 2'b01) begin
        if(PEG_Yvec_45__ap_ready) begin
          if(PEG_Yvec_45__ap_done) begin
            PEG_Yvec_45__state <= 2'b10;
          end else begin
            PEG_Yvec_45__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_45__state == 2'b11) begin
        if(PEG_Yvec_45__ap_done) begin
          PEG_Yvec_45__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_45__state == 2'b10) begin
        if(PEG_Yvec_45__ap_done_global__q0) begin
          PEG_Yvec_45__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_45__ap_start = (PEG_Yvec_45__state == 2'b01);
  assign PEG_Yvec_46__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_46__is_done__q0 = (PEG_Yvec_46__state == 2'b10);
  assign PEG_Yvec_46__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_46__state <= 2'b00;
    end else begin
      if(PEG_Yvec_46__state == 2'b00) begin
        if(PEG_Yvec_46__ap_start_global__q0) begin
          PEG_Yvec_46__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_46__state == 2'b01) begin
        if(PEG_Yvec_46__ap_ready) begin
          if(PEG_Yvec_46__ap_done) begin
            PEG_Yvec_46__state <= 2'b10;
          end else begin
            PEG_Yvec_46__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_46__state == 2'b11) begin
        if(PEG_Yvec_46__ap_done) begin
          PEG_Yvec_46__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_46__state == 2'b10) begin
        if(PEG_Yvec_46__ap_done_global__q0) begin
          PEG_Yvec_46__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_46__ap_start = (PEG_Yvec_46__state == 2'b01);
  assign PEG_Yvec_47__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_47__is_done__q0 = (PEG_Yvec_47__state == 2'b10);
  assign PEG_Yvec_47__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_47__state <= 2'b00;
    end else begin
      if(PEG_Yvec_47__state == 2'b00) begin
        if(PEG_Yvec_47__ap_start_global__q0) begin
          PEG_Yvec_47__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_47__state == 2'b01) begin
        if(PEG_Yvec_47__ap_ready) begin
          if(PEG_Yvec_47__ap_done) begin
            PEG_Yvec_47__state <= 2'b10;
          end else begin
            PEG_Yvec_47__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_47__state == 2'b11) begin
        if(PEG_Yvec_47__ap_done) begin
          PEG_Yvec_47__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_47__state == 2'b10) begin
        if(PEG_Yvec_47__ap_done_global__q0) begin
          PEG_Yvec_47__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_47__ap_start = (PEG_Yvec_47__state == 2'b01);
  assign PEG_Yvec_48__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_48__is_done__q0 = (PEG_Yvec_48__state == 2'b10);
  assign PEG_Yvec_48__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_48__state <= 2'b00;
    end else begin
      if(PEG_Yvec_48__state == 2'b00) begin
        if(PEG_Yvec_48__ap_start_global__q0) begin
          PEG_Yvec_48__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_48__state == 2'b01) begin
        if(PEG_Yvec_48__ap_ready) begin
          if(PEG_Yvec_48__ap_done) begin
            PEG_Yvec_48__state <= 2'b10;
          end else begin
            PEG_Yvec_48__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_48__state == 2'b11) begin
        if(PEG_Yvec_48__ap_done) begin
          PEG_Yvec_48__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_48__state == 2'b10) begin
        if(PEG_Yvec_48__ap_done_global__q0) begin
          PEG_Yvec_48__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_48__ap_start = (PEG_Yvec_48__state == 2'b01);
  assign PEG_Yvec_49__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_49__is_done__q0 = (PEG_Yvec_49__state == 2'b10);
  assign PEG_Yvec_49__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_49__state <= 2'b00;
    end else begin
      if(PEG_Yvec_49__state == 2'b00) begin
        if(PEG_Yvec_49__ap_start_global__q0) begin
          PEG_Yvec_49__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_49__state == 2'b01) begin
        if(PEG_Yvec_49__ap_ready) begin
          if(PEG_Yvec_49__ap_done) begin
            PEG_Yvec_49__state <= 2'b10;
          end else begin
            PEG_Yvec_49__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_49__state == 2'b11) begin
        if(PEG_Yvec_49__ap_done) begin
          PEG_Yvec_49__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_49__state == 2'b10) begin
        if(PEG_Yvec_49__ap_done_global__q0) begin
          PEG_Yvec_49__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_49__ap_start = (PEG_Yvec_49__state == 2'b01);
  assign PEG_Yvec_50__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_50__is_done__q0 = (PEG_Yvec_50__state == 2'b10);
  assign PEG_Yvec_50__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_50__state <= 2'b00;
    end else begin
      if(PEG_Yvec_50__state == 2'b00) begin
        if(PEG_Yvec_50__ap_start_global__q0) begin
          PEG_Yvec_50__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_50__state == 2'b01) begin
        if(PEG_Yvec_50__ap_ready) begin
          if(PEG_Yvec_50__ap_done) begin
            PEG_Yvec_50__state <= 2'b10;
          end else begin
            PEG_Yvec_50__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_50__state == 2'b11) begin
        if(PEG_Yvec_50__ap_done) begin
          PEG_Yvec_50__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_50__state == 2'b10) begin
        if(PEG_Yvec_50__ap_done_global__q0) begin
          PEG_Yvec_50__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_50__ap_start = (PEG_Yvec_50__state == 2'b01);
  assign PEG_Yvec_51__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_51__is_done__q0 = (PEG_Yvec_51__state == 2'b10);
  assign PEG_Yvec_51__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_51__state <= 2'b00;
    end else begin
      if(PEG_Yvec_51__state == 2'b00) begin
        if(PEG_Yvec_51__ap_start_global__q0) begin
          PEG_Yvec_51__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_51__state == 2'b01) begin
        if(PEG_Yvec_51__ap_ready) begin
          if(PEG_Yvec_51__ap_done) begin
            PEG_Yvec_51__state <= 2'b10;
          end else begin
            PEG_Yvec_51__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_51__state == 2'b11) begin
        if(PEG_Yvec_51__ap_done) begin
          PEG_Yvec_51__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_51__state == 2'b10) begin
        if(PEG_Yvec_51__ap_done_global__q0) begin
          PEG_Yvec_51__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_51__ap_start = (PEG_Yvec_51__state == 2'b01);
  assign PEG_Yvec_52__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_52__is_done__q0 = (PEG_Yvec_52__state == 2'b10);
  assign PEG_Yvec_52__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_52__state <= 2'b00;
    end else begin
      if(PEG_Yvec_52__state == 2'b00) begin
        if(PEG_Yvec_52__ap_start_global__q0) begin
          PEG_Yvec_52__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_52__state == 2'b01) begin
        if(PEG_Yvec_52__ap_ready) begin
          if(PEG_Yvec_52__ap_done) begin
            PEG_Yvec_52__state <= 2'b10;
          end else begin
            PEG_Yvec_52__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_52__state == 2'b11) begin
        if(PEG_Yvec_52__ap_done) begin
          PEG_Yvec_52__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_52__state == 2'b10) begin
        if(PEG_Yvec_52__ap_done_global__q0) begin
          PEG_Yvec_52__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_52__ap_start = (PEG_Yvec_52__state == 2'b01);
  assign PEG_Yvec_53__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_53__is_done__q0 = (PEG_Yvec_53__state == 2'b10);
  assign PEG_Yvec_53__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_53__state <= 2'b00;
    end else begin
      if(PEG_Yvec_53__state == 2'b00) begin
        if(PEG_Yvec_53__ap_start_global__q0) begin
          PEG_Yvec_53__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_53__state == 2'b01) begin
        if(PEG_Yvec_53__ap_ready) begin
          if(PEG_Yvec_53__ap_done) begin
            PEG_Yvec_53__state <= 2'b10;
          end else begin
            PEG_Yvec_53__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_53__state == 2'b11) begin
        if(PEG_Yvec_53__ap_done) begin
          PEG_Yvec_53__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_53__state == 2'b10) begin
        if(PEG_Yvec_53__ap_done_global__q0) begin
          PEG_Yvec_53__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_53__ap_start = (PEG_Yvec_53__state == 2'b01);
  assign PEG_Yvec_54__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_54__is_done__q0 = (PEG_Yvec_54__state == 2'b10);
  assign PEG_Yvec_54__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_54__state <= 2'b00;
    end else begin
      if(PEG_Yvec_54__state == 2'b00) begin
        if(PEG_Yvec_54__ap_start_global__q0) begin
          PEG_Yvec_54__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_54__state == 2'b01) begin
        if(PEG_Yvec_54__ap_ready) begin
          if(PEG_Yvec_54__ap_done) begin
            PEG_Yvec_54__state <= 2'b10;
          end else begin
            PEG_Yvec_54__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_54__state == 2'b11) begin
        if(PEG_Yvec_54__ap_done) begin
          PEG_Yvec_54__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_54__state == 2'b10) begin
        if(PEG_Yvec_54__ap_done_global__q0) begin
          PEG_Yvec_54__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_54__ap_start = (PEG_Yvec_54__state == 2'b01);
  assign PEG_Yvec_55__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_55__is_done__q0 = (PEG_Yvec_55__state == 2'b10);
  assign PEG_Yvec_55__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_55__state <= 2'b00;
    end else begin
      if(PEG_Yvec_55__state == 2'b00) begin
        if(PEG_Yvec_55__ap_start_global__q0) begin
          PEG_Yvec_55__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_55__state == 2'b01) begin
        if(PEG_Yvec_55__ap_ready) begin
          if(PEG_Yvec_55__ap_done) begin
            PEG_Yvec_55__state <= 2'b10;
          end else begin
            PEG_Yvec_55__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_55__state == 2'b11) begin
        if(PEG_Yvec_55__ap_done) begin
          PEG_Yvec_55__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_55__state == 2'b10) begin
        if(PEG_Yvec_55__ap_done_global__q0) begin
          PEG_Yvec_55__state <= 2'b00;
        end 
      end 
    end
  end
  assign PEG_Yvec_55__ap_start = (PEG_Yvec_55__state == 2'b01);
  assign black_hole_float_v16_0__ap_start_global__q0 = ap_start__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      black_hole_float_v16_0__ap_start <= 1'b0;
    end else if(black_hole_float_v16_0__ap_start_global__q0) begin
      black_hole_float_v16_0__ap_start <= 1'b1;
    end 
  end
  assign black_hole_int_0__ap_start_global__q0 = ap_start__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      black_hole_int_0__ap_start <= 1'b0;
    end else if(black_hole_int_0__ap_start_global__q0) begin
      black_hole_int_0__ap_start <= 1'b1;
    end 
  end
  assign read_A_0__ap_start_global__q0 = ap_start__q0;
  assign read_A_0__is_done__q0 = (read_A_0__state == 2'b10);
  assign read_A_0__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_0__state <= 2'b00;
    end else begin
      if(read_A_0__state == 2'b00) begin
        if(read_A_0__ap_start_global__q0) begin
          read_A_0__state <= 2'b01;
        end 
      end 
      if(read_A_0__state == 2'b01) begin
        if(read_A_0__ap_ready) begin
          if(read_A_0__ap_done) begin
            read_A_0__state <= 2'b10;
          end else begin
            read_A_0__state <= 2'b11;
          end
        end 
      end 
      if(read_A_0__state == 2'b11) begin
        if(read_A_0__ap_done) begin
          read_A_0__state <= 2'b10;
        end 
      end 
      if(read_A_0__state == 2'b10) begin
        if(read_A_0__ap_done_global__q0) begin
          read_A_0__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_0__ap_start = (read_A_0__state == 2'b01);
  assign read_A_1__ap_start_global__q0 = ap_start__q0;
  assign read_A_1__is_done__q0 = (read_A_1__state == 2'b10);
  assign read_A_1__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_1__state <= 2'b00;
    end else begin
      if(read_A_1__state == 2'b00) begin
        if(read_A_1__ap_start_global__q0) begin
          read_A_1__state <= 2'b01;
        end 
      end 
      if(read_A_1__state == 2'b01) begin
        if(read_A_1__ap_ready) begin
          if(read_A_1__ap_done) begin
            read_A_1__state <= 2'b10;
          end else begin
            read_A_1__state <= 2'b11;
          end
        end 
      end 
      if(read_A_1__state == 2'b11) begin
        if(read_A_1__ap_done) begin
          read_A_1__state <= 2'b10;
        end 
      end 
      if(read_A_1__state == 2'b10) begin
        if(read_A_1__ap_done_global__q0) begin
          read_A_1__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_1__ap_start = (read_A_1__state == 2'b01);
  assign read_A_2__ap_start_global__q0 = ap_start__q0;
  assign read_A_2__is_done__q0 = (read_A_2__state == 2'b10);
  assign read_A_2__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_2__state <= 2'b00;
    end else begin
      if(read_A_2__state == 2'b00) begin
        if(read_A_2__ap_start_global__q0) begin
          read_A_2__state <= 2'b01;
        end 
      end 
      if(read_A_2__state == 2'b01) begin
        if(read_A_2__ap_ready) begin
          if(read_A_2__ap_done) begin
            read_A_2__state <= 2'b10;
          end else begin
            read_A_2__state <= 2'b11;
          end
        end 
      end 
      if(read_A_2__state == 2'b11) begin
        if(read_A_2__ap_done) begin
          read_A_2__state <= 2'b10;
        end 
      end 
      if(read_A_2__state == 2'b10) begin
        if(read_A_2__ap_done_global__q0) begin
          read_A_2__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_2__ap_start = (read_A_2__state == 2'b01);
  assign read_A_3__ap_start_global__q0 = ap_start__q0;
  assign read_A_3__is_done__q0 = (read_A_3__state == 2'b10);
  assign read_A_3__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_3__state <= 2'b00;
    end else begin
      if(read_A_3__state == 2'b00) begin
        if(read_A_3__ap_start_global__q0) begin
          read_A_3__state <= 2'b01;
        end 
      end 
      if(read_A_3__state == 2'b01) begin
        if(read_A_3__ap_ready) begin
          if(read_A_3__ap_done) begin
            read_A_3__state <= 2'b10;
          end else begin
            read_A_3__state <= 2'b11;
          end
        end 
      end 
      if(read_A_3__state == 2'b11) begin
        if(read_A_3__ap_done) begin
          read_A_3__state <= 2'b10;
        end 
      end 
      if(read_A_3__state == 2'b10) begin
        if(read_A_3__ap_done_global__q0) begin
          read_A_3__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_3__ap_start = (read_A_3__state == 2'b01);
  assign read_A_4__ap_start_global__q0 = ap_start__q0;
  assign read_A_4__is_done__q0 = (read_A_4__state == 2'b10);
  assign read_A_4__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_4__state <= 2'b00;
    end else begin
      if(read_A_4__state == 2'b00) begin
        if(read_A_4__ap_start_global__q0) begin
          read_A_4__state <= 2'b01;
        end 
      end 
      if(read_A_4__state == 2'b01) begin
        if(read_A_4__ap_ready) begin
          if(read_A_4__ap_done) begin
            read_A_4__state <= 2'b10;
          end else begin
            read_A_4__state <= 2'b11;
          end
        end 
      end 
      if(read_A_4__state == 2'b11) begin
        if(read_A_4__ap_done) begin
          read_A_4__state <= 2'b10;
        end 
      end 
      if(read_A_4__state == 2'b10) begin
        if(read_A_4__ap_done_global__q0) begin
          read_A_4__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_4__ap_start = (read_A_4__state == 2'b01);
  assign read_A_5__ap_start_global__q0 = ap_start__q0;
  assign read_A_5__is_done__q0 = (read_A_5__state == 2'b10);
  assign read_A_5__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_5__state <= 2'b00;
    end else begin
      if(read_A_5__state == 2'b00) begin
        if(read_A_5__ap_start_global__q0) begin
          read_A_5__state <= 2'b01;
        end 
      end 
      if(read_A_5__state == 2'b01) begin
        if(read_A_5__ap_ready) begin
          if(read_A_5__ap_done) begin
            read_A_5__state <= 2'b10;
          end else begin
            read_A_5__state <= 2'b11;
          end
        end 
      end 
      if(read_A_5__state == 2'b11) begin
        if(read_A_5__ap_done) begin
          read_A_5__state <= 2'b10;
        end 
      end 
      if(read_A_5__state == 2'b10) begin
        if(read_A_5__ap_done_global__q0) begin
          read_A_5__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_5__ap_start = (read_A_5__state == 2'b01);
  assign read_A_6__ap_start_global__q0 = ap_start__q0;
  assign read_A_6__is_done__q0 = (read_A_6__state == 2'b10);
  assign read_A_6__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_6__state <= 2'b00;
    end else begin
      if(read_A_6__state == 2'b00) begin
        if(read_A_6__ap_start_global__q0) begin
          read_A_6__state <= 2'b01;
        end 
      end 
      if(read_A_6__state == 2'b01) begin
        if(read_A_6__ap_ready) begin
          if(read_A_6__ap_done) begin
            read_A_6__state <= 2'b10;
          end else begin
            read_A_6__state <= 2'b11;
          end
        end 
      end 
      if(read_A_6__state == 2'b11) begin
        if(read_A_6__ap_done) begin
          read_A_6__state <= 2'b10;
        end 
      end 
      if(read_A_6__state == 2'b10) begin
        if(read_A_6__ap_done_global__q0) begin
          read_A_6__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_6__ap_start = (read_A_6__state == 2'b01);
  assign read_A_7__ap_start_global__q0 = ap_start__q0;
  assign read_A_7__is_done__q0 = (read_A_7__state == 2'b10);
  assign read_A_7__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_7__state <= 2'b00;
    end else begin
      if(read_A_7__state == 2'b00) begin
        if(read_A_7__ap_start_global__q0) begin
          read_A_7__state <= 2'b01;
        end 
      end 
      if(read_A_7__state == 2'b01) begin
        if(read_A_7__ap_ready) begin
          if(read_A_7__ap_done) begin
            read_A_7__state <= 2'b10;
          end else begin
            read_A_7__state <= 2'b11;
          end
        end 
      end 
      if(read_A_7__state == 2'b11) begin
        if(read_A_7__ap_done) begin
          read_A_7__state <= 2'b10;
        end 
      end 
      if(read_A_7__state == 2'b10) begin
        if(read_A_7__ap_done_global__q0) begin
          read_A_7__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_7__ap_start = (read_A_7__state == 2'b01);
  assign read_A_8__ap_start_global__q0 = ap_start__q0;
  assign read_A_8__is_done__q0 = (read_A_8__state == 2'b10);
  assign read_A_8__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_8__state <= 2'b00;
    end else begin
      if(read_A_8__state == 2'b00) begin
        if(read_A_8__ap_start_global__q0) begin
          read_A_8__state <= 2'b01;
        end 
      end 
      if(read_A_8__state == 2'b01) begin
        if(read_A_8__ap_ready) begin
          if(read_A_8__ap_done) begin
            read_A_8__state <= 2'b10;
          end else begin
            read_A_8__state <= 2'b11;
          end
        end 
      end 
      if(read_A_8__state == 2'b11) begin
        if(read_A_8__ap_done) begin
          read_A_8__state <= 2'b10;
        end 
      end 
      if(read_A_8__state == 2'b10) begin
        if(read_A_8__ap_done_global__q0) begin
          read_A_8__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_8__ap_start = (read_A_8__state == 2'b01);
  assign read_A_9__ap_start_global__q0 = ap_start__q0;
  assign read_A_9__is_done__q0 = (read_A_9__state == 2'b10);
  assign read_A_9__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_9__state <= 2'b00;
    end else begin
      if(read_A_9__state == 2'b00) begin
        if(read_A_9__ap_start_global__q0) begin
          read_A_9__state <= 2'b01;
        end 
      end 
      if(read_A_9__state == 2'b01) begin
        if(read_A_9__ap_ready) begin
          if(read_A_9__ap_done) begin
            read_A_9__state <= 2'b10;
          end else begin
            read_A_9__state <= 2'b11;
          end
        end 
      end 
      if(read_A_9__state == 2'b11) begin
        if(read_A_9__ap_done) begin
          read_A_9__state <= 2'b10;
        end 
      end 
      if(read_A_9__state == 2'b10) begin
        if(read_A_9__ap_done_global__q0) begin
          read_A_9__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_9__ap_start = (read_A_9__state == 2'b01);
  assign read_A_10__ap_start_global__q0 = ap_start__q0;
  assign read_A_10__is_done__q0 = (read_A_10__state == 2'b10);
  assign read_A_10__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_10__state <= 2'b00;
    end else begin
      if(read_A_10__state == 2'b00) begin
        if(read_A_10__ap_start_global__q0) begin
          read_A_10__state <= 2'b01;
        end 
      end 
      if(read_A_10__state == 2'b01) begin
        if(read_A_10__ap_ready) begin
          if(read_A_10__ap_done) begin
            read_A_10__state <= 2'b10;
          end else begin
            read_A_10__state <= 2'b11;
          end
        end 
      end 
      if(read_A_10__state == 2'b11) begin
        if(read_A_10__ap_done) begin
          read_A_10__state <= 2'b10;
        end 
      end 
      if(read_A_10__state == 2'b10) begin
        if(read_A_10__ap_done_global__q0) begin
          read_A_10__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_10__ap_start = (read_A_10__state == 2'b01);
  assign read_A_11__ap_start_global__q0 = ap_start__q0;
  assign read_A_11__is_done__q0 = (read_A_11__state == 2'b10);
  assign read_A_11__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_11__state <= 2'b00;
    end else begin
      if(read_A_11__state == 2'b00) begin
        if(read_A_11__ap_start_global__q0) begin
          read_A_11__state <= 2'b01;
        end 
      end 
      if(read_A_11__state == 2'b01) begin
        if(read_A_11__ap_ready) begin
          if(read_A_11__ap_done) begin
            read_A_11__state <= 2'b10;
          end else begin
            read_A_11__state <= 2'b11;
          end
        end 
      end 
      if(read_A_11__state == 2'b11) begin
        if(read_A_11__ap_done) begin
          read_A_11__state <= 2'b10;
        end 
      end 
      if(read_A_11__state == 2'b10) begin
        if(read_A_11__ap_done_global__q0) begin
          read_A_11__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_11__ap_start = (read_A_11__state == 2'b01);
  assign read_A_12__ap_start_global__q0 = ap_start__q0;
  assign read_A_12__is_done__q0 = (read_A_12__state == 2'b10);
  assign read_A_12__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_12__state <= 2'b00;
    end else begin
      if(read_A_12__state == 2'b00) begin
        if(read_A_12__ap_start_global__q0) begin
          read_A_12__state <= 2'b01;
        end 
      end 
      if(read_A_12__state == 2'b01) begin
        if(read_A_12__ap_ready) begin
          if(read_A_12__ap_done) begin
            read_A_12__state <= 2'b10;
          end else begin
            read_A_12__state <= 2'b11;
          end
        end 
      end 
      if(read_A_12__state == 2'b11) begin
        if(read_A_12__ap_done) begin
          read_A_12__state <= 2'b10;
        end 
      end 
      if(read_A_12__state == 2'b10) begin
        if(read_A_12__ap_done_global__q0) begin
          read_A_12__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_12__ap_start = (read_A_12__state == 2'b01);
  assign read_A_13__ap_start_global__q0 = ap_start__q0;
  assign read_A_13__is_done__q0 = (read_A_13__state == 2'b10);
  assign read_A_13__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_13__state <= 2'b00;
    end else begin
      if(read_A_13__state == 2'b00) begin
        if(read_A_13__ap_start_global__q0) begin
          read_A_13__state <= 2'b01;
        end 
      end 
      if(read_A_13__state == 2'b01) begin
        if(read_A_13__ap_ready) begin
          if(read_A_13__ap_done) begin
            read_A_13__state <= 2'b10;
          end else begin
            read_A_13__state <= 2'b11;
          end
        end 
      end 
      if(read_A_13__state == 2'b11) begin
        if(read_A_13__ap_done) begin
          read_A_13__state <= 2'b10;
        end 
      end 
      if(read_A_13__state == 2'b10) begin
        if(read_A_13__ap_done_global__q0) begin
          read_A_13__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_13__ap_start = (read_A_13__state == 2'b01);
  assign read_A_14__ap_start_global__q0 = ap_start__q0;
  assign read_A_14__is_done__q0 = (read_A_14__state == 2'b10);
  assign read_A_14__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_14__state <= 2'b00;
    end else begin
      if(read_A_14__state == 2'b00) begin
        if(read_A_14__ap_start_global__q0) begin
          read_A_14__state <= 2'b01;
        end 
      end 
      if(read_A_14__state == 2'b01) begin
        if(read_A_14__ap_ready) begin
          if(read_A_14__ap_done) begin
            read_A_14__state <= 2'b10;
          end else begin
            read_A_14__state <= 2'b11;
          end
        end 
      end 
      if(read_A_14__state == 2'b11) begin
        if(read_A_14__ap_done) begin
          read_A_14__state <= 2'b10;
        end 
      end 
      if(read_A_14__state == 2'b10) begin
        if(read_A_14__ap_done_global__q0) begin
          read_A_14__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_14__ap_start = (read_A_14__state == 2'b01);
  assign read_A_15__ap_start_global__q0 = ap_start__q0;
  assign read_A_15__is_done__q0 = (read_A_15__state == 2'b10);
  assign read_A_15__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_15__state <= 2'b00;
    end else begin
      if(read_A_15__state == 2'b00) begin
        if(read_A_15__ap_start_global__q0) begin
          read_A_15__state <= 2'b01;
        end 
      end 
      if(read_A_15__state == 2'b01) begin
        if(read_A_15__ap_ready) begin
          if(read_A_15__ap_done) begin
            read_A_15__state <= 2'b10;
          end else begin
            read_A_15__state <= 2'b11;
          end
        end 
      end 
      if(read_A_15__state == 2'b11) begin
        if(read_A_15__ap_done) begin
          read_A_15__state <= 2'b10;
        end 
      end 
      if(read_A_15__state == 2'b10) begin
        if(read_A_15__ap_done_global__q0) begin
          read_A_15__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_15__ap_start = (read_A_15__state == 2'b01);
  assign read_A_16__ap_start_global__q0 = ap_start__q0;
  assign read_A_16__is_done__q0 = (read_A_16__state == 2'b10);
  assign read_A_16__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_16__state <= 2'b00;
    end else begin
      if(read_A_16__state == 2'b00) begin
        if(read_A_16__ap_start_global__q0) begin
          read_A_16__state <= 2'b01;
        end 
      end 
      if(read_A_16__state == 2'b01) begin
        if(read_A_16__ap_ready) begin
          if(read_A_16__ap_done) begin
            read_A_16__state <= 2'b10;
          end else begin
            read_A_16__state <= 2'b11;
          end
        end 
      end 
      if(read_A_16__state == 2'b11) begin
        if(read_A_16__ap_done) begin
          read_A_16__state <= 2'b10;
        end 
      end 
      if(read_A_16__state == 2'b10) begin
        if(read_A_16__ap_done_global__q0) begin
          read_A_16__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_16__ap_start = (read_A_16__state == 2'b01);
  assign read_A_17__ap_start_global__q0 = ap_start__q0;
  assign read_A_17__is_done__q0 = (read_A_17__state == 2'b10);
  assign read_A_17__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_17__state <= 2'b00;
    end else begin
      if(read_A_17__state == 2'b00) begin
        if(read_A_17__ap_start_global__q0) begin
          read_A_17__state <= 2'b01;
        end 
      end 
      if(read_A_17__state == 2'b01) begin
        if(read_A_17__ap_ready) begin
          if(read_A_17__ap_done) begin
            read_A_17__state <= 2'b10;
          end else begin
            read_A_17__state <= 2'b11;
          end
        end 
      end 
      if(read_A_17__state == 2'b11) begin
        if(read_A_17__ap_done) begin
          read_A_17__state <= 2'b10;
        end 
      end 
      if(read_A_17__state == 2'b10) begin
        if(read_A_17__ap_done_global__q0) begin
          read_A_17__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_17__ap_start = (read_A_17__state == 2'b01);
  assign read_A_18__ap_start_global__q0 = ap_start__q0;
  assign read_A_18__is_done__q0 = (read_A_18__state == 2'b10);
  assign read_A_18__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_18__state <= 2'b00;
    end else begin
      if(read_A_18__state == 2'b00) begin
        if(read_A_18__ap_start_global__q0) begin
          read_A_18__state <= 2'b01;
        end 
      end 
      if(read_A_18__state == 2'b01) begin
        if(read_A_18__ap_ready) begin
          if(read_A_18__ap_done) begin
            read_A_18__state <= 2'b10;
          end else begin
            read_A_18__state <= 2'b11;
          end
        end 
      end 
      if(read_A_18__state == 2'b11) begin
        if(read_A_18__ap_done) begin
          read_A_18__state <= 2'b10;
        end 
      end 
      if(read_A_18__state == 2'b10) begin
        if(read_A_18__ap_done_global__q0) begin
          read_A_18__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_18__ap_start = (read_A_18__state == 2'b01);
  assign read_A_19__ap_start_global__q0 = ap_start__q0;
  assign read_A_19__is_done__q0 = (read_A_19__state == 2'b10);
  assign read_A_19__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_19__state <= 2'b00;
    end else begin
      if(read_A_19__state == 2'b00) begin
        if(read_A_19__ap_start_global__q0) begin
          read_A_19__state <= 2'b01;
        end 
      end 
      if(read_A_19__state == 2'b01) begin
        if(read_A_19__ap_ready) begin
          if(read_A_19__ap_done) begin
            read_A_19__state <= 2'b10;
          end else begin
            read_A_19__state <= 2'b11;
          end
        end 
      end 
      if(read_A_19__state == 2'b11) begin
        if(read_A_19__ap_done) begin
          read_A_19__state <= 2'b10;
        end 
      end 
      if(read_A_19__state == 2'b10) begin
        if(read_A_19__ap_done_global__q0) begin
          read_A_19__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_19__ap_start = (read_A_19__state == 2'b01);
  assign read_A_20__ap_start_global__q0 = ap_start__q0;
  assign read_A_20__is_done__q0 = (read_A_20__state == 2'b10);
  assign read_A_20__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_20__state <= 2'b00;
    end else begin
      if(read_A_20__state == 2'b00) begin
        if(read_A_20__ap_start_global__q0) begin
          read_A_20__state <= 2'b01;
        end 
      end 
      if(read_A_20__state == 2'b01) begin
        if(read_A_20__ap_ready) begin
          if(read_A_20__ap_done) begin
            read_A_20__state <= 2'b10;
          end else begin
            read_A_20__state <= 2'b11;
          end
        end 
      end 
      if(read_A_20__state == 2'b11) begin
        if(read_A_20__ap_done) begin
          read_A_20__state <= 2'b10;
        end 
      end 
      if(read_A_20__state == 2'b10) begin
        if(read_A_20__ap_done_global__q0) begin
          read_A_20__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_20__ap_start = (read_A_20__state == 2'b01);
  assign read_A_21__ap_start_global__q0 = ap_start__q0;
  assign read_A_21__is_done__q0 = (read_A_21__state == 2'b10);
  assign read_A_21__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_21__state <= 2'b00;
    end else begin
      if(read_A_21__state == 2'b00) begin
        if(read_A_21__ap_start_global__q0) begin
          read_A_21__state <= 2'b01;
        end 
      end 
      if(read_A_21__state == 2'b01) begin
        if(read_A_21__ap_ready) begin
          if(read_A_21__ap_done) begin
            read_A_21__state <= 2'b10;
          end else begin
            read_A_21__state <= 2'b11;
          end
        end 
      end 
      if(read_A_21__state == 2'b11) begin
        if(read_A_21__ap_done) begin
          read_A_21__state <= 2'b10;
        end 
      end 
      if(read_A_21__state == 2'b10) begin
        if(read_A_21__ap_done_global__q0) begin
          read_A_21__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_21__ap_start = (read_A_21__state == 2'b01);
  assign read_A_22__ap_start_global__q0 = ap_start__q0;
  assign read_A_22__is_done__q0 = (read_A_22__state == 2'b10);
  assign read_A_22__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_22__state <= 2'b00;
    end else begin
      if(read_A_22__state == 2'b00) begin
        if(read_A_22__ap_start_global__q0) begin
          read_A_22__state <= 2'b01;
        end 
      end 
      if(read_A_22__state == 2'b01) begin
        if(read_A_22__ap_ready) begin
          if(read_A_22__ap_done) begin
            read_A_22__state <= 2'b10;
          end else begin
            read_A_22__state <= 2'b11;
          end
        end 
      end 
      if(read_A_22__state == 2'b11) begin
        if(read_A_22__ap_done) begin
          read_A_22__state <= 2'b10;
        end 
      end 
      if(read_A_22__state == 2'b10) begin
        if(read_A_22__ap_done_global__q0) begin
          read_A_22__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_22__ap_start = (read_A_22__state == 2'b01);
  assign read_A_23__ap_start_global__q0 = ap_start__q0;
  assign read_A_23__is_done__q0 = (read_A_23__state == 2'b10);
  assign read_A_23__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_23__state <= 2'b00;
    end else begin
      if(read_A_23__state == 2'b00) begin
        if(read_A_23__ap_start_global__q0) begin
          read_A_23__state <= 2'b01;
        end 
      end 
      if(read_A_23__state == 2'b01) begin
        if(read_A_23__ap_ready) begin
          if(read_A_23__ap_done) begin
            read_A_23__state <= 2'b10;
          end else begin
            read_A_23__state <= 2'b11;
          end
        end 
      end 
      if(read_A_23__state == 2'b11) begin
        if(read_A_23__ap_done) begin
          read_A_23__state <= 2'b10;
        end 
      end 
      if(read_A_23__state == 2'b10) begin
        if(read_A_23__ap_done_global__q0) begin
          read_A_23__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_23__ap_start = (read_A_23__state == 2'b01);
  assign read_A_24__ap_start_global__q0 = ap_start__q0;
  assign read_A_24__is_done__q0 = (read_A_24__state == 2'b10);
  assign read_A_24__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_24__state <= 2'b00;
    end else begin
      if(read_A_24__state == 2'b00) begin
        if(read_A_24__ap_start_global__q0) begin
          read_A_24__state <= 2'b01;
        end 
      end 
      if(read_A_24__state == 2'b01) begin
        if(read_A_24__ap_ready) begin
          if(read_A_24__ap_done) begin
            read_A_24__state <= 2'b10;
          end else begin
            read_A_24__state <= 2'b11;
          end
        end 
      end 
      if(read_A_24__state == 2'b11) begin
        if(read_A_24__ap_done) begin
          read_A_24__state <= 2'b10;
        end 
      end 
      if(read_A_24__state == 2'b10) begin
        if(read_A_24__ap_done_global__q0) begin
          read_A_24__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_24__ap_start = (read_A_24__state == 2'b01);
  assign read_A_25__ap_start_global__q0 = ap_start__q0;
  assign read_A_25__is_done__q0 = (read_A_25__state == 2'b10);
  assign read_A_25__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_25__state <= 2'b00;
    end else begin
      if(read_A_25__state == 2'b00) begin
        if(read_A_25__ap_start_global__q0) begin
          read_A_25__state <= 2'b01;
        end 
      end 
      if(read_A_25__state == 2'b01) begin
        if(read_A_25__ap_ready) begin
          if(read_A_25__ap_done) begin
            read_A_25__state <= 2'b10;
          end else begin
            read_A_25__state <= 2'b11;
          end
        end 
      end 
      if(read_A_25__state == 2'b11) begin
        if(read_A_25__ap_done) begin
          read_A_25__state <= 2'b10;
        end 
      end 
      if(read_A_25__state == 2'b10) begin
        if(read_A_25__ap_done_global__q0) begin
          read_A_25__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_25__ap_start = (read_A_25__state == 2'b01);
  assign read_A_26__ap_start_global__q0 = ap_start__q0;
  assign read_A_26__is_done__q0 = (read_A_26__state == 2'b10);
  assign read_A_26__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_26__state <= 2'b00;
    end else begin
      if(read_A_26__state == 2'b00) begin
        if(read_A_26__ap_start_global__q0) begin
          read_A_26__state <= 2'b01;
        end 
      end 
      if(read_A_26__state == 2'b01) begin
        if(read_A_26__ap_ready) begin
          if(read_A_26__ap_done) begin
            read_A_26__state <= 2'b10;
          end else begin
            read_A_26__state <= 2'b11;
          end
        end 
      end 
      if(read_A_26__state == 2'b11) begin
        if(read_A_26__ap_done) begin
          read_A_26__state <= 2'b10;
        end 
      end 
      if(read_A_26__state == 2'b10) begin
        if(read_A_26__ap_done_global__q0) begin
          read_A_26__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_26__ap_start = (read_A_26__state == 2'b01);
  assign read_A_27__ap_start_global__q0 = ap_start__q0;
  assign read_A_27__is_done__q0 = (read_A_27__state == 2'b10);
  assign read_A_27__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_27__state <= 2'b00;
    end else begin
      if(read_A_27__state == 2'b00) begin
        if(read_A_27__ap_start_global__q0) begin
          read_A_27__state <= 2'b01;
        end 
      end 
      if(read_A_27__state == 2'b01) begin
        if(read_A_27__ap_ready) begin
          if(read_A_27__ap_done) begin
            read_A_27__state <= 2'b10;
          end else begin
            read_A_27__state <= 2'b11;
          end
        end 
      end 
      if(read_A_27__state == 2'b11) begin
        if(read_A_27__ap_done) begin
          read_A_27__state <= 2'b10;
        end 
      end 
      if(read_A_27__state == 2'b10) begin
        if(read_A_27__ap_done_global__q0) begin
          read_A_27__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_27__ap_start = (read_A_27__state == 2'b01);
  assign read_A_28__ap_start_global__q0 = ap_start__q0;
  assign read_A_28__is_done__q0 = (read_A_28__state == 2'b10);
  assign read_A_28__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_28__state <= 2'b00;
    end else begin
      if(read_A_28__state == 2'b00) begin
        if(read_A_28__ap_start_global__q0) begin
          read_A_28__state <= 2'b01;
        end 
      end 
      if(read_A_28__state == 2'b01) begin
        if(read_A_28__ap_ready) begin
          if(read_A_28__ap_done) begin
            read_A_28__state <= 2'b10;
          end else begin
            read_A_28__state <= 2'b11;
          end
        end 
      end 
      if(read_A_28__state == 2'b11) begin
        if(read_A_28__ap_done) begin
          read_A_28__state <= 2'b10;
        end 
      end 
      if(read_A_28__state == 2'b10) begin
        if(read_A_28__ap_done_global__q0) begin
          read_A_28__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_28__ap_start = (read_A_28__state == 2'b01);
  assign read_A_29__ap_start_global__q0 = ap_start__q0;
  assign read_A_29__is_done__q0 = (read_A_29__state == 2'b10);
  assign read_A_29__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_29__state <= 2'b00;
    end else begin
      if(read_A_29__state == 2'b00) begin
        if(read_A_29__ap_start_global__q0) begin
          read_A_29__state <= 2'b01;
        end 
      end 
      if(read_A_29__state == 2'b01) begin
        if(read_A_29__ap_ready) begin
          if(read_A_29__ap_done) begin
            read_A_29__state <= 2'b10;
          end else begin
            read_A_29__state <= 2'b11;
          end
        end 
      end 
      if(read_A_29__state == 2'b11) begin
        if(read_A_29__ap_done) begin
          read_A_29__state <= 2'b10;
        end 
      end 
      if(read_A_29__state == 2'b10) begin
        if(read_A_29__ap_done_global__q0) begin
          read_A_29__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_29__ap_start = (read_A_29__state == 2'b01);
  assign read_A_30__ap_start_global__q0 = ap_start__q0;
  assign read_A_30__is_done__q0 = (read_A_30__state == 2'b10);
  assign read_A_30__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_30__state <= 2'b00;
    end else begin
      if(read_A_30__state == 2'b00) begin
        if(read_A_30__ap_start_global__q0) begin
          read_A_30__state <= 2'b01;
        end 
      end 
      if(read_A_30__state == 2'b01) begin
        if(read_A_30__ap_ready) begin
          if(read_A_30__ap_done) begin
            read_A_30__state <= 2'b10;
          end else begin
            read_A_30__state <= 2'b11;
          end
        end 
      end 
      if(read_A_30__state == 2'b11) begin
        if(read_A_30__ap_done) begin
          read_A_30__state <= 2'b10;
        end 
      end 
      if(read_A_30__state == 2'b10) begin
        if(read_A_30__ap_done_global__q0) begin
          read_A_30__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_30__ap_start = (read_A_30__state == 2'b01);
  assign read_A_31__ap_start_global__q0 = ap_start__q0;
  assign read_A_31__is_done__q0 = (read_A_31__state == 2'b10);
  assign read_A_31__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_31__state <= 2'b00;
    end else begin
      if(read_A_31__state == 2'b00) begin
        if(read_A_31__ap_start_global__q0) begin
          read_A_31__state <= 2'b01;
        end 
      end 
      if(read_A_31__state == 2'b01) begin
        if(read_A_31__ap_ready) begin
          if(read_A_31__ap_done) begin
            read_A_31__state <= 2'b10;
          end else begin
            read_A_31__state <= 2'b11;
          end
        end 
      end 
      if(read_A_31__state == 2'b11) begin
        if(read_A_31__ap_done) begin
          read_A_31__state <= 2'b10;
        end 
      end 
      if(read_A_31__state == 2'b10) begin
        if(read_A_31__ap_done_global__q0) begin
          read_A_31__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_31__ap_start = (read_A_31__state == 2'b01);
  assign read_A_32__ap_start_global__q0 = ap_start__q0;
  assign read_A_32__is_done__q0 = (read_A_32__state == 2'b10);
  assign read_A_32__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_32__state <= 2'b00;
    end else begin
      if(read_A_32__state == 2'b00) begin
        if(read_A_32__ap_start_global__q0) begin
          read_A_32__state <= 2'b01;
        end 
      end 
      if(read_A_32__state == 2'b01) begin
        if(read_A_32__ap_ready) begin
          if(read_A_32__ap_done) begin
            read_A_32__state <= 2'b10;
          end else begin
            read_A_32__state <= 2'b11;
          end
        end 
      end 
      if(read_A_32__state == 2'b11) begin
        if(read_A_32__ap_done) begin
          read_A_32__state <= 2'b10;
        end 
      end 
      if(read_A_32__state == 2'b10) begin
        if(read_A_32__ap_done_global__q0) begin
          read_A_32__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_32__ap_start = (read_A_32__state == 2'b01);
  assign read_A_33__ap_start_global__q0 = ap_start__q0;
  assign read_A_33__is_done__q0 = (read_A_33__state == 2'b10);
  assign read_A_33__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_33__state <= 2'b00;
    end else begin
      if(read_A_33__state == 2'b00) begin
        if(read_A_33__ap_start_global__q0) begin
          read_A_33__state <= 2'b01;
        end 
      end 
      if(read_A_33__state == 2'b01) begin
        if(read_A_33__ap_ready) begin
          if(read_A_33__ap_done) begin
            read_A_33__state <= 2'b10;
          end else begin
            read_A_33__state <= 2'b11;
          end
        end 
      end 
      if(read_A_33__state == 2'b11) begin
        if(read_A_33__ap_done) begin
          read_A_33__state <= 2'b10;
        end 
      end 
      if(read_A_33__state == 2'b10) begin
        if(read_A_33__ap_done_global__q0) begin
          read_A_33__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_33__ap_start = (read_A_33__state == 2'b01);
  assign read_A_34__ap_start_global__q0 = ap_start__q0;
  assign read_A_34__is_done__q0 = (read_A_34__state == 2'b10);
  assign read_A_34__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_34__state <= 2'b00;
    end else begin
      if(read_A_34__state == 2'b00) begin
        if(read_A_34__ap_start_global__q0) begin
          read_A_34__state <= 2'b01;
        end 
      end 
      if(read_A_34__state == 2'b01) begin
        if(read_A_34__ap_ready) begin
          if(read_A_34__ap_done) begin
            read_A_34__state <= 2'b10;
          end else begin
            read_A_34__state <= 2'b11;
          end
        end 
      end 
      if(read_A_34__state == 2'b11) begin
        if(read_A_34__ap_done) begin
          read_A_34__state <= 2'b10;
        end 
      end 
      if(read_A_34__state == 2'b10) begin
        if(read_A_34__ap_done_global__q0) begin
          read_A_34__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_34__ap_start = (read_A_34__state == 2'b01);
  assign read_A_35__ap_start_global__q0 = ap_start__q0;
  assign read_A_35__is_done__q0 = (read_A_35__state == 2'b10);
  assign read_A_35__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_35__state <= 2'b00;
    end else begin
      if(read_A_35__state == 2'b00) begin
        if(read_A_35__ap_start_global__q0) begin
          read_A_35__state <= 2'b01;
        end 
      end 
      if(read_A_35__state == 2'b01) begin
        if(read_A_35__ap_ready) begin
          if(read_A_35__ap_done) begin
            read_A_35__state <= 2'b10;
          end else begin
            read_A_35__state <= 2'b11;
          end
        end 
      end 
      if(read_A_35__state == 2'b11) begin
        if(read_A_35__ap_done) begin
          read_A_35__state <= 2'b10;
        end 
      end 
      if(read_A_35__state == 2'b10) begin
        if(read_A_35__ap_done_global__q0) begin
          read_A_35__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_35__ap_start = (read_A_35__state == 2'b01);
  assign read_A_36__ap_start_global__q0 = ap_start__q0;
  assign read_A_36__is_done__q0 = (read_A_36__state == 2'b10);
  assign read_A_36__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_36__state <= 2'b00;
    end else begin
      if(read_A_36__state == 2'b00) begin
        if(read_A_36__ap_start_global__q0) begin
          read_A_36__state <= 2'b01;
        end 
      end 
      if(read_A_36__state == 2'b01) begin
        if(read_A_36__ap_ready) begin
          if(read_A_36__ap_done) begin
            read_A_36__state <= 2'b10;
          end else begin
            read_A_36__state <= 2'b11;
          end
        end 
      end 
      if(read_A_36__state == 2'b11) begin
        if(read_A_36__ap_done) begin
          read_A_36__state <= 2'b10;
        end 
      end 
      if(read_A_36__state == 2'b10) begin
        if(read_A_36__ap_done_global__q0) begin
          read_A_36__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_36__ap_start = (read_A_36__state == 2'b01);
  assign read_A_37__ap_start_global__q0 = ap_start__q0;
  assign read_A_37__is_done__q0 = (read_A_37__state == 2'b10);
  assign read_A_37__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_37__state <= 2'b00;
    end else begin
      if(read_A_37__state == 2'b00) begin
        if(read_A_37__ap_start_global__q0) begin
          read_A_37__state <= 2'b01;
        end 
      end 
      if(read_A_37__state == 2'b01) begin
        if(read_A_37__ap_ready) begin
          if(read_A_37__ap_done) begin
            read_A_37__state <= 2'b10;
          end else begin
            read_A_37__state <= 2'b11;
          end
        end 
      end 
      if(read_A_37__state == 2'b11) begin
        if(read_A_37__ap_done) begin
          read_A_37__state <= 2'b10;
        end 
      end 
      if(read_A_37__state == 2'b10) begin
        if(read_A_37__ap_done_global__q0) begin
          read_A_37__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_37__ap_start = (read_A_37__state == 2'b01);
  assign read_A_38__ap_start_global__q0 = ap_start__q0;
  assign read_A_38__is_done__q0 = (read_A_38__state == 2'b10);
  assign read_A_38__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_38__state <= 2'b00;
    end else begin
      if(read_A_38__state == 2'b00) begin
        if(read_A_38__ap_start_global__q0) begin
          read_A_38__state <= 2'b01;
        end 
      end 
      if(read_A_38__state == 2'b01) begin
        if(read_A_38__ap_ready) begin
          if(read_A_38__ap_done) begin
            read_A_38__state <= 2'b10;
          end else begin
            read_A_38__state <= 2'b11;
          end
        end 
      end 
      if(read_A_38__state == 2'b11) begin
        if(read_A_38__ap_done) begin
          read_A_38__state <= 2'b10;
        end 
      end 
      if(read_A_38__state == 2'b10) begin
        if(read_A_38__ap_done_global__q0) begin
          read_A_38__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_38__ap_start = (read_A_38__state == 2'b01);
  assign read_A_39__ap_start_global__q0 = ap_start__q0;
  assign read_A_39__is_done__q0 = (read_A_39__state == 2'b10);
  assign read_A_39__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_39__state <= 2'b00;
    end else begin
      if(read_A_39__state == 2'b00) begin
        if(read_A_39__ap_start_global__q0) begin
          read_A_39__state <= 2'b01;
        end 
      end 
      if(read_A_39__state == 2'b01) begin
        if(read_A_39__ap_ready) begin
          if(read_A_39__ap_done) begin
            read_A_39__state <= 2'b10;
          end else begin
            read_A_39__state <= 2'b11;
          end
        end 
      end 
      if(read_A_39__state == 2'b11) begin
        if(read_A_39__ap_done) begin
          read_A_39__state <= 2'b10;
        end 
      end 
      if(read_A_39__state == 2'b10) begin
        if(read_A_39__ap_done_global__q0) begin
          read_A_39__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_39__ap_start = (read_A_39__state == 2'b01);
  assign read_A_40__ap_start_global__q0 = ap_start__q0;
  assign read_A_40__is_done__q0 = (read_A_40__state == 2'b10);
  assign read_A_40__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_40__state <= 2'b00;
    end else begin
      if(read_A_40__state == 2'b00) begin
        if(read_A_40__ap_start_global__q0) begin
          read_A_40__state <= 2'b01;
        end 
      end 
      if(read_A_40__state == 2'b01) begin
        if(read_A_40__ap_ready) begin
          if(read_A_40__ap_done) begin
            read_A_40__state <= 2'b10;
          end else begin
            read_A_40__state <= 2'b11;
          end
        end 
      end 
      if(read_A_40__state == 2'b11) begin
        if(read_A_40__ap_done) begin
          read_A_40__state <= 2'b10;
        end 
      end 
      if(read_A_40__state == 2'b10) begin
        if(read_A_40__ap_done_global__q0) begin
          read_A_40__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_40__ap_start = (read_A_40__state == 2'b01);
  assign read_A_41__ap_start_global__q0 = ap_start__q0;
  assign read_A_41__is_done__q0 = (read_A_41__state == 2'b10);
  assign read_A_41__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_41__state <= 2'b00;
    end else begin
      if(read_A_41__state == 2'b00) begin
        if(read_A_41__ap_start_global__q0) begin
          read_A_41__state <= 2'b01;
        end 
      end 
      if(read_A_41__state == 2'b01) begin
        if(read_A_41__ap_ready) begin
          if(read_A_41__ap_done) begin
            read_A_41__state <= 2'b10;
          end else begin
            read_A_41__state <= 2'b11;
          end
        end 
      end 
      if(read_A_41__state == 2'b11) begin
        if(read_A_41__ap_done) begin
          read_A_41__state <= 2'b10;
        end 
      end 
      if(read_A_41__state == 2'b10) begin
        if(read_A_41__ap_done_global__q0) begin
          read_A_41__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_41__ap_start = (read_A_41__state == 2'b01);
  assign read_A_42__ap_start_global__q0 = ap_start__q0;
  assign read_A_42__is_done__q0 = (read_A_42__state == 2'b10);
  assign read_A_42__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_42__state <= 2'b00;
    end else begin
      if(read_A_42__state == 2'b00) begin
        if(read_A_42__ap_start_global__q0) begin
          read_A_42__state <= 2'b01;
        end 
      end 
      if(read_A_42__state == 2'b01) begin
        if(read_A_42__ap_ready) begin
          if(read_A_42__ap_done) begin
            read_A_42__state <= 2'b10;
          end else begin
            read_A_42__state <= 2'b11;
          end
        end 
      end 
      if(read_A_42__state == 2'b11) begin
        if(read_A_42__ap_done) begin
          read_A_42__state <= 2'b10;
        end 
      end 
      if(read_A_42__state == 2'b10) begin
        if(read_A_42__ap_done_global__q0) begin
          read_A_42__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_42__ap_start = (read_A_42__state == 2'b01);
  assign read_A_43__ap_start_global__q0 = ap_start__q0;
  assign read_A_43__is_done__q0 = (read_A_43__state == 2'b10);
  assign read_A_43__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_43__state <= 2'b00;
    end else begin
      if(read_A_43__state == 2'b00) begin
        if(read_A_43__ap_start_global__q0) begin
          read_A_43__state <= 2'b01;
        end 
      end 
      if(read_A_43__state == 2'b01) begin
        if(read_A_43__ap_ready) begin
          if(read_A_43__ap_done) begin
            read_A_43__state <= 2'b10;
          end else begin
            read_A_43__state <= 2'b11;
          end
        end 
      end 
      if(read_A_43__state == 2'b11) begin
        if(read_A_43__ap_done) begin
          read_A_43__state <= 2'b10;
        end 
      end 
      if(read_A_43__state == 2'b10) begin
        if(read_A_43__ap_done_global__q0) begin
          read_A_43__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_43__ap_start = (read_A_43__state == 2'b01);
  assign read_A_44__ap_start_global__q0 = ap_start__q0;
  assign read_A_44__is_done__q0 = (read_A_44__state == 2'b10);
  assign read_A_44__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_44__state <= 2'b00;
    end else begin
      if(read_A_44__state == 2'b00) begin
        if(read_A_44__ap_start_global__q0) begin
          read_A_44__state <= 2'b01;
        end 
      end 
      if(read_A_44__state == 2'b01) begin
        if(read_A_44__ap_ready) begin
          if(read_A_44__ap_done) begin
            read_A_44__state <= 2'b10;
          end else begin
            read_A_44__state <= 2'b11;
          end
        end 
      end 
      if(read_A_44__state == 2'b11) begin
        if(read_A_44__ap_done) begin
          read_A_44__state <= 2'b10;
        end 
      end 
      if(read_A_44__state == 2'b10) begin
        if(read_A_44__ap_done_global__q0) begin
          read_A_44__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_44__ap_start = (read_A_44__state == 2'b01);
  assign read_A_45__ap_start_global__q0 = ap_start__q0;
  assign read_A_45__is_done__q0 = (read_A_45__state == 2'b10);
  assign read_A_45__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_45__state <= 2'b00;
    end else begin
      if(read_A_45__state == 2'b00) begin
        if(read_A_45__ap_start_global__q0) begin
          read_A_45__state <= 2'b01;
        end 
      end 
      if(read_A_45__state == 2'b01) begin
        if(read_A_45__ap_ready) begin
          if(read_A_45__ap_done) begin
            read_A_45__state <= 2'b10;
          end else begin
            read_A_45__state <= 2'b11;
          end
        end 
      end 
      if(read_A_45__state == 2'b11) begin
        if(read_A_45__ap_done) begin
          read_A_45__state <= 2'b10;
        end 
      end 
      if(read_A_45__state == 2'b10) begin
        if(read_A_45__ap_done_global__q0) begin
          read_A_45__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_45__ap_start = (read_A_45__state == 2'b01);
  assign read_A_46__ap_start_global__q0 = ap_start__q0;
  assign read_A_46__is_done__q0 = (read_A_46__state == 2'b10);
  assign read_A_46__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_46__state <= 2'b00;
    end else begin
      if(read_A_46__state == 2'b00) begin
        if(read_A_46__ap_start_global__q0) begin
          read_A_46__state <= 2'b01;
        end 
      end 
      if(read_A_46__state == 2'b01) begin
        if(read_A_46__ap_ready) begin
          if(read_A_46__ap_done) begin
            read_A_46__state <= 2'b10;
          end else begin
            read_A_46__state <= 2'b11;
          end
        end 
      end 
      if(read_A_46__state == 2'b11) begin
        if(read_A_46__ap_done) begin
          read_A_46__state <= 2'b10;
        end 
      end 
      if(read_A_46__state == 2'b10) begin
        if(read_A_46__ap_done_global__q0) begin
          read_A_46__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_46__ap_start = (read_A_46__state == 2'b01);
  assign read_A_47__ap_start_global__q0 = ap_start__q0;
  assign read_A_47__is_done__q0 = (read_A_47__state == 2'b10);
  assign read_A_47__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_47__state <= 2'b00;
    end else begin
      if(read_A_47__state == 2'b00) begin
        if(read_A_47__ap_start_global__q0) begin
          read_A_47__state <= 2'b01;
        end 
      end 
      if(read_A_47__state == 2'b01) begin
        if(read_A_47__ap_ready) begin
          if(read_A_47__ap_done) begin
            read_A_47__state <= 2'b10;
          end else begin
            read_A_47__state <= 2'b11;
          end
        end 
      end 
      if(read_A_47__state == 2'b11) begin
        if(read_A_47__ap_done) begin
          read_A_47__state <= 2'b10;
        end 
      end 
      if(read_A_47__state == 2'b10) begin
        if(read_A_47__ap_done_global__q0) begin
          read_A_47__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_47__ap_start = (read_A_47__state == 2'b01);
  assign read_A_48__ap_start_global__q0 = ap_start__q0;
  assign read_A_48__is_done__q0 = (read_A_48__state == 2'b10);
  assign read_A_48__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_48__state <= 2'b00;
    end else begin
      if(read_A_48__state == 2'b00) begin
        if(read_A_48__ap_start_global__q0) begin
          read_A_48__state <= 2'b01;
        end 
      end 
      if(read_A_48__state == 2'b01) begin
        if(read_A_48__ap_ready) begin
          if(read_A_48__ap_done) begin
            read_A_48__state <= 2'b10;
          end else begin
            read_A_48__state <= 2'b11;
          end
        end 
      end 
      if(read_A_48__state == 2'b11) begin
        if(read_A_48__ap_done) begin
          read_A_48__state <= 2'b10;
        end 
      end 
      if(read_A_48__state == 2'b10) begin
        if(read_A_48__ap_done_global__q0) begin
          read_A_48__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_48__ap_start = (read_A_48__state == 2'b01);
  assign read_A_49__ap_start_global__q0 = ap_start__q0;
  assign read_A_49__is_done__q0 = (read_A_49__state == 2'b10);
  assign read_A_49__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_49__state <= 2'b00;
    end else begin
      if(read_A_49__state == 2'b00) begin
        if(read_A_49__ap_start_global__q0) begin
          read_A_49__state <= 2'b01;
        end 
      end 
      if(read_A_49__state == 2'b01) begin
        if(read_A_49__ap_ready) begin
          if(read_A_49__ap_done) begin
            read_A_49__state <= 2'b10;
          end else begin
            read_A_49__state <= 2'b11;
          end
        end 
      end 
      if(read_A_49__state == 2'b11) begin
        if(read_A_49__ap_done) begin
          read_A_49__state <= 2'b10;
        end 
      end 
      if(read_A_49__state == 2'b10) begin
        if(read_A_49__ap_done_global__q0) begin
          read_A_49__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_49__ap_start = (read_A_49__state == 2'b01);
  assign read_A_50__ap_start_global__q0 = ap_start__q0;
  assign read_A_50__is_done__q0 = (read_A_50__state == 2'b10);
  assign read_A_50__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_50__state <= 2'b00;
    end else begin
      if(read_A_50__state == 2'b00) begin
        if(read_A_50__ap_start_global__q0) begin
          read_A_50__state <= 2'b01;
        end 
      end 
      if(read_A_50__state == 2'b01) begin
        if(read_A_50__ap_ready) begin
          if(read_A_50__ap_done) begin
            read_A_50__state <= 2'b10;
          end else begin
            read_A_50__state <= 2'b11;
          end
        end 
      end 
      if(read_A_50__state == 2'b11) begin
        if(read_A_50__ap_done) begin
          read_A_50__state <= 2'b10;
        end 
      end 
      if(read_A_50__state == 2'b10) begin
        if(read_A_50__ap_done_global__q0) begin
          read_A_50__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_50__ap_start = (read_A_50__state == 2'b01);
  assign read_A_51__ap_start_global__q0 = ap_start__q0;
  assign read_A_51__is_done__q0 = (read_A_51__state == 2'b10);
  assign read_A_51__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_51__state <= 2'b00;
    end else begin
      if(read_A_51__state == 2'b00) begin
        if(read_A_51__ap_start_global__q0) begin
          read_A_51__state <= 2'b01;
        end 
      end 
      if(read_A_51__state == 2'b01) begin
        if(read_A_51__ap_ready) begin
          if(read_A_51__ap_done) begin
            read_A_51__state <= 2'b10;
          end else begin
            read_A_51__state <= 2'b11;
          end
        end 
      end 
      if(read_A_51__state == 2'b11) begin
        if(read_A_51__ap_done) begin
          read_A_51__state <= 2'b10;
        end 
      end 
      if(read_A_51__state == 2'b10) begin
        if(read_A_51__ap_done_global__q0) begin
          read_A_51__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_51__ap_start = (read_A_51__state == 2'b01);
  assign read_A_52__ap_start_global__q0 = ap_start__q0;
  assign read_A_52__is_done__q0 = (read_A_52__state == 2'b10);
  assign read_A_52__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_52__state <= 2'b00;
    end else begin
      if(read_A_52__state == 2'b00) begin
        if(read_A_52__ap_start_global__q0) begin
          read_A_52__state <= 2'b01;
        end 
      end 
      if(read_A_52__state == 2'b01) begin
        if(read_A_52__ap_ready) begin
          if(read_A_52__ap_done) begin
            read_A_52__state <= 2'b10;
          end else begin
            read_A_52__state <= 2'b11;
          end
        end 
      end 
      if(read_A_52__state == 2'b11) begin
        if(read_A_52__ap_done) begin
          read_A_52__state <= 2'b10;
        end 
      end 
      if(read_A_52__state == 2'b10) begin
        if(read_A_52__ap_done_global__q0) begin
          read_A_52__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_52__ap_start = (read_A_52__state == 2'b01);
  assign read_A_53__ap_start_global__q0 = ap_start__q0;
  assign read_A_53__is_done__q0 = (read_A_53__state == 2'b10);
  assign read_A_53__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_53__state <= 2'b00;
    end else begin
      if(read_A_53__state == 2'b00) begin
        if(read_A_53__ap_start_global__q0) begin
          read_A_53__state <= 2'b01;
        end 
      end 
      if(read_A_53__state == 2'b01) begin
        if(read_A_53__ap_ready) begin
          if(read_A_53__ap_done) begin
            read_A_53__state <= 2'b10;
          end else begin
            read_A_53__state <= 2'b11;
          end
        end 
      end 
      if(read_A_53__state == 2'b11) begin
        if(read_A_53__ap_done) begin
          read_A_53__state <= 2'b10;
        end 
      end 
      if(read_A_53__state == 2'b10) begin
        if(read_A_53__ap_done_global__q0) begin
          read_A_53__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_53__ap_start = (read_A_53__state == 2'b01);
  assign read_A_54__ap_start_global__q0 = ap_start__q0;
  assign read_A_54__is_done__q0 = (read_A_54__state == 2'b10);
  assign read_A_54__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_54__state <= 2'b00;
    end else begin
      if(read_A_54__state == 2'b00) begin
        if(read_A_54__ap_start_global__q0) begin
          read_A_54__state <= 2'b01;
        end 
      end 
      if(read_A_54__state == 2'b01) begin
        if(read_A_54__ap_ready) begin
          if(read_A_54__ap_done) begin
            read_A_54__state <= 2'b10;
          end else begin
            read_A_54__state <= 2'b11;
          end
        end 
      end 
      if(read_A_54__state == 2'b11) begin
        if(read_A_54__ap_done) begin
          read_A_54__state <= 2'b10;
        end 
      end 
      if(read_A_54__state == 2'b10) begin
        if(read_A_54__ap_done_global__q0) begin
          read_A_54__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_54__ap_start = (read_A_54__state == 2'b01);
  assign read_A_55__ap_start_global__q0 = ap_start__q0;
  assign read_A_55__is_done__q0 = (read_A_55__state == 2'b10);
  assign read_A_55__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_55__state <= 2'b00;
    end else begin
      if(read_A_55__state == 2'b00) begin
        if(read_A_55__ap_start_global__q0) begin
          read_A_55__state <= 2'b01;
        end 
      end 
      if(read_A_55__state == 2'b01) begin
        if(read_A_55__ap_ready) begin
          if(read_A_55__ap_done) begin
            read_A_55__state <= 2'b10;
          end else begin
            read_A_55__state <= 2'b11;
          end
        end 
      end 
      if(read_A_55__state == 2'b11) begin
        if(read_A_55__ap_done) begin
          read_A_55__state <= 2'b10;
        end 
      end 
      if(read_A_55__state == 2'b10) begin
        if(read_A_55__ap_done_global__q0) begin
          read_A_55__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_A_55__ap_start = (read_A_55__state == 2'b01);
  assign read_X_0__ap_start_global__q0 = ap_start__q0;
  assign read_X_0__is_done__q0 = (read_X_0__state == 2'b10);
  assign read_X_0__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_X_0__state <= 2'b00;
    end else begin
      if(read_X_0__state == 2'b00) begin
        if(read_X_0__ap_start_global__q0) begin
          read_X_0__state <= 2'b01;
        end 
      end 
      if(read_X_0__state == 2'b01) begin
        if(read_X_0__ap_ready) begin
          if(read_X_0__ap_done) begin
            read_X_0__state <= 2'b10;
          end else begin
            read_X_0__state <= 2'b11;
          end
        end 
      end 
      if(read_X_0__state == 2'b11) begin
        if(read_X_0__ap_done) begin
          read_X_0__state <= 2'b10;
        end 
      end 
      if(read_X_0__state == 2'b10) begin
        if(read_X_0__ap_done_global__q0) begin
          read_X_0__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_X_0__ap_start = (read_X_0__state == 2'b01);
  assign read_Y_0__ap_start_global__q0 = ap_start__q0;
  assign read_Y_0__is_done__q0 = (read_Y_0__state == 2'b10);
  assign read_Y_0__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_Y_0__state <= 2'b00;
    end else begin
      if(read_Y_0__state == 2'b00) begin
        if(read_Y_0__ap_start_global__q0) begin
          read_Y_0__state <= 2'b01;
        end 
      end 
      if(read_Y_0__state == 2'b01) begin
        if(read_Y_0__ap_ready) begin
          if(read_Y_0__ap_done) begin
            read_Y_0__state <= 2'b10;
          end else begin
            read_Y_0__state <= 2'b11;
          end
        end 
      end 
      if(read_Y_0__state == 2'b11) begin
        if(read_Y_0__ap_done) begin
          read_Y_0__state <= 2'b10;
        end 
      end 
      if(read_Y_0__state == 2'b10) begin
        if(read_Y_0__ap_done_global__q0) begin
          read_Y_0__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_Y_0__ap_start = (read_Y_0__state == 2'b01);
  assign read_edge_list_ptr_0__ap_start_global__q0 = ap_start__q0;
  assign read_edge_list_ptr_0__is_done__q0 = (read_edge_list_ptr_0__state == 2'b10);
  assign read_edge_list_ptr_0__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_edge_list_ptr_0__state <= 2'b00;
    end else begin
      if(read_edge_list_ptr_0__state == 2'b00) begin
        if(read_edge_list_ptr_0__ap_start_global__q0) begin
          read_edge_list_ptr_0__state <= 2'b01;
        end 
      end 
      if(read_edge_list_ptr_0__state == 2'b01) begin
        if(read_edge_list_ptr_0__ap_ready) begin
          if(read_edge_list_ptr_0__ap_done) begin
            read_edge_list_ptr_0__state <= 2'b10;
          end else begin
            read_edge_list_ptr_0__state <= 2'b11;
          end
        end 
      end 
      if(read_edge_list_ptr_0__state == 2'b11) begin
        if(read_edge_list_ptr_0__ap_done) begin
          read_edge_list_ptr_0__state <= 2'b10;
        end 
      end 
      if(read_edge_list_ptr_0__state == 2'b10) begin
        if(read_edge_list_ptr_0__ap_done_global__q0) begin
          read_edge_list_ptr_0__state <= 2'b00;
        end 
      end 
    end
  end
  assign read_edge_list_ptr_0__ap_start = (read_edge_list_ptr_0__state == 2'b01);
  assign write_Y_0__ap_start_global__q0 = ap_start__q0;
  assign write_Y_0__is_done__q0 = (write_Y_0__state == 2'b10);
  assign write_Y_0__ap_done_global__q0 = ap_done__q0;
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      write_Y_0__state <= 2'b00;
    end else begin
      if(write_Y_0__state == 2'b00) begin
        if(write_Y_0__ap_start_global__q0) begin
          write_Y_0__state <= 2'b01;
        end 
      end 
      if(write_Y_0__state == 2'b01) begin
        if(write_Y_0__ap_ready) begin
          if(write_Y_0__ap_done) begin
            write_Y_0__state <= 2'b10;
          end else begin
            write_Y_0__state <= 2'b11;
          end
        end 
      end 
      if(write_Y_0__state == 2'b11) begin
        if(write_Y_0__ap_done) begin
          write_Y_0__state <= 2'b10;
        end 
      end 
      if(write_Y_0__state == 2'b10) begin
        if(write_Y_0__ap_done_global__q0) begin
          write_Y_0__state <= 2'b00;
        end 
      end 
    end
  end
  assign write_Y_0__ap_start = (write_Y_0__state == 2'b01);
  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      tapa_state <= 2'b00;
    end else begin
      case(tapa_state)
        2'b00: begin
          if(ap_start__q0) begin
            tapa_state <= 2'b01;
          end 
        end
        2'b01: begin
          if(Arbiter_Y_0__is_done__q0 && Arbiter_Y_1__is_done__q0 && Arbiter_Y_2__is_done__q0 && Arbiter_Y_3__is_done__q0 && Arbiter_Y_4__is_done__q0 && Arbiter_Y_5__is_done__q0 && Arbiter_Y_6__is_done__q0 && Arbiter_Y_7__is_done__q0 && FloatvMultConst_0__is_done__q0 && FloatvMultConst_1__is_done__q0 && PEG_Xvec_0__is_done__q0 && PEG_Xvec_1__is_done__q0 && PEG_Xvec_2__is_done__q0 && PEG_Xvec_3__is_done__q0 && PEG_Xvec_4__is_done__q0 && PEG_Xvec_5__is_done__q0 && PEG_Xvec_6__is_done__q0 && PEG_Xvec_7__is_done__q0 && PEG_Xvec_8__is_done__q0 && PEG_Xvec_9__is_done__q0 && PEG_Xvec_10__is_done__q0 && PEG_Xvec_11__is_done__q0 && PEG_Xvec_12__is_done__q0 && PEG_Xvec_13__is_done__q0 && PEG_Xvec_14__is_done__q0 && PEG_Xvec_15__is_done__q0 && PEG_Xvec_16__is_done__q0 && PEG_Xvec_17__is_done__q0 && PEG_Xvec_18__is_done__q0 && PEG_Xvec_19__is_done__q0 && PEG_Xvec_20__is_done__q0 && PEG_Xvec_21__is_done__q0 && PEG_Xvec_22__is_done__q0 && PEG_Xvec_23__is_done__q0 && PEG_Xvec_24__is_done__q0 && PEG_Xvec_25__is_done__q0 && PEG_Xvec_26__is_done__q0 && PEG_Xvec_27__is_done__q0 && PEG_Xvec_28__is_done__q0 && PEG_Xvec_29__is_done__q0 && PEG_Xvec_30__is_done__q0 && PEG_Xvec_31__is_done__q0 && PEG_Xvec_32__is_done__q0 && PEG_Xvec_33__is_done__q0 && PEG_Xvec_34__is_done__q0 && PEG_Xvec_35__is_done__q0 && PEG_Xvec_36__is_done__q0 && PEG_Xvec_37__is_done__q0 && PEG_Xvec_38__is_done__q0 && PEG_Xvec_39__is_done__q0 && PEG_Xvec_40__is_done__q0 && PEG_Xvec_41__is_done__q0 && PEG_Xvec_42__is_done__q0 && PEG_Xvec_43__is_done__q0 && PEG_Xvec_44__is_done__q0 && PEG_Xvec_45__is_done__q0 && PEG_Xvec_46__is_done__q0 && PEG_Xvec_47__is_done__q0 && PEG_Xvec_48__is_done__q0 && PEG_Xvec_49__is_done__q0 && PEG_Xvec_50__is_done__q0 && PEG_Xvec_51__is_done__q0 && PEG_Xvec_52__is_done__q0 && PEG_Xvec_53__is_done__q0 && PEG_Xvec_54__is_done__q0 && PEG_Xvec_55__is_done__q0 && PEG_Yvec_0__is_done__q0 && PEG_Yvec_1__is_done__q0 && PEG_Yvec_2__is_done__q0 && PEG_Yvec_3__is_done__q0 && PEG_Yvec_4__is_done__q0 && PEG_Yvec_5__is_done__q0 && PEG_Yvec_6__is_done__q0 && PEG_Yvec_7__is_done__q0 && PEG_Yvec_8__is_done__q0 && PEG_Yvec_9__is_done__q0 && PEG_Yvec_10__is_done__q0 && PEG_Yvec_11__is_done__q0 && PEG_Yvec_12__is_done__q0 && PEG_Yvec_13__is_done__q0 && PEG_Yvec_14__is_done__q0 && PEG_Yvec_15__is_done__q0 && PEG_Yvec_16__is_done__q0 && PEG_Yvec_17__is_done__q0 && PEG_Yvec_18__is_done__q0 && PEG_Yvec_19__is_done__q0 && PEG_Yvec_20__is_done__q0 && PEG_Yvec_21__is_done__q0 && PEG_Yvec_22__is_done__q0 && PEG_Yvec_23__is_done__q0 && PEG_Yvec_24__is_done__q0 && PEG_Yvec_25__is_done__q0 && PEG_Yvec_26__is_done__q0 && PEG_Yvec_27__is_done__q0 && PEG_Yvec_28__is_done__q0 && PEG_Yvec_29__is_done__q0 && PEG_Yvec_30__is_done__q0 && PEG_Yvec_31__is_done__q0 && PEG_Yvec_32__is_done__q0 && PEG_Yvec_33__is_done__q0 && PEG_Yvec_34__is_done__q0 && PEG_Yvec_35__is_done__q0 && PEG_Yvec_36__is_done__q0 && PEG_Yvec_37__is_done__q0 && PEG_Yvec_38__is_done__q0 && PEG_Yvec_39__is_done__q0 && PEG_Yvec_40__is_done__q0 && PEG_Yvec_41__is_done__q0 && PEG_Yvec_42__is_done__q0 && PEG_Yvec_43__is_done__q0 && PEG_Yvec_44__is_done__q0 && PEG_Yvec_45__is_done__q0 && PEG_Yvec_46__is_done__q0 && PEG_Yvec_47__is_done__q0 && PEG_Yvec_48__is_done__q0 && PEG_Yvec_49__is_done__q0 && PEG_Yvec_50__is_done__q0 && PEG_Yvec_51__is_done__q0 && PEG_Yvec_52__is_done__q0 && PEG_Yvec_53__is_done__q0 && PEG_Yvec_54__is_done__q0 && PEG_Yvec_55__is_done__q0 && read_A_0__is_done__q0 && read_A_1__is_done__q0 && read_A_2__is_done__q0 && read_A_3__is_done__q0 && read_A_4__is_done__q0 && read_A_5__is_done__q0 && read_A_6__is_done__q0 && read_A_7__is_done__q0 && read_A_8__is_done__q0 && read_A_9__is_done__q0 && read_A_10__is_done__q0 && read_A_11__is_done__q0 && read_A_12__is_done__q0 && read_A_13__is_done__q0 && read_A_14__is_done__q0 && read_A_15__is_done__q0 && read_A_16__is_done__q0 && read_A_17__is_done__q0 && read_A_18__is_done__q0 && read_A_19__is_done__q0 && read_A_20__is_done__q0 && read_A_21__is_done__q0 && read_A_22__is_done__q0 && read_A_23__is_done__q0 && read_A_24__is_done__q0 && read_A_25__is_done__q0 && read_A_26__is_done__q0 && read_A_27__is_done__q0 && read_A_28__is_done__q0 && read_A_29__is_done__q0 && read_A_30__is_done__q0 && read_A_31__is_done__q0 && read_A_32__is_done__q0 && read_A_33__is_done__q0 && read_A_34__is_done__q0 && read_A_35__is_done__q0 && read_A_36__is_done__q0 && read_A_37__is_done__q0 && read_A_38__is_done__q0 && read_A_39__is_done__q0 && read_A_40__is_done__q0 && read_A_41__is_done__q0 && read_A_42__is_done__q0 && read_A_43__is_done__q0 && read_A_44__is_done__q0 && read_A_45__is_done__q0 && read_A_46__is_done__q0 && read_A_47__is_done__q0 && read_A_48__is_done__q0 && read_A_49__is_done__q0 && read_A_50__is_done__q0 && read_A_51__is_done__q0 && read_A_52__is_done__q0 && read_A_53__is_done__q0 && read_A_54__is_done__q0 && read_A_55__is_done__q0 && read_X_0__is_done__q0 && read_Y_0__is_done__q0 && read_edge_list_ptr_0__is_done__q0 && write_Y_0__is_done__q0) begin
            tapa_state <= 2'b10;
          end 
        end
        2'b10: begin
          tapa_state <= 2'b00;
          countdown <= 1'd0;
        end
        2'b11: begin
          if(countdown == 1'd0) begin
            tapa_state <= 2'b00;
          end else begin
            countdown <= (countdown - 1'd1);
          end
        end
      endcase
    end
  end
  assign ap_idle = (tapa_state == 2'b00);
  assign ap_done = ap_done__q0;
  assign ap_ready = ap_done__q0;
  assign ap_start__q0 = ap_start;
  assign ap_done__q0 = (tapa_state == 2'b10);
endmodule