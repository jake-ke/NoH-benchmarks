`timescale 1 ns / 1 ps
 
(* CORE_GENERATION_INFO = "jacobi3d_kernel_jacobi3d_kernel,hls_ip_2023_2_2,{HLS_INPUT_TYPE=cxx,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=0,HLS_INPUT_PART=xcvp1802-lsvc4072-2MP-e-S,HLS_INPUT_CLOCK=3.330000,HLS_INPUT_ARCH=others,HLS_SYN_CLOCK=1.000000,HLS_SYN_LAT=0,HLS_SYN_TPT=none,HLS_SYN_MEM=0,HLS_SYN_DSP=0,HLS_SYN_FF=246,HLS_SYN_LUT=424,HLS_VERSION=2023_2_2}" *)module __rs_jacobi3d_kernel_aux #(
    parameter C_S_AXI_CONTROL_DATA_WIDTH  = 32,
    parameter C_S_AXI_CONTROL_ADDR_WIDTH  = 6,
    parameter C_S_AXI_DATA_WIDTH          = 32,
    parameter C_S_AXI_CONTROL_WSTRB_WIDTH = 4,
    parameter C_S_AXI_WSTRB_WIDTH         = 4
) (
    input wire                                           s_axi_control_AWVALID,
    output wire                                          s_axi_control_AWREADY,
    input wire  [    (C_S_AXI_CONTROL_ADDR_WIDTH - 1):0] s_axi_control_AWADDR,
    input wire                                           s_axi_control_WVALID,
    output wire                                          s_axi_control_WREADY,
    input wire  [    (C_S_AXI_CONTROL_DATA_WIDTH - 1):0] s_axi_control_WDATA,
    input wire  [   (C_S_AXI_CONTROL_WSTRB_WIDTH - 1):0] s_axi_control_WSTRB,
    input wire                                           s_axi_control_ARVALID,
    output wire                                          s_axi_control_ARREADY,
    input wire  [    (C_S_AXI_CONTROL_ADDR_WIDTH - 1):0] s_axi_control_ARADDR,
    output wire                                          s_axi_control_RVALID,
    input wire                                           s_axi_control_RREADY,
    output wire [    (C_S_AXI_CONTROL_DATA_WIDTH - 1):0] s_axi_control_RDATA,
    output wire [                                   1:0] s_axi_control_RRESP,
    output wire                                          s_axi_control_BVALID,
    input wire                                           s_axi_control_BREADY,
    output wire [                                   1:0] s_axi_control_BRESP,
    input wire                                           ap_clk,
    input wire                                           ap_rst_n,
    output wire                                          interrupt,
    output wire [                                  63:0] m_axi_bank_0_t1_ARADDR,
    output wire [                                   1:0] m_axi_bank_0_t1_ARBURST,
    output wire [                                   3:0] m_axi_bank_0_t1_ARCACHE,
    output wire [                                   0:0] m_axi_bank_0_t1_ARID,
    output wire [                                   7:0] m_axi_bank_0_t1_ARLEN,
    output wire                                          m_axi_bank_0_t1_ARLOCK,
    output wire [                                   2:0] m_axi_bank_0_t1_ARPROT,
    output wire [                                   3:0] m_axi_bank_0_t1_ARQOS,
    input wire                                           m_axi_bank_0_t1_ARREADY,
    output wire [                                   2:0] m_axi_bank_0_t1_ARSIZE,
    output wire                                          m_axi_bank_0_t1_ARVALID,
    output wire [                                  63:0] m_axi_bank_0_t1_AWADDR,
    output wire [                                   1:0] m_axi_bank_0_t1_AWBURST,
    output wire [                                   3:0] m_axi_bank_0_t1_AWCACHE,
    output wire [                                   0:0] m_axi_bank_0_t1_AWID,
    output wire [                                   7:0] m_axi_bank_0_t1_AWLEN,
    output wire                                          m_axi_bank_0_t1_AWLOCK,
    output wire [                                   2:0] m_axi_bank_0_t1_AWPROT,
    output wire [                                   3:0] m_axi_bank_0_t1_AWQOS,
    input wire                                           m_axi_bank_0_t1_AWREADY,
    output wire [                                   2:0] m_axi_bank_0_t1_AWSIZE,
    output wire                                          m_axi_bank_0_t1_AWVALID,
    input wire  [                                   0:0] m_axi_bank_0_t1_BID,
    output wire                                          m_axi_bank_0_t1_BREADY,
    input wire  [                                   1:0] m_axi_bank_0_t1_BRESP,
    input wire                                           m_axi_bank_0_t1_BVALID,
    input wire  [                                 511:0] m_axi_bank_0_t1_RDATA,
    input wire  [                                   0:0] m_axi_bank_0_t1_RID,
    input wire                                           m_axi_bank_0_t1_RLAST,
    output wire                                          m_axi_bank_0_t1_RREADY,
    input wire  [                                   1:0] m_axi_bank_0_t1_RRESP,
    input wire                                           m_axi_bank_0_t1_RVALID,
    output wire [                                 511:0] m_axi_bank_0_t1_WDATA,
    output wire                                          m_axi_bank_0_t1_WLAST,
    input wire                                           m_axi_bank_0_t1_WREADY,
    output wire [                                  63:0] m_axi_bank_0_t1_WSTRB,
    output wire                                          m_axi_bank_0_t1_WVALID,
    output wire [                                  63:0] m_axi_bank_1_t0_ARADDR,
    output wire [                                   1:0] m_axi_bank_1_t0_ARBURST,
    output wire [                                   3:0] m_axi_bank_1_t0_ARCACHE,
    output wire [                                   0:0] m_axi_bank_1_t0_ARID,
    output wire [                                   7:0] m_axi_bank_1_t0_ARLEN,
    output wire                                          m_axi_bank_1_t0_ARLOCK,
    output wire [                                   2:0] m_axi_bank_1_t0_ARPROT,
    output wire [                                   3:0] m_axi_bank_1_t0_ARQOS,
    input wire                                           m_axi_bank_1_t0_ARREADY,
    output wire [                                   2:0] m_axi_bank_1_t0_ARSIZE,
    output wire                                          m_axi_bank_1_t0_ARVALID,
    output wire [                                  63:0] m_axi_bank_1_t0_AWADDR,
    output wire [                                   1:0] m_axi_bank_1_t0_AWBURST,
    output wire [                                   3:0] m_axi_bank_1_t0_AWCACHE,
    output wire [                                   0:0] m_axi_bank_1_t0_AWID,
    output wire [                                   7:0] m_axi_bank_1_t0_AWLEN,
    output wire                                          m_axi_bank_1_t0_AWLOCK,
    output wire [                                   2:0] m_axi_bank_1_t0_AWPROT,
    output wire [                                   3:0] m_axi_bank_1_t0_AWQOS,
    input wire                                           m_axi_bank_1_t0_AWREADY,
    output wire [                                   2:0] m_axi_bank_1_t0_AWSIZE,
    output wire                                          m_axi_bank_1_t0_AWVALID,
    input wire  [                                   0:0] m_axi_bank_1_t0_BID,
    output wire                                          m_axi_bank_1_t0_BREADY,
    input wire  [                                   1:0] m_axi_bank_1_t0_BRESP,
    input wire                                           m_axi_bank_1_t0_BVALID,
    input wire  [                                 511:0] m_axi_bank_1_t0_RDATA,
    input wire  [                                   0:0] m_axi_bank_1_t0_RID,
    input wire                                           m_axi_bank_1_t0_RLAST,
    output wire                                          m_axi_bank_1_t0_RREADY,
    input wire  [                                   1:0] m_axi_bank_1_t0_RRESP,
    input wire                                           m_axi_bank_1_t0_RVALID,
    output wire [                                 511:0] m_axi_bank_1_t0_WDATA,
    output wire                                          m_axi_bank_1_t0_WLAST,
    input wire                                           m_axi_bank_1_t0_WREADY,
    output wire [                                  63:0] m_axi_bank_1_t0_WSTRB,
    output wire                                          m_axi_bank_1_t0_WVALID,
    output wire                                          control_s_axi_U_ACLK,
    output wire                                          control_s_axi_U_ACLK_EN,
    output wire [    (C_S_AXI_CONTROL_ADDR_WIDTH - 1):0] control_s_axi_U_ARADDR,
    output wire                                          control_s_axi_U_ARESET,
    input wire                                           control_s_axi_U_ARREADY,
    output wire                                          control_s_axi_U_ARVALID,
    output wire [    (C_S_AXI_CONTROL_ADDR_WIDTH - 1):0] control_s_axi_U_AWADDR,
    input wire                                           control_s_axi_U_AWREADY,
    output wire                                          control_s_axi_U_AWVALID,
    output wire                                          control_s_axi_U_BREADY,
    input wire  [                                   1:0] control_s_axi_U_BRESP,
    input wire                                           control_s_axi_U_BVALID,
    input wire  [    (C_S_AXI_CONTROL_DATA_WIDTH - 1):0] control_s_axi_U_RDATA,
    output wire                                          control_s_axi_U_RREADY,
    input wire  [                                   1:0] control_s_axi_U_RRESP,
    input wire                                           control_s_axi_U_RVALID,
    output wire [    (C_S_AXI_CONTROL_DATA_WIDTH - 1):0] control_s_axi_U_WDATA,
    input wire                                           control_s_axi_U_WREADY,
    output wire [(C_S_AXI_CONTROL_DATA_WIDTH / 8 - 1):0] control_s_axi_U_WSTRB,
    output wire                                          control_s_axi_U_WVALID,
    output wire                                          control_s_axi_U_ap_done,
    output wire                                          control_s_axi_U_ap_idle,
    output wire                                          control_s_axi_U_ap_ready,
    input wire                                           control_s_axi_U_ap_start,
    input wire  [                                  63:0] control_s_axi_U_bank_0_t1,
    input wire  [                                  63:0] control_s_axi_U_bank_1_t0,
    input wire  [                                  63:0] control_s_axi_U_coalesced_data_num,
    input wire                                           control_s_axi_U_interrupt,
    output wire                                          bank_0_t1_buf_clk,
    output wire [                                 512:0] bank_0_t1_buf_if_din,
    input wire  [                                 512:0] bank_0_t1_buf_if_dout,
    input wire                                           bank_0_t1_buf_if_empty_n,
    input wire                                           bank_0_t1_buf_if_full_n,
    output wire                                          bank_0_t1_buf_if_read,
    output wire                                          bank_0_t1_buf_if_read_ce,
    output wire                                          bank_0_t1_buf_if_write,
    output wire                                          bank_0_t1_buf_if_write_ce,
    output wire                                          bank_0_t1_buf_reset,
    output wire                                          bank_1_t0_buf_clk,
    output wire [                                 512:0] bank_1_t0_buf_if_din,
    input wire  [                                 512:0] bank_1_t0_buf_if_dout,
    input wire                                           bank_1_t0_buf_if_empty_n,
    input wire                                           bank_1_t0_buf_if_full_n,
    output wire                                          bank_1_t0_buf_if_read,
    output wire                                          bank_1_t0_buf_if_read_ce,
    output wire                                          bank_1_t0_buf_if_write,
    output wire                                          bank_1_t0_buf_if_write_ce,
    output wire                                          bank_1_t0_buf_reset,
    output wire                                          from_t0_to_t0_bank_1_clk,
    output wire [                                 512:0] from_t0_to_t0_bank_1_if_din,
    input wire  [                                 512:0] from_t0_to_t0_bank_1_if_dout,
    input wire                                           from_t0_to_t0_bank_1_if_empty_n,
    input wire                                           from_t0_to_t0_bank_1_if_full_n,
    output wire                                          from_t0_to_t0_bank_1_if_read,
    output wire                                          from_t0_to_t0_bank_1_if_read_ce,
    output wire                                          from_t0_to_t0_bank_1_if_write,
    output wire                                          from_t0_to_t0_bank_1_if_write_ce,
    output wire                                          from_t0_to_t0_bank_1_reset,
    output wire                                          from_t1_bank_0_to_t1_iter1_clk,
    output wire [                                 512:0] from_t1_bank_0_to_t1_iter1_if_din,
    input wire  [                                 512:0] from_t1_bank_0_to_t1_iter1_if_dout,
    input wire                                           from_t1_bank_0_to_t1_iter1_if_empty_n,
    input wire                                           from_t1_bank_0_to_t1_iter1_if_full_n,
    output wire                                          from_t1_bank_0_to_t1_iter1_if_read,
    output wire                                          from_t1_bank_0_to_t1_iter1_if_read_ce,
    output wire                                          from_t1_bank_0_to_t1_iter1_if_write,
    output wire                                          from_t1_bank_0_to_t1_iter1_if_write_ce,
    output wire                                          from_t1_bank_0_to_t1_iter1_reset,
    output wire                                          from_t1_iter100_to_t1_iter101_clk,
    output wire [                                 512:0] from_t1_iter100_to_t1_iter101_if_din,
    input wire  [                                 512:0] from_t1_iter100_to_t1_iter101_if_dout,
    input wire                                           from_t1_iter100_to_t1_iter101_if_empty_n,
    input wire                                           from_t1_iter100_to_t1_iter101_if_full_n,
    output wire                                          from_t1_iter100_to_t1_iter101_if_read,
    output wire                                          from_t1_iter100_to_t1_iter101_if_read_ce,
    output wire                                          from_t1_iter100_to_t1_iter101_if_write,
    output wire                                          from_t1_iter100_to_t1_iter101_if_write_ce,
    output wire                                          from_t1_iter100_to_t1_iter101_reset,
    output wire                                          from_t1_iter101_to_t1_iter102_clk,
    output wire [                                 512:0] from_t1_iter101_to_t1_iter102_if_din,
    input wire  [                                 512:0] from_t1_iter101_to_t1_iter102_if_dout,
    input wire                                           from_t1_iter101_to_t1_iter102_if_empty_n,
    input wire                                           from_t1_iter101_to_t1_iter102_if_full_n,
    output wire                                          from_t1_iter101_to_t1_iter102_if_read,
    output wire                                          from_t1_iter101_to_t1_iter102_if_read_ce,
    output wire                                          from_t1_iter101_to_t1_iter102_if_write,
    output wire                                          from_t1_iter101_to_t1_iter102_if_write_ce,
    output wire                                          from_t1_iter101_to_t1_iter102_reset,
    output wire                                          from_t1_iter102_to_t1_iter103_clk,
    output wire [                                 512:0] from_t1_iter102_to_t1_iter103_if_din,
    input wire  [                                 512:0] from_t1_iter102_to_t1_iter103_if_dout,
    input wire                                           from_t1_iter102_to_t1_iter103_if_empty_n,
    input wire                                           from_t1_iter102_to_t1_iter103_if_full_n,
    output wire                                          from_t1_iter102_to_t1_iter103_if_read,
    output wire                                          from_t1_iter102_to_t1_iter103_if_read_ce,
    output wire                                          from_t1_iter102_to_t1_iter103_if_write,
    output wire                                          from_t1_iter102_to_t1_iter103_if_write_ce,
    output wire                                          from_t1_iter102_to_t1_iter103_reset,
    output wire                                          from_t1_iter103_to_t1_iter104_clk,
    output wire [                                 512:0] from_t1_iter103_to_t1_iter104_if_din,
    input wire  [                                 512:0] from_t1_iter103_to_t1_iter104_if_dout,
    input wire                                           from_t1_iter103_to_t1_iter104_if_empty_n,
    input wire                                           from_t1_iter103_to_t1_iter104_if_full_n,
    output wire                                          from_t1_iter103_to_t1_iter104_if_read,
    output wire                                          from_t1_iter103_to_t1_iter104_if_read_ce,
    output wire                                          from_t1_iter103_to_t1_iter104_if_write,
    output wire                                          from_t1_iter103_to_t1_iter104_if_write_ce,
    output wire                                          from_t1_iter103_to_t1_iter104_reset,
    output wire                                          from_t1_iter104_to_t1_iter105_clk,
    output wire [                                 512:0] from_t1_iter104_to_t1_iter105_if_din,
    input wire  [                                 512:0] from_t1_iter104_to_t1_iter105_if_dout,
    input wire                                           from_t1_iter104_to_t1_iter105_if_empty_n,
    input wire                                           from_t1_iter104_to_t1_iter105_if_full_n,
    output wire                                          from_t1_iter104_to_t1_iter105_if_read,
    output wire                                          from_t1_iter104_to_t1_iter105_if_read_ce,
    output wire                                          from_t1_iter104_to_t1_iter105_if_write,
    output wire                                          from_t1_iter104_to_t1_iter105_if_write_ce,
    output wire                                          from_t1_iter104_to_t1_iter105_reset,
    output wire                                          from_t1_iter105_to_t1_iter106_clk,
    output wire [                                 512:0] from_t1_iter105_to_t1_iter106_if_din,
    input wire  [                                 512:0] from_t1_iter105_to_t1_iter106_if_dout,
    input wire                                           from_t1_iter105_to_t1_iter106_if_empty_n,
    input wire                                           from_t1_iter105_to_t1_iter106_if_full_n,
    output wire                                          from_t1_iter105_to_t1_iter106_if_read,
    output wire                                          from_t1_iter105_to_t1_iter106_if_read_ce,
    output wire                                          from_t1_iter105_to_t1_iter106_if_write,
    output wire                                          from_t1_iter105_to_t1_iter106_if_write_ce,
    output wire                                          from_t1_iter105_to_t1_iter106_reset,
    output wire                                          from_t1_iter106_to_t1_iter107_clk,
    output wire [                                 512:0] from_t1_iter106_to_t1_iter107_if_din,
    input wire  [                                 512:0] from_t1_iter106_to_t1_iter107_if_dout,
    input wire                                           from_t1_iter106_to_t1_iter107_if_empty_n,
    input wire                                           from_t1_iter106_to_t1_iter107_if_full_n,
    output wire                                          from_t1_iter106_to_t1_iter107_if_read,
    output wire                                          from_t1_iter106_to_t1_iter107_if_read_ce,
    output wire                                          from_t1_iter106_to_t1_iter107_if_write,
    output wire                                          from_t1_iter106_to_t1_iter107_if_write_ce,
    output wire                                          from_t1_iter106_to_t1_iter107_reset,
    output wire                                          from_t1_iter107_to_t1_iter108_clk,
    output wire [                                 512:0] from_t1_iter107_to_t1_iter108_if_din,
    input wire  [                                 512:0] from_t1_iter107_to_t1_iter108_if_dout,
    input wire                                           from_t1_iter107_to_t1_iter108_if_empty_n,
    input wire                                           from_t1_iter107_to_t1_iter108_if_full_n,
    output wire                                          from_t1_iter107_to_t1_iter108_if_read,
    output wire                                          from_t1_iter107_to_t1_iter108_if_read_ce,
    output wire                                          from_t1_iter107_to_t1_iter108_if_write,
    output wire                                          from_t1_iter107_to_t1_iter108_if_write_ce,
    output wire                                          from_t1_iter107_to_t1_iter108_reset,
    output wire                                          from_t1_iter108_to_t0_clk,
    output wire [                                 512:0] from_t1_iter108_to_t0_if_din,
    input wire  [                                 512:0] from_t1_iter108_to_t0_if_dout,
    input wire                                           from_t1_iter108_to_t0_if_empty_n,
    input wire                                           from_t1_iter108_to_t0_if_full_n,
    output wire                                          from_t1_iter108_to_t0_if_read,
    output wire                                          from_t1_iter108_to_t0_if_read_ce,
    output wire                                          from_t1_iter108_to_t0_if_write,
    output wire                                          from_t1_iter108_to_t0_if_write_ce,
    output wire                                          from_t1_iter108_to_t0_reset,
    output wire                                          from_t1_iter10_to_t1_iter11_clk,
    output wire [                                 512:0] from_t1_iter10_to_t1_iter11_if_din,
    input wire  [                                 512:0] from_t1_iter10_to_t1_iter11_if_dout,
    input wire                                           from_t1_iter10_to_t1_iter11_if_empty_n,
    input wire                                           from_t1_iter10_to_t1_iter11_if_full_n,
    output wire                                          from_t1_iter10_to_t1_iter11_if_read,
    output wire                                          from_t1_iter10_to_t1_iter11_if_read_ce,
    output wire                                          from_t1_iter10_to_t1_iter11_if_write,
    output wire                                          from_t1_iter10_to_t1_iter11_if_write_ce,
    output wire                                          from_t1_iter10_to_t1_iter11_reset,
    output wire                                          from_t1_iter11_to_t1_iter12_clk,
    output wire [                                 512:0] from_t1_iter11_to_t1_iter12_if_din,
    input wire  [                                 512:0] from_t1_iter11_to_t1_iter12_if_dout,
    input wire                                           from_t1_iter11_to_t1_iter12_if_empty_n,
    input wire                                           from_t1_iter11_to_t1_iter12_if_full_n,
    output wire                                          from_t1_iter11_to_t1_iter12_if_read,
    output wire                                          from_t1_iter11_to_t1_iter12_if_read_ce,
    output wire                                          from_t1_iter11_to_t1_iter12_if_write,
    output wire                                          from_t1_iter11_to_t1_iter12_if_write_ce,
    output wire                                          from_t1_iter11_to_t1_iter12_reset,
    output wire                                          from_t1_iter12_to_t1_iter13_clk,
    output wire [                                 512:0] from_t1_iter12_to_t1_iter13_if_din,
    input wire  [                                 512:0] from_t1_iter12_to_t1_iter13_if_dout,
    input wire                                           from_t1_iter12_to_t1_iter13_if_empty_n,
    input wire                                           from_t1_iter12_to_t1_iter13_if_full_n,
    output wire                                          from_t1_iter12_to_t1_iter13_if_read,
    output wire                                          from_t1_iter12_to_t1_iter13_if_read_ce,
    output wire                                          from_t1_iter12_to_t1_iter13_if_write,
    output wire                                          from_t1_iter12_to_t1_iter13_if_write_ce,
    output wire                                          from_t1_iter12_to_t1_iter13_reset,
    output wire                                          from_t1_iter13_to_t1_iter14_clk,
    output wire [                                 512:0] from_t1_iter13_to_t1_iter14_if_din,
    input wire  [                                 512:0] from_t1_iter13_to_t1_iter14_if_dout,
    input wire                                           from_t1_iter13_to_t1_iter14_if_empty_n,
    input wire                                           from_t1_iter13_to_t1_iter14_if_full_n,
    output wire                                          from_t1_iter13_to_t1_iter14_if_read,
    output wire                                          from_t1_iter13_to_t1_iter14_if_read_ce,
    output wire                                          from_t1_iter13_to_t1_iter14_if_write,
    output wire                                          from_t1_iter13_to_t1_iter14_if_write_ce,
    output wire                                          from_t1_iter13_to_t1_iter14_reset,
    output wire                                          from_t1_iter14_to_t1_iter15_clk,
    output wire [                                 512:0] from_t1_iter14_to_t1_iter15_if_din,
    input wire  [                                 512:0] from_t1_iter14_to_t1_iter15_if_dout,
    input wire                                           from_t1_iter14_to_t1_iter15_if_empty_n,
    input wire                                           from_t1_iter14_to_t1_iter15_if_full_n,
    output wire                                          from_t1_iter14_to_t1_iter15_if_read,
    output wire                                          from_t1_iter14_to_t1_iter15_if_read_ce,
    output wire                                          from_t1_iter14_to_t1_iter15_if_write,
    output wire                                          from_t1_iter14_to_t1_iter15_if_write_ce,
    output wire                                          from_t1_iter14_to_t1_iter15_reset,
    output wire                                          from_t1_iter15_to_t1_iter16_clk,
    output wire [                                 512:0] from_t1_iter15_to_t1_iter16_if_din,
    input wire  [                                 512:0] from_t1_iter15_to_t1_iter16_if_dout,
    input wire                                           from_t1_iter15_to_t1_iter16_if_empty_n,
    input wire                                           from_t1_iter15_to_t1_iter16_if_full_n,
    output wire                                          from_t1_iter15_to_t1_iter16_if_read,
    output wire                                          from_t1_iter15_to_t1_iter16_if_read_ce,
    output wire                                          from_t1_iter15_to_t1_iter16_if_write,
    output wire                                          from_t1_iter15_to_t1_iter16_if_write_ce,
    output wire                                          from_t1_iter15_to_t1_iter16_reset,
    output wire                                          from_t1_iter16_to_t1_iter17_clk,
    output wire [                                 512:0] from_t1_iter16_to_t1_iter17_if_din,
    input wire  [                                 512:0] from_t1_iter16_to_t1_iter17_if_dout,
    input wire                                           from_t1_iter16_to_t1_iter17_if_empty_n,
    input wire                                           from_t1_iter16_to_t1_iter17_if_full_n,
    output wire                                          from_t1_iter16_to_t1_iter17_if_read,
    output wire                                          from_t1_iter16_to_t1_iter17_if_read_ce,
    output wire                                          from_t1_iter16_to_t1_iter17_if_write,
    output wire                                          from_t1_iter16_to_t1_iter17_if_write_ce,
    output wire                                          from_t1_iter16_to_t1_iter17_reset,
    output wire                                          from_t1_iter17_to_t1_iter18_clk,
    output wire [                                 512:0] from_t1_iter17_to_t1_iter18_if_din,
    input wire  [                                 512:0] from_t1_iter17_to_t1_iter18_if_dout,
    input wire                                           from_t1_iter17_to_t1_iter18_if_empty_n,
    input wire                                           from_t1_iter17_to_t1_iter18_if_full_n,
    output wire                                          from_t1_iter17_to_t1_iter18_if_read,
    output wire                                          from_t1_iter17_to_t1_iter18_if_read_ce,
    output wire                                          from_t1_iter17_to_t1_iter18_if_write,
    output wire                                          from_t1_iter17_to_t1_iter18_if_write_ce,
    output wire                                          from_t1_iter17_to_t1_iter18_reset,
    output wire                                          from_t1_iter18_to_t1_iter19_clk,
    output wire [                                 512:0] from_t1_iter18_to_t1_iter19_if_din,
    input wire  [                                 512:0] from_t1_iter18_to_t1_iter19_if_dout,
    input wire                                           from_t1_iter18_to_t1_iter19_if_empty_n,
    input wire                                           from_t1_iter18_to_t1_iter19_if_full_n,
    output wire                                          from_t1_iter18_to_t1_iter19_if_read,
    output wire                                          from_t1_iter18_to_t1_iter19_if_read_ce,
    output wire                                          from_t1_iter18_to_t1_iter19_if_write,
    output wire                                          from_t1_iter18_to_t1_iter19_if_write_ce,
    output wire                                          from_t1_iter18_to_t1_iter19_reset,
    output wire                                          from_t1_iter19_to_t1_iter20_clk,
    output wire [                                 512:0] from_t1_iter19_to_t1_iter20_if_din,
    input wire  [                                 512:0] from_t1_iter19_to_t1_iter20_if_dout,
    input wire                                           from_t1_iter19_to_t1_iter20_if_empty_n,
    input wire                                           from_t1_iter19_to_t1_iter20_if_full_n,
    output wire                                          from_t1_iter19_to_t1_iter20_if_read,
    output wire                                          from_t1_iter19_to_t1_iter20_if_read_ce,
    output wire                                          from_t1_iter19_to_t1_iter20_if_write,
    output wire                                          from_t1_iter19_to_t1_iter20_if_write_ce,
    output wire                                          from_t1_iter19_to_t1_iter20_reset,
    output wire                                          from_t1_iter1_to_t1_iter2_clk,
    output wire [                                 512:0] from_t1_iter1_to_t1_iter2_if_din,
    input wire  [                                 512:0] from_t1_iter1_to_t1_iter2_if_dout,
    input wire                                           from_t1_iter1_to_t1_iter2_if_empty_n,
    input wire                                           from_t1_iter1_to_t1_iter2_if_full_n,
    output wire                                          from_t1_iter1_to_t1_iter2_if_read,
    output wire                                          from_t1_iter1_to_t1_iter2_if_read_ce,
    output wire                                          from_t1_iter1_to_t1_iter2_if_write,
    output wire                                          from_t1_iter1_to_t1_iter2_if_write_ce,
    output wire                                          from_t1_iter1_to_t1_iter2_reset,
    output wire                                          from_t1_iter20_to_t1_iter21_clk,
    output wire [                                 512:0] from_t1_iter20_to_t1_iter21_if_din,
    input wire  [                                 512:0] from_t1_iter20_to_t1_iter21_if_dout,
    input wire                                           from_t1_iter20_to_t1_iter21_if_empty_n,
    input wire                                           from_t1_iter20_to_t1_iter21_if_full_n,
    output wire                                          from_t1_iter20_to_t1_iter21_if_read,
    output wire                                          from_t1_iter20_to_t1_iter21_if_read_ce,
    output wire                                          from_t1_iter20_to_t1_iter21_if_write,
    output wire                                          from_t1_iter20_to_t1_iter21_if_write_ce,
    output wire                                          from_t1_iter20_to_t1_iter21_reset,
    output wire                                          from_t1_iter21_to_t1_iter22_clk,
    output wire [                                 512:0] from_t1_iter21_to_t1_iter22_if_din,
    input wire  [                                 512:0] from_t1_iter21_to_t1_iter22_if_dout,
    input wire                                           from_t1_iter21_to_t1_iter22_if_empty_n,
    input wire                                           from_t1_iter21_to_t1_iter22_if_full_n,
    output wire                                          from_t1_iter21_to_t1_iter22_if_read,
    output wire                                          from_t1_iter21_to_t1_iter22_if_read_ce,
    output wire                                          from_t1_iter21_to_t1_iter22_if_write,
    output wire                                          from_t1_iter21_to_t1_iter22_if_write_ce,
    output wire                                          from_t1_iter21_to_t1_iter22_reset,
    output wire                                          from_t1_iter22_to_t1_iter23_clk,
    output wire [                                 512:0] from_t1_iter22_to_t1_iter23_if_din,
    input wire  [                                 512:0] from_t1_iter22_to_t1_iter23_if_dout,
    input wire                                           from_t1_iter22_to_t1_iter23_if_empty_n,
    input wire                                           from_t1_iter22_to_t1_iter23_if_full_n,
    output wire                                          from_t1_iter22_to_t1_iter23_if_read,
    output wire                                          from_t1_iter22_to_t1_iter23_if_read_ce,
    output wire                                          from_t1_iter22_to_t1_iter23_if_write,
    output wire                                          from_t1_iter22_to_t1_iter23_if_write_ce,
    output wire                                          from_t1_iter22_to_t1_iter23_reset,
    output wire                                          from_t1_iter23_to_t1_iter24_clk,
    output wire [                                 512:0] from_t1_iter23_to_t1_iter24_if_din,
    input wire  [                                 512:0] from_t1_iter23_to_t1_iter24_if_dout,
    input wire                                           from_t1_iter23_to_t1_iter24_if_empty_n,
    input wire                                           from_t1_iter23_to_t1_iter24_if_full_n,
    output wire                                          from_t1_iter23_to_t1_iter24_if_read,
    output wire                                          from_t1_iter23_to_t1_iter24_if_read_ce,
    output wire                                          from_t1_iter23_to_t1_iter24_if_write,
    output wire                                          from_t1_iter23_to_t1_iter24_if_write_ce,
    output wire                                          from_t1_iter23_to_t1_iter24_reset,
    output wire                                          from_t1_iter24_to_t1_iter25_clk,
    output wire [                                 512:0] from_t1_iter24_to_t1_iter25_if_din,
    input wire  [                                 512:0] from_t1_iter24_to_t1_iter25_if_dout,
    input wire                                           from_t1_iter24_to_t1_iter25_if_empty_n,
    input wire                                           from_t1_iter24_to_t1_iter25_if_full_n,
    output wire                                          from_t1_iter24_to_t1_iter25_if_read,
    output wire                                          from_t1_iter24_to_t1_iter25_if_read_ce,
    output wire                                          from_t1_iter24_to_t1_iter25_if_write,
    output wire                                          from_t1_iter24_to_t1_iter25_if_write_ce,
    output wire                                          from_t1_iter24_to_t1_iter25_reset,
    output wire                                          from_t1_iter25_to_t1_iter26_clk,
    output wire [                                 512:0] from_t1_iter25_to_t1_iter26_if_din,
    input wire  [                                 512:0] from_t1_iter25_to_t1_iter26_if_dout,
    input wire                                           from_t1_iter25_to_t1_iter26_if_empty_n,
    input wire                                           from_t1_iter25_to_t1_iter26_if_full_n,
    output wire                                          from_t1_iter25_to_t1_iter26_if_read,
    output wire                                          from_t1_iter25_to_t1_iter26_if_read_ce,
    output wire                                          from_t1_iter25_to_t1_iter26_if_write,
    output wire                                          from_t1_iter25_to_t1_iter26_if_write_ce,
    output wire                                          from_t1_iter25_to_t1_iter26_reset,
    output wire                                          from_t1_iter26_to_t1_iter27_clk,
    output wire [                                 512:0] from_t1_iter26_to_t1_iter27_if_din,
    input wire  [                                 512:0] from_t1_iter26_to_t1_iter27_if_dout,
    input wire                                           from_t1_iter26_to_t1_iter27_if_empty_n,
    input wire                                           from_t1_iter26_to_t1_iter27_if_full_n,
    output wire                                          from_t1_iter26_to_t1_iter27_if_read,
    output wire                                          from_t1_iter26_to_t1_iter27_if_read_ce,
    output wire                                          from_t1_iter26_to_t1_iter27_if_write,
    output wire                                          from_t1_iter26_to_t1_iter27_if_write_ce,
    output wire                                          from_t1_iter26_to_t1_iter27_reset,
    output wire                                          from_t1_iter27_to_t1_iter28_clk,
    output wire [                                 512:0] from_t1_iter27_to_t1_iter28_if_din,
    input wire  [                                 512:0] from_t1_iter27_to_t1_iter28_if_dout,
    input wire                                           from_t1_iter27_to_t1_iter28_if_empty_n,
    input wire                                           from_t1_iter27_to_t1_iter28_if_full_n,
    output wire                                          from_t1_iter27_to_t1_iter28_if_read,
    output wire                                          from_t1_iter27_to_t1_iter28_if_read_ce,
    output wire                                          from_t1_iter27_to_t1_iter28_if_write,
    output wire                                          from_t1_iter27_to_t1_iter28_if_write_ce,
    output wire                                          from_t1_iter27_to_t1_iter28_reset,
    output wire                                          from_t1_iter28_to_t1_iter29_clk,
    output wire [                                 512:0] from_t1_iter28_to_t1_iter29_if_din,
    input wire  [                                 512:0] from_t1_iter28_to_t1_iter29_if_dout,
    input wire                                           from_t1_iter28_to_t1_iter29_if_empty_n,
    input wire                                           from_t1_iter28_to_t1_iter29_if_full_n,
    output wire                                          from_t1_iter28_to_t1_iter29_if_read,
    output wire                                          from_t1_iter28_to_t1_iter29_if_read_ce,
    output wire                                          from_t1_iter28_to_t1_iter29_if_write,
    output wire                                          from_t1_iter28_to_t1_iter29_if_write_ce,
    output wire                                          from_t1_iter28_to_t1_iter29_reset,
    output wire                                          from_t1_iter29_to_t1_iter30_clk,
    output wire [                                 512:0] from_t1_iter29_to_t1_iter30_if_din,
    input wire  [                                 512:0] from_t1_iter29_to_t1_iter30_if_dout,
    input wire                                           from_t1_iter29_to_t1_iter30_if_empty_n,
    input wire                                           from_t1_iter29_to_t1_iter30_if_full_n,
    output wire                                          from_t1_iter29_to_t1_iter30_if_read,
    output wire                                          from_t1_iter29_to_t1_iter30_if_read_ce,
    output wire                                          from_t1_iter29_to_t1_iter30_if_write,
    output wire                                          from_t1_iter29_to_t1_iter30_if_write_ce,
    output wire                                          from_t1_iter29_to_t1_iter30_reset,
    output wire                                          from_t1_iter2_to_t1_iter3_clk,
    output wire [                                 512:0] from_t1_iter2_to_t1_iter3_if_din,
    input wire  [                                 512:0] from_t1_iter2_to_t1_iter3_if_dout,
    input wire                                           from_t1_iter2_to_t1_iter3_if_empty_n,
    input wire                                           from_t1_iter2_to_t1_iter3_if_full_n,
    output wire                                          from_t1_iter2_to_t1_iter3_if_read,
    output wire                                          from_t1_iter2_to_t1_iter3_if_read_ce,
    output wire                                          from_t1_iter2_to_t1_iter3_if_write,
    output wire                                          from_t1_iter2_to_t1_iter3_if_write_ce,
    output wire                                          from_t1_iter2_to_t1_iter3_reset,
    output wire                                          from_t1_iter30_to_t1_iter31_clk,
    output wire [                                 512:0] from_t1_iter30_to_t1_iter31_if_din,
    input wire  [                                 512:0] from_t1_iter30_to_t1_iter31_if_dout,
    input wire                                           from_t1_iter30_to_t1_iter31_if_empty_n,
    input wire                                           from_t1_iter30_to_t1_iter31_if_full_n,
    output wire                                          from_t1_iter30_to_t1_iter31_if_read,
    output wire                                          from_t1_iter30_to_t1_iter31_if_read_ce,
    output wire                                          from_t1_iter30_to_t1_iter31_if_write,
    output wire                                          from_t1_iter30_to_t1_iter31_if_write_ce,
    output wire                                          from_t1_iter30_to_t1_iter31_reset,
    output wire                                          from_t1_iter31_to_t1_iter32_clk,
    output wire [                                 512:0] from_t1_iter31_to_t1_iter32_if_din,
    input wire  [                                 512:0] from_t1_iter31_to_t1_iter32_if_dout,
    input wire                                           from_t1_iter31_to_t1_iter32_if_empty_n,
    input wire                                           from_t1_iter31_to_t1_iter32_if_full_n,
    output wire                                          from_t1_iter31_to_t1_iter32_if_read,
    output wire                                          from_t1_iter31_to_t1_iter32_if_read_ce,
    output wire                                          from_t1_iter31_to_t1_iter32_if_write,
    output wire                                          from_t1_iter31_to_t1_iter32_if_write_ce,
    output wire                                          from_t1_iter31_to_t1_iter32_reset,
    output wire                                          from_t1_iter32_to_t1_iter33_clk,
    output wire [                                 512:0] from_t1_iter32_to_t1_iter33_if_din,
    input wire  [                                 512:0] from_t1_iter32_to_t1_iter33_if_dout,
    input wire                                           from_t1_iter32_to_t1_iter33_if_empty_n,
    input wire                                           from_t1_iter32_to_t1_iter33_if_full_n,
    output wire                                          from_t1_iter32_to_t1_iter33_if_read,
    output wire                                          from_t1_iter32_to_t1_iter33_if_read_ce,
    output wire                                          from_t1_iter32_to_t1_iter33_if_write,
    output wire                                          from_t1_iter32_to_t1_iter33_if_write_ce,
    output wire                                          from_t1_iter32_to_t1_iter33_reset,
    output wire                                          from_t1_iter33_to_t1_iter34_clk,
    output wire [                                 512:0] from_t1_iter33_to_t1_iter34_if_din,
    input wire  [                                 512:0] from_t1_iter33_to_t1_iter34_if_dout,
    input wire                                           from_t1_iter33_to_t1_iter34_if_empty_n,
    input wire                                           from_t1_iter33_to_t1_iter34_if_full_n,
    output wire                                          from_t1_iter33_to_t1_iter34_if_read,
    output wire                                          from_t1_iter33_to_t1_iter34_if_read_ce,
    output wire                                          from_t1_iter33_to_t1_iter34_if_write,
    output wire                                          from_t1_iter33_to_t1_iter34_if_write_ce,
    output wire                                          from_t1_iter33_to_t1_iter34_reset,
    output wire                                          from_t1_iter34_to_t1_iter35_clk,
    output wire [                                 512:0] from_t1_iter34_to_t1_iter35_if_din,
    input wire  [                                 512:0] from_t1_iter34_to_t1_iter35_if_dout,
    input wire                                           from_t1_iter34_to_t1_iter35_if_empty_n,
    input wire                                           from_t1_iter34_to_t1_iter35_if_full_n,
    output wire                                          from_t1_iter34_to_t1_iter35_if_read,
    output wire                                          from_t1_iter34_to_t1_iter35_if_read_ce,
    output wire                                          from_t1_iter34_to_t1_iter35_if_write,
    output wire                                          from_t1_iter34_to_t1_iter35_if_write_ce,
    output wire                                          from_t1_iter34_to_t1_iter35_reset,
    output wire                                          from_t1_iter35_to_t1_iter36_clk,
    output wire [                                 512:0] from_t1_iter35_to_t1_iter36_if_din,
    input wire  [                                 512:0] from_t1_iter35_to_t1_iter36_if_dout,
    input wire                                           from_t1_iter35_to_t1_iter36_if_empty_n,
    input wire                                           from_t1_iter35_to_t1_iter36_if_full_n,
    output wire                                          from_t1_iter35_to_t1_iter36_if_read,
    output wire                                          from_t1_iter35_to_t1_iter36_if_read_ce,
    output wire                                          from_t1_iter35_to_t1_iter36_if_write,
    output wire                                          from_t1_iter35_to_t1_iter36_if_write_ce,
    output wire                                          from_t1_iter35_to_t1_iter36_reset,
    output wire                                          from_t1_iter36_to_t1_iter37_clk,
    output wire [                                 512:0] from_t1_iter36_to_t1_iter37_if_din,
    input wire  [                                 512:0] from_t1_iter36_to_t1_iter37_if_dout,
    input wire                                           from_t1_iter36_to_t1_iter37_if_empty_n,
    input wire                                           from_t1_iter36_to_t1_iter37_if_full_n,
    output wire                                          from_t1_iter36_to_t1_iter37_if_read,
    output wire                                          from_t1_iter36_to_t1_iter37_if_read_ce,
    output wire                                          from_t1_iter36_to_t1_iter37_if_write,
    output wire                                          from_t1_iter36_to_t1_iter37_if_write_ce,
    output wire                                          from_t1_iter36_to_t1_iter37_reset,
    output wire                                          from_t1_iter37_to_t1_iter38_clk,
    output wire [                                 512:0] from_t1_iter37_to_t1_iter38_if_din,
    input wire  [                                 512:0] from_t1_iter37_to_t1_iter38_if_dout,
    input wire                                           from_t1_iter37_to_t1_iter38_if_empty_n,
    input wire                                           from_t1_iter37_to_t1_iter38_if_full_n,
    output wire                                          from_t1_iter37_to_t1_iter38_if_read,
    output wire                                          from_t1_iter37_to_t1_iter38_if_read_ce,
    output wire                                          from_t1_iter37_to_t1_iter38_if_write,
    output wire                                          from_t1_iter37_to_t1_iter38_if_write_ce,
    output wire                                          from_t1_iter37_to_t1_iter38_reset,
    output wire                                          from_t1_iter38_to_t1_iter39_clk,
    output wire [                                 512:0] from_t1_iter38_to_t1_iter39_if_din,
    input wire  [                                 512:0] from_t1_iter38_to_t1_iter39_if_dout,
    input wire                                           from_t1_iter38_to_t1_iter39_if_empty_n,
    input wire                                           from_t1_iter38_to_t1_iter39_if_full_n,
    output wire                                          from_t1_iter38_to_t1_iter39_if_read,
    output wire                                          from_t1_iter38_to_t1_iter39_if_read_ce,
    output wire                                          from_t1_iter38_to_t1_iter39_if_write,
    output wire                                          from_t1_iter38_to_t1_iter39_if_write_ce,
    output wire                                          from_t1_iter38_to_t1_iter39_reset,
    output wire                                          from_t1_iter39_to_t1_iter40_clk,
    output wire [                                 512:0] from_t1_iter39_to_t1_iter40_if_din,
    input wire  [                                 512:0] from_t1_iter39_to_t1_iter40_if_dout,
    input wire                                           from_t1_iter39_to_t1_iter40_if_empty_n,
    input wire                                           from_t1_iter39_to_t1_iter40_if_full_n,
    output wire                                          from_t1_iter39_to_t1_iter40_if_read,
    output wire                                          from_t1_iter39_to_t1_iter40_if_read_ce,
    output wire                                          from_t1_iter39_to_t1_iter40_if_write,
    output wire                                          from_t1_iter39_to_t1_iter40_if_write_ce,
    output wire                                          from_t1_iter39_to_t1_iter40_reset,
    output wire                                          from_t1_iter3_to_t1_iter4_clk,
    output wire [                                 512:0] from_t1_iter3_to_t1_iter4_if_din,
    input wire  [                                 512:0] from_t1_iter3_to_t1_iter4_if_dout,
    input wire                                           from_t1_iter3_to_t1_iter4_if_empty_n,
    input wire                                           from_t1_iter3_to_t1_iter4_if_full_n,
    output wire                                          from_t1_iter3_to_t1_iter4_if_read,
    output wire                                          from_t1_iter3_to_t1_iter4_if_read_ce,
    output wire                                          from_t1_iter3_to_t1_iter4_if_write,
    output wire                                          from_t1_iter3_to_t1_iter4_if_write_ce,
    output wire                                          from_t1_iter3_to_t1_iter4_reset,
    output wire                                          from_t1_iter40_to_t1_iter41_clk,
    output wire [                                 512:0] from_t1_iter40_to_t1_iter41_if_din,
    input wire  [                                 512:0] from_t1_iter40_to_t1_iter41_if_dout,
    input wire                                           from_t1_iter40_to_t1_iter41_if_empty_n,
    input wire                                           from_t1_iter40_to_t1_iter41_if_full_n,
    output wire                                          from_t1_iter40_to_t1_iter41_if_read,
    output wire                                          from_t1_iter40_to_t1_iter41_if_read_ce,
    output wire                                          from_t1_iter40_to_t1_iter41_if_write,
    output wire                                          from_t1_iter40_to_t1_iter41_if_write_ce,
    output wire                                          from_t1_iter40_to_t1_iter41_reset,
    output wire                                          from_t1_iter41_to_t1_iter42_clk,
    output wire [                                 512:0] from_t1_iter41_to_t1_iter42_if_din,
    input wire  [                                 512:0] from_t1_iter41_to_t1_iter42_if_dout,
    input wire                                           from_t1_iter41_to_t1_iter42_if_empty_n,
    input wire                                           from_t1_iter41_to_t1_iter42_if_full_n,
    output wire                                          from_t1_iter41_to_t1_iter42_if_read,
    output wire                                          from_t1_iter41_to_t1_iter42_if_read_ce,
    output wire                                          from_t1_iter41_to_t1_iter42_if_write,
    output wire                                          from_t1_iter41_to_t1_iter42_if_write_ce,
    output wire                                          from_t1_iter41_to_t1_iter42_reset,
    output wire                                          from_t1_iter42_to_t1_iter43_clk,
    output wire [                                 512:0] from_t1_iter42_to_t1_iter43_if_din,
    input wire  [                                 512:0] from_t1_iter42_to_t1_iter43_if_dout,
    input wire                                           from_t1_iter42_to_t1_iter43_if_empty_n,
    input wire                                           from_t1_iter42_to_t1_iter43_if_full_n,
    output wire                                          from_t1_iter42_to_t1_iter43_if_read,
    output wire                                          from_t1_iter42_to_t1_iter43_if_read_ce,
    output wire                                          from_t1_iter42_to_t1_iter43_if_write,
    output wire                                          from_t1_iter42_to_t1_iter43_if_write_ce,
    output wire                                          from_t1_iter42_to_t1_iter43_reset,
    output wire                                          from_t1_iter43_to_t1_iter44_clk,
    output wire [                                 512:0] from_t1_iter43_to_t1_iter44_if_din,
    input wire  [                                 512:0] from_t1_iter43_to_t1_iter44_if_dout,
    input wire                                           from_t1_iter43_to_t1_iter44_if_empty_n,
    input wire                                           from_t1_iter43_to_t1_iter44_if_full_n,
    output wire                                          from_t1_iter43_to_t1_iter44_if_read,
    output wire                                          from_t1_iter43_to_t1_iter44_if_read_ce,
    output wire                                          from_t1_iter43_to_t1_iter44_if_write,
    output wire                                          from_t1_iter43_to_t1_iter44_if_write_ce,
    output wire                                          from_t1_iter43_to_t1_iter44_reset,
    output wire                                          from_t1_iter44_to_t1_iter45_clk,
    output wire [                                 512:0] from_t1_iter44_to_t1_iter45_if_din,
    input wire  [                                 512:0] from_t1_iter44_to_t1_iter45_if_dout,
    input wire                                           from_t1_iter44_to_t1_iter45_if_empty_n,
    input wire                                           from_t1_iter44_to_t1_iter45_if_full_n,
    output wire                                          from_t1_iter44_to_t1_iter45_if_read,
    output wire                                          from_t1_iter44_to_t1_iter45_if_read_ce,
    output wire                                          from_t1_iter44_to_t1_iter45_if_write,
    output wire                                          from_t1_iter44_to_t1_iter45_if_write_ce,
    output wire                                          from_t1_iter44_to_t1_iter45_reset,
    output wire                                          from_t1_iter45_to_t1_iter46_clk,
    output wire [                                 512:0] from_t1_iter45_to_t1_iter46_if_din,
    input wire  [                                 512:0] from_t1_iter45_to_t1_iter46_if_dout,
    input wire                                           from_t1_iter45_to_t1_iter46_if_empty_n,
    input wire                                           from_t1_iter45_to_t1_iter46_if_full_n,
    output wire                                          from_t1_iter45_to_t1_iter46_if_read,
    output wire                                          from_t1_iter45_to_t1_iter46_if_read_ce,
    output wire                                          from_t1_iter45_to_t1_iter46_if_write,
    output wire                                          from_t1_iter45_to_t1_iter46_if_write_ce,
    output wire                                          from_t1_iter45_to_t1_iter46_reset,
    output wire                                          from_t1_iter46_to_t1_iter47_clk,
    output wire [                                 512:0] from_t1_iter46_to_t1_iter47_if_din,
    input wire  [                                 512:0] from_t1_iter46_to_t1_iter47_if_dout,
    input wire                                           from_t1_iter46_to_t1_iter47_if_empty_n,
    input wire                                           from_t1_iter46_to_t1_iter47_if_full_n,
    output wire                                          from_t1_iter46_to_t1_iter47_if_read,
    output wire                                          from_t1_iter46_to_t1_iter47_if_read_ce,
    output wire                                          from_t1_iter46_to_t1_iter47_if_write,
    output wire                                          from_t1_iter46_to_t1_iter47_if_write_ce,
    output wire                                          from_t1_iter46_to_t1_iter47_reset,
    output wire                                          from_t1_iter47_to_t1_iter48_clk,
    output wire [                                 512:0] from_t1_iter47_to_t1_iter48_if_din,
    input wire  [                                 512:0] from_t1_iter47_to_t1_iter48_if_dout,
    input wire                                           from_t1_iter47_to_t1_iter48_if_empty_n,
    input wire                                           from_t1_iter47_to_t1_iter48_if_full_n,
    output wire                                          from_t1_iter47_to_t1_iter48_if_read,
    output wire                                          from_t1_iter47_to_t1_iter48_if_read_ce,
    output wire                                          from_t1_iter47_to_t1_iter48_if_write,
    output wire                                          from_t1_iter47_to_t1_iter48_if_write_ce,
    output wire                                          from_t1_iter47_to_t1_iter48_reset,
    output wire                                          from_t1_iter48_to_t1_iter49_clk,
    output wire [                                 512:0] from_t1_iter48_to_t1_iter49_if_din,
    input wire  [                                 512:0] from_t1_iter48_to_t1_iter49_if_dout,
    input wire                                           from_t1_iter48_to_t1_iter49_if_empty_n,
    input wire                                           from_t1_iter48_to_t1_iter49_if_full_n,
    output wire                                          from_t1_iter48_to_t1_iter49_if_read,
    output wire                                          from_t1_iter48_to_t1_iter49_if_read_ce,
    output wire                                          from_t1_iter48_to_t1_iter49_if_write,
    output wire                                          from_t1_iter48_to_t1_iter49_if_write_ce,
    output wire                                          from_t1_iter48_to_t1_iter49_reset,
    output wire                                          from_t1_iter49_to_t1_iter50_clk,
    output wire [                                 512:0] from_t1_iter49_to_t1_iter50_if_din,
    input wire  [                                 512:0] from_t1_iter49_to_t1_iter50_if_dout,
    input wire                                           from_t1_iter49_to_t1_iter50_if_empty_n,
    input wire                                           from_t1_iter49_to_t1_iter50_if_full_n,
    output wire                                          from_t1_iter49_to_t1_iter50_if_read,
    output wire                                          from_t1_iter49_to_t1_iter50_if_read_ce,
    output wire                                          from_t1_iter49_to_t1_iter50_if_write,
    output wire                                          from_t1_iter49_to_t1_iter50_if_write_ce,
    output wire                                          from_t1_iter49_to_t1_iter50_reset,
    output wire                                          from_t1_iter4_to_t1_iter5_clk,
    output wire [                                 512:0] from_t1_iter4_to_t1_iter5_if_din,
    input wire  [                                 512:0] from_t1_iter4_to_t1_iter5_if_dout,
    input wire                                           from_t1_iter4_to_t1_iter5_if_empty_n,
    input wire                                           from_t1_iter4_to_t1_iter5_if_full_n,
    output wire                                          from_t1_iter4_to_t1_iter5_if_read,
    output wire                                          from_t1_iter4_to_t1_iter5_if_read_ce,
    output wire                                          from_t1_iter4_to_t1_iter5_if_write,
    output wire                                          from_t1_iter4_to_t1_iter5_if_write_ce,
    output wire                                          from_t1_iter4_to_t1_iter5_reset,
    output wire                                          from_t1_iter50_to_t1_iter51_clk,
    output wire [                                 512:0] from_t1_iter50_to_t1_iter51_if_din,
    input wire  [                                 512:0] from_t1_iter50_to_t1_iter51_if_dout,
    input wire                                           from_t1_iter50_to_t1_iter51_if_empty_n,
    input wire                                           from_t1_iter50_to_t1_iter51_if_full_n,
    output wire                                          from_t1_iter50_to_t1_iter51_if_read,
    output wire                                          from_t1_iter50_to_t1_iter51_if_read_ce,
    output wire                                          from_t1_iter50_to_t1_iter51_if_write,
    output wire                                          from_t1_iter50_to_t1_iter51_if_write_ce,
    output wire                                          from_t1_iter50_to_t1_iter51_reset,
    output wire                                          from_t1_iter51_to_t1_iter52_clk,
    output wire [                                 512:0] from_t1_iter51_to_t1_iter52_if_din,
    input wire  [                                 512:0] from_t1_iter51_to_t1_iter52_if_dout,
    input wire                                           from_t1_iter51_to_t1_iter52_if_empty_n,
    input wire                                           from_t1_iter51_to_t1_iter52_if_full_n,
    output wire                                          from_t1_iter51_to_t1_iter52_if_read,
    output wire                                          from_t1_iter51_to_t1_iter52_if_read_ce,
    output wire                                          from_t1_iter51_to_t1_iter52_if_write,
    output wire                                          from_t1_iter51_to_t1_iter52_if_write_ce,
    output wire                                          from_t1_iter51_to_t1_iter52_reset,
    output wire                                          from_t1_iter52_to_t1_iter53_clk,
    output wire [                                 512:0] from_t1_iter52_to_t1_iter53_if_din,
    input wire  [                                 512:0] from_t1_iter52_to_t1_iter53_if_dout,
    input wire                                           from_t1_iter52_to_t1_iter53_if_empty_n,
    input wire                                           from_t1_iter52_to_t1_iter53_if_full_n,
    output wire                                          from_t1_iter52_to_t1_iter53_if_read,
    output wire                                          from_t1_iter52_to_t1_iter53_if_read_ce,
    output wire                                          from_t1_iter52_to_t1_iter53_if_write,
    output wire                                          from_t1_iter52_to_t1_iter53_if_write_ce,
    output wire                                          from_t1_iter52_to_t1_iter53_reset,
    output wire                                          from_t1_iter53_to_t1_iter54_clk,
    output wire [                                 512:0] from_t1_iter53_to_t1_iter54_if_din,
    input wire  [                                 512:0] from_t1_iter53_to_t1_iter54_if_dout,
    input wire                                           from_t1_iter53_to_t1_iter54_if_empty_n,
    input wire                                           from_t1_iter53_to_t1_iter54_if_full_n,
    output wire                                          from_t1_iter53_to_t1_iter54_if_read,
    output wire                                          from_t1_iter53_to_t1_iter54_if_read_ce,
    output wire                                          from_t1_iter53_to_t1_iter54_if_write,
    output wire                                          from_t1_iter53_to_t1_iter54_if_write_ce,
    output wire                                          from_t1_iter53_to_t1_iter54_reset,
    output wire                                          from_t1_iter54_to_t1_iter55_clk,
    output wire [                                 512:0] from_t1_iter54_to_t1_iter55_if_din,
    input wire  [                                 512:0] from_t1_iter54_to_t1_iter55_if_dout,
    input wire                                           from_t1_iter54_to_t1_iter55_if_empty_n,
    input wire                                           from_t1_iter54_to_t1_iter55_if_full_n,
    output wire                                          from_t1_iter54_to_t1_iter55_if_read,
    output wire                                          from_t1_iter54_to_t1_iter55_if_read_ce,
    output wire                                          from_t1_iter54_to_t1_iter55_if_write,
    output wire                                          from_t1_iter54_to_t1_iter55_if_write_ce,
    output wire                                          from_t1_iter54_to_t1_iter55_reset,
    output wire                                          from_t1_iter55_to_t1_iter56_clk,
    output wire [                                 512:0] from_t1_iter55_to_t1_iter56_if_din,
    input wire  [                                 512:0] from_t1_iter55_to_t1_iter56_if_dout,
    input wire                                           from_t1_iter55_to_t1_iter56_if_empty_n,
    input wire                                           from_t1_iter55_to_t1_iter56_if_full_n,
    output wire                                          from_t1_iter55_to_t1_iter56_if_read,
    output wire                                          from_t1_iter55_to_t1_iter56_if_read_ce,
    output wire                                          from_t1_iter55_to_t1_iter56_if_write,
    output wire                                          from_t1_iter55_to_t1_iter56_if_write_ce,
    output wire                                          from_t1_iter55_to_t1_iter56_reset,
    output wire                                          from_t1_iter56_to_t1_iter57_clk,
    output wire [                                 512:0] from_t1_iter56_to_t1_iter57_if_din,
    input wire  [                                 512:0] from_t1_iter56_to_t1_iter57_if_dout,
    input wire                                           from_t1_iter56_to_t1_iter57_if_empty_n,
    input wire                                           from_t1_iter56_to_t1_iter57_if_full_n,
    output wire                                          from_t1_iter56_to_t1_iter57_if_read,
    output wire                                          from_t1_iter56_to_t1_iter57_if_read_ce,
    output wire                                          from_t1_iter56_to_t1_iter57_if_write,
    output wire                                          from_t1_iter56_to_t1_iter57_if_write_ce,
    output wire                                          from_t1_iter56_to_t1_iter57_reset,
    output wire                                          from_t1_iter57_to_t1_iter58_clk,
    output wire [                                 512:0] from_t1_iter57_to_t1_iter58_if_din,
    input wire  [                                 512:0] from_t1_iter57_to_t1_iter58_if_dout,
    input wire                                           from_t1_iter57_to_t1_iter58_if_empty_n,
    input wire                                           from_t1_iter57_to_t1_iter58_if_full_n,
    output wire                                          from_t1_iter57_to_t1_iter58_if_read,
    output wire                                          from_t1_iter57_to_t1_iter58_if_read_ce,
    output wire                                          from_t1_iter57_to_t1_iter58_if_write,
    output wire                                          from_t1_iter57_to_t1_iter58_if_write_ce,
    output wire                                          from_t1_iter57_to_t1_iter58_reset,
    output wire                                          from_t1_iter58_to_t1_iter59_clk,
    output wire [                                 512:0] from_t1_iter58_to_t1_iter59_if_din,
    input wire  [                                 512:0] from_t1_iter58_to_t1_iter59_if_dout,
    input wire                                           from_t1_iter58_to_t1_iter59_if_empty_n,
    input wire                                           from_t1_iter58_to_t1_iter59_if_full_n,
    output wire                                          from_t1_iter58_to_t1_iter59_if_read,
    output wire                                          from_t1_iter58_to_t1_iter59_if_read_ce,
    output wire                                          from_t1_iter58_to_t1_iter59_if_write,
    output wire                                          from_t1_iter58_to_t1_iter59_if_write_ce,
    output wire                                          from_t1_iter58_to_t1_iter59_reset,
    output wire                                          from_t1_iter59_to_t1_iter60_clk,
    output wire [                                 512:0] from_t1_iter59_to_t1_iter60_if_din,
    input wire  [                                 512:0] from_t1_iter59_to_t1_iter60_if_dout,
    input wire                                           from_t1_iter59_to_t1_iter60_if_empty_n,
    input wire                                           from_t1_iter59_to_t1_iter60_if_full_n,
    output wire                                          from_t1_iter59_to_t1_iter60_if_read,
    output wire                                          from_t1_iter59_to_t1_iter60_if_read_ce,
    output wire                                          from_t1_iter59_to_t1_iter60_if_write,
    output wire                                          from_t1_iter59_to_t1_iter60_if_write_ce,
    output wire                                          from_t1_iter59_to_t1_iter60_reset,
    output wire                                          from_t1_iter5_to_t1_iter6_clk,
    output wire [                                 512:0] from_t1_iter5_to_t1_iter6_if_din,
    input wire  [                                 512:0] from_t1_iter5_to_t1_iter6_if_dout,
    input wire                                           from_t1_iter5_to_t1_iter6_if_empty_n,
    input wire                                           from_t1_iter5_to_t1_iter6_if_full_n,
    output wire                                          from_t1_iter5_to_t1_iter6_if_read,
    output wire                                          from_t1_iter5_to_t1_iter6_if_read_ce,
    output wire                                          from_t1_iter5_to_t1_iter6_if_write,
    output wire                                          from_t1_iter5_to_t1_iter6_if_write_ce,
    output wire                                          from_t1_iter5_to_t1_iter6_reset,
    output wire                                          from_t1_iter60_to_t1_iter61_clk,
    output wire [                                 512:0] from_t1_iter60_to_t1_iter61_if_din,
    input wire  [                                 512:0] from_t1_iter60_to_t1_iter61_if_dout,
    input wire                                           from_t1_iter60_to_t1_iter61_if_empty_n,
    input wire                                           from_t1_iter60_to_t1_iter61_if_full_n,
    output wire                                          from_t1_iter60_to_t1_iter61_if_read,
    output wire                                          from_t1_iter60_to_t1_iter61_if_read_ce,
    output wire                                          from_t1_iter60_to_t1_iter61_if_write,
    output wire                                          from_t1_iter60_to_t1_iter61_if_write_ce,
    output wire                                          from_t1_iter60_to_t1_iter61_reset,
    output wire                                          from_t1_iter61_to_t1_iter62_clk,
    output wire [                                 512:0] from_t1_iter61_to_t1_iter62_if_din,
    input wire  [                                 512:0] from_t1_iter61_to_t1_iter62_if_dout,
    input wire                                           from_t1_iter61_to_t1_iter62_if_empty_n,
    input wire                                           from_t1_iter61_to_t1_iter62_if_full_n,
    output wire                                          from_t1_iter61_to_t1_iter62_if_read,
    output wire                                          from_t1_iter61_to_t1_iter62_if_read_ce,
    output wire                                          from_t1_iter61_to_t1_iter62_if_write,
    output wire                                          from_t1_iter61_to_t1_iter62_if_write_ce,
    output wire                                          from_t1_iter61_to_t1_iter62_reset,
    output wire                                          from_t1_iter62_to_t1_iter63_clk,
    output wire [                                 512:0] from_t1_iter62_to_t1_iter63_if_din,
    input wire  [                                 512:0] from_t1_iter62_to_t1_iter63_if_dout,
    input wire                                           from_t1_iter62_to_t1_iter63_if_empty_n,
    input wire                                           from_t1_iter62_to_t1_iter63_if_full_n,
    output wire                                          from_t1_iter62_to_t1_iter63_if_read,
    output wire                                          from_t1_iter62_to_t1_iter63_if_read_ce,
    output wire                                          from_t1_iter62_to_t1_iter63_if_write,
    output wire                                          from_t1_iter62_to_t1_iter63_if_write_ce,
    output wire                                          from_t1_iter62_to_t1_iter63_reset,
    output wire                                          from_t1_iter63_to_t1_iter64_clk,
    output wire [                                 512:0] from_t1_iter63_to_t1_iter64_if_din,
    input wire  [                                 512:0] from_t1_iter63_to_t1_iter64_if_dout,
    input wire                                           from_t1_iter63_to_t1_iter64_if_empty_n,
    input wire                                           from_t1_iter63_to_t1_iter64_if_full_n,
    output wire                                          from_t1_iter63_to_t1_iter64_if_read,
    output wire                                          from_t1_iter63_to_t1_iter64_if_read_ce,
    output wire                                          from_t1_iter63_to_t1_iter64_if_write,
    output wire                                          from_t1_iter63_to_t1_iter64_if_write_ce,
    output wire                                          from_t1_iter63_to_t1_iter64_reset,
    output wire                                          from_t1_iter64_to_t1_iter65_clk,
    output wire [                                 512:0] from_t1_iter64_to_t1_iter65_if_din,
    input wire  [                                 512:0] from_t1_iter64_to_t1_iter65_if_dout,
    input wire                                           from_t1_iter64_to_t1_iter65_if_empty_n,
    input wire                                           from_t1_iter64_to_t1_iter65_if_full_n,
    output wire                                          from_t1_iter64_to_t1_iter65_if_read,
    output wire                                          from_t1_iter64_to_t1_iter65_if_read_ce,
    output wire                                          from_t1_iter64_to_t1_iter65_if_write,
    output wire                                          from_t1_iter64_to_t1_iter65_if_write_ce,
    output wire                                          from_t1_iter64_to_t1_iter65_reset,
    output wire                                          from_t1_iter65_to_t1_iter66_clk,
    output wire [                                 512:0] from_t1_iter65_to_t1_iter66_if_din,
    input wire  [                                 512:0] from_t1_iter65_to_t1_iter66_if_dout,
    input wire                                           from_t1_iter65_to_t1_iter66_if_empty_n,
    input wire                                           from_t1_iter65_to_t1_iter66_if_full_n,
    output wire                                          from_t1_iter65_to_t1_iter66_if_read,
    output wire                                          from_t1_iter65_to_t1_iter66_if_read_ce,
    output wire                                          from_t1_iter65_to_t1_iter66_if_write,
    output wire                                          from_t1_iter65_to_t1_iter66_if_write_ce,
    output wire                                          from_t1_iter65_to_t1_iter66_reset,
    output wire                                          from_t1_iter66_to_t1_iter67_clk,
    output wire [                                 512:0] from_t1_iter66_to_t1_iter67_if_din,
    input wire  [                                 512:0] from_t1_iter66_to_t1_iter67_if_dout,
    input wire                                           from_t1_iter66_to_t1_iter67_if_empty_n,
    input wire                                           from_t1_iter66_to_t1_iter67_if_full_n,
    output wire                                          from_t1_iter66_to_t1_iter67_if_read,
    output wire                                          from_t1_iter66_to_t1_iter67_if_read_ce,
    output wire                                          from_t1_iter66_to_t1_iter67_if_write,
    output wire                                          from_t1_iter66_to_t1_iter67_if_write_ce,
    output wire                                          from_t1_iter66_to_t1_iter67_reset,
    output wire                                          from_t1_iter67_to_t1_iter68_clk,
    output wire [                                 512:0] from_t1_iter67_to_t1_iter68_if_din,
    input wire  [                                 512:0] from_t1_iter67_to_t1_iter68_if_dout,
    input wire                                           from_t1_iter67_to_t1_iter68_if_empty_n,
    input wire                                           from_t1_iter67_to_t1_iter68_if_full_n,
    output wire                                          from_t1_iter67_to_t1_iter68_if_read,
    output wire                                          from_t1_iter67_to_t1_iter68_if_read_ce,
    output wire                                          from_t1_iter67_to_t1_iter68_if_write,
    output wire                                          from_t1_iter67_to_t1_iter68_if_write_ce,
    output wire                                          from_t1_iter67_to_t1_iter68_reset,
    output wire                                          from_t1_iter68_to_t1_iter69_clk,
    output wire [                                 512:0] from_t1_iter68_to_t1_iter69_if_din,
    input wire  [                                 512:0] from_t1_iter68_to_t1_iter69_if_dout,
    input wire                                           from_t1_iter68_to_t1_iter69_if_empty_n,
    input wire                                           from_t1_iter68_to_t1_iter69_if_full_n,
    output wire                                          from_t1_iter68_to_t1_iter69_if_read,
    output wire                                          from_t1_iter68_to_t1_iter69_if_read_ce,
    output wire                                          from_t1_iter68_to_t1_iter69_if_write,
    output wire                                          from_t1_iter68_to_t1_iter69_if_write_ce,
    output wire                                          from_t1_iter68_to_t1_iter69_reset,
    output wire                                          from_t1_iter69_to_t1_iter70_clk,
    output wire [                                 512:0] from_t1_iter69_to_t1_iter70_if_din,
    input wire  [                                 512:0] from_t1_iter69_to_t1_iter70_if_dout,
    input wire                                           from_t1_iter69_to_t1_iter70_if_empty_n,
    input wire                                           from_t1_iter69_to_t1_iter70_if_full_n,
    output wire                                          from_t1_iter69_to_t1_iter70_if_read,
    output wire                                          from_t1_iter69_to_t1_iter70_if_read_ce,
    output wire                                          from_t1_iter69_to_t1_iter70_if_write,
    output wire                                          from_t1_iter69_to_t1_iter70_if_write_ce,
    output wire                                          from_t1_iter69_to_t1_iter70_reset,
    output wire                                          from_t1_iter6_to_t1_iter7_clk,
    output wire [                                 512:0] from_t1_iter6_to_t1_iter7_if_din,
    input wire  [                                 512:0] from_t1_iter6_to_t1_iter7_if_dout,
    input wire                                           from_t1_iter6_to_t1_iter7_if_empty_n,
    input wire                                           from_t1_iter6_to_t1_iter7_if_full_n,
    output wire                                          from_t1_iter6_to_t1_iter7_if_read,
    output wire                                          from_t1_iter6_to_t1_iter7_if_read_ce,
    output wire                                          from_t1_iter6_to_t1_iter7_if_write,
    output wire                                          from_t1_iter6_to_t1_iter7_if_write_ce,
    output wire                                          from_t1_iter6_to_t1_iter7_reset,
    output wire                                          from_t1_iter70_to_t1_iter71_clk,
    output wire [                                 512:0] from_t1_iter70_to_t1_iter71_if_din,
    input wire  [                                 512:0] from_t1_iter70_to_t1_iter71_if_dout,
    input wire                                           from_t1_iter70_to_t1_iter71_if_empty_n,
    input wire                                           from_t1_iter70_to_t1_iter71_if_full_n,
    output wire                                          from_t1_iter70_to_t1_iter71_if_read,
    output wire                                          from_t1_iter70_to_t1_iter71_if_read_ce,
    output wire                                          from_t1_iter70_to_t1_iter71_if_write,
    output wire                                          from_t1_iter70_to_t1_iter71_if_write_ce,
    output wire                                          from_t1_iter70_to_t1_iter71_reset,
    output wire                                          from_t1_iter71_to_t1_iter72_clk,
    output wire [                                 512:0] from_t1_iter71_to_t1_iter72_if_din,
    input wire  [                                 512:0] from_t1_iter71_to_t1_iter72_if_dout,
    input wire                                           from_t1_iter71_to_t1_iter72_if_empty_n,
    input wire                                           from_t1_iter71_to_t1_iter72_if_full_n,
    output wire                                          from_t1_iter71_to_t1_iter72_if_read,
    output wire                                          from_t1_iter71_to_t1_iter72_if_read_ce,
    output wire                                          from_t1_iter71_to_t1_iter72_if_write,
    output wire                                          from_t1_iter71_to_t1_iter72_if_write_ce,
    output wire                                          from_t1_iter71_to_t1_iter72_reset,
    output wire                                          from_t1_iter72_to_t1_iter73_clk,
    output wire [                                 512:0] from_t1_iter72_to_t1_iter73_if_din,
    input wire  [                                 512:0] from_t1_iter72_to_t1_iter73_if_dout,
    input wire                                           from_t1_iter72_to_t1_iter73_if_empty_n,
    input wire                                           from_t1_iter72_to_t1_iter73_if_full_n,
    output wire                                          from_t1_iter72_to_t1_iter73_if_read,
    output wire                                          from_t1_iter72_to_t1_iter73_if_read_ce,
    output wire                                          from_t1_iter72_to_t1_iter73_if_write,
    output wire                                          from_t1_iter72_to_t1_iter73_if_write_ce,
    output wire                                          from_t1_iter72_to_t1_iter73_reset,
    output wire                                          from_t1_iter73_to_t1_iter74_clk,
    output wire [                                 512:0] from_t1_iter73_to_t1_iter74_if_din,
    input wire  [                                 512:0] from_t1_iter73_to_t1_iter74_if_dout,
    input wire                                           from_t1_iter73_to_t1_iter74_if_empty_n,
    input wire                                           from_t1_iter73_to_t1_iter74_if_full_n,
    output wire                                          from_t1_iter73_to_t1_iter74_if_read,
    output wire                                          from_t1_iter73_to_t1_iter74_if_read_ce,
    output wire                                          from_t1_iter73_to_t1_iter74_if_write,
    output wire                                          from_t1_iter73_to_t1_iter74_if_write_ce,
    output wire                                          from_t1_iter73_to_t1_iter74_reset,
    output wire                                          from_t1_iter74_to_t1_iter75_clk,
    output wire [                                 512:0] from_t1_iter74_to_t1_iter75_if_din,
    input wire  [                                 512:0] from_t1_iter74_to_t1_iter75_if_dout,
    input wire                                           from_t1_iter74_to_t1_iter75_if_empty_n,
    input wire                                           from_t1_iter74_to_t1_iter75_if_full_n,
    output wire                                          from_t1_iter74_to_t1_iter75_if_read,
    output wire                                          from_t1_iter74_to_t1_iter75_if_read_ce,
    output wire                                          from_t1_iter74_to_t1_iter75_if_write,
    output wire                                          from_t1_iter74_to_t1_iter75_if_write_ce,
    output wire                                          from_t1_iter74_to_t1_iter75_reset,
    output wire                                          from_t1_iter75_to_t1_iter76_clk,
    output wire [                                 512:0] from_t1_iter75_to_t1_iter76_if_din,
    input wire  [                                 512:0] from_t1_iter75_to_t1_iter76_if_dout,
    input wire                                           from_t1_iter75_to_t1_iter76_if_empty_n,
    input wire                                           from_t1_iter75_to_t1_iter76_if_full_n,
    output wire                                          from_t1_iter75_to_t1_iter76_if_read,
    output wire                                          from_t1_iter75_to_t1_iter76_if_read_ce,
    output wire                                          from_t1_iter75_to_t1_iter76_if_write,
    output wire                                          from_t1_iter75_to_t1_iter76_if_write_ce,
    output wire                                          from_t1_iter75_to_t1_iter76_reset,
    output wire                                          from_t1_iter76_to_t1_iter77_clk,
    output wire [                                 512:0] from_t1_iter76_to_t1_iter77_if_din,
    input wire  [                                 512:0] from_t1_iter76_to_t1_iter77_if_dout,
    input wire                                           from_t1_iter76_to_t1_iter77_if_empty_n,
    input wire                                           from_t1_iter76_to_t1_iter77_if_full_n,
    output wire                                          from_t1_iter76_to_t1_iter77_if_read,
    output wire                                          from_t1_iter76_to_t1_iter77_if_read_ce,
    output wire                                          from_t1_iter76_to_t1_iter77_if_write,
    output wire                                          from_t1_iter76_to_t1_iter77_if_write_ce,
    output wire                                          from_t1_iter76_to_t1_iter77_reset,
    output wire                                          from_t1_iter77_to_t1_iter78_clk,
    output wire [                                 512:0] from_t1_iter77_to_t1_iter78_if_din,
    input wire  [                                 512:0] from_t1_iter77_to_t1_iter78_if_dout,
    input wire                                           from_t1_iter77_to_t1_iter78_if_empty_n,
    input wire                                           from_t1_iter77_to_t1_iter78_if_full_n,
    output wire                                          from_t1_iter77_to_t1_iter78_if_read,
    output wire                                          from_t1_iter77_to_t1_iter78_if_read_ce,
    output wire                                          from_t1_iter77_to_t1_iter78_if_write,
    output wire                                          from_t1_iter77_to_t1_iter78_if_write_ce,
    output wire                                          from_t1_iter77_to_t1_iter78_reset,
    output wire                                          from_t1_iter78_to_t1_iter79_clk,
    output wire [                                 512:0] from_t1_iter78_to_t1_iter79_if_din,
    input wire  [                                 512:0] from_t1_iter78_to_t1_iter79_if_dout,
    input wire                                           from_t1_iter78_to_t1_iter79_if_empty_n,
    input wire                                           from_t1_iter78_to_t1_iter79_if_full_n,
    output wire                                          from_t1_iter78_to_t1_iter79_if_read,
    output wire                                          from_t1_iter78_to_t1_iter79_if_read_ce,
    output wire                                          from_t1_iter78_to_t1_iter79_if_write,
    output wire                                          from_t1_iter78_to_t1_iter79_if_write_ce,
    output wire                                          from_t1_iter78_to_t1_iter79_reset,
    output wire                                          from_t1_iter79_to_t1_iter80_clk,
    output wire [                                 512:0] from_t1_iter79_to_t1_iter80_if_din,
    input wire  [                                 512:0] from_t1_iter79_to_t1_iter80_if_dout,
    input wire                                           from_t1_iter79_to_t1_iter80_if_empty_n,
    input wire                                           from_t1_iter79_to_t1_iter80_if_full_n,
    output wire                                          from_t1_iter79_to_t1_iter80_if_read,
    output wire                                          from_t1_iter79_to_t1_iter80_if_read_ce,
    output wire                                          from_t1_iter79_to_t1_iter80_if_write,
    output wire                                          from_t1_iter79_to_t1_iter80_if_write_ce,
    output wire                                          from_t1_iter79_to_t1_iter80_reset,
    output wire                                          from_t1_iter7_to_t1_iter8_clk,
    output wire [                                 512:0] from_t1_iter7_to_t1_iter8_if_din,
    input wire  [                                 512:0] from_t1_iter7_to_t1_iter8_if_dout,
    input wire                                           from_t1_iter7_to_t1_iter8_if_empty_n,
    input wire                                           from_t1_iter7_to_t1_iter8_if_full_n,
    output wire                                          from_t1_iter7_to_t1_iter8_if_read,
    output wire                                          from_t1_iter7_to_t1_iter8_if_read_ce,
    output wire                                          from_t1_iter7_to_t1_iter8_if_write,
    output wire                                          from_t1_iter7_to_t1_iter8_if_write_ce,
    output wire                                          from_t1_iter7_to_t1_iter8_reset,
    output wire                                          from_t1_iter80_to_t1_iter81_clk,
    output wire [                                 512:0] from_t1_iter80_to_t1_iter81_if_din,
    input wire  [                                 512:0] from_t1_iter80_to_t1_iter81_if_dout,
    input wire                                           from_t1_iter80_to_t1_iter81_if_empty_n,
    input wire                                           from_t1_iter80_to_t1_iter81_if_full_n,
    output wire                                          from_t1_iter80_to_t1_iter81_if_read,
    output wire                                          from_t1_iter80_to_t1_iter81_if_read_ce,
    output wire                                          from_t1_iter80_to_t1_iter81_if_write,
    output wire                                          from_t1_iter80_to_t1_iter81_if_write_ce,
    output wire                                          from_t1_iter80_to_t1_iter81_reset,
    output wire                                          from_t1_iter81_to_t1_iter82_clk,
    output wire [                                 512:0] from_t1_iter81_to_t1_iter82_if_din,
    input wire  [                                 512:0] from_t1_iter81_to_t1_iter82_if_dout,
    input wire                                           from_t1_iter81_to_t1_iter82_if_empty_n,
    input wire                                           from_t1_iter81_to_t1_iter82_if_full_n,
    output wire                                          from_t1_iter81_to_t1_iter82_if_read,
    output wire                                          from_t1_iter81_to_t1_iter82_if_read_ce,
    output wire                                          from_t1_iter81_to_t1_iter82_if_write,
    output wire                                          from_t1_iter81_to_t1_iter82_if_write_ce,
    output wire                                          from_t1_iter81_to_t1_iter82_reset,
    output wire                                          from_t1_iter82_to_t1_iter83_clk,
    output wire [                                 512:0] from_t1_iter82_to_t1_iter83_if_din,
    input wire  [                                 512:0] from_t1_iter82_to_t1_iter83_if_dout,
    input wire                                           from_t1_iter82_to_t1_iter83_if_empty_n,
    input wire                                           from_t1_iter82_to_t1_iter83_if_full_n,
    output wire                                          from_t1_iter82_to_t1_iter83_if_read,
    output wire                                          from_t1_iter82_to_t1_iter83_if_read_ce,
    output wire                                          from_t1_iter82_to_t1_iter83_if_write,
    output wire                                          from_t1_iter82_to_t1_iter83_if_write_ce,
    output wire                                          from_t1_iter82_to_t1_iter83_reset,
    output wire                                          from_t1_iter83_to_t1_iter84_clk,
    output wire [                                 512:0] from_t1_iter83_to_t1_iter84_if_din,
    input wire  [                                 512:0] from_t1_iter83_to_t1_iter84_if_dout,
    input wire                                           from_t1_iter83_to_t1_iter84_if_empty_n,
    input wire                                           from_t1_iter83_to_t1_iter84_if_full_n,
    output wire                                          from_t1_iter83_to_t1_iter84_if_read,
    output wire                                          from_t1_iter83_to_t1_iter84_if_read_ce,
    output wire                                          from_t1_iter83_to_t1_iter84_if_write,
    output wire                                          from_t1_iter83_to_t1_iter84_if_write_ce,
    output wire                                          from_t1_iter83_to_t1_iter84_reset,
    output wire                                          from_t1_iter84_to_t1_iter85_clk,
    output wire [                                 512:0] from_t1_iter84_to_t1_iter85_if_din,
    input wire  [                                 512:0] from_t1_iter84_to_t1_iter85_if_dout,
    input wire                                           from_t1_iter84_to_t1_iter85_if_empty_n,
    input wire                                           from_t1_iter84_to_t1_iter85_if_full_n,
    output wire                                          from_t1_iter84_to_t1_iter85_if_read,
    output wire                                          from_t1_iter84_to_t1_iter85_if_read_ce,
    output wire                                          from_t1_iter84_to_t1_iter85_if_write,
    output wire                                          from_t1_iter84_to_t1_iter85_if_write_ce,
    output wire                                          from_t1_iter84_to_t1_iter85_reset,
    output wire                                          from_t1_iter85_to_t1_iter86_clk,
    output wire [                                 512:0] from_t1_iter85_to_t1_iter86_if_din,
    input wire  [                                 512:0] from_t1_iter85_to_t1_iter86_if_dout,
    input wire                                           from_t1_iter85_to_t1_iter86_if_empty_n,
    input wire                                           from_t1_iter85_to_t1_iter86_if_full_n,
    output wire                                          from_t1_iter85_to_t1_iter86_if_read,
    output wire                                          from_t1_iter85_to_t1_iter86_if_read_ce,
    output wire                                          from_t1_iter85_to_t1_iter86_if_write,
    output wire                                          from_t1_iter85_to_t1_iter86_if_write_ce,
    output wire                                          from_t1_iter85_to_t1_iter86_reset,
    output wire                                          from_t1_iter86_to_t1_iter87_clk,
    output wire [                                 512:0] from_t1_iter86_to_t1_iter87_if_din,
    input wire  [                                 512:0] from_t1_iter86_to_t1_iter87_if_dout,
    input wire                                           from_t1_iter86_to_t1_iter87_if_empty_n,
    input wire                                           from_t1_iter86_to_t1_iter87_if_full_n,
    output wire                                          from_t1_iter86_to_t1_iter87_if_read,
    output wire                                          from_t1_iter86_to_t1_iter87_if_read_ce,
    output wire                                          from_t1_iter86_to_t1_iter87_if_write,
    output wire                                          from_t1_iter86_to_t1_iter87_if_write_ce,
    output wire                                          from_t1_iter86_to_t1_iter87_reset,
    output wire                                          from_t1_iter87_to_t1_iter88_clk,
    output wire [                                 512:0] from_t1_iter87_to_t1_iter88_if_din,
    input wire  [                                 512:0] from_t1_iter87_to_t1_iter88_if_dout,
    input wire                                           from_t1_iter87_to_t1_iter88_if_empty_n,
    input wire                                           from_t1_iter87_to_t1_iter88_if_full_n,
    output wire                                          from_t1_iter87_to_t1_iter88_if_read,
    output wire                                          from_t1_iter87_to_t1_iter88_if_read_ce,
    output wire                                          from_t1_iter87_to_t1_iter88_if_write,
    output wire                                          from_t1_iter87_to_t1_iter88_if_write_ce,
    output wire                                          from_t1_iter87_to_t1_iter88_reset,
    output wire                                          from_t1_iter88_to_t1_iter89_clk,
    output wire [                                 512:0] from_t1_iter88_to_t1_iter89_if_din,
    input wire  [                                 512:0] from_t1_iter88_to_t1_iter89_if_dout,
    input wire                                           from_t1_iter88_to_t1_iter89_if_empty_n,
    input wire                                           from_t1_iter88_to_t1_iter89_if_full_n,
    output wire                                          from_t1_iter88_to_t1_iter89_if_read,
    output wire                                          from_t1_iter88_to_t1_iter89_if_read_ce,
    output wire                                          from_t1_iter88_to_t1_iter89_if_write,
    output wire                                          from_t1_iter88_to_t1_iter89_if_write_ce,
    output wire                                          from_t1_iter88_to_t1_iter89_reset,
    output wire                                          from_t1_iter89_to_t1_iter90_clk,
    output wire [                                 512:0] from_t1_iter89_to_t1_iter90_if_din,
    input wire  [                                 512:0] from_t1_iter89_to_t1_iter90_if_dout,
    input wire                                           from_t1_iter89_to_t1_iter90_if_empty_n,
    input wire                                           from_t1_iter89_to_t1_iter90_if_full_n,
    output wire                                          from_t1_iter89_to_t1_iter90_if_read,
    output wire                                          from_t1_iter89_to_t1_iter90_if_read_ce,
    output wire                                          from_t1_iter89_to_t1_iter90_if_write,
    output wire                                          from_t1_iter89_to_t1_iter90_if_write_ce,
    output wire                                          from_t1_iter89_to_t1_iter90_reset,
    output wire                                          from_t1_iter8_to_t1_iter9_clk,
    output wire [                                 512:0] from_t1_iter8_to_t1_iter9_if_din,
    input wire  [                                 512:0] from_t1_iter8_to_t1_iter9_if_dout,
    input wire                                           from_t1_iter8_to_t1_iter9_if_empty_n,
    input wire                                           from_t1_iter8_to_t1_iter9_if_full_n,
    output wire                                          from_t1_iter8_to_t1_iter9_if_read,
    output wire                                          from_t1_iter8_to_t1_iter9_if_read_ce,
    output wire                                          from_t1_iter8_to_t1_iter9_if_write,
    output wire                                          from_t1_iter8_to_t1_iter9_if_write_ce,
    output wire                                          from_t1_iter8_to_t1_iter9_reset,
    output wire                                          from_t1_iter90_to_t1_iter91_clk,
    output wire [                                 512:0] from_t1_iter90_to_t1_iter91_if_din,
    input wire  [                                 512:0] from_t1_iter90_to_t1_iter91_if_dout,
    input wire                                           from_t1_iter90_to_t1_iter91_if_empty_n,
    input wire                                           from_t1_iter90_to_t1_iter91_if_full_n,
    output wire                                          from_t1_iter90_to_t1_iter91_if_read,
    output wire                                          from_t1_iter90_to_t1_iter91_if_read_ce,
    output wire                                          from_t1_iter90_to_t1_iter91_if_write,
    output wire                                          from_t1_iter90_to_t1_iter91_if_write_ce,
    output wire                                          from_t1_iter90_to_t1_iter91_reset,
    output wire                                          from_t1_iter91_to_t1_iter92_clk,
    output wire [                                 512:0] from_t1_iter91_to_t1_iter92_if_din,
    input wire  [                                 512:0] from_t1_iter91_to_t1_iter92_if_dout,
    input wire                                           from_t1_iter91_to_t1_iter92_if_empty_n,
    input wire                                           from_t1_iter91_to_t1_iter92_if_full_n,
    output wire                                          from_t1_iter91_to_t1_iter92_if_read,
    output wire                                          from_t1_iter91_to_t1_iter92_if_read_ce,
    output wire                                          from_t1_iter91_to_t1_iter92_if_write,
    output wire                                          from_t1_iter91_to_t1_iter92_if_write_ce,
    output wire                                          from_t1_iter91_to_t1_iter92_reset,
    output wire                                          from_t1_iter92_to_t1_iter93_clk,
    output wire [                                 512:0] from_t1_iter92_to_t1_iter93_if_din,
    input wire  [                                 512:0] from_t1_iter92_to_t1_iter93_if_dout,
    input wire                                           from_t1_iter92_to_t1_iter93_if_empty_n,
    input wire                                           from_t1_iter92_to_t1_iter93_if_full_n,
    output wire                                          from_t1_iter92_to_t1_iter93_if_read,
    output wire                                          from_t1_iter92_to_t1_iter93_if_read_ce,
    output wire                                          from_t1_iter92_to_t1_iter93_if_write,
    output wire                                          from_t1_iter92_to_t1_iter93_if_write_ce,
    output wire                                          from_t1_iter92_to_t1_iter93_reset,
    output wire                                          from_t1_iter93_to_t1_iter94_clk,
    output wire [                                 512:0] from_t1_iter93_to_t1_iter94_if_din,
    input wire  [                                 512:0] from_t1_iter93_to_t1_iter94_if_dout,
    input wire                                           from_t1_iter93_to_t1_iter94_if_empty_n,
    input wire                                           from_t1_iter93_to_t1_iter94_if_full_n,
    output wire                                          from_t1_iter93_to_t1_iter94_if_read,
    output wire                                          from_t1_iter93_to_t1_iter94_if_read_ce,
    output wire                                          from_t1_iter93_to_t1_iter94_if_write,
    output wire                                          from_t1_iter93_to_t1_iter94_if_write_ce,
    output wire                                          from_t1_iter93_to_t1_iter94_reset,
    output wire                                          from_t1_iter94_to_t1_iter95_clk,
    output wire [                                 512:0] from_t1_iter94_to_t1_iter95_if_din,
    input wire  [                                 512:0] from_t1_iter94_to_t1_iter95_if_dout,
    input wire                                           from_t1_iter94_to_t1_iter95_if_empty_n,
    input wire                                           from_t1_iter94_to_t1_iter95_if_full_n,
    output wire                                          from_t1_iter94_to_t1_iter95_if_read,
    output wire                                          from_t1_iter94_to_t1_iter95_if_read_ce,
    output wire                                          from_t1_iter94_to_t1_iter95_if_write,
    output wire                                          from_t1_iter94_to_t1_iter95_if_write_ce,
    output wire                                          from_t1_iter94_to_t1_iter95_reset,
    output wire                                          from_t1_iter95_to_t1_iter96_clk,
    output wire [                                 512:0] from_t1_iter95_to_t1_iter96_if_din,
    input wire  [                                 512:0] from_t1_iter95_to_t1_iter96_if_dout,
    input wire                                           from_t1_iter95_to_t1_iter96_if_empty_n,
    input wire                                           from_t1_iter95_to_t1_iter96_if_full_n,
    output wire                                          from_t1_iter95_to_t1_iter96_if_read,
    output wire                                          from_t1_iter95_to_t1_iter96_if_read_ce,
    output wire                                          from_t1_iter95_to_t1_iter96_if_write,
    output wire                                          from_t1_iter95_to_t1_iter96_if_write_ce,
    output wire                                          from_t1_iter95_to_t1_iter96_reset,
    output wire                                          from_t1_iter96_to_t1_iter97_clk,
    output wire [                                 512:0] from_t1_iter96_to_t1_iter97_if_din,
    input wire  [                                 512:0] from_t1_iter96_to_t1_iter97_if_dout,
    input wire                                           from_t1_iter96_to_t1_iter97_if_empty_n,
    input wire                                           from_t1_iter96_to_t1_iter97_if_full_n,
    output wire                                          from_t1_iter96_to_t1_iter97_if_read,
    output wire                                          from_t1_iter96_to_t1_iter97_if_read_ce,
    output wire                                          from_t1_iter96_to_t1_iter97_if_write,
    output wire                                          from_t1_iter96_to_t1_iter97_if_write_ce,
    output wire                                          from_t1_iter96_to_t1_iter97_reset,
    output wire                                          from_t1_iter97_to_t1_iter98_clk,
    output wire [                                 512:0] from_t1_iter97_to_t1_iter98_if_din,
    input wire  [                                 512:0] from_t1_iter97_to_t1_iter98_if_dout,
    input wire                                           from_t1_iter97_to_t1_iter98_if_empty_n,
    input wire                                           from_t1_iter97_to_t1_iter98_if_full_n,
    output wire                                          from_t1_iter97_to_t1_iter98_if_read,
    output wire                                          from_t1_iter97_to_t1_iter98_if_read_ce,
    output wire                                          from_t1_iter97_to_t1_iter98_if_write,
    output wire                                          from_t1_iter97_to_t1_iter98_if_write_ce,
    output wire                                          from_t1_iter97_to_t1_iter98_reset,
    output wire                                          from_t1_iter98_to_t1_iter99_clk,
    output wire [                                 512:0] from_t1_iter98_to_t1_iter99_if_din,
    input wire  [                                 512:0] from_t1_iter98_to_t1_iter99_if_dout,
    input wire                                           from_t1_iter98_to_t1_iter99_if_empty_n,
    input wire                                           from_t1_iter98_to_t1_iter99_if_full_n,
    output wire                                          from_t1_iter98_to_t1_iter99_if_read,
    output wire                                          from_t1_iter98_to_t1_iter99_if_read_ce,
    output wire                                          from_t1_iter98_to_t1_iter99_if_write,
    output wire                                          from_t1_iter98_to_t1_iter99_if_write_ce,
    output wire                                          from_t1_iter98_to_t1_iter99_reset,
    output wire                                          from_t1_iter99_to_t1_iter100_clk,
    output wire [                                 512:0] from_t1_iter99_to_t1_iter100_if_din,
    input wire  [                                 512:0] from_t1_iter99_to_t1_iter100_if_dout,
    input wire                                           from_t1_iter99_to_t1_iter100_if_empty_n,
    input wire                                           from_t1_iter99_to_t1_iter100_if_full_n,
    output wire                                          from_t1_iter99_to_t1_iter100_if_read,
    output wire                                          from_t1_iter99_to_t1_iter100_if_read_ce,
    output wire                                          from_t1_iter99_to_t1_iter100_if_write,
    output wire                                          from_t1_iter99_to_t1_iter100_if_write_ce,
    output wire                                          from_t1_iter99_to_t1_iter100_reset,
    output wire                                          from_t1_iter9_to_t1_iter10_clk,
    output wire [                                 512:0] from_t1_iter9_to_t1_iter10_if_din,
    input wire  [                                 512:0] from_t1_iter9_to_t1_iter10_if_dout,
    input wire                                           from_t1_iter9_to_t1_iter10_if_empty_n,
    input wire                                           from_t1_iter9_to_t1_iter10_if_full_n,
    output wire                                          from_t1_iter9_to_t1_iter10_if_read,
    output wire                                          from_t1_iter9_to_t1_iter10_if_read_ce,
    output wire                                          from_t1_iter9_to_t1_iter10_if_write,
    output wire                                          from_t1_iter9_to_t1_iter10_if_write_ce,
    output wire                                          from_t1_iter9_to_t1_iter10_reset,
    output wire                                          BurstRead_floatx16_0_ap_clk,
    input wire                                           BurstRead_floatx16_0_ap_done,
    input wire                                           BurstRead_floatx16_0_ap_idle,
    input wire                                           BurstRead_floatx16_0_ap_ready,
    output wire                                          BurstRead_floatx16_0_ap_rst_n,
    output wire                                          BurstRead_floatx16_0_ap_start,
    input wire  [                                 512:0] BurstRead_floatx16_0_dest_din,
    output wire                                          BurstRead_floatx16_0_dest_full_n,
    input wire                                           BurstRead_floatx16_0_dest_write,
    output wire [                                  63:0] BurstRead_floatx16_0_n,
    output wire [                                  63:0] BurstRead_floatx16_0_src_read_addr_offset,
    input wire  [                                  63:0] BurstRead_floatx16_0_src_read_addr_s_din,
    output wire                                          BurstRead_floatx16_0_src_read_addr_s_full_n,
    input wire                                           BurstRead_floatx16_0_src_read_addr_s_write,
    output wire [                                 512:0] BurstRead_floatx16_0_src_read_data_peek_dout,
    output wire                                          BurstRead_floatx16_0_src_read_data_peek_empty_n,
    input wire                                           BurstRead_floatx16_0_src_read_data_peek_read,
    output wire [                                 512:0] BurstRead_floatx16_0_src_read_data_s_dout,
    output wire                                          BurstRead_floatx16_0_src_read_data_s_empty_n,
    input wire                                           BurstRead_floatx16_0_src_read_data_s_read,
    output wire [                                  63:0] BurstRead_floatx16_0_src_write_addr_offset,
    input wire  [                                  63:0] BurstRead_floatx16_0_src_write_addr_s_din,
    output wire                                          BurstRead_floatx16_0_src_write_addr_s_full_n,
    input wire                                           BurstRead_floatx16_0_src_write_addr_s_write,
    input wire  [                                 512:0] BurstRead_floatx16_0_src_write_data_din,
    output wire                                          BurstRead_floatx16_0_src_write_data_full_n,
    input wire                                           BurstRead_floatx16_0_src_write_data_write,
    output wire [                                   8:0] BurstRead_floatx16_0_src_write_resp_peek_dout,
    output wire                                          BurstRead_floatx16_0_src_write_resp_peek_empty_n,
    input wire                                           BurstRead_floatx16_0_src_write_resp_peek_read,
    output wire [                                   8:0] BurstRead_floatx16_0_src_write_resp_s_dout,
    output wire                                          BurstRead_floatx16_0_src_write_resp_s_empty_n,
    input wire                                           BurstRead_floatx16_0_src_write_resp_s_read,
    output wire                                          BurstWrite_floatx16_0_ap_clk,
    input wire                                           BurstWrite_floatx16_0_ap_done,
    input wire                                           BurstWrite_floatx16_0_ap_idle,
    input wire                                           BurstWrite_floatx16_0_ap_ready,
    output wire                                          BurstWrite_floatx16_0_ap_rst_n,
    output wire                                          BurstWrite_floatx16_0_ap_start,
    output wire [                                  63:0] BurstWrite_floatx16_0_dest_read_addr_offset,
    input wire  [                                  63:0] BurstWrite_floatx16_0_dest_read_addr_s_din,
    output wire                                          BurstWrite_floatx16_0_dest_read_addr_s_full_n,
    input wire                                           BurstWrite_floatx16_0_dest_read_addr_s_write,
    output wire [                                 512:0] BurstWrite_floatx16_0_dest_read_data_peek_dout,
    output wire                                          BurstWrite_floatx16_0_dest_read_data_peek_empty_n,
    input wire                                           BurstWrite_floatx16_0_dest_read_data_peek_read,
    output wire [                                 512:0] BurstWrite_floatx16_0_dest_read_data_s_dout,
    output wire                                          BurstWrite_floatx16_0_dest_read_data_s_empty_n,
    input wire                                           BurstWrite_floatx16_0_dest_read_data_s_read,
    output wire [                                  63:0] BurstWrite_floatx16_0_dest_write_addr_offset,
    input wire  [                                  63:0] BurstWrite_floatx16_0_dest_write_addr_s_din,
    output wire                                          BurstWrite_floatx16_0_dest_write_addr_s_full_n,
    input wire                                           BurstWrite_floatx16_0_dest_write_addr_s_write,
    input wire  [                                 512:0] BurstWrite_floatx16_0_dest_write_data_din,
    output wire                                          BurstWrite_floatx16_0_dest_write_data_full_n,
    input wire                                           BurstWrite_floatx16_0_dest_write_data_write,
    output wire [                                   8:0] BurstWrite_floatx16_0_dest_write_resp_peek_dout,
    output wire                                          BurstWrite_floatx16_0_dest_write_resp_peek_empty_n,
    input wire                                           BurstWrite_floatx16_0_dest_write_resp_peek_read,
    output wire [                                   8:0] BurstWrite_floatx16_0_dest_write_resp_s_dout,
    output wire                                          BurstWrite_floatx16_0_dest_write_resp_s_empty_n,
    input wire                                           BurstWrite_floatx16_0_dest_write_resp_s_read,
    output wire [                                  63:0] BurstWrite_floatx16_0_n,
    output wire [                                 512:0] BurstWrite_floatx16_0_src_peek_dout,
    output wire                                          BurstWrite_floatx16_0_src_peek_empty_n,
    input wire                                           BurstWrite_floatx16_0_src_peek_read,
    output wire [                                 512:0] BurstWrite_floatx16_0_src_s_dout,
    output wire                                          BurstWrite_floatx16_0_src_s_empty_n,
    input wire                                           BurstWrite_floatx16_0_src_s_read,
    output wire                                          Module0Func_0_ap_clk,
    input wire                                           Module0Func_0_ap_done,
    input wire                                           Module0Func_0_ap_idle,
    input wire                                           Module0Func_0_ap_ready,
    output wire                                          Module0Func_0_ap_rst_n,
    output wire                                          Module0Func_0_ap_start,
    output wire [                                 512:0] Module0Func_0_dram_t1_bank_0_fifo_peek_dout,
    output wire                                          Module0Func_0_dram_t1_bank_0_fifo_peek_empty_n,
    input wire                                           Module0Func_0_dram_t1_bank_0_fifo_peek_read,
    output wire [                                 512:0] Module0Func_0_dram_t1_bank_0_fifo_s_dout,
    output wire                                          Module0Func_0_dram_t1_bank_0_fifo_s_empty_n,
    input wire                                           Module0Func_0_dram_t1_bank_0_fifo_s_read,
    input wire  [                                 512:0] Module0Func_0_fifo_st_0_din,
    output wire                                          Module0Func_0_fifo_st_0_full_n,
    input wire                                           Module0Func_0_fifo_st_0_write,
    output wire                                          Module1Func_0_ap_clk,
    input wire                                           Module1Func_0_ap_done,
    input wire                                           Module1Func_0_ap_idle,
    input wire                                           Module1Func_0_ap_ready,
    output wire                                          Module1Func_0_ap_rst_n,
    output wire                                          Module1Func_0_ap_start,
    output wire [                                 512:0] Module1Func_0_fifo_ld_0_peek_dout,
    output wire                                          Module1Func_0_fifo_ld_0_peek_empty_n,
    input wire                                           Module1Func_0_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module1Func_0_fifo_ld_0_s_dout,
    output wire                                          Module1Func_0_fifo_ld_0_s_empty_n,
    input wire                                           Module1Func_0_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module1Func_0_fifo_st_0_din,
    output wire                                          Module1Func_0_fifo_st_0_full_n,
    input wire                                           Module1Func_0_fifo_st_0_write,
    output wire                                          Module2Func_0_ap_clk,
    input wire                                           Module2Func_0_ap_done,
    input wire                                           Module2Func_0_ap_idle,
    input wire                                           Module2Func_0_ap_ready,
    output wire                                          Module2Func_0_ap_rst_n,
    output wire                                          Module2Func_0_ap_start,
    output wire [                                 512:0] Module2Func_0_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_0_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_0_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_0_fifo_ld_0_s_dout,
    output wire                                          Module2Func_0_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_0_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_0_fifo_st_0_din,
    output wire                                          Module2Func_0_fifo_st_0_full_n,
    input wire                                           Module2Func_0_fifo_st_0_write,
    output wire                                          Module2Func_1_ap_clk,
    input wire                                           Module2Func_1_ap_done,
    input wire                                           Module2Func_1_ap_idle,
    input wire                                           Module2Func_1_ap_ready,
    output wire                                          Module2Func_1_ap_rst_n,
    output wire                                          Module2Func_1_ap_start,
    output wire [                                 512:0] Module2Func_1_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_1_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_1_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_1_fifo_ld_0_s_dout,
    output wire                                          Module2Func_1_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_1_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_1_fifo_st_0_din,
    output wire                                          Module2Func_1_fifo_st_0_full_n,
    input wire                                           Module2Func_1_fifo_st_0_write,
    output wire                                          Module2Func_2_ap_clk,
    input wire                                           Module2Func_2_ap_done,
    input wire                                           Module2Func_2_ap_idle,
    input wire                                           Module2Func_2_ap_ready,
    output wire                                          Module2Func_2_ap_rst_n,
    output wire                                          Module2Func_2_ap_start,
    output wire [                                 512:0] Module2Func_2_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_2_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_2_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_2_fifo_ld_0_s_dout,
    output wire                                          Module2Func_2_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_2_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_2_fifo_st_0_din,
    output wire                                          Module2Func_2_fifo_st_0_full_n,
    input wire                                           Module2Func_2_fifo_st_0_write,
    output wire                                          Module2Func_3_ap_clk,
    input wire                                           Module2Func_3_ap_done,
    input wire                                           Module2Func_3_ap_idle,
    input wire                                           Module2Func_3_ap_ready,
    output wire                                          Module2Func_3_ap_rst_n,
    output wire                                          Module2Func_3_ap_start,
    output wire [                                 512:0] Module2Func_3_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_3_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_3_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_3_fifo_ld_0_s_dout,
    output wire                                          Module2Func_3_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_3_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_3_fifo_st_0_din,
    output wire                                          Module2Func_3_fifo_st_0_full_n,
    input wire                                           Module2Func_3_fifo_st_0_write,
    output wire                                          Module2Func_4_ap_clk,
    input wire                                           Module2Func_4_ap_done,
    input wire                                           Module2Func_4_ap_idle,
    input wire                                           Module2Func_4_ap_ready,
    output wire                                          Module2Func_4_ap_rst_n,
    output wire                                          Module2Func_4_ap_start,
    output wire [                                 512:0] Module2Func_4_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_4_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_4_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_4_fifo_ld_0_s_dout,
    output wire                                          Module2Func_4_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_4_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_4_fifo_st_0_din,
    output wire                                          Module2Func_4_fifo_st_0_full_n,
    input wire                                           Module2Func_4_fifo_st_0_write,
    output wire                                          Module2Func_5_ap_clk,
    input wire                                           Module2Func_5_ap_done,
    input wire                                           Module2Func_5_ap_idle,
    input wire                                           Module2Func_5_ap_ready,
    output wire                                          Module2Func_5_ap_rst_n,
    output wire                                          Module2Func_5_ap_start,
    output wire [                                 512:0] Module2Func_5_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_5_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_5_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_5_fifo_ld_0_s_dout,
    output wire                                          Module2Func_5_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_5_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_5_fifo_st_0_din,
    output wire                                          Module2Func_5_fifo_st_0_full_n,
    input wire                                           Module2Func_5_fifo_st_0_write,
    output wire                                          Module2Func_6_ap_clk,
    input wire                                           Module2Func_6_ap_done,
    input wire                                           Module2Func_6_ap_idle,
    input wire                                           Module2Func_6_ap_ready,
    output wire                                          Module2Func_6_ap_rst_n,
    output wire                                          Module2Func_6_ap_start,
    output wire [                                 512:0] Module2Func_6_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_6_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_6_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_6_fifo_ld_0_s_dout,
    output wire                                          Module2Func_6_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_6_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_6_fifo_st_0_din,
    output wire                                          Module2Func_6_fifo_st_0_full_n,
    input wire                                           Module2Func_6_fifo_st_0_write,
    output wire                                          Module2Func_7_ap_clk,
    input wire                                           Module2Func_7_ap_done,
    input wire                                           Module2Func_7_ap_idle,
    input wire                                           Module2Func_7_ap_ready,
    output wire                                          Module2Func_7_ap_rst_n,
    output wire                                          Module2Func_7_ap_start,
    output wire [                                 512:0] Module2Func_7_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_7_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_7_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_7_fifo_ld_0_s_dout,
    output wire                                          Module2Func_7_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_7_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_7_fifo_st_0_din,
    output wire                                          Module2Func_7_fifo_st_0_full_n,
    input wire                                           Module2Func_7_fifo_st_0_write,
    output wire                                          Module2Func_8_ap_clk,
    input wire                                           Module2Func_8_ap_done,
    input wire                                           Module2Func_8_ap_idle,
    input wire                                           Module2Func_8_ap_ready,
    output wire                                          Module2Func_8_ap_rst_n,
    output wire                                          Module2Func_8_ap_start,
    output wire [                                 512:0] Module2Func_8_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_8_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_8_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_8_fifo_ld_0_s_dout,
    output wire                                          Module2Func_8_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_8_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_8_fifo_st_0_din,
    output wire                                          Module2Func_8_fifo_st_0_full_n,
    input wire                                           Module2Func_8_fifo_st_0_write,
    output wire                                          Module2Func_9_ap_clk,
    input wire                                           Module2Func_9_ap_done,
    input wire                                           Module2Func_9_ap_idle,
    input wire                                           Module2Func_9_ap_ready,
    output wire                                          Module2Func_9_ap_rst_n,
    output wire                                          Module2Func_9_ap_start,
    output wire [                                 512:0] Module2Func_9_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_9_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_9_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_9_fifo_ld_0_s_dout,
    output wire                                          Module2Func_9_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_9_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_9_fifo_st_0_din,
    output wire                                          Module2Func_9_fifo_st_0_full_n,
    input wire                                           Module2Func_9_fifo_st_0_write,
    output wire                                          Module2Func_10_ap_clk,
    input wire                                           Module2Func_10_ap_done,
    input wire                                           Module2Func_10_ap_idle,
    input wire                                           Module2Func_10_ap_ready,
    output wire                                          Module2Func_10_ap_rst_n,
    output wire                                          Module2Func_10_ap_start,
    output wire [                                 512:0] Module2Func_10_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_10_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_10_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_10_fifo_ld_0_s_dout,
    output wire                                          Module2Func_10_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_10_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_10_fifo_st_0_din,
    output wire                                          Module2Func_10_fifo_st_0_full_n,
    input wire                                           Module2Func_10_fifo_st_0_write,
    output wire                                          Module2Func_11_ap_clk,
    input wire                                           Module2Func_11_ap_done,
    input wire                                           Module2Func_11_ap_idle,
    input wire                                           Module2Func_11_ap_ready,
    output wire                                          Module2Func_11_ap_rst_n,
    output wire                                          Module2Func_11_ap_start,
    output wire [                                 512:0] Module2Func_11_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_11_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_11_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_11_fifo_ld_0_s_dout,
    output wire                                          Module2Func_11_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_11_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_11_fifo_st_0_din,
    output wire                                          Module2Func_11_fifo_st_0_full_n,
    input wire                                           Module2Func_11_fifo_st_0_write,
    output wire                                          Module2Func_12_ap_clk,
    input wire                                           Module2Func_12_ap_done,
    input wire                                           Module2Func_12_ap_idle,
    input wire                                           Module2Func_12_ap_ready,
    output wire                                          Module2Func_12_ap_rst_n,
    output wire                                          Module2Func_12_ap_start,
    output wire [                                 512:0] Module2Func_12_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_12_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_12_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_12_fifo_ld_0_s_dout,
    output wire                                          Module2Func_12_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_12_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_12_fifo_st_0_din,
    output wire                                          Module2Func_12_fifo_st_0_full_n,
    input wire                                           Module2Func_12_fifo_st_0_write,
    output wire                                          Module2Func_13_ap_clk,
    input wire                                           Module2Func_13_ap_done,
    input wire                                           Module2Func_13_ap_idle,
    input wire                                           Module2Func_13_ap_ready,
    output wire                                          Module2Func_13_ap_rst_n,
    output wire                                          Module2Func_13_ap_start,
    output wire [                                 512:0] Module2Func_13_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_13_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_13_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_13_fifo_ld_0_s_dout,
    output wire                                          Module2Func_13_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_13_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_13_fifo_st_0_din,
    output wire                                          Module2Func_13_fifo_st_0_full_n,
    input wire                                           Module2Func_13_fifo_st_0_write,
    output wire                                          Module2Func_14_ap_clk,
    input wire                                           Module2Func_14_ap_done,
    input wire                                           Module2Func_14_ap_idle,
    input wire                                           Module2Func_14_ap_ready,
    output wire                                          Module2Func_14_ap_rst_n,
    output wire                                          Module2Func_14_ap_start,
    output wire [                                 512:0] Module2Func_14_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_14_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_14_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_14_fifo_ld_0_s_dout,
    output wire                                          Module2Func_14_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_14_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_14_fifo_st_0_din,
    output wire                                          Module2Func_14_fifo_st_0_full_n,
    input wire                                           Module2Func_14_fifo_st_0_write,
    output wire                                          Module2Func_15_ap_clk,
    input wire                                           Module2Func_15_ap_done,
    input wire                                           Module2Func_15_ap_idle,
    input wire                                           Module2Func_15_ap_ready,
    output wire                                          Module2Func_15_ap_rst_n,
    output wire                                          Module2Func_15_ap_start,
    output wire [                                 512:0] Module2Func_15_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_15_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_15_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_15_fifo_ld_0_s_dout,
    output wire                                          Module2Func_15_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_15_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_15_fifo_st_0_din,
    output wire                                          Module2Func_15_fifo_st_0_full_n,
    input wire                                           Module2Func_15_fifo_st_0_write,
    output wire                                          Module2Func_16_ap_clk,
    input wire                                           Module2Func_16_ap_done,
    input wire                                           Module2Func_16_ap_idle,
    input wire                                           Module2Func_16_ap_ready,
    output wire                                          Module2Func_16_ap_rst_n,
    output wire                                          Module2Func_16_ap_start,
    output wire [                                 512:0] Module2Func_16_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_16_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_16_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_16_fifo_ld_0_s_dout,
    output wire                                          Module2Func_16_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_16_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_16_fifo_st_0_din,
    output wire                                          Module2Func_16_fifo_st_0_full_n,
    input wire                                           Module2Func_16_fifo_st_0_write,
    output wire                                          Module2Func_17_ap_clk,
    input wire                                           Module2Func_17_ap_done,
    input wire                                           Module2Func_17_ap_idle,
    input wire                                           Module2Func_17_ap_ready,
    output wire                                          Module2Func_17_ap_rst_n,
    output wire                                          Module2Func_17_ap_start,
    output wire [                                 512:0] Module2Func_17_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_17_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_17_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_17_fifo_ld_0_s_dout,
    output wire                                          Module2Func_17_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_17_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_17_fifo_st_0_din,
    output wire                                          Module2Func_17_fifo_st_0_full_n,
    input wire                                           Module2Func_17_fifo_st_0_write,
    output wire                                          Module2Func_18_ap_clk,
    input wire                                           Module2Func_18_ap_done,
    input wire                                           Module2Func_18_ap_idle,
    input wire                                           Module2Func_18_ap_ready,
    output wire                                          Module2Func_18_ap_rst_n,
    output wire                                          Module2Func_18_ap_start,
    output wire [                                 512:0] Module2Func_18_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_18_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_18_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_18_fifo_ld_0_s_dout,
    output wire                                          Module2Func_18_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_18_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_18_fifo_st_0_din,
    output wire                                          Module2Func_18_fifo_st_0_full_n,
    input wire                                           Module2Func_18_fifo_st_0_write,
    output wire                                          Module2Func_19_ap_clk,
    input wire                                           Module2Func_19_ap_done,
    input wire                                           Module2Func_19_ap_idle,
    input wire                                           Module2Func_19_ap_ready,
    output wire                                          Module2Func_19_ap_rst_n,
    output wire                                          Module2Func_19_ap_start,
    output wire [                                 512:0] Module2Func_19_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_19_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_19_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_19_fifo_ld_0_s_dout,
    output wire                                          Module2Func_19_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_19_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_19_fifo_st_0_din,
    output wire                                          Module2Func_19_fifo_st_0_full_n,
    input wire                                           Module2Func_19_fifo_st_0_write,
    output wire                                          Module2Func_20_ap_clk,
    input wire                                           Module2Func_20_ap_done,
    input wire                                           Module2Func_20_ap_idle,
    input wire                                           Module2Func_20_ap_ready,
    output wire                                          Module2Func_20_ap_rst_n,
    output wire                                          Module2Func_20_ap_start,
    output wire [                                 512:0] Module2Func_20_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_20_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_20_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_20_fifo_ld_0_s_dout,
    output wire                                          Module2Func_20_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_20_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_20_fifo_st_0_din,
    output wire                                          Module2Func_20_fifo_st_0_full_n,
    input wire                                           Module2Func_20_fifo_st_0_write,
    output wire                                          Module2Func_21_ap_clk,
    input wire                                           Module2Func_21_ap_done,
    input wire                                           Module2Func_21_ap_idle,
    input wire                                           Module2Func_21_ap_ready,
    output wire                                          Module2Func_21_ap_rst_n,
    output wire                                          Module2Func_21_ap_start,
    output wire [                                 512:0] Module2Func_21_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_21_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_21_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_21_fifo_ld_0_s_dout,
    output wire                                          Module2Func_21_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_21_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_21_fifo_st_0_din,
    output wire                                          Module2Func_21_fifo_st_0_full_n,
    input wire                                           Module2Func_21_fifo_st_0_write,
    output wire                                          Module2Func_22_ap_clk,
    input wire                                           Module2Func_22_ap_done,
    input wire                                           Module2Func_22_ap_idle,
    input wire                                           Module2Func_22_ap_ready,
    output wire                                          Module2Func_22_ap_rst_n,
    output wire                                          Module2Func_22_ap_start,
    output wire [                                 512:0] Module2Func_22_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_22_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_22_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_22_fifo_ld_0_s_dout,
    output wire                                          Module2Func_22_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_22_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_22_fifo_st_0_din,
    output wire                                          Module2Func_22_fifo_st_0_full_n,
    input wire                                           Module2Func_22_fifo_st_0_write,
    output wire                                          Module2Func_23_ap_clk,
    input wire                                           Module2Func_23_ap_done,
    input wire                                           Module2Func_23_ap_idle,
    input wire                                           Module2Func_23_ap_ready,
    output wire                                          Module2Func_23_ap_rst_n,
    output wire                                          Module2Func_23_ap_start,
    output wire [                                 512:0] Module2Func_23_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_23_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_23_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_23_fifo_ld_0_s_dout,
    output wire                                          Module2Func_23_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_23_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_23_fifo_st_0_din,
    output wire                                          Module2Func_23_fifo_st_0_full_n,
    input wire                                           Module2Func_23_fifo_st_0_write,
    output wire                                          Module2Func_24_ap_clk,
    input wire                                           Module2Func_24_ap_done,
    input wire                                           Module2Func_24_ap_idle,
    input wire                                           Module2Func_24_ap_ready,
    output wire                                          Module2Func_24_ap_rst_n,
    output wire                                          Module2Func_24_ap_start,
    output wire [                                 512:0] Module2Func_24_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_24_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_24_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_24_fifo_ld_0_s_dout,
    output wire                                          Module2Func_24_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_24_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_24_fifo_st_0_din,
    output wire                                          Module2Func_24_fifo_st_0_full_n,
    input wire                                           Module2Func_24_fifo_st_0_write,
    output wire                                          Module2Func_25_ap_clk,
    input wire                                           Module2Func_25_ap_done,
    input wire                                           Module2Func_25_ap_idle,
    input wire                                           Module2Func_25_ap_ready,
    output wire                                          Module2Func_25_ap_rst_n,
    output wire                                          Module2Func_25_ap_start,
    output wire [                                 512:0] Module2Func_25_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_25_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_25_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_25_fifo_ld_0_s_dout,
    output wire                                          Module2Func_25_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_25_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_25_fifo_st_0_din,
    output wire                                          Module2Func_25_fifo_st_0_full_n,
    input wire                                           Module2Func_25_fifo_st_0_write,
    output wire                                          Module2Func_26_ap_clk,
    input wire                                           Module2Func_26_ap_done,
    input wire                                           Module2Func_26_ap_idle,
    input wire                                           Module2Func_26_ap_ready,
    output wire                                          Module2Func_26_ap_rst_n,
    output wire                                          Module2Func_26_ap_start,
    output wire [                                 512:0] Module2Func_26_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_26_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_26_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_26_fifo_ld_0_s_dout,
    output wire                                          Module2Func_26_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_26_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_26_fifo_st_0_din,
    output wire                                          Module2Func_26_fifo_st_0_full_n,
    input wire                                           Module2Func_26_fifo_st_0_write,
    output wire                                          Module2Func_27_ap_clk,
    input wire                                           Module2Func_27_ap_done,
    input wire                                           Module2Func_27_ap_idle,
    input wire                                           Module2Func_27_ap_ready,
    output wire                                          Module2Func_27_ap_rst_n,
    output wire                                          Module2Func_27_ap_start,
    output wire [                                 512:0] Module2Func_27_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_27_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_27_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_27_fifo_ld_0_s_dout,
    output wire                                          Module2Func_27_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_27_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_27_fifo_st_0_din,
    output wire                                          Module2Func_27_fifo_st_0_full_n,
    input wire                                           Module2Func_27_fifo_st_0_write,
    output wire                                          Module2Func_28_ap_clk,
    input wire                                           Module2Func_28_ap_done,
    input wire                                           Module2Func_28_ap_idle,
    input wire                                           Module2Func_28_ap_ready,
    output wire                                          Module2Func_28_ap_rst_n,
    output wire                                          Module2Func_28_ap_start,
    output wire [                                 512:0] Module2Func_28_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_28_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_28_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_28_fifo_ld_0_s_dout,
    output wire                                          Module2Func_28_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_28_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_28_fifo_st_0_din,
    output wire                                          Module2Func_28_fifo_st_0_full_n,
    input wire                                           Module2Func_28_fifo_st_0_write,
    output wire                                          Module2Func_29_ap_clk,
    input wire                                           Module2Func_29_ap_done,
    input wire                                           Module2Func_29_ap_idle,
    input wire                                           Module2Func_29_ap_ready,
    output wire                                          Module2Func_29_ap_rst_n,
    output wire                                          Module2Func_29_ap_start,
    output wire [                                 512:0] Module2Func_29_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_29_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_29_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_29_fifo_ld_0_s_dout,
    output wire                                          Module2Func_29_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_29_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_29_fifo_st_0_din,
    output wire                                          Module2Func_29_fifo_st_0_full_n,
    input wire                                           Module2Func_29_fifo_st_0_write,
    output wire                                          Module2Func_30_ap_clk,
    input wire                                           Module2Func_30_ap_done,
    input wire                                           Module2Func_30_ap_idle,
    input wire                                           Module2Func_30_ap_ready,
    output wire                                          Module2Func_30_ap_rst_n,
    output wire                                          Module2Func_30_ap_start,
    output wire [                                 512:0] Module2Func_30_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_30_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_30_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_30_fifo_ld_0_s_dout,
    output wire                                          Module2Func_30_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_30_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_30_fifo_st_0_din,
    output wire                                          Module2Func_30_fifo_st_0_full_n,
    input wire                                           Module2Func_30_fifo_st_0_write,
    output wire                                          Module2Func_31_ap_clk,
    input wire                                           Module2Func_31_ap_done,
    input wire                                           Module2Func_31_ap_idle,
    input wire                                           Module2Func_31_ap_ready,
    output wire                                          Module2Func_31_ap_rst_n,
    output wire                                          Module2Func_31_ap_start,
    output wire [                                 512:0] Module2Func_31_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_31_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_31_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_31_fifo_ld_0_s_dout,
    output wire                                          Module2Func_31_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_31_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_31_fifo_st_0_din,
    output wire                                          Module2Func_31_fifo_st_0_full_n,
    input wire                                           Module2Func_31_fifo_st_0_write,
    output wire                                          Module2Func_32_ap_clk,
    input wire                                           Module2Func_32_ap_done,
    input wire                                           Module2Func_32_ap_idle,
    input wire                                           Module2Func_32_ap_ready,
    output wire                                          Module2Func_32_ap_rst_n,
    output wire                                          Module2Func_32_ap_start,
    output wire [                                 512:0] Module2Func_32_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_32_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_32_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_32_fifo_ld_0_s_dout,
    output wire                                          Module2Func_32_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_32_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_32_fifo_st_0_din,
    output wire                                          Module2Func_32_fifo_st_0_full_n,
    input wire                                           Module2Func_32_fifo_st_0_write,
    output wire                                          Module2Func_33_ap_clk,
    input wire                                           Module2Func_33_ap_done,
    input wire                                           Module2Func_33_ap_idle,
    input wire                                           Module2Func_33_ap_ready,
    output wire                                          Module2Func_33_ap_rst_n,
    output wire                                          Module2Func_33_ap_start,
    output wire [                                 512:0] Module2Func_33_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_33_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_33_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_33_fifo_ld_0_s_dout,
    output wire                                          Module2Func_33_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_33_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_33_fifo_st_0_din,
    output wire                                          Module2Func_33_fifo_st_0_full_n,
    input wire                                           Module2Func_33_fifo_st_0_write,
    output wire                                          Module2Func_34_ap_clk,
    input wire                                           Module2Func_34_ap_done,
    input wire                                           Module2Func_34_ap_idle,
    input wire                                           Module2Func_34_ap_ready,
    output wire                                          Module2Func_34_ap_rst_n,
    output wire                                          Module2Func_34_ap_start,
    output wire [                                 512:0] Module2Func_34_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_34_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_34_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_34_fifo_ld_0_s_dout,
    output wire                                          Module2Func_34_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_34_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_34_fifo_st_0_din,
    output wire                                          Module2Func_34_fifo_st_0_full_n,
    input wire                                           Module2Func_34_fifo_st_0_write,
    output wire                                          Module2Func_35_ap_clk,
    input wire                                           Module2Func_35_ap_done,
    input wire                                           Module2Func_35_ap_idle,
    input wire                                           Module2Func_35_ap_ready,
    output wire                                          Module2Func_35_ap_rst_n,
    output wire                                          Module2Func_35_ap_start,
    output wire [                                 512:0] Module2Func_35_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_35_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_35_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_35_fifo_ld_0_s_dout,
    output wire                                          Module2Func_35_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_35_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_35_fifo_st_0_din,
    output wire                                          Module2Func_35_fifo_st_0_full_n,
    input wire                                           Module2Func_35_fifo_st_0_write,
    output wire                                          Module2Func_36_ap_clk,
    input wire                                           Module2Func_36_ap_done,
    input wire                                           Module2Func_36_ap_idle,
    input wire                                           Module2Func_36_ap_ready,
    output wire                                          Module2Func_36_ap_rst_n,
    output wire                                          Module2Func_36_ap_start,
    output wire [                                 512:0] Module2Func_36_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_36_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_36_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_36_fifo_ld_0_s_dout,
    output wire                                          Module2Func_36_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_36_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_36_fifo_st_0_din,
    output wire                                          Module2Func_36_fifo_st_0_full_n,
    input wire                                           Module2Func_36_fifo_st_0_write,
    output wire                                          Module2Func_37_ap_clk,
    input wire                                           Module2Func_37_ap_done,
    input wire                                           Module2Func_37_ap_idle,
    input wire                                           Module2Func_37_ap_ready,
    output wire                                          Module2Func_37_ap_rst_n,
    output wire                                          Module2Func_37_ap_start,
    output wire [                                 512:0] Module2Func_37_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_37_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_37_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_37_fifo_ld_0_s_dout,
    output wire                                          Module2Func_37_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_37_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_37_fifo_st_0_din,
    output wire                                          Module2Func_37_fifo_st_0_full_n,
    input wire                                           Module2Func_37_fifo_st_0_write,
    output wire                                          Module2Func_38_ap_clk,
    input wire                                           Module2Func_38_ap_done,
    input wire                                           Module2Func_38_ap_idle,
    input wire                                           Module2Func_38_ap_ready,
    output wire                                          Module2Func_38_ap_rst_n,
    output wire                                          Module2Func_38_ap_start,
    output wire [                                 512:0] Module2Func_38_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_38_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_38_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_38_fifo_ld_0_s_dout,
    output wire                                          Module2Func_38_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_38_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_38_fifo_st_0_din,
    output wire                                          Module2Func_38_fifo_st_0_full_n,
    input wire                                           Module2Func_38_fifo_st_0_write,
    output wire                                          Module2Func_39_ap_clk,
    input wire                                           Module2Func_39_ap_done,
    input wire                                           Module2Func_39_ap_idle,
    input wire                                           Module2Func_39_ap_ready,
    output wire                                          Module2Func_39_ap_rst_n,
    output wire                                          Module2Func_39_ap_start,
    output wire [                                 512:0] Module2Func_39_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_39_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_39_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_39_fifo_ld_0_s_dout,
    output wire                                          Module2Func_39_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_39_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_39_fifo_st_0_din,
    output wire                                          Module2Func_39_fifo_st_0_full_n,
    input wire                                           Module2Func_39_fifo_st_0_write,
    output wire                                          Module2Func_40_ap_clk,
    input wire                                           Module2Func_40_ap_done,
    input wire                                           Module2Func_40_ap_idle,
    input wire                                           Module2Func_40_ap_ready,
    output wire                                          Module2Func_40_ap_rst_n,
    output wire                                          Module2Func_40_ap_start,
    output wire [                                 512:0] Module2Func_40_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_40_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_40_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_40_fifo_ld_0_s_dout,
    output wire                                          Module2Func_40_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_40_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_40_fifo_st_0_din,
    output wire                                          Module2Func_40_fifo_st_0_full_n,
    input wire                                           Module2Func_40_fifo_st_0_write,
    output wire                                          Module2Func_41_ap_clk,
    input wire                                           Module2Func_41_ap_done,
    input wire                                           Module2Func_41_ap_idle,
    input wire                                           Module2Func_41_ap_ready,
    output wire                                          Module2Func_41_ap_rst_n,
    output wire                                          Module2Func_41_ap_start,
    output wire [                                 512:0] Module2Func_41_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_41_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_41_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_41_fifo_ld_0_s_dout,
    output wire                                          Module2Func_41_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_41_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_41_fifo_st_0_din,
    output wire                                          Module2Func_41_fifo_st_0_full_n,
    input wire                                           Module2Func_41_fifo_st_0_write,
    output wire                                          Module2Func_42_ap_clk,
    input wire                                           Module2Func_42_ap_done,
    input wire                                           Module2Func_42_ap_idle,
    input wire                                           Module2Func_42_ap_ready,
    output wire                                          Module2Func_42_ap_rst_n,
    output wire                                          Module2Func_42_ap_start,
    output wire [                                 512:0] Module2Func_42_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_42_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_42_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_42_fifo_ld_0_s_dout,
    output wire                                          Module2Func_42_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_42_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_42_fifo_st_0_din,
    output wire                                          Module2Func_42_fifo_st_0_full_n,
    input wire                                           Module2Func_42_fifo_st_0_write,
    output wire                                          Module2Func_43_ap_clk,
    input wire                                           Module2Func_43_ap_done,
    input wire                                           Module2Func_43_ap_idle,
    input wire                                           Module2Func_43_ap_ready,
    output wire                                          Module2Func_43_ap_rst_n,
    output wire                                          Module2Func_43_ap_start,
    output wire [                                 512:0] Module2Func_43_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_43_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_43_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_43_fifo_ld_0_s_dout,
    output wire                                          Module2Func_43_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_43_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_43_fifo_st_0_din,
    output wire                                          Module2Func_43_fifo_st_0_full_n,
    input wire                                           Module2Func_43_fifo_st_0_write,
    output wire                                          Module2Func_44_ap_clk,
    input wire                                           Module2Func_44_ap_done,
    input wire                                           Module2Func_44_ap_idle,
    input wire                                           Module2Func_44_ap_ready,
    output wire                                          Module2Func_44_ap_rst_n,
    output wire                                          Module2Func_44_ap_start,
    output wire [                                 512:0] Module2Func_44_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_44_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_44_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_44_fifo_ld_0_s_dout,
    output wire                                          Module2Func_44_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_44_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_44_fifo_st_0_din,
    output wire                                          Module2Func_44_fifo_st_0_full_n,
    input wire                                           Module2Func_44_fifo_st_0_write,
    output wire                                          Module2Func_45_ap_clk,
    input wire                                           Module2Func_45_ap_done,
    input wire                                           Module2Func_45_ap_idle,
    input wire                                           Module2Func_45_ap_ready,
    output wire                                          Module2Func_45_ap_rst_n,
    output wire                                          Module2Func_45_ap_start,
    output wire [                                 512:0] Module2Func_45_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_45_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_45_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_45_fifo_ld_0_s_dout,
    output wire                                          Module2Func_45_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_45_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_45_fifo_st_0_din,
    output wire                                          Module2Func_45_fifo_st_0_full_n,
    input wire                                           Module2Func_45_fifo_st_0_write,
    output wire                                          Module2Func_46_ap_clk,
    input wire                                           Module2Func_46_ap_done,
    input wire                                           Module2Func_46_ap_idle,
    input wire                                           Module2Func_46_ap_ready,
    output wire                                          Module2Func_46_ap_rst_n,
    output wire                                          Module2Func_46_ap_start,
    output wire [                                 512:0] Module2Func_46_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_46_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_46_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_46_fifo_ld_0_s_dout,
    output wire                                          Module2Func_46_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_46_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_46_fifo_st_0_din,
    output wire                                          Module2Func_46_fifo_st_0_full_n,
    input wire                                           Module2Func_46_fifo_st_0_write,
    output wire                                          Module2Func_47_ap_clk,
    input wire                                           Module2Func_47_ap_done,
    input wire                                           Module2Func_47_ap_idle,
    input wire                                           Module2Func_47_ap_ready,
    output wire                                          Module2Func_47_ap_rst_n,
    output wire                                          Module2Func_47_ap_start,
    output wire [                                 512:0] Module2Func_47_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_47_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_47_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_47_fifo_ld_0_s_dout,
    output wire                                          Module2Func_47_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_47_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_47_fifo_st_0_din,
    output wire                                          Module2Func_47_fifo_st_0_full_n,
    input wire                                           Module2Func_47_fifo_st_0_write,
    output wire                                          Module2Func_48_ap_clk,
    input wire                                           Module2Func_48_ap_done,
    input wire                                           Module2Func_48_ap_idle,
    input wire                                           Module2Func_48_ap_ready,
    output wire                                          Module2Func_48_ap_rst_n,
    output wire                                          Module2Func_48_ap_start,
    output wire [                                 512:0] Module2Func_48_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_48_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_48_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_48_fifo_ld_0_s_dout,
    output wire                                          Module2Func_48_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_48_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_48_fifo_st_0_din,
    output wire                                          Module2Func_48_fifo_st_0_full_n,
    input wire                                           Module2Func_48_fifo_st_0_write,
    output wire                                          Module2Func_49_ap_clk,
    input wire                                           Module2Func_49_ap_done,
    input wire                                           Module2Func_49_ap_idle,
    input wire                                           Module2Func_49_ap_ready,
    output wire                                          Module2Func_49_ap_rst_n,
    output wire                                          Module2Func_49_ap_start,
    output wire [                                 512:0] Module2Func_49_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_49_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_49_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_49_fifo_ld_0_s_dout,
    output wire                                          Module2Func_49_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_49_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_49_fifo_st_0_din,
    output wire                                          Module2Func_49_fifo_st_0_full_n,
    input wire                                           Module2Func_49_fifo_st_0_write,
    output wire                                          Module2Func_50_ap_clk,
    input wire                                           Module2Func_50_ap_done,
    input wire                                           Module2Func_50_ap_idle,
    input wire                                           Module2Func_50_ap_ready,
    output wire                                          Module2Func_50_ap_rst_n,
    output wire                                          Module2Func_50_ap_start,
    output wire [                                 512:0] Module2Func_50_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_50_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_50_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_50_fifo_ld_0_s_dout,
    output wire                                          Module2Func_50_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_50_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_50_fifo_st_0_din,
    output wire                                          Module2Func_50_fifo_st_0_full_n,
    input wire                                           Module2Func_50_fifo_st_0_write,
    output wire                                          Module2Func_51_ap_clk,
    input wire                                           Module2Func_51_ap_done,
    input wire                                           Module2Func_51_ap_idle,
    input wire                                           Module2Func_51_ap_ready,
    output wire                                          Module2Func_51_ap_rst_n,
    output wire                                          Module2Func_51_ap_start,
    output wire [                                 512:0] Module2Func_51_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_51_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_51_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_51_fifo_ld_0_s_dout,
    output wire                                          Module2Func_51_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_51_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_51_fifo_st_0_din,
    output wire                                          Module2Func_51_fifo_st_0_full_n,
    input wire                                           Module2Func_51_fifo_st_0_write,
    output wire                                          Module2Func_52_ap_clk,
    input wire                                           Module2Func_52_ap_done,
    input wire                                           Module2Func_52_ap_idle,
    input wire                                           Module2Func_52_ap_ready,
    output wire                                          Module2Func_52_ap_rst_n,
    output wire                                          Module2Func_52_ap_start,
    output wire [                                 512:0] Module2Func_52_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_52_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_52_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_52_fifo_ld_0_s_dout,
    output wire                                          Module2Func_52_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_52_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_52_fifo_st_0_din,
    output wire                                          Module2Func_52_fifo_st_0_full_n,
    input wire                                           Module2Func_52_fifo_st_0_write,
    output wire                                          Module2Func_53_ap_clk,
    input wire                                           Module2Func_53_ap_done,
    input wire                                           Module2Func_53_ap_idle,
    input wire                                           Module2Func_53_ap_ready,
    output wire                                          Module2Func_53_ap_rst_n,
    output wire                                          Module2Func_53_ap_start,
    output wire [                                 512:0] Module2Func_53_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_53_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_53_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_53_fifo_ld_0_s_dout,
    output wire                                          Module2Func_53_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_53_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_53_fifo_st_0_din,
    output wire                                          Module2Func_53_fifo_st_0_full_n,
    input wire                                           Module2Func_53_fifo_st_0_write,
    output wire                                          Module2Func_54_ap_clk,
    input wire                                           Module2Func_54_ap_done,
    input wire                                           Module2Func_54_ap_idle,
    input wire                                           Module2Func_54_ap_ready,
    output wire                                          Module2Func_54_ap_rst_n,
    output wire                                          Module2Func_54_ap_start,
    output wire [                                 512:0] Module2Func_54_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_54_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_54_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_54_fifo_ld_0_s_dout,
    output wire                                          Module2Func_54_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_54_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_54_fifo_st_0_din,
    output wire                                          Module2Func_54_fifo_st_0_full_n,
    input wire                                           Module2Func_54_fifo_st_0_write,
    output wire                                          Module2Func_55_ap_clk,
    input wire                                           Module2Func_55_ap_done,
    input wire                                           Module2Func_55_ap_idle,
    input wire                                           Module2Func_55_ap_ready,
    output wire                                          Module2Func_55_ap_rst_n,
    output wire                                          Module2Func_55_ap_start,
    output wire [                                 512:0] Module2Func_55_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_55_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_55_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_55_fifo_ld_0_s_dout,
    output wire                                          Module2Func_55_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_55_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_55_fifo_st_0_din,
    output wire                                          Module2Func_55_fifo_st_0_full_n,
    input wire                                           Module2Func_55_fifo_st_0_write,
    output wire                                          Module2Func_56_ap_clk,
    input wire                                           Module2Func_56_ap_done,
    input wire                                           Module2Func_56_ap_idle,
    input wire                                           Module2Func_56_ap_ready,
    output wire                                          Module2Func_56_ap_rst_n,
    output wire                                          Module2Func_56_ap_start,
    output wire [                                 512:0] Module2Func_56_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_56_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_56_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_56_fifo_ld_0_s_dout,
    output wire                                          Module2Func_56_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_56_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_56_fifo_st_0_din,
    output wire                                          Module2Func_56_fifo_st_0_full_n,
    input wire                                           Module2Func_56_fifo_st_0_write,
    output wire                                          Module2Func_57_ap_clk,
    input wire                                           Module2Func_57_ap_done,
    input wire                                           Module2Func_57_ap_idle,
    input wire                                           Module2Func_57_ap_ready,
    output wire                                          Module2Func_57_ap_rst_n,
    output wire                                          Module2Func_57_ap_start,
    output wire [                                 512:0] Module2Func_57_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_57_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_57_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_57_fifo_ld_0_s_dout,
    output wire                                          Module2Func_57_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_57_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_57_fifo_st_0_din,
    output wire                                          Module2Func_57_fifo_st_0_full_n,
    input wire                                           Module2Func_57_fifo_st_0_write,
    output wire                                          Module2Func_58_ap_clk,
    input wire                                           Module2Func_58_ap_done,
    input wire                                           Module2Func_58_ap_idle,
    input wire                                           Module2Func_58_ap_ready,
    output wire                                          Module2Func_58_ap_rst_n,
    output wire                                          Module2Func_58_ap_start,
    output wire [                                 512:0] Module2Func_58_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_58_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_58_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_58_fifo_ld_0_s_dout,
    output wire                                          Module2Func_58_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_58_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_58_fifo_st_0_din,
    output wire                                          Module2Func_58_fifo_st_0_full_n,
    input wire                                           Module2Func_58_fifo_st_0_write,
    output wire                                          Module2Func_59_ap_clk,
    input wire                                           Module2Func_59_ap_done,
    input wire                                           Module2Func_59_ap_idle,
    input wire                                           Module2Func_59_ap_ready,
    output wire                                          Module2Func_59_ap_rst_n,
    output wire                                          Module2Func_59_ap_start,
    output wire [                                 512:0] Module2Func_59_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_59_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_59_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_59_fifo_ld_0_s_dout,
    output wire                                          Module2Func_59_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_59_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_59_fifo_st_0_din,
    output wire                                          Module2Func_59_fifo_st_0_full_n,
    input wire                                           Module2Func_59_fifo_st_0_write,
    output wire                                          Module2Func_60_ap_clk,
    input wire                                           Module2Func_60_ap_done,
    input wire                                           Module2Func_60_ap_idle,
    input wire                                           Module2Func_60_ap_ready,
    output wire                                          Module2Func_60_ap_rst_n,
    output wire                                          Module2Func_60_ap_start,
    output wire [                                 512:0] Module2Func_60_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_60_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_60_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_60_fifo_ld_0_s_dout,
    output wire                                          Module2Func_60_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_60_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_60_fifo_st_0_din,
    output wire                                          Module2Func_60_fifo_st_0_full_n,
    input wire                                           Module2Func_60_fifo_st_0_write,
    output wire                                          Module2Func_61_ap_clk,
    input wire                                           Module2Func_61_ap_done,
    input wire                                           Module2Func_61_ap_idle,
    input wire                                           Module2Func_61_ap_ready,
    output wire                                          Module2Func_61_ap_rst_n,
    output wire                                          Module2Func_61_ap_start,
    output wire [                                 512:0] Module2Func_61_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_61_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_61_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_61_fifo_ld_0_s_dout,
    output wire                                          Module2Func_61_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_61_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_61_fifo_st_0_din,
    output wire                                          Module2Func_61_fifo_st_0_full_n,
    input wire                                           Module2Func_61_fifo_st_0_write,
    output wire                                          Module2Func_62_ap_clk,
    input wire                                           Module2Func_62_ap_done,
    input wire                                           Module2Func_62_ap_idle,
    input wire                                           Module2Func_62_ap_ready,
    output wire                                          Module2Func_62_ap_rst_n,
    output wire                                          Module2Func_62_ap_start,
    output wire [                                 512:0] Module2Func_62_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_62_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_62_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_62_fifo_ld_0_s_dout,
    output wire                                          Module2Func_62_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_62_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_62_fifo_st_0_din,
    output wire                                          Module2Func_62_fifo_st_0_full_n,
    input wire                                           Module2Func_62_fifo_st_0_write,
    output wire                                          Module2Func_63_ap_clk,
    input wire                                           Module2Func_63_ap_done,
    input wire                                           Module2Func_63_ap_idle,
    input wire                                           Module2Func_63_ap_ready,
    output wire                                          Module2Func_63_ap_rst_n,
    output wire                                          Module2Func_63_ap_start,
    output wire [                                 512:0] Module2Func_63_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_63_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_63_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_63_fifo_ld_0_s_dout,
    output wire                                          Module2Func_63_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_63_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_63_fifo_st_0_din,
    output wire                                          Module2Func_63_fifo_st_0_full_n,
    input wire                                           Module2Func_63_fifo_st_0_write,
    output wire                                          Module2Func_64_ap_clk,
    input wire                                           Module2Func_64_ap_done,
    input wire                                           Module2Func_64_ap_idle,
    input wire                                           Module2Func_64_ap_ready,
    output wire                                          Module2Func_64_ap_rst_n,
    output wire                                          Module2Func_64_ap_start,
    output wire [                                 512:0] Module2Func_64_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_64_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_64_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_64_fifo_ld_0_s_dout,
    output wire                                          Module2Func_64_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_64_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_64_fifo_st_0_din,
    output wire                                          Module2Func_64_fifo_st_0_full_n,
    input wire                                           Module2Func_64_fifo_st_0_write,
    output wire                                          Module2Func_65_ap_clk,
    input wire                                           Module2Func_65_ap_done,
    input wire                                           Module2Func_65_ap_idle,
    input wire                                           Module2Func_65_ap_ready,
    output wire                                          Module2Func_65_ap_rst_n,
    output wire                                          Module2Func_65_ap_start,
    output wire [                                 512:0] Module2Func_65_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_65_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_65_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_65_fifo_ld_0_s_dout,
    output wire                                          Module2Func_65_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_65_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_65_fifo_st_0_din,
    output wire                                          Module2Func_65_fifo_st_0_full_n,
    input wire                                           Module2Func_65_fifo_st_0_write,
    output wire                                          Module2Func_66_ap_clk,
    input wire                                           Module2Func_66_ap_done,
    input wire                                           Module2Func_66_ap_idle,
    input wire                                           Module2Func_66_ap_ready,
    output wire                                          Module2Func_66_ap_rst_n,
    output wire                                          Module2Func_66_ap_start,
    output wire [                                 512:0] Module2Func_66_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_66_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_66_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_66_fifo_ld_0_s_dout,
    output wire                                          Module2Func_66_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_66_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_66_fifo_st_0_din,
    output wire                                          Module2Func_66_fifo_st_0_full_n,
    input wire                                           Module2Func_66_fifo_st_0_write,
    output wire                                          Module2Func_67_ap_clk,
    input wire                                           Module2Func_67_ap_done,
    input wire                                           Module2Func_67_ap_idle,
    input wire                                           Module2Func_67_ap_ready,
    output wire                                          Module2Func_67_ap_rst_n,
    output wire                                          Module2Func_67_ap_start,
    output wire [                                 512:0] Module2Func_67_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_67_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_67_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_67_fifo_ld_0_s_dout,
    output wire                                          Module2Func_67_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_67_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_67_fifo_st_0_din,
    output wire                                          Module2Func_67_fifo_st_0_full_n,
    input wire                                           Module2Func_67_fifo_st_0_write,
    output wire                                          Module2Func_68_ap_clk,
    input wire                                           Module2Func_68_ap_done,
    input wire                                           Module2Func_68_ap_idle,
    input wire                                           Module2Func_68_ap_ready,
    output wire                                          Module2Func_68_ap_rst_n,
    output wire                                          Module2Func_68_ap_start,
    output wire [                                 512:0] Module2Func_68_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_68_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_68_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_68_fifo_ld_0_s_dout,
    output wire                                          Module2Func_68_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_68_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_68_fifo_st_0_din,
    output wire                                          Module2Func_68_fifo_st_0_full_n,
    input wire                                           Module2Func_68_fifo_st_0_write,
    output wire                                          Module2Func_69_ap_clk,
    input wire                                           Module2Func_69_ap_done,
    input wire                                           Module2Func_69_ap_idle,
    input wire                                           Module2Func_69_ap_ready,
    output wire                                          Module2Func_69_ap_rst_n,
    output wire                                          Module2Func_69_ap_start,
    output wire [                                 512:0] Module2Func_69_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_69_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_69_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_69_fifo_ld_0_s_dout,
    output wire                                          Module2Func_69_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_69_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_69_fifo_st_0_din,
    output wire                                          Module2Func_69_fifo_st_0_full_n,
    input wire                                           Module2Func_69_fifo_st_0_write,
    output wire                                          Module2Func_70_ap_clk,
    input wire                                           Module2Func_70_ap_done,
    input wire                                           Module2Func_70_ap_idle,
    input wire                                           Module2Func_70_ap_ready,
    output wire                                          Module2Func_70_ap_rst_n,
    output wire                                          Module2Func_70_ap_start,
    output wire [                                 512:0] Module2Func_70_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_70_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_70_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_70_fifo_ld_0_s_dout,
    output wire                                          Module2Func_70_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_70_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_70_fifo_st_0_din,
    output wire                                          Module2Func_70_fifo_st_0_full_n,
    input wire                                           Module2Func_70_fifo_st_0_write,
    output wire                                          Module2Func_71_ap_clk,
    input wire                                           Module2Func_71_ap_done,
    input wire                                           Module2Func_71_ap_idle,
    input wire                                           Module2Func_71_ap_ready,
    output wire                                          Module2Func_71_ap_rst_n,
    output wire                                          Module2Func_71_ap_start,
    output wire [                                 512:0] Module2Func_71_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_71_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_71_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_71_fifo_ld_0_s_dout,
    output wire                                          Module2Func_71_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_71_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_71_fifo_st_0_din,
    output wire                                          Module2Func_71_fifo_st_0_full_n,
    input wire                                           Module2Func_71_fifo_st_0_write,
    output wire                                          Module2Func_72_ap_clk,
    input wire                                           Module2Func_72_ap_done,
    input wire                                           Module2Func_72_ap_idle,
    input wire                                           Module2Func_72_ap_ready,
    output wire                                          Module2Func_72_ap_rst_n,
    output wire                                          Module2Func_72_ap_start,
    output wire [                                 512:0] Module2Func_72_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_72_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_72_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_72_fifo_ld_0_s_dout,
    output wire                                          Module2Func_72_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_72_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_72_fifo_st_0_din,
    output wire                                          Module2Func_72_fifo_st_0_full_n,
    input wire                                           Module2Func_72_fifo_st_0_write,
    output wire                                          Module2Func_73_ap_clk,
    input wire                                           Module2Func_73_ap_done,
    input wire                                           Module2Func_73_ap_idle,
    input wire                                           Module2Func_73_ap_ready,
    output wire                                          Module2Func_73_ap_rst_n,
    output wire                                          Module2Func_73_ap_start,
    output wire [                                 512:0] Module2Func_73_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_73_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_73_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_73_fifo_ld_0_s_dout,
    output wire                                          Module2Func_73_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_73_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_73_fifo_st_0_din,
    output wire                                          Module2Func_73_fifo_st_0_full_n,
    input wire                                           Module2Func_73_fifo_st_0_write,
    output wire                                          Module2Func_74_ap_clk,
    input wire                                           Module2Func_74_ap_done,
    input wire                                           Module2Func_74_ap_idle,
    input wire                                           Module2Func_74_ap_ready,
    output wire                                          Module2Func_74_ap_rst_n,
    output wire                                          Module2Func_74_ap_start,
    output wire [                                 512:0] Module2Func_74_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_74_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_74_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_74_fifo_ld_0_s_dout,
    output wire                                          Module2Func_74_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_74_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_74_fifo_st_0_din,
    output wire                                          Module2Func_74_fifo_st_0_full_n,
    input wire                                           Module2Func_74_fifo_st_0_write,
    output wire                                          Module2Func_75_ap_clk,
    input wire                                           Module2Func_75_ap_done,
    input wire                                           Module2Func_75_ap_idle,
    input wire                                           Module2Func_75_ap_ready,
    output wire                                          Module2Func_75_ap_rst_n,
    output wire                                          Module2Func_75_ap_start,
    output wire [                                 512:0] Module2Func_75_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_75_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_75_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_75_fifo_ld_0_s_dout,
    output wire                                          Module2Func_75_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_75_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_75_fifo_st_0_din,
    output wire                                          Module2Func_75_fifo_st_0_full_n,
    input wire                                           Module2Func_75_fifo_st_0_write,
    output wire                                          Module2Func_76_ap_clk,
    input wire                                           Module2Func_76_ap_done,
    input wire                                           Module2Func_76_ap_idle,
    input wire                                           Module2Func_76_ap_ready,
    output wire                                          Module2Func_76_ap_rst_n,
    output wire                                          Module2Func_76_ap_start,
    output wire [                                 512:0] Module2Func_76_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_76_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_76_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_76_fifo_ld_0_s_dout,
    output wire                                          Module2Func_76_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_76_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_76_fifo_st_0_din,
    output wire                                          Module2Func_76_fifo_st_0_full_n,
    input wire                                           Module2Func_76_fifo_st_0_write,
    output wire                                          Module2Func_77_ap_clk,
    input wire                                           Module2Func_77_ap_done,
    input wire                                           Module2Func_77_ap_idle,
    input wire                                           Module2Func_77_ap_ready,
    output wire                                          Module2Func_77_ap_rst_n,
    output wire                                          Module2Func_77_ap_start,
    output wire [                                 512:0] Module2Func_77_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_77_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_77_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_77_fifo_ld_0_s_dout,
    output wire                                          Module2Func_77_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_77_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_77_fifo_st_0_din,
    output wire                                          Module2Func_77_fifo_st_0_full_n,
    input wire                                           Module2Func_77_fifo_st_0_write,
    output wire                                          Module2Func_78_ap_clk,
    input wire                                           Module2Func_78_ap_done,
    input wire                                           Module2Func_78_ap_idle,
    input wire                                           Module2Func_78_ap_ready,
    output wire                                          Module2Func_78_ap_rst_n,
    output wire                                          Module2Func_78_ap_start,
    output wire [                                 512:0] Module2Func_78_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_78_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_78_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_78_fifo_ld_0_s_dout,
    output wire                                          Module2Func_78_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_78_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_78_fifo_st_0_din,
    output wire                                          Module2Func_78_fifo_st_0_full_n,
    input wire                                           Module2Func_78_fifo_st_0_write,
    output wire                                          Module2Func_79_ap_clk,
    input wire                                           Module2Func_79_ap_done,
    input wire                                           Module2Func_79_ap_idle,
    input wire                                           Module2Func_79_ap_ready,
    output wire                                          Module2Func_79_ap_rst_n,
    output wire                                          Module2Func_79_ap_start,
    output wire [                                 512:0] Module2Func_79_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_79_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_79_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_79_fifo_ld_0_s_dout,
    output wire                                          Module2Func_79_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_79_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_79_fifo_st_0_din,
    output wire                                          Module2Func_79_fifo_st_0_full_n,
    input wire                                           Module2Func_79_fifo_st_0_write,
    output wire                                          Module2Func_80_ap_clk,
    input wire                                           Module2Func_80_ap_done,
    input wire                                           Module2Func_80_ap_idle,
    input wire                                           Module2Func_80_ap_ready,
    output wire                                          Module2Func_80_ap_rst_n,
    output wire                                          Module2Func_80_ap_start,
    output wire [                                 512:0] Module2Func_80_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_80_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_80_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_80_fifo_ld_0_s_dout,
    output wire                                          Module2Func_80_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_80_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_80_fifo_st_0_din,
    output wire                                          Module2Func_80_fifo_st_0_full_n,
    input wire                                           Module2Func_80_fifo_st_0_write,
    output wire                                          Module2Func_81_ap_clk,
    input wire                                           Module2Func_81_ap_done,
    input wire                                           Module2Func_81_ap_idle,
    input wire                                           Module2Func_81_ap_ready,
    output wire                                          Module2Func_81_ap_rst_n,
    output wire                                          Module2Func_81_ap_start,
    output wire [                                 512:0] Module2Func_81_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_81_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_81_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_81_fifo_ld_0_s_dout,
    output wire                                          Module2Func_81_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_81_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_81_fifo_st_0_din,
    output wire                                          Module2Func_81_fifo_st_0_full_n,
    input wire                                           Module2Func_81_fifo_st_0_write,
    output wire                                          Module2Func_82_ap_clk,
    input wire                                           Module2Func_82_ap_done,
    input wire                                           Module2Func_82_ap_idle,
    input wire                                           Module2Func_82_ap_ready,
    output wire                                          Module2Func_82_ap_rst_n,
    output wire                                          Module2Func_82_ap_start,
    output wire [                                 512:0] Module2Func_82_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_82_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_82_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_82_fifo_ld_0_s_dout,
    output wire                                          Module2Func_82_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_82_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_82_fifo_st_0_din,
    output wire                                          Module2Func_82_fifo_st_0_full_n,
    input wire                                           Module2Func_82_fifo_st_0_write,
    output wire                                          Module2Func_83_ap_clk,
    input wire                                           Module2Func_83_ap_done,
    input wire                                           Module2Func_83_ap_idle,
    input wire                                           Module2Func_83_ap_ready,
    output wire                                          Module2Func_83_ap_rst_n,
    output wire                                          Module2Func_83_ap_start,
    output wire [                                 512:0] Module2Func_83_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_83_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_83_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_83_fifo_ld_0_s_dout,
    output wire                                          Module2Func_83_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_83_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_83_fifo_st_0_din,
    output wire                                          Module2Func_83_fifo_st_0_full_n,
    input wire                                           Module2Func_83_fifo_st_0_write,
    output wire                                          Module2Func_84_ap_clk,
    input wire                                           Module2Func_84_ap_done,
    input wire                                           Module2Func_84_ap_idle,
    input wire                                           Module2Func_84_ap_ready,
    output wire                                          Module2Func_84_ap_rst_n,
    output wire                                          Module2Func_84_ap_start,
    output wire [                                 512:0] Module2Func_84_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_84_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_84_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_84_fifo_ld_0_s_dout,
    output wire                                          Module2Func_84_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_84_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_84_fifo_st_0_din,
    output wire                                          Module2Func_84_fifo_st_0_full_n,
    input wire                                           Module2Func_84_fifo_st_0_write,
    output wire                                          Module2Func_85_ap_clk,
    input wire                                           Module2Func_85_ap_done,
    input wire                                           Module2Func_85_ap_idle,
    input wire                                           Module2Func_85_ap_ready,
    output wire                                          Module2Func_85_ap_rst_n,
    output wire                                          Module2Func_85_ap_start,
    output wire [                                 512:0] Module2Func_85_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_85_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_85_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_85_fifo_ld_0_s_dout,
    output wire                                          Module2Func_85_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_85_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_85_fifo_st_0_din,
    output wire                                          Module2Func_85_fifo_st_0_full_n,
    input wire                                           Module2Func_85_fifo_st_0_write,
    output wire                                          Module2Func_86_ap_clk,
    input wire                                           Module2Func_86_ap_done,
    input wire                                           Module2Func_86_ap_idle,
    input wire                                           Module2Func_86_ap_ready,
    output wire                                          Module2Func_86_ap_rst_n,
    output wire                                          Module2Func_86_ap_start,
    output wire [                                 512:0] Module2Func_86_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_86_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_86_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_86_fifo_ld_0_s_dout,
    output wire                                          Module2Func_86_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_86_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_86_fifo_st_0_din,
    output wire                                          Module2Func_86_fifo_st_0_full_n,
    input wire                                           Module2Func_86_fifo_st_0_write,
    output wire                                          Module2Func_87_ap_clk,
    input wire                                           Module2Func_87_ap_done,
    input wire                                           Module2Func_87_ap_idle,
    input wire                                           Module2Func_87_ap_ready,
    output wire                                          Module2Func_87_ap_rst_n,
    output wire                                          Module2Func_87_ap_start,
    output wire [                                 512:0] Module2Func_87_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_87_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_87_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_87_fifo_ld_0_s_dout,
    output wire                                          Module2Func_87_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_87_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_87_fifo_st_0_din,
    output wire                                          Module2Func_87_fifo_st_0_full_n,
    input wire                                           Module2Func_87_fifo_st_0_write,
    output wire                                          Module2Func_88_ap_clk,
    input wire                                           Module2Func_88_ap_done,
    input wire                                           Module2Func_88_ap_idle,
    input wire                                           Module2Func_88_ap_ready,
    output wire                                          Module2Func_88_ap_rst_n,
    output wire                                          Module2Func_88_ap_start,
    output wire [                                 512:0] Module2Func_88_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_88_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_88_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_88_fifo_ld_0_s_dout,
    output wire                                          Module2Func_88_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_88_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_88_fifo_st_0_din,
    output wire                                          Module2Func_88_fifo_st_0_full_n,
    input wire                                           Module2Func_88_fifo_st_0_write,
    output wire                                          Module2Func_89_ap_clk,
    input wire                                           Module2Func_89_ap_done,
    input wire                                           Module2Func_89_ap_idle,
    input wire                                           Module2Func_89_ap_ready,
    output wire                                          Module2Func_89_ap_rst_n,
    output wire                                          Module2Func_89_ap_start,
    output wire [                                 512:0] Module2Func_89_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_89_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_89_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_89_fifo_ld_0_s_dout,
    output wire                                          Module2Func_89_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_89_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_89_fifo_st_0_din,
    output wire                                          Module2Func_89_fifo_st_0_full_n,
    input wire                                           Module2Func_89_fifo_st_0_write,
    output wire                                          Module2Func_90_ap_clk,
    input wire                                           Module2Func_90_ap_done,
    input wire                                           Module2Func_90_ap_idle,
    input wire                                           Module2Func_90_ap_ready,
    output wire                                          Module2Func_90_ap_rst_n,
    output wire                                          Module2Func_90_ap_start,
    output wire [                                 512:0] Module2Func_90_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_90_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_90_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_90_fifo_ld_0_s_dout,
    output wire                                          Module2Func_90_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_90_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_90_fifo_st_0_din,
    output wire                                          Module2Func_90_fifo_st_0_full_n,
    input wire                                           Module2Func_90_fifo_st_0_write,
    output wire                                          Module2Func_91_ap_clk,
    input wire                                           Module2Func_91_ap_done,
    input wire                                           Module2Func_91_ap_idle,
    input wire                                           Module2Func_91_ap_ready,
    output wire                                          Module2Func_91_ap_rst_n,
    output wire                                          Module2Func_91_ap_start,
    output wire [                                 512:0] Module2Func_91_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_91_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_91_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_91_fifo_ld_0_s_dout,
    output wire                                          Module2Func_91_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_91_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_91_fifo_st_0_din,
    output wire                                          Module2Func_91_fifo_st_0_full_n,
    input wire                                           Module2Func_91_fifo_st_0_write,
    output wire                                          Module2Func_92_ap_clk,
    input wire                                           Module2Func_92_ap_done,
    input wire                                           Module2Func_92_ap_idle,
    input wire                                           Module2Func_92_ap_ready,
    output wire                                          Module2Func_92_ap_rst_n,
    output wire                                          Module2Func_92_ap_start,
    output wire [                                 512:0] Module2Func_92_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_92_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_92_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_92_fifo_ld_0_s_dout,
    output wire                                          Module2Func_92_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_92_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_92_fifo_st_0_din,
    output wire                                          Module2Func_92_fifo_st_0_full_n,
    input wire                                           Module2Func_92_fifo_st_0_write,
    output wire                                          Module2Func_93_ap_clk,
    input wire                                           Module2Func_93_ap_done,
    input wire                                           Module2Func_93_ap_idle,
    input wire                                           Module2Func_93_ap_ready,
    output wire                                          Module2Func_93_ap_rst_n,
    output wire                                          Module2Func_93_ap_start,
    output wire [                                 512:0] Module2Func_93_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_93_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_93_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_93_fifo_ld_0_s_dout,
    output wire                                          Module2Func_93_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_93_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_93_fifo_st_0_din,
    output wire                                          Module2Func_93_fifo_st_0_full_n,
    input wire                                           Module2Func_93_fifo_st_0_write,
    output wire                                          Module2Func_94_ap_clk,
    input wire                                           Module2Func_94_ap_done,
    input wire                                           Module2Func_94_ap_idle,
    input wire                                           Module2Func_94_ap_ready,
    output wire                                          Module2Func_94_ap_rst_n,
    output wire                                          Module2Func_94_ap_start,
    output wire [                                 512:0] Module2Func_94_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_94_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_94_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_94_fifo_ld_0_s_dout,
    output wire                                          Module2Func_94_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_94_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_94_fifo_st_0_din,
    output wire                                          Module2Func_94_fifo_st_0_full_n,
    input wire                                           Module2Func_94_fifo_st_0_write,
    output wire                                          Module2Func_95_ap_clk,
    input wire                                           Module2Func_95_ap_done,
    input wire                                           Module2Func_95_ap_idle,
    input wire                                           Module2Func_95_ap_ready,
    output wire                                          Module2Func_95_ap_rst_n,
    output wire                                          Module2Func_95_ap_start,
    output wire [                                 512:0] Module2Func_95_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_95_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_95_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_95_fifo_ld_0_s_dout,
    output wire                                          Module2Func_95_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_95_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_95_fifo_st_0_din,
    output wire                                          Module2Func_95_fifo_st_0_full_n,
    input wire                                           Module2Func_95_fifo_st_0_write,
    output wire                                          Module2Func_96_ap_clk,
    input wire                                           Module2Func_96_ap_done,
    input wire                                           Module2Func_96_ap_idle,
    input wire                                           Module2Func_96_ap_ready,
    output wire                                          Module2Func_96_ap_rst_n,
    output wire                                          Module2Func_96_ap_start,
    output wire [                                 512:0] Module2Func_96_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_96_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_96_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_96_fifo_ld_0_s_dout,
    output wire                                          Module2Func_96_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_96_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_96_fifo_st_0_din,
    output wire                                          Module2Func_96_fifo_st_0_full_n,
    input wire                                           Module2Func_96_fifo_st_0_write,
    output wire                                          Module2Func_97_ap_clk,
    input wire                                           Module2Func_97_ap_done,
    input wire                                           Module2Func_97_ap_idle,
    input wire                                           Module2Func_97_ap_ready,
    output wire                                          Module2Func_97_ap_rst_n,
    output wire                                          Module2Func_97_ap_start,
    output wire [                                 512:0] Module2Func_97_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_97_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_97_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_97_fifo_ld_0_s_dout,
    output wire                                          Module2Func_97_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_97_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_97_fifo_st_0_din,
    output wire                                          Module2Func_97_fifo_st_0_full_n,
    input wire                                           Module2Func_97_fifo_st_0_write,
    output wire                                          Module2Func_98_ap_clk,
    input wire                                           Module2Func_98_ap_done,
    input wire                                           Module2Func_98_ap_idle,
    input wire                                           Module2Func_98_ap_ready,
    output wire                                          Module2Func_98_ap_rst_n,
    output wire                                          Module2Func_98_ap_start,
    output wire [                                 512:0] Module2Func_98_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_98_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_98_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_98_fifo_ld_0_s_dout,
    output wire                                          Module2Func_98_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_98_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_98_fifo_st_0_din,
    output wire                                          Module2Func_98_fifo_st_0_full_n,
    input wire                                           Module2Func_98_fifo_st_0_write,
    output wire                                          Module2Func_99_ap_clk,
    input wire                                           Module2Func_99_ap_done,
    input wire                                           Module2Func_99_ap_idle,
    input wire                                           Module2Func_99_ap_ready,
    output wire                                          Module2Func_99_ap_rst_n,
    output wire                                          Module2Func_99_ap_start,
    output wire [                                 512:0] Module2Func_99_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_99_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_99_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_99_fifo_ld_0_s_dout,
    output wire                                          Module2Func_99_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_99_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_99_fifo_st_0_din,
    output wire                                          Module2Func_99_fifo_st_0_full_n,
    input wire                                           Module2Func_99_fifo_st_0_write,
    output wire                                          Module2Func_100_ap_clk,
    input wire                                           Module2Func_100_ap_done,
    input wire                                           Module2Func_100_ap_idle,
    input wire                                           Module2Func_100_ap_ready,
    output wire                                          Module2Func_100_ap_rst_n,
    output wire                                          Module2Func_100_ap_start,
    output wire [                                 512:0] Module2Func_100_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_100_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_100_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_100_fifo_ld_0_s_dout,
    output wire                                          Module2Func_100_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_100_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_100_fifo_st_0_din,
    output wire                                          Module2Func_100_fifo_st_0_full_n,
    input wire                                           Module2Func_100_fifo_st_0_write,
    output wire                                          Module2Func_101_ap_clk,
    input wire                                           Module2Func_101_ap_done,
    input wire                                           Module2Func_101_ap_idle,
    input wire                                           Module2Func_101_ap_ready,
    output wire                                          Module2Func_101_ap_rst_n,
    output wire                                          Module2Func_101_ap_start,
    output wire [                                 512:0] Module2Func_101_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_101_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_101_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_101_fifo_ld_0_s_dout,
    output wire                                          Module2Func_101_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_101_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_101_fifo_st_0_din,
    output wire                                          Module2Func_101_fifo_st_0_full_n,
    input wire                                           Module2Func_101_fifo_st_0_write,
    output wire                                          Module2Func_102_ap_clk,
    input wire                                           Module2Func_102_ap_done,
    input wire                                           Module2Func_102_ap_idle,
    input wire                                           Module2Func_102_ap_ready,
    output wire                                          Module2Func_102_ap_rst_n,
    output wire                                          Module2Func_102_ap_start,
    output wire [                                 512:0] Module2Func_102_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_102_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_102_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_102_fifo_ld_0_s_dout,
    output wire                                          Module2Func_102_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_102_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_102_fifo_st_0_din,
    output wire                                          Module2Func_102_fifo_st_0_full_n,
    input wire                                           Module2Func_102_fifo_st_0_write,
    output wire                                          Module2Func_103_ap_clk,
    input wire                                           Module2Func_103_ap_done,
    input wire                                           Module2Func_103_ap_idle,
    input wire                                           Module2Func_103_ap_ready,
    output wire                                          Module2Func_103_ap_rst_n,
    output wire                                          Module2Func_103_ap_start,
    output wire [                                 512:0] Module2Func_103_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_103_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_103_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_103_fifo_ld_0_s_dout,
    output wire                                          Module2Func_103_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_103_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_103_fifo_st_0_din,
    output wire                                          Module2Func_103_fifo_st_0_full_n,
    input wire                                           Module2Func_103_fifo_st_0_write,
    output wire                                          Module2Func_104_ap_clk,
    input wire                                           Module2Func_104_ap_done,
    input wire                                           Module2Func_104_ap_idle,
    input wire                                           Module2Func_104_ap_ready,
    output wire                                          Module2Func_104_ap_rst_n,
    output wire                                          Module2Func_104_ap_start,
    output wire [                                 512:0] Module2Func_104_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_104_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_104_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_104_fifo_ld_0_s_dout,
    output wire                                          Module2Func_104_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_104_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_104_fifo_st_0_din,
    output wire                                          Module2Func_104_fifo_st_0_full_n,
    input wire                                           Module2Func_104_fifo_st_0_write,
    output wire                                          Module2Func_105_ap_clk,
    input wire                                           Module2Func_105_ap_done,
    input wire                                           Module2Func_105_ap_idle,
    input wire                                           Module2Func_105_ap_ready,
    output wire                                          Module2Func_105_ap_rst_n,
    output wire                                          Module2Func_105_ap_start,
    output wire [                                 512:0] Module2Func_105_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_105_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_105_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_105_fifo_ld_0_s_dout,
    output wire                                          Module2Func_105_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_105_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_105_fifo_st_0_din,
    output wire                                          Module2Func_105_fifo_st_0_full_n,
    input wire                                           Module2Func_105_fifo_st_0_write,
    output wire                                          Module2Func_106_ap_clk,
    input wire                                           Module2Func_106_ap_done,
    input wire                                           Module2Func_106_ap_idle,
    input wire                                           Module2Func_106_ap_ready,
    output wire                                          Module2Func_106_ap_rst_n,
    output wire                                          Module2Func_106_ap_start,
    output wire [                                 512:0] Module2Func_106_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_106_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_106_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_106_fifo_ld_0_s_dout,
    output wire                                          Module2Func_106_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_106_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_106_fifo_st_0_din,
    output wire                                          Module2Func_106_fifo_st_0_full_n,
    input wire                                           Module2Func_106_fifo_st_0_write,
    output wire                                          Module2Func_107_ap_clk,
    input wire                                           Module2Func_107_ap_done,
    input wire                                           Module2Func_107_ap_idle,
    input wire                                           Module2Func_107_ap_ready,
    output wire                                          Module2Func_107_ap_rst_n,
    output wire                                          Module2Func_107_ap_start,
    output wire [                                 512:0] Module2Func_107_fifo_ld_0_peek_dout,
    output wire                                          Module2Func_107_fifo_ld_0_peek_empty_n,
    input wire                                           Module2Func_107_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module2Func_107_fifo_ld_0_s_dout,
    output wire                                          Module2Func_107_fifo_ld_0_s_empty_n,
    input wire                                           Module2Func_107_fifo_ld_0_s_read,
    input wire  [                                 512:0] Module2Func_107_fifo_st_0_din,
    output wire                                          Module2Func_107_fifo_st_0_full_n,
    input wire                                           Module2Func_107_fifo_st_0_write,
    output wire                                          Module3Func_0_ap_clk,
    input wire                                           Module3Func_0_ap_done,
    input wire                                           Module3Func_0_ap_idle,
    input wire                                           Module3Func_0_ap_ready,
    output wire                                          Module3Func_0_ap_rst_n,
    output wire                                          Module3Func_0_ap_start,
    input wire  [                                 512:0] Module3Func_0_dram_t0_bank_1_fifo_din,
    output wire                                          Module3Func_0_dram_t0_bank_1_fifo_full_n,
    input wire                                           Module3Func_0_dram_t0_bank_1_fifo_write,
    output wire [                                 512:0] Module3Func_0_fifo_ld_0_peek_dout,
    output wire                                          Module3Func_0_fifo_ld_0_peek_empty_n,
    input wire                                           Module3Func_0_fifo_ld_0_peek_read,
    output wire [                                 512:0] Module3Func_0_fifo_ld_0_s_dout,
    output wire                                          Module3Func_0_fifo_ld_0_s_empty_n,
    input wire                                           Module3Func_0_fifo_ld_0_s_read,
    output wire                                          bank_0_t1__m_axi_clk,
    input wire  [                                  63:0] bank_0_t1__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] bank_0_t1__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] bank_0_t1__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] bank_0_t1__m_axi_m_axi_ARID,
    input wire  [                                   7:0] bank_0_t1__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] bank_0_t1__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] bank_0_t1__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] bank_0_t1__m_axi_m_axi_ARQOS,
    output wire                                          bank_0_t1__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] bank_0_t1__m_axi_m_axi_ARSIZE,
    input wire                                           bank_0_t1__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] bank_0_t1__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] bank_0_t1__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] bank_0_t1__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] bank_0_t1__m_axi_m_axi_AWID,
    input wire  [                                   7:0] bank_0_t1__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] bank_0_t1__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] bank_0_t1__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] bank_0_t1__m_axi_m_axi_AWQOS,
    output wire                                          bank_0_t1__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] bank_0_t1__m_axi_m_axi_AWSIZE,
    input wire                                           bank_0_t1__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] bank_0_t1__m_axi_m_axi_BID,
    input wire                                           bank_0_t1__m_axi_m_axi_BREADY,
    output wire [                                   1:0] bank_0_t1__m_axi_m_axi_BRESP,
    output wire                                          bank_0_t1__m_axi_m_axi_BVALID,
    output wire [                                 511:0] bank_0_t1__m_axi_m_axi_RDATA,
    output wire [                                   0:0] bank_0_t1__m_axi_m_axi_RID,
    output wire                                          bank_0_t1__m_axi_m_axi_RLAST,
    input wire                                           bank_0_t1__m_axi_m_axi_RREADY,
    output wire [                                   1:0] bank_0_t1__m_axi_m_axi_RRESP,
    output wire                                          bank_0_t1__m_axi_m_axi_RVALID,
    input wire  [                                 511:0] bank_0_t1__m_axi_m_axi_WDATA,
    input wire                                           bank_0_t1__m_axi_m_axi_WLAST,
    output wire                                          bank_0_t1__m_axi_m_axi_WREADY,
    input wire  [                                  63:0] bank_0_t1__m_axi_m_axi_WSTRB,
    input wire                                           bank_0_t1__m_axi_m_axi_WVALID,
    output wire [                                  63:0] bank_0_t1__m_axi_read_addr_din,
    input wire                                           bank_0_t1__m_axi_read_addr_full_n,
    output wire                                          bank_0_t1__m_axi_read_addr_write,
    input wire  [                                 511:0] bank_0_t1__m_axi_read_data_dout,
    input wire                                           bank_0_t1__m_axi_read_data_empty_n,
    output wire                                          bank_0_t1__m_axi_read_data_read,
    output wire                                          bank_0_t1__m_axi_rst,
    output wire [                                  63:0] bank_0_t1__m_axi_write_addr_din,
    input wire                                           bank_0_t1__m_axi_write_addr_full_n,
    output wire                                          bank_0_t1__m_axi_write_addr_write,
    output wire [                                 511:0] bank_0_t1__m_axi_write_data_din,
    input wire                                           bank_0_t1__m_axi_write_data_full_n,
    output wire                                          bank_0_t1__m_axi_write_data_write,
    input wire  [                                   7:0] bank_0_t1__m_axi_write_resp_dout,
    input wire                                           bank_0_t1__m_axi_write_resp_empty_n,
    output wire                                          bank_0_t1__m_axi_write_resp_read,
    output wire                                          bank_1_t0__m_axi_clk,
    input wire  [                                  63:0] bank_1_t0__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] bank_1_t0__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] bank_1_t0__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] bank_1_t0__m_axi_m_axi_ARID,
    input wire  [                                   7:0] bank_1_t0__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] bank_1_t0__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] bank_1_t0__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] bank_1_t0__m_axi_m_axi_ARQOS,
    output wire                                          bank_1_t0__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] bank_1_t0__m_axi_m_axi_ARSIZE,
    input wire                                           bank_1_t0__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] bank_1_t0__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] bank_1_t0__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] bank_1_t0__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] bank_1_t0__m_axi_m_axi_AWID,
    input wire  [                                   7:0] bank_1_t0__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] bank_1_t0__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] bank_1_t0__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] bank_1_t0__m_axi_m_axi_AWQOS,
    output wire                                          bank_1_t0__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] bank_1_t0__m_axi_m_axi_AWSIZE,
    input wire                                           bank_1_t0__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] bank_1_t0__m_axi_m_axi_BID,
    input wire                                           bank_1_t0__m_axi_m_axi_BREADY,
    output wire [                                   1:0] bank_1_t0__m_axi_m_axi_BRESP,
    output wire                                          bank_1_t0__m_axi_m_axi_BVALID,
    output wire [                                 511:0] bank_1_t0__m_axi_m_axi_RDATA,
    output wire [                                   0:0] bank_1_t0__m_axi_m_axi_RID,
    output wire                                          bank_1_t0__m_axi_m_axi_RLAST,
    input wire                                           bank_1_t0__m_axi_m_axi_RREADY,
    output wire [                                   1:0] bank_1_t0__m_axi_m_axi_RRESP,
    output wire                                          bank_1_t0__m_axi_m_axi_RVALID,
    input wire  [                                 511:0] bank_1_t0__m_axi_m_axi_WDATA,
    input wire                                           bank_1_t0__m_axi_m_axi_WLAST,
    output wire                                          bank_1_t0__m_axi_m_axi_WREADY,
    input wire  [                                  63:0] bank_1_t0__m_axi_m_axi_WSTRB,
    input wire                                           bank_1_t0__m_axi_m_axi_WVALID,
    output wire [                                  63:0] bank_1_t0__m_axi_read_addr_din,
    input wire                                           bank_1_t0__m_axi_read_addr_full_n,
    output wire                                          bank_1_t0__m_axi_read_addr_write,
    input wire  [                                 511:0] bank_1_t0__m_axi_read_data_dout,
    input wire                                           bank_1_t0__m_axi_read_data_empty_n,
    output wire                                          bank_1_t0__m_axi_read_data_read,
    output wire                                          bank_1_t0__m_axi_rst,
    output wire [                                  63:0] bank_1_t0__m_axi_write_addr_din,
    input wire                                           bank_1_t0__m_axi_write_addr_full_n,
    output wire                                          bank_1_t0__m_axi_write_addr_write,
    output wire [                                 511:0] bank_1_t0__m_axi_write_data_din,
    input wire                                           bank_1_t0__m_axi_write_data_full_n,
    output wire                                          bank_1_t0__m_axi_write_data_write,
    input wire  [                                   7:0] bank_1_t0__m_axi_write_resp_dout,
    input wire                                           bank_1_t0__m_axi_write_resp_empty_n,
    output wire                                          bank_1_t0__m_axi_write_resp_read,
    input wire  [                                  63:0] __tapa_fsm_unit_BurstRead_floatx16_0___bank_0_t1__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_BurstRead_floatx16_0___coalesced_data_num__q0,
    output wire                                          __tapa_fsm_unit_BurstRead_floatx16_0__ap_done,
    output wire                                          __tapa_fsm_unit_BurstRead_floatx16_0__ap_idle,
    output wire                                          __tapa_fsm_unit_BurstRead_floatx16_0__ap_ready,
    input wire                                           __tapa_fsm_unit_BurstRead_floatx16_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_BurstWrite_floatx16_0___bank_1_t0__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_BurstWrite_floatx16_0___coalesced_data_num__q0,
    output wire                                          __tapa_fsm_unit_BurstWrite_floatx16_0__ap_done,
    output wire                                          __tapa_fsm_unit_BurstWrite_floatx16_0__ap_idle,
    output wire                                          __tapa_fsm_unit_BurstWrite_floatx16_0__ap_ready,
    input wire                                           __tapa_fsm_unit_BurstWrite_floatx16_0__ap_start,
    input wire                                           __tapa_fsm_unit_Module0Func_0__ap_start,
    input wire                                           __tapa_fsm_unit_Module1Func_0__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_0__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_100__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_101__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_102__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_103__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_104__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_105__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_106__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_107__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_10__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_11__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_12__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_13__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_14__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_15__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_16__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_17__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_18__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_19__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_1__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_20__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_21__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_22__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_23__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_24__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_25__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_26__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_27__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_28__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_29__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_2__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_30__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_31__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_32__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_33__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_34__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_35__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_36__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_37__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_38__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_39__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_3__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_40__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_41__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_42__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_43__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_44__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_45__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_46__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_47__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_48__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_49__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_4__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_50__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_51__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_52__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_53__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_54__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_55__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_56__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_57__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_58__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_59__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_5__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_60__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_61__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_62__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_63__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_64__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_65__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_66__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_67__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_68__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_69__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_6__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_70__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_71__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_72__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_73__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_74__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_75__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_76__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_77__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_78__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_79__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_7__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_80__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_81__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_82__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_83__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_84__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_85__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_86__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_87__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_88__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_89__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_8__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_90__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_91__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_92__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_93__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_94__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_95__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_96__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_97__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_98__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_99__ap_start,
    input wire                                           __tapa_fsm_unit_Module2Func_9__ap_start,
    input wire                                           __tapa_fsm_unit_Module3Func_0__ap_start,
    output wire                                          __tapa_fsm_unit_ap_clk,
    input wire                                           __tapa_fsm_unit_ap_done,
    input wire                                           __tapa_fsm_unit_ap_idle,
    input wire                                           __tapa_fsm_unit_ap_ready,
    output wire                                          __tapa_fsm_unit_ap_rst_n,
    output wire                                          __tapa_fsm_unit_ap_start,
    output wire [                                  63:0] __tapa_fsm_unit_bank_0_t1,
    output wire [                                  63:0] __tapa_fsm_unit_bank_1_t0,
    output wire [                                  63:0] __tapa_fsm_unit_coalesced_data_num
);
  wire ap_start;
  wire [63:0] bank_1_t0;
  wire [63:0] bank_0_t1;
  wire [63:0] coalesced_data_num;
  wire [512:0] bank_0_t1_buf__dout;
  wire bank_0_t1_buf__empty_n;
  wire bank_0_t1_buf__read;
  wire [512:0] bank_0_t1_buf__din;
  wire bank_0_t1_buf__full_n;
  wire bank_0_t1_buf__write;
  wire [512:0] bank_1_t0_buf__dout;
  wire bank_1_t0_buf__empty_n;
  wire bank_1_t0_buf__read;
  wire [512:0] bank_1_t0_buf__din;
  wire bank_1_t0_buf__full_n;
  wire bank_1_t0_buf__write;
  wire [512:0] from_t0_to_t0_bank_1__dout;
  wire from_t0_to_t0_bank_1__empty_n;
  wire from_t0_to_t0_bank_1__read;
  wire [512:0] from_t0_to_t0_bank_1__din;
  wire from_t0_to_t0_bank_1__full_n;
  wire from_t0_to_t0_bank_1__write;
  wire [512:0] from_t1_bank_0_to_t1_iter1__dout;
  wire from_t1_bank_0_to_t1_iter1__empty_n;
  wire from_t1_bank_0_to_t1_iter1__read;
  wire [512:0] from_t1_bank_0_to_t1_iter1__din;
  wire from_t1_bank_0_to_t1_iter1__full_n;
  wire from_t1_bank_0_to_t1_iter1__write;
  wire [512:0] from_t1_iter100_to_t1_iter101__dout;
  wire from_t1_iter100_to_t1_iter101__empty_n;
  wire from_t1_iter100_to_t1_iter101__read;
  wire [512:0] from_t1_iter100_to_t1_iter101__din;
  wire from_t1_iter100_to_t1_iter101__full_n;
  wire from_t1_iter100_to_t1_iter101__write;
  wire [512:0] from_t1_iter101_to_t1_iter102__dout;
  wire from_t1_iter101_to_t1_iter102__empty_n;
  wire from_t1_iter101_to_t1_iter102__read;
  wire [512:0] from_t1_iter101_to_t1_iter102__din;
  wire from_t1_iter101_to_t1_iter102__full_n;
  wire from_t1_iter101_to_t1_iter102__write;
  wire [512:0] from_t1_iter102_to_t1_iter103__dout;
  wire from_t1_iter102_to_t1_iter103__empty_n;
  wire from_t1_iter102_to_t1_iter103__read;
  wire [512:0] from_t1_iter102_to_t1_iter103__din;
  wire from_t1_iter102_to_t1_iter103__full_n;
  wire from_t1_iter102_to_t1_iter103__write;
  wire [512:0] from_t1_iter103_to_t1_iter104__dout;
  wire from_t1_iter103_to_t1_iter104__empty_n;
  wire from_t1_iter103_to_t1_iter104__read;
  wire [512:0] from_t1_iter103_to_t1_iter104__din;
  wire from_t1_iter103_to_t1_iter104__full_n;
  wire from_t1_iter103_to_t1_iter104__write;
  wire [512:0] from_t1_iter104_to_t1_iter105__dout;
  wire from_t1_iter104_to_t1_iter105__empty_n;
  wire from_t1_iter104_to_t1_iter105__read;
  wire [512:0] from_t1_iter104_to_t1_iter105__din;
  wire from_t1_iter104_to_t1_iter105__full_n;
  wire from_t1_iter104_to_t1_iter105__write;
  wire [512:0] from_t1_iter105_to_t1_iter106__dout;
  wire from_t1_iter105_to_t1_iter106__empty_n;
  wire from_t1_iter105_to_t1_iter106__read;
  wire [512:0] from_t1_iter105_to_t1_iter106__din;
  wire from_t1_iter105_to_t1_iter106__full_n;
  wire from_t1_iter105_to_t1_iter106__write;
  wire [512:0] from_t1_iter106_to_t1_iter107__dout;
  wire from_t1_iter106_to_t1_iter107__empty_n;
  wire from_t1_iter106_to_t1_iter107__read;
  wire [512:0] from_t1_iter106_to_t1_iter107__din;
  wire from_t1_iter106_to_t1_iter107__full_n;
  wire from_t1_iter106_to_t1_iter107__write;
  wire [512:0] from_t1_iter107_to_t1_iter108__dout;
  wire from_t1_iter107_to_t1_iter108__empty_n;
  wire from_t1_iter107_to_t1_iter108__read;
  wire [512:0] from_t1_iter107_to_t1_iter108__din;
  wire from_t1_iter107_to_t1_iter108__full_n;
  wire from_t1_iter107_to_t1_iter108__write;
  wire [512:0] from_t1_iter108_to_t0__dout;
  wire from_t1_iter108_to_t0__empty_n;
  wire from_t1_iter108_to_t0__read;
  wire [512:0] from_t1_iter108_to_t0__din;
  wire from_t1_iter108_to_t0__full_n;
  wire from_t1_iter108_to_t0__write;
  wire [512:0] from_t1_iter10_to_t1_iter11__dout;
  wire from_t1_iter10_to_t1_iter11__empty_n;
  wire from_t1_iter10_to_t1_iter11__read;
  wire [512:0] from_t1_iter10_to_t1_iter11__din;
  wire from_t1_iter10_to_t1_iter11__full_n;
  wire from_t1_iter10_to_t1_iter11__write;
  wire [512:0] from_t1_iter11_to_t1_iter12__dout;
  wire from_t1_iter11_to_t1_iter12__empty_n;
  wire from_t1_iter11_to_t1_iter12__read;
  wire [512:0] from_t1_iter11_to_t1_iter12__din;
  wire from_t1_iter11_to_t1_iter12__full_n;
  wire from_t1_iter11_to_t1_iter12__write;
  wire [512:0] from_t1_iter12_to_t1_iter13__dout;
  wire from_t1_iter12_to_t1_iter13__empty_n;
  wire from_t1_iter12_to_t1_iter13__read;
  wire [512:0] from_t1_iter12_to_t1_iter13__din;
  wire from_t1_iter12_to_t1_iter13__full_n;
  wire from_t1_iter12_to_t1_iter13__write;
  wire [512:0] from_t1_iter13_to_t1_iter14__dout;
  wire from_t1_iter13_to_t1_iter14__empty_n;
  wire from_t1_iter13_to_t1_iter14__read;
  wire [512:0] from_t1_iter13_to_t1_iter14__din;
  wire from_t1_iter13_to_t1_iter14__full_n;
  wire from_t1_iter13_to_t1_iter14__write;
  wire [512:0] from_t1_iter14_to_t1_iter15__dout;
  wire from_t1_iter14_to_t1_iter15__empty_n;
  wire from_t1_iter14_to_t1_iter15__read;
  wire [512:0] from_t1_iter14_to_t1_iter15__din;
  wire from_t1_iter14_to_t1_iter15__full_n;
  wire from_t1_iter14_to_t1_iter15__write;
  wire [512:0] from_t1_iter15_to_t1_iter16__dout;
  wire from_t1_iter15_to_t1_iter16__empty_n;
  wire from_t1_iter15_to_t1_iter16__read;
  wire [512:0] from_t1_iter15_to_t1_iter16__din;
  wire from_t1_iter15_to_t1_iter16__full_n;
  wire from_t1_iter15_to_t1_iter16__write;
  wire [512:0] from_t1_iter16_to_t1_iter17__dout;
  wire from_t1_iter16_to_t1_iter17__empty_n;
  wire from_t1_iter16_to_t1_iter17__read;
  wire [512:0] from_t1_iter16_to_t1_iter17__din;
  wire from_t1_iter16_to_t1_iter17__full_n;
  wire from_t1_iter16_to_t1_iter17__write;
  wire [512:0] from_t1_iter17_to_t1_iter18__dout;
  wire from_t1_iter17_to_t1_iter18__empty_n;
  wire from_t1_iter17_to_t1_iter18__read;
  wire [512:0] from_t1_iter17_to_t1_iter18__din;
  wire from_t1_iter17_to_t1_iter18__full_n;
  wire from_t1_iter17_to_t1_iter18__write;
  wire [512:0] from_t1_iter18_to_t1_iter19__dout;
  wire from_t1_iter18_to_t1_iter19__empty_n;
  wire from_t1_iter18_to_t1_iter19__read;
  wire [512:0] from_t1_iter18_to_t1_iter19__din;
  wire from_t1_iter18_to_t1_iter19__full_n;
  wire from_t1_iter18_to_t1_iter19__write;
  wire [512:0] from_t1_iter19_to_t1_iter20__dout;
  wire from_t1_iter19_to_t1_iter20__empty_n;
  wire from_t1_iter19_to_t1_iter20__read;
  wire [512:0] from_t1_iter19_to_t1_iter20__din;
  wire from_t1_iter19_to_t1_iter20__full_n;
  wire from_t1_iter19_to_t1_iter20__write;
  wire [512:0] from_t1_iter1_to_t1_iter2__dout;
  wire from_t1_iter1_to_t1_iter2__empty_n;
  wire from_t1_iter1_to_t1_iter2__read;
  wire [512:0] from_t1_iter1_to_t1_iter2__din;
  wire from_t1_iter1_to_t1_iter2__full_n;
  wire from_t1_iter1_to_t1_iter2__write;
  wire [512:0] from_t1_iter20_to_t1_iter21__dout;
  wire from_t1_iter20_to_t1_iter21__empty_n;
  wire from_t1_iter20_to_t1_iter21__read;
  wire [512:0] from_t1_iter20_to_t1_iter21__din;
  wire from_t1_iter20_to_t1_iter21__full_n;
  wire from_t1_iter20_to_t1_iter21__write;
  wire [512:0] from_t1_iter21_to_t1_iter22__dout;
  wire from_t1_iter21_to_t1_iter22__empty_n;
  wire from_t1_iter21_to_t1_iter22__read;
  wire [512:0] from_t1_iter21_to_t1_iter22__din;
  wire from_t1_iter21_to_t1_iter22__full_n;
  wire from_t1_iter21_to_t1_iter22__write;
  wire [512:0] from_t1_iter22_to_t1_iter23__dout;
  wire from_t1_iter22_to_t1_iter23__empty_n;
  wire from_t1_iter22_to_t1_iter23__read;
  wire [512:0] from_t1_iter22_to_t1_iter23__din;
  wire from_t1_iter22_to_t1_iter23__full_n;
  wire from_t1_iter22_to_t1_iter23__write;
  wire [512:0] from_t1_iter23_to_t1_iter24__dout;
  wire from_t1_iter23_to_t1_iter24__empty_n;
  wire from_t1_iter23_to_t1_iter24__read;
  wire [512:0] from_t1_iter23_to_t1_iter24__din;
  wire from_t1_iter23_to_t1_iter24__full_n;
  wire from_t1_iter23_to_t1_iter24__write;
  wire [512:0] from_t1_iter24_to_t1_iter25__dout;
  wire from_t1_iter24_to_t1_iter25__empty_n;
  wire from_t1_iter24_to_t1_iter25__read;
  wire [512:0] from_t1_iter24_to_t1_iter25__din;
  wire from_t1_iter24_to_t1_iter25__full_n;
  wire from_t1_iter24_to_t1_iter25__write;
  wire [512:0] from_t1_iter25_to_t1_iter26__dout;
  wire from_t1_iter25_to_t1_iter26__empty_n;
  wire from_t1_iter25_to_t1_iter26__read;
  wire [512:0] from_t1_iter25_to_t1_iter26__din;
  wire from_t1_iter25_to_t1_iter26__full_n;
  wire from_t1_iter25_to_t1_iter26__write;
  wire [512:0] from_t1_iter26_to_t1_iter27__dout;
  wire from_t1_iter26_to_t1_iter27__empty_n;
  wire from_t1_iter26_to_t1_iter27__read;
  wire [512:0] from_t1_iter26_to_t1_iter27__din;
  wire from_t1_iter26_to_t1_iter27__full_n;
  wire from_t1_iter26_to_t1_iter27__write;
  wire [512:0] from_t1_iter27_to_t1_iter28__dout;
  wire from_t1_iter27_to_t1_iter28__empty_n;
  wire from_t1_iter27_to_t1_iter28__read;
  wire [512:0] from_t1_iter27_to_t1_iter28__din;
  wire from_t1_iter27_to_t1_iter28__full_n;
  wire from_t1_iter27_to_t1_iter28__write;
  wire [512:0] from_t1_iter28_to_t1_iter29__dout;
  wire from_t1_iter28_to_t1_iter29__empty_n;
  wire from_t1_iter28_to_t1_iter29__read;
  wire [512:0] from_t1_iter28_to_t1_iter29__din;
  wire from_t1_iter28_to_t1_iter29__full_n;
  wire from_t1_iter28_to_t1_iter29__write;
  wire [512:0] from_t1_iter29_to_t1_iter30__dout;
  wire from_t1_iter29_to_t1_iter30__empty_n;
  wire from_t1_iter29_to_t1_iter30__read;
  wire [512:0] from_t1_iter29_to_t1_iter30__din;
  wire from_t1_iter29_to_t1_iter30__full_n;
  wire from_t1_iter29_to_t1_iter30__write;
  wire [512:0] from_t1_iter2_to_t1_iter3__dout;
  wire from_t1_iter2_to_t1_iter3__empty_n;
  wire from_t1_iter2_to_t1_iter3__read;
  wire [512:0] from_t1_iter2_to_t1_iter3__din;
  wire from_t1_iter2_to_t1_iter3__full_n;
  wire from_t1_iter2_to_t1_iter3__write;
  wire [512:0] from_t1_iter30_to_t1_iter31__dout;
  wire from_t1_iter30_to_t1_iter31__empty_n;
  wire from_t1_iter30_to_t1_iter31__read;
  wire [512:0] from_t1_iter30_to_t1_iter31__din;
  wire from_t1_iter30_to_t1_iter31__full_n;
  wire from_t1_iter30_to_t1_iter31__write;
  wire [512:0] from_t1_iter31_to_t1_iter32__dout;
  wire from_t1_iter31_to_t1_iter32__empty_n;
  wire from_t1_iter31_to_t1_iter32__read;
  wire [512:0] from_t1_iter31_to_t1_iter32__din;
  wire from_t1_iter31_to_t1_iter32__full_n;
  wire from_t1_iter31_to_t1_iter32__write;
  wire [512:0] from_t1_iter32_to_t1_iter33__dout;
  wire from_t1_iter32_to_t1_iter33__empty_n;
  wire from_t1_iter32_to_t1_iter33__read;
  wire [512:0] from_t1_iter32_to_t1_iter33__din;
  wire from_t1_iter32_to_t1_iter33__full_n;
  wire from_t1_iter32_to_t1_iter33__write;
  wire [512:0] from_t1_iter33_to_t1_iter34__dout;
  wire from_t1_iter33_to_t1_iter34__empty_n;
  wire from_t1_iter33_to_t1_iter34__read;
  wire [512:0] from_t1_iter33_to_t1_iter34__din;
  wire from_t1_iter33_to_t1_iter34__full_n;
  wire from_t1_iter33_to_t1_iter34__write;
  wire [512:0] from_t1_iter34_to_t1_iter35__dout;
  wire from_t1_iter34_to_t1_iter35__empty_n;
  wire from_t1_iter34_to_t1_iter35__read;
  wire [512:0] from_t1_iter34_to_t1_iter35__din;
  wire from_t1_iter34_to_t1_iter35__full_n;
  wire from_t1_iter34_to_t1_iter35__write;
  wire [512:0] from_t1_iter35_to_t1_iter36__dout;
  wire from_t1_iter35_to_t1_iter36__empty_n;
  wire from_t1_iter35_to_t1_iter36__read;
  wire [512:0] from_t1_iter35_to_t1_iter36__din;
  wire from_t1_iter35_to_t1_iter36__full_n;
  wire from_t1_iter35_to_t1_iter36__write;
  wire [512:0] from_t1_iter36_to_t1_iter37__dout;
  wire from_t1_iter36_to_t1_iter37__empty_n;
  wire from_t1_iter36_to_t1_iter37__read;
  wire [512:0] from_t1_iter36_to_t1_iter37__din;
  wire from_t1_iter36_to_t1_iter37__full_n;
  wire from_t1_iter36_to_t1_iter37__write;
  wire [512:0] from_t1_iter37_to_t1_iter38__dout;
  wire from_t1_iter37_to_t1_iter38__empty_n;
  wire from_t1_iter37_to_t1_iter38__read;
  wire [512:0] from_t1_iter37_to_t1_iter38__din;
  wire from_t1_iter37_to_t1_iter38__full_n;
  wire from_t1_iter37_to_t1_iter38__write;
  wire [512:0] from_t1_iter38_to_t1_iter39__dout;
  wire from_t1_iter38_to_t1_iter39__empty_n;
  wire from_t1_iter38_to_t1_iter39__read;
  wire [512:0] from_t1_iter38_to_t1_iter39__din;
  wire from_t1_iter38_to_t1_iter39__full_n;
  wire from_t1_iter38_to_t1_iter39__write;
  wire [512:0] from_t1_iter39_to_t1_iter40__dout;
  wire from_t1_iter39_to_t1_iter40__empty_n;
  wire from_t1_iter39_to_t1_iter40__read;
  wire [512:0] from_t1_iter39_to_t1_iter40__din;
  wire from_t1_iter39_to_t1_iter40__full_n;
  wire from_t1_iter39_to_t1_iter40__write;
  wire [512:0] from_t1_iter3_to_t1_iter4__dout;
  wire from_t1_iter3_to_t1_iter4__empty_n;
  wire from_t1_iter3_to_t1_iter4__read;
  wire [512:0] from_t1_iter3_to_t1_iter4__din;
  wire from_t1_iter3_to_t1_iter4__full_n;
  wire from_t1_iter3_to_t1_iter4__write;
  wire [512:0] from_t1_iter40_to_t1_iter41__dout;
  wire from_t1_iter40_to_t1_iter41__empty_n;
  wire from_t1_iter40_to_t1_iter41__read;
  wire [512:0] from_t1_iter40_to_t1_iter41__din;
  wire from_t1_iter40_to_t1_iter41__full_n;
  wire from_t1_iter40_to_t1_iter41__write;
  wire [512:0] from_t1_iter41_to_t1_iter42__dout;
  wire from_t1_iter41_to_t1_iter42__empty_n;
  wire from_t1_iter41_to_t1_iter42__read;
  wire [512:0] from_t1_iter41_to_t1_iter42__din;
  wire from_t1_iter41_to_t1_iter42__full_n;
  wire from_t1_iter41_to_t1_iter42__write;
  wire [512:0] from_t1_iter42_to_t1_iter43__dout;
  wire from_t1_iter42_to_t1_iter43__empty_n;
  wire from_t1_iter42_to_t1_iter43__read;
  wire [512:0] from_t1_iter42_to_t1_iter43__din;
  wire from_t1_iter42_to_t1_iter43__full_n;
  wire from_t1_iter42_to_t1_iter43__write;
  wire [512:0] from_t1_iter43_to_t1_iter44__dout;
  wire from_t1_iter43_to_t1_iter44__empty_n;
  wire from_t1_iter43_to_t1_iter44__read;
  wire [512:0] from_t1_iter43_to_t1_iter44__din;
  wire from_t1_iter43_to_t1_iter44__full_n;
  wire from_t1_iter43_to_t1_iter44__write;
  wire [512:0] from_t1_iter44_to_t1_iter45__dout;
  wire from_t1_iter44_to_t1_iter45__empty_n;
  wire from_t1_iter44_to_t1_iter45__read;
  wire [512:0] from_t1_iter44_to_t1_iter45__din;
  wire from_t1_iter44_to_t1_iter45__full_n;
  wire from_t1_iter44_to_t1_iter45__write;
  wire [512:0] from_t1_iter45_to_t1_iter46__dout;
  wire from_t1_iter45_to_t1_iter46__empty_n;
  wire from_t1_iter45_to_t1_iter46__read;
  wire [512:0] from_t1_iter45_to_t1_iter46__din;
  wire from_t1_iter45_to_t1_iter46__full_n;
  wire from_t1_iter45_to_t1_iter46__write;
  wire [512:0] from_t1_iter46_to_t1_iter47__dout;
  wire from_t1_iter46_to_t1_iter47__empty_n;
  wire from_t1_iter46_to_t1_iter47__read;
  wire [512:0] from_t1_iter46_to_t1_iter47__din;
  wire from_t1_iter46_to_t1_iter47__full_n;
  wire from_t1_iter46_to_t1_iter47__write;
  wire [512:0] from_t1_iter47_to_t1_iter48__dout;
  wire from_t1_iter47_to_t1_iter48__empty_n;
  wire from_t1_iter47_to_t1_iter48__read;
  wire [512:0] from_t1_iter47_to_t1_iter48__din;
  wire from_t1_iter47_to_t1_iter48__full_n;
  wire from_t1_iter47_to_t1_iter48__write;
  wire [512:0] from_t1_iter48_to_t1_iter49__dout;
  wire from_t1_iter48_to_t1_iter49__empty_n;
  wire from_t1_iter48_to_t1_iter49__read;
  wire [512:0] from_t1_iter48_to_t1_iter49__din;
  wire from_t1_iter48_to_t1_iter49__full_n;
  wire from_t1_iter48_to_t1_iter49__write;
  wire [512:0] from_t1_iter49_to_t1_iter50__dout;
  wire from_t1_iter49_to_t1_iter50__empty_n;
  wire from_t1_iter49_to_t1_iter50__read;
  wire [512:0] from_t1_iter49_to_t1_iter50__din;
  wire from_t1_iter49_to_t1_iter50__full_n;
  wire from_t1_iter49_to_t1_iter50__write;
  wire [512:0] from_t1_iter4_to_t1_iter5__dout;
  wire from_t1_iter4_to_t1_iter5__empty_n;
  wire from_t1_iter4_to_t1_iter5__read;
  wire [512:0] from_t1_iter4_to_t1_iter5__din;
  wire from_t1_iter4_to_t1_iter5__full_n;
  wire from_t1_iter4_to_t1_iter5__write;
  wire [512:0] from_t1_iter50_to_t1_iter51__dout;
  wire from_t1_iter50_to_t1_iter51__empty_n;
  wire from_t1_iter50_to_t1_iter51__read;
  wire [512:0] from_t1_iter50_to_t1_iter51__din;
  wire from_t1_iter50_to_t1_iter51__full_n;
  wire from_t1_iter50_to_t1_iter51__write;
  wire [512:0] from_t1_iter51_to_t1_iter52__dout;
  wire from_t1_iter51_to_t1_iter52__empty_n;
  wire from_t1_iter51_to_t1_iter52__read;
  wire [512:0] from_t1_iter51_to_t1_iter52__din;
  wire from_t1_iter51_to_t1_iter52__full_n;
  wire from_t1_iter51_to_t1_iter52__write;
  wire [512:0] from_t1_iter52_to_t1_iter53__dout;
  wire from_t1_iter52_to_t1_iter53__empty_n;
  wire from_t1_iter52_to_t1_iter53__read;
  wire [512:0] from_t1_iter52_to_t1_iter53__din;
  wire from_t1_iter52_to_t1_iter53__full_n;
  wire from_t1_iter52_to_t1_iter53__write;
  wire [512:0] from_t1_iter53_to_t1_iter54__dout;
  wire from_t1_iter53_to_t1_iter54__empty_n;
  wire from_t1_iter53_to_t1_iter54__read;
  wire [512:0] from_t1_iter53_to_t1_iter54__din;
  wire from_t1_iter53_to_t1_iter54__full_n;
  wire from_t1_iter53_to_t1_iter54__write;
  wire [512:0] from_t1_iter54_to_t1_iter55__dout;
  wire from_t1_iter54_to_t1_iter55__empty_n;
  wire from_t1_iter54_to_t1_iter55__read;
  wire [512:0] from_t1_iter54_to_t1_iter55__din;
  wire from_t1_iter54_to_t1_iter55__full_n;
  wire from_t1_iter54_to_t1_iter55__write;
  wire [512:0] from_t1_iter55_to_t1_iter56__dout;
  wire from_t1_iter55_to_t1_iter56__empty_n;
  wire from_t1_iter55_to_t1_iter56__read;
  wire [512:0] from_t1_iter55_to_t1_iter56__din;
  wire from_t1_iter55_to_t1_iter56__full_n;
  wire from_t1_iter55_to_t1_iter56__write;
  wire [512:0] from_t1_iter56_to_t1_iter57__dout;
  wire from_t1_iter56_to_t1_iter57__empty_n;
  wire from_t1_iter56_to_t1_iter57__read;
  wire [512:0] from_t1_iter56_to_t1_iter57__din;
  wire from_t1_iter56_to_t1_iter57__full_n;
  wire from_t1_iter56_to_t1_iter57__write;
  wire [512:0] from_t1_iter57_to_t1_iter58__dout;
  wire from_t1_iter57_to_t1_iter58__empty_n;
  wire from_t1_iter57_to_t1_iter58__read;
  wire [512:0] from_t1_iter57_to_t1_iter58__din;
  wire from_t1_iter57_to_t1_iter58__full_n;
  wire from_t1_iter57_to_t1_iter58__write;
  wire [512:0] from_t1_iter58_to_t1_iter59__dout;
  wire from_t1_iter58_to_t1_iter59__empty_n;
  wire from_t1_iter58_to_t1_iter59__read;
  wire [512:0] from_t1_iter58_to_t1_iter59__din;
  wire from_t1_iter58_to_t1_iter59__full_n;
  wire from_t1_iter58_to_t1_iter59__write;
  wire [512:0] from_t1_iter59_to_t1_iter60__dout;
  wire from_t1_iter59_to_t1_iter60__empty_n;
  wire from_t1_iter59_to_t1_iter60__read;
  wire [512:0] from_t1_iter59_to_t1_iter60__din;
  wire from_t1_iter59_to_t1_iter60__full_n;
  wire from_t1_iter59_to_t1_iter60__write;
  wire [512:0] from_t1_iter5_to_t1_iter6__dout;
  wire from_t1_iter5_to_t1_iter6__empty_n;
  wire from_t1_iter5_to_t1_iter6__read;
  wire [512:0] from_t1_iter5_to_t1_iter6__din;
  wire from_t1_iter5_to_t1_iter6__full_n;
  wire from_t1_iter5_to_t1_iter6__write;
  wire [512:0] from_t1_iter60_to_t1_iter61__dout;
  wire from_t1_iter60_to_t1_iter61__empty_n;
  wire from_t1_iter60_to_t1_iter61__read;
  wire [512:0] from_t1_iter60_to_t1_iter61__din;
  wire from_t1_iter60_to_t1_iter61__full_n;
  wire from_t1_iter60_to_t1_iter61__write;
  wire [512:0] from_t1_iter61_to_t1_iter62__dout;
  wire from_t1_iter61_to_t1_iter62__empty_n;
  wire from_t1_iter61_to_t1_iter62__read;
  wire [512:0] from_t1_iter61_to_t1_iter62__din;
  wire from_t1_iter61_to_t1_iter62__full_n;
  wire from_t1_iter61_to_t1_iter62__write;
  wire [512:0] from_t1_iter62_to_t1_iter63__dout;
  wire from_t1_iter62_to_t1_iter63__empty_n;
  wire from_t1_iter62_to_t1_iter63__read;
  wire [512:0] from_t1_iter62_to_t1_iter63__din;
  wire from_t1_iter62_to_t1_iter63__full_n;
  wire from_t1_iter62_to_t1_iter63__write;
  wire [512:0] from_t1_iter63_to_t1_iter64__dout;
  wire from_t1_iter63_to_t1_iter64__empty_n;
  wire from_t1_iter63_to_t1_iter64__read;
  wire [512:0] from_t1_iter63_to_t1_iter64__din;
  wire from_t1_iter63_to_t1_iter64__full_n;
  wire from_t1_iter63_to_t1_iter64__write;
  wire [512:0] from_t1_iter64_to_t1_iter65__dout;
  wire from_t1_iter64_to_t1_iter65__empty_n;
  wire from_t1_iter64_to_t1_iter65__read;
  wire [512:0] from_t1_iter64_to_t1_iter65__din;
  wire from_t1_iter64_to_t1_iter65__full_n;
  wire from_t1_iter64_to_t1_iter65__write;
  wire [512:0] from_t1_iter65_to_t1_iter66__dout;
  wire from_t1_iter65_to_t1_iter66__empty_n;
  wire from_t1_iter65_to_t1_iter66__read;
  wire [512:0] from_t1_iter65_to_t1_iter66__din;
  wire from_t1_iter65_to_t1_iter66__full_n;
  wire from_t1_iter65_to_t1_iter66__write;
  wire [512:0] from_t1_iter66_to_t1_iter67__dout;
  wire from_t1_iter66_to_t1_iter67__empty_n;
  wire from_t1_iter66_to_t1_iter67__read;
  wire [512:0] from_t1_iter66_to_t1_iter67__din;
  wire from_t1_iter66_to_t1_iter67__full_n;
  wire from_t1_iter66_to_t1_iter67__write;
  wire [512:0] from_t1_iter67_to_t1_iter68__dout;
  wire from_t1_iter67_to_t1_iter68__empty_n;
  wire from_t1_iter67_to_t1_iter68__read;
  wire [512:0] from_t1_iter67_to_t1_iter68__din;
  wire from_t1_iter67_to_t1_iter68__full_n;
  wire from_t1_iter67_to_t1_iter68__write;
  wire [512:0] from_t1_iter68_to_t1_iter69__dout;
  wire from_t1_iter68_to_t1_iter69__empty_n;
  wire from_t1_iter68_to_t1_iter69__read;
  wire [512:0] from_t1_iter68_to_t1_iter69__din;
  wire from_t1_iter68_to_t1_iter69__full_n;
  wire from_t1_iter68_to_t1_iter69__write;
  wire [512:0] from_t1_iter69_to_t1_iter70__dout;
  wire from_t1_iter69_to_t1_iter70__empty_n;
  wire from_t1_iter69_to_t1_iter70__read;
  wire [512:0] from_t1_iter69_to_t1_iter70__din;
  wire from_t1_iter69_to_t1_iter70__full_n;
  wire from_t1_iter69_to_t1_iter70__write;
  wire [512:0] from_t1_iter6_to_t1_iter7__dout;
  wire from_t1_iter6_to_t1_iter7__empty_n;
  wire from_t1_iter6_to_t1_iter7__read;
  wire [512:0] from_t1_iter6_to_t1_iter7__din;
  wire from_t1_iter6_to_t1_iter7__full_n;
  wire from_t1_iter6_to_t1_iter7__write;
  wire [512:0] from_t1_iter70_to_t1_iter71__dout;
  wire from_t1_iter70_to_t1_iter71__empty_n;
  wire from_t1_iter70_to_t1_iter71__read;
  wire [512:0] from_t1_iter70_to_t1_iter71__din;
  wire from_t1_iter70_to_t1_iter71__full_n;
  wire from_t1_iter70_to_t1_iter71__write;
  wire [512:0] from_t1_iter71_to_t1_iter72__dout;
  wire from_t1_iter71_to_t1_iter72__empty_n;
  wire from_t1_iter71_to_t1_iter72__read;
  wire [512:0] from_t1_iter71_to_t1_iter72__din;
  wire from_t1_iter71_to_t1_iter72__full_n;
  wire from_t1_iter71_to_t1_iter72__write;
  wire [512:0] from_t1_iter72_to_t1_iter73__dout;
  wire from_t1_iter72_to_t1_iter73__empty_n;
  wire from_t1_iter72_to_t1_iter73__read;
  wire [512:0] from_t1_iter72_to_t1_iter73__din;
  wire from_t1_iter72_to_t1_iter73__full_n;
  wire from_t1_iter72_to_t1_iter73__write;
  wire [512:0] from_t1_iter73_to_t1_iter74__dout;
  wire from_t1_iter73_to_t1_iter74__empty_n;
  wire from_t1_iter73_to_t1_iter74__read;
  wire [512:0] from_t1_iter73_to_t1_iter74__din;
  wire from_t1_iter73_to_t1_iter74__full_n;
  wire from_t1_iter73_to_t1_iter74__write;
  wire [512:0] from_t1_iter74_to_t1_iter75__dout;
  wire from_t1_iter74_to_t1_iter75__empty_n;
  wire from_t1_iter74_to_t1_iter75__read;
  wire [512:0] from_t1_iter74_to_t1_iter75__din;
  wire from_t1_iter74_to_t1_iter75__full_n;
  wire from_t1_iter74_to_t1_iter75__write;
  wire [512:0] from_t1_iter75_to_t1_iter76__dout;
  wire from_t1_iter75_to_t1_iter76__empty_n;
  wire from_t1_iter75_to_t1_iter76__read;
  wire [512:0] from_t1_iter75_to_t1_iter76__din;
  wire from_t1_iter75_to_t1_iter76__full_n;
  wire from_t1_iter75_to_t1_iter76__write;
  wire [512:0] from_t1_iter76_to_t1_iter77__dout;
  wire from_t1_iter76_to_t1_iter77__empty_n;
  wire from_t1_iter76_to_t1_iter77__read;
  wire [512:0] from_t1_iter76_to_t1_iter77__din;
  wire from_t1_iter76_to_t1_iter77__full_n;
  wire from_t1_iter76_to_t1_iter77__write;
  wire [512:0] from_t1_iter77_to_t1_iter78__dout;
  wire from_t1_iter77_to_t1_iter78__empty_n;
  wire from_t1_iter77_to_t1_iter78__read;
  wire [512:0] from_t1_iter77_to_t1_iter78__din;
  wire from_t1_iter77_to_t1_iter78__full_n;
  wire from_t1_iter77_to_t1_iter78__write;
  wire [512:0] from_t1_iter78_to_t1_iter79__dout;
  wire from_t1_iter78_to_t1_iter79__empty_n;
  wire from_t1_iter78_to_t1_iter79__read;
  wire [512:0] from_t1_iter78_to_t1_iter79__din;
  wire from_t1_iter78_to_t1_iter79__full_n;
  wire from_t1_iter78_to_t1_iter79__write;
  wire [512:0] from_t1_iter79_to_t1_iter80__dout;
  wire from_t1_iter79_to_t1_iter80__empty_n;
  wire from_t1_iter79_to_t1_iter80__read;
  wire [512:0] from_t1_iter79_to_t1_iter80__din;
  wire from_t1_iter79_to_t1_iter80__full_n;
  wire from_t1_iter79_to_t1_iter80__write;
  wire [512:0] from_t1_iter7_to_t1_iter8__dout;
  wire from_t1_iter7_to_t1_iter8__empty_n;
  wire from_t1_iter7_to_t1_iter8__read;
  wire [512:0] from_t1_iter7_to_t1_iter8__din;
  wire from_t1_iter7_to_t1_iter8__full_n;
  wire from_t1_iter7_to_t1_iter8__write;
  wire [512:0] from_t1_iter80_to_t1_iter81__dout;
  wire from_t1_iter80_to_t1_iter81__empty_n;
  wire from_t1_iter80_to_t1_iter81__read;
  wire [512:0] from_t1_iter80_to_t1_iter81__din;
  wire from_t1_iter80_to_t1_iter81__full_n;
  wire from_t1_iter80_to_t1_iter81__write;
  wire [512:0] from_t1_iter81_to_t1_iter82__dout;
  wire from_t1_iter81_to_t1_iter82__empty_n;
  wire from_t1_iter81_to_t1_iter82__read;
  wire [512:0] from_t1_iter81_to_t1_iter82__din;
  wire from_t1_iter81_to_t1_iter82__full_n;
  wire from_t1_iter81_to_t1_iter82__write;
  wire [512:0] from_t1_iter82_to_t1_iter83__dout;
  wire from_t1_iter82_to_t1_iter83__empty_n;
  wire from_t1_iter82_to_t1_iter83__read;
  wire [512:0] from_t1_iter82_to_t1_iter83__din;
  wire from_t1_iter82_to_t1_iter83__full_n;
  wire from_t1_iter82_to_t1_iter83__write;
  wire [512:0] from_t1_iter83_to_t1_iter84__dout;
  wire from_t1_iter83_to_t1_iter84__empty_n;
  wire from_t1_iter83_to_t1_iter84__read;
  wire [512:0] from_t1_iter83_to_t1_iter84__din;
  wire from_t1_iter83_to_t1_iter84__full_n;
  wire from_t1_iter83_to_t1_iter84__write;
  wire [512:0] from_t1_iter84_to_t1_iter85__dout;
  wire from_t1_iter84_to_t1_iter85__empty_n;
  wire from_t1_iter84_to_t1_iter85__read;
  wire [512:0] from_t1_iter84_to_t1_iter85__din;
  wire from_t1_iter84_to_t1_iter85__full_n;
  wire from_t1_iter84_to_t1_iter85__write;
  wire [512:0] from_t1_iter85_to_t1_iter86__dout;
  wire from_t1_iter85_to_t1_iter86__empty_n;
  wire from_t1_iter85_to_t1_iter86__read;
  wire [512:0] from_t1_iter85_to_t1_iter86__din;
  wire from_t1_iter85_to_t1_iter86__full_n;
  wire from_t1_iter85_to_t1_iter86__write;
  wire [512:0] from_t1_iter86_to_t1_iter87__dout;
  wire from_t1_iter86_to_t1_iter87__empty_n;
  wire from_t1_iter86_to_t1_iter87__read;
  wire [512:0] from_t1_iter86_to_t1_iter87__din;
  wire from_t1_iter86_to_t1_iter87__full_n;
  wire from_t1_iter86_to_t1_iter87__write;
  wire [512:0] from_t1_iter87_to_t1_iter88__dout;
  wire from_t1_iter87_to_t1_iter88__empty_n;
  wire from_t1_iter87_to_t1_iter88__read;
  wire [512:0] from_t1_iter87_to_t1_iter88__din;
  wire from_t1_iter87_to_t1_iter88__full_n;
  wire from_t1_iter87_to_t1_iter88__write;
  wire [512:0] from_t1_iter88_to_t1_iter89__dout;
  wire from_t1_iter88_to_t1_iter89__empty_n;
  wire from_t1_iter88_to_t1_iter89__read;
  wire [512:0] from_t1_iter88_to_t1_iter89__din;
  wire from_t1_iter88_to_t1_iter89__full_n;
  wire from_t1_iter88_to_t1_iter89__write;
  wire [512:0] from_t1_iter89_to_t1_iter90__dout;
  wire from_t1_iter89_to_t1_iter90__empty_n;
  wire from_t1_iter89_to_t1_iter90__read;
  wire [512:0] from_t1_iter89_to_t1_iter90__din;
  wire from_t1_iter89_to_t1_iter90__full_n;
  wire from_t1_iter89_to_t1_iter90__write;
  wire [512:0] from_t1_iter8_to_t1_iter9__dout;
  wire from_t1_iter8_to_t1_iter9__empty_n;
  wire from_t1_iter8_to_t1_iter9__read;
  wire [512:0] from_t1_iter8_to_t1_iter9__din;
  wire from_t1_iter8_to_t1_iter9__full_n;
  wire from_t1_iter8_to_t1_iter9__write;
  wire [512:0] from_t1_iter90_to_t1_iter91__dout;
  wire from_t1_iter90_to_t1_iter91__empty_n;
  wire from_t1_iter90_to_t1_iter91__read;
  wire [512:0] from_t1_iter90_to_t1_iter91__din;
  wire from_t1_iter90_to_t1_iter91__full_n;
  wire from_t1_iter90_to_t1_iter91__write;
  wire [512:0] from_t1_iter91_to_t1_iter92__dout;
  wire from_t1_iter91_to_t1_iter92__empty_n;
  wire from_t1_iter91_to_t1_iter92__read;
  wire [512:0] from_t1_iter91_to_t1_iter92__din;
  wire from_t1_iter91_to_t1_iter92__full_n;
  wire from_t1_iter91_to_t1_iter92__write;
  wire [512:0] from_t1_iter92_to_t1_iter93__dout;
  wire from_t1_iter92_to_t1_iter93__empty_n;
  wire from_t1_iter92_to_t1_iter93__read;
  wire [512:0] from_t1_iter92_to_t1_iter93__din;
  wire from_t1_iter92_to_t1_iter93__full_n;
  wire from_t1_iter92_to_t1_iter93__write;
  wire [512:0] from_t1_iter93_to_t1_iter94__dout;
  wire from_t1_iter93_to_t1_iter94__empty_n;
  wire from_t1_iter93_to_t1_iter94__read;
  wire [512:0] from_t1_iter93_to_t1_iter94__din;
  wire from_t1_iter93_to_t1_iter94__full_n;
  wire from_t1_iter93_to_t1_iter94__write;
  wire [512:0] from_t1_iter94_to_t1_iter95__dout;
  wire from_t1_iter94_to_t1_iter95__empty_n;
  wire from_t1_iter94_to_t1_iter95__read;
  wire [512:0] from_t1_iter94_to_t1_iter95__din;
  wire from_t1_iter94_to_t1_iter95__full_n;
  wire from_t1_iter94_to_t1_iter95__write;
  wire [512:0] from_t1_iter95_to_t1_iter96__dout;
  wire from_t1_iter95_to_t1_iter96__empty_n;
  wire from_t1_iter95_to_t1_iter96__read;
  wire [512:0] from_t1_iter95_to_t1_iter96__din;
  wire from_t1_iter95_to_t1_iter96__full_n;
  wire from_t1_iter95_to_t1_iter96__write;
  wire [512:0] from_t1_iter96_to_t1_iter97__dout;
  wire from_t1_iter96_to_t1_iter97__empty_n;
  wire from_t1_iter96_to_t1_iter97__read;
  wire [512:0] from_t1_iter96_to_t1_iter97__din;
  wire from_t1_iter96_to_t1_iter97__full_n;
  wire from_t1_iter96_to_t1_iter97__write;
  wire [512:0] from_t1_iter97_to_t1_iter98__dout;
  wire from_t1_iter97_to_t1_iter98__empty_n;
  wire from_t1_iter97_to_t1_iter98__read;
  wire [512:0] from_t1_iter97_to_t1_iter98__din;
  wire from_t1_iter97_to_t1_iter98__full_n;
  wire from_t1_iter97_to_t1_iter98__write;
  wire [512:0] from_t1_iter98_to_t1_iter99__dout;
  wire from_t1_iter98_to_t1_iter99__empty_n;
  wire from_t1_iter98_to_t1_iter99__read;
  wire [512:0] from_t1_iter98_to_t1_iter99__din;
  wire from_t1_iter98_to_t1_iter99__full_n;
  wire from_t1_iter98_to_t1_iter99__write;
  wire [512:0] from_t1_iter99_to_t1_iter100__dout;
  wire from_t1_iter99_to_t1_iter100__empty_n;
  wire from_t1_iter99_to_t1_iter100__read;
  wire [512:0] from_t1_iter99_to_t1_iter100__din;
  wire from_t1_iter99_to_t1_iter100__full_n;
  wire from_t1_iter99_to_t1_iter100__write;
  wire [512:0] from_t1_iter9_to_t1_iter10__dout;
  wire from_t1_iter9_to_t1_iter10__empty_n;
  wire from_t1_iter9_to_t1_iter10__read;
  wire [512:0] from_t1_iter9_to_t1_iter10__din;
  wire from_t1_iter9_to_t1_iter10__full_n;
  wire from_t1_iter9_to_t1_iter10__write;
  wire [63:0] BurstRead_floatx16_0___bank_0_t1__q0;
  wire [63:0] bank_0_t1_read_addr__din;
  wire bank_0_t1_read_addr__full_n;
  wire bank_0_t1_read_addr__write;
  wire [511:0] bank_0_t1_read_data__dout;
  wire bank_0_t1_read_data__empty_n;
  wire bank_0_t1_read_data__read;
  wire [63:0] bank_0_t1_write_addr__din;
  wire bank_0_t1_write_addr__full_n;
  wire bank_0_t1_write_addr__write;
  wire [511:0] bank_0_t1_write_data__din;
  wire bank_0_t1_write_data__full_n;
  wire bank_0_t1_write_data__write;
  wire [7:0] bank_0_t1_write_resp__dout;
  wire bank_0_t1_write_resp__empty_n;
  wire bank_0_t1_write_resp__read;
  wire [63:0] BurstRead_floatx16_0___coalesced_data_num__q0;
  wire BurstRead_floatx16_0__ap_start;
  wire BurstRead_floatx16_0__ap_ready;
  wire BurstRead_floatx16_0__ap_done;
  wire BurstRead_floatx16_0__ap_idle;
  wire [63:0] BurstWrite_floatx16_0___bank_1_t0__q0;
  wire [63:0] bank_1_t0_read_addr__din;
  wire bank_1_t0_read_addr__full_n;
  wire bank_1_t0_read_addr__write;
  wire [511:0] bank_1_t0_read_data__dout;
  wire bank_1_t0_read_data__empty_n;
  wire bank_1_t0_read_data__read;
  wire [63:0] bank_1_t0_write_addr__din;
  wire bank_1_t0_write_addr__full_n;
  wire bank_1_t0_write_addr__write;
  wire [511:0] bank_1_t0_write_data__din;
  wire bank_1_t0_write_data__full_n;
  wire bank_1_t0_write_data__write;
  wire [7:0] bank_1_t0_write_resp__dout;
  wire bank_1_t0_write_resp__empty_n;
  wire bank_1_t0_write_resp__read;
  wire [63:0] BurstWrite_floatx16_0___coalesced_data_num__q0;
  wire BurstWrite_floatx16_0__ap_start;
  wire BurstWrite_floatx16_0__ap_ready;
  wire BurstWrite_floatx16_0__ap_done;
  wire BurstWrite_floatx16_0__ap_idle;
  wire Module0Func_0__ap_start;
  wire Module1Func_0__ap_start;
  wire Module2Func_0__ap_start;
  wire Module2Func_1__ap_start;
  wire Module2Func_2__ap_start;
  wire Module2Func_3__ap_start;
  wire Module2Func_4__ap_start;
  wire Module2Func_5__ap_start;
  wire Module2Func_6__ap_start;
  wire Module2Func_7__ap_start;
  wire Module2Func_8__ap_start;
  wire Module2Func_9__ap_start;
  wire Module2Func_10__ap_start;
  wire Module2Func_11__ap_start;
  wire Module2Func_12__ap_start;
  wire Module2Func_13__ap_start;
  wire Module2Func_14__ap_start;
  wire Module2Func_15__ap_start;
  wire Module2Func_16__ap_start;
  wire Module2Func_17__ap_start;
  wire Module2Func_18__ap_start;
  wire Module2Func_19__ap_start;
  wire Module2Func_20__ap_start;
  wire Module2Func_21__ap_start;
  wire Module2Func_22__ap_start;
  wire Module2Func_23__ap_start;
  wire Module2Func_24__ap_start;
  wire Module2Func_25__ap_start;
  wire Module2Func_26__ap_start;
  wire Module2Func_27__ap_start;
  wire Module2Func_28__ap_start;
  wire Module2Func_29__ap_start;
  wire Module2Func_30__ap_start;
  wire Module2Func_31__ap_start;
  wire Module2Func_32__ap_start;
  wire Module2Func_33__ap_start;
  wire Module2Func_34__ap_start;
  wire Module2Func_35__ap_start;
  wire Module2Func_36__ap_start;
  wire Module2Func_37__ap_start;
  wire Module2Func_38__ap_start;
  wire Module2Func_39__ap_start;
  wire Module2Func_40__ap_start;
  wire Module2Func_41__ap_start;
  wire Module2Func_42__ap_start;
  wire Module2Func_43__ap_start;
  wire Module2Func_44__ap_start;
  wire Module2Func_45__ap_start;
  wire Module2Func_46__ap_start;
  wire Module2Func_47__ap_start;
  wire Module2Func_48__ap_start;
  wire Module2Func_49__ap_start;
  wire Module2Func_50__ap_start;
  wire Module2Func_51__ap_start;
  wire Module2Func_52__ap_start;
  wire Module2Func_53__ap_start;
  wire Module2Func_54__ap_start;
  wire Module2Func_55__ap_start;
  wire Module2Func_56__ap_start;
  wire Module2Func_57__ap_start;
  wire Module2Func_58__ap_start;
  wire Module2Func_59__ap_start;
  wire Module2Func_60__ap_start;
  wire Module2Func_61__ap_start;
  wire Module2Func_62__ap_start;
  wire Module2Func_63__ap_start;
  wire Module2Func_64__ap_start;
  wire Module2Func_65__ap_start;
  wire Module2Func_66__ap_start;
  wire Module2Func_67__ap_start;
  wire Module2Func_68__ap_start;
  wire Module2Func_69__ap_start;
  wire Module2Func_70__ap_start;
  wire Module2Func_71__ap_start;
  wire Module2Func_72__ap_start;
  wire Module2Func_73__ap_start;
  wire Module2Func_74__ap_start;
  wire Module2Func_75__ap_start;
  wire Module2Func_76__ap_start;
  wire Module2Func_77__ap_start;
  wire Module2Func_78__ap_start;
  wire Module2Func_79__ap_start;
  wire Module2Func_80__ap_start;
  wire Module2Func_81__ap_start;
  wire Module2Func_82__ap_start;
  wire Module2Func_83__ap_start;
  wire Module2Func_84__ap_start;
  wire Module2Func_85__ap_start;
  wire Module2Func_86__ap_start;
  wire Module2Func_87__ap_start;
  wire Module2Func_88__ap_start;
  wire Module2Func_89__ap_start;
  wire Module2Func_90__ap_start;
  wire Module2Func_91__ap_start;
  wire Module2Func_92__ap_start;
  wire Module2Func_93__ap_start;
  wire Module2Func_94__ap_start;
  wire Module2Func_95__ap_start;
  wire Module2Func_96__ap_start;
  wire Module2Func_97__ap_start;
  wire Module2Func_98__ap_start;
  wire Module2Func_99__ap_start;
  wire Module2Func_100__ap_start;
  wire Module2Func_101__ap_start;
  wire Module2Func_102__ap_start;
  wire Module2Func_103__ap_start;
  wire Module2Func_104__ap_start;
  wire Module2Func_105__ap_start;
  wire Module2Func_106__ap_start;
  wire Module2Func_107__ap_start;
  wire Module3Func_0__ap_start;
  wire ap_rst_n_inv;
  wire ap_done;
  wire ap_idle;
  wire ap_ready;
  assign ap_rst_n_inv = (~ap_rst_n);
  assign control_s_axi_U_ACLK = ap_clk;
  assign control_s_axi_U_ACLK_EN = 1'b1;
  assign control_s_axi_U_ARADDR = s_axi_control_ARADDR;
  assign control_s_axi_U_ARESET = ap_rst_n_inv;
  assign s_axi_control_ARREADY = control_s_axi_U_ARREADY;
  assign control_s_axi_U_ARVALID = s_axi_control_ARVALID;
  assign control_s_axi_U_AWADDR = s_axi_control_AWADDR;
  assign s_axi_control_AWREADY = control_s_axi_U_AWREADY;
  assign control_s_axi_U_AWVALID = s_axi_control_AWVALID;
  assign control_s_axi_U_BREADY = s_axi_control_BREADY;
  assign s_axi_control_BRESP = control_s_axi_U_BRESP;
  assign s_axi_control_BVALID = control_s_axi_U_BVALID;
  assign s_axi_control_RDATA = control_s_axi_U_RDATA;
  assign control_s_axi_U_RREADY = s_axi_control_RREADY;
  assign s_axi_control_RRESP = control_s_axi_U_RRESP;
  assign s_axi_control_RVALID = control_s_axi_U_RVALID;
  assign control_s_axi_U_WDATA = s_axi_control_WDATA;
  assign s_axi_control_WREADY = control_s_axi_U_WREADY;
  assign control_s_axi_U_WSTRB = s_axi_control_WSTRB;
  assign control_s_axi_U_WVALID = s_axi_control_WVALID;
  assign control_s_axi_U_ap_done = ap_done;
  assign control_s_axi_U_ap_idle = ap_idle;
  assign control_s_axi_U_ap_ready = ap_ready;
  assign ap_start = control_s_axi_U_ap_start;
  assign bank_0_t1 = control_s_axi_U_bank_0_t1;
  assign bank_1_t0 = control_s_axi_U_bank_1_t0;
  assign coalesced_data_num = control_s_axi_U_coalesced_data_num;
  assign interrupt = control_s_axi_U_interrupt;
  assign bank_0_t1_buf_clk = ap_clk;
  assign bank_0_t1_buf_if_din = bank_0_t1_buf__din;
  assign bank_0_t1_buf__dout = bank_0_t1_buf_if_dout;
  assign bank_0_t1_buf__empty_n = bank_0_t1_buf_if_empty_n;
  assign bank_0_t1_buf__full_n = bank_0_t1_buf_if_full_n;
  assign bank_0_t1_buf_if_read = bank_0_t1_buf__read;
  assign bank_0_t1_buf_if_read_ce = 1'b1;
  assign bank_0_t1_buf_if_write = bank_0_t1_buf__write;
  assign bank_0_t1_buf_if_write_ce = 1'b1;
  assign bank_0_t1_buf_reset = ~ ap_rst_n;
  assign bank_1_t0_buf_clk = ap_clk;
  assign bank_1_t0_buf_if_din = bank_1_t0_buf__din;
  assign bank_1_t0_buf__dout = bank_1_t0_buf_if_dout;
  assign bank_1_t0_buf__empty_n = bank_1_t0_buf_if_empty_n;
  assign bank_1_t0_buf__full_n = bank_1_t0_buf_if_full_n;
  assign bank_1_t0_buf_if_read = bank_1_t0_buf__read;
  assign bank_1_t0_buf_if_read_ce = 1'b1;
  assign bank_1_t0_buf_if_write = bank_1_t0_buf__write;
  assign bank_1_t0_buf_if_write_ce = 1'b1;
  assign bank_1_t0_buf_reset = ~ ap_rst_n;
  assign from_t0_to_t0_bank_1_clk = ap_clk;
  assign from_t0_to_t0_bank_1_if_din = from_t0_to_t0_bank_1__din;
  assign from_t0_to_t0_bank_1__dout = from_t0_to_t0_bank_1_if_dout;
  assign from_t0_to_t0_bank_1__empty_n = from_t0_to_t0_bank_1_if_empty_n;
  assign from_t0_to_t0_bank_1__full_n = from_t0_to_t0_bank_1_if_full_n;
  assign from_t0_to_t0_bank_1_if_read = from_t0_to_t0_bank_1__read;
  assign from_t0_to_t0_bank_1_if_read_ce = 1'b1;
  assign from_t0_to_t0_bank_1_if_write = from_t0_to_t0_bank_1__write;
  assign from_t0_to_t0_bank_1_if_write_ce = 1'b1;
  assign from_t0_to_t0_bank_1_reset = ~ ap_rst_n;
  assign from_t1_bank_0_to_t1_iter1_clk = ap_clk;
  assign from_t1_bank_0_to_t1_iter1_if_din = from_t1_bank_0_to_t1_iter1__din;
  assign from_t1_bank_0_to_t1_iter1__dout = from_t1_bank_0_to_t1_iter1_if_dout;
  assign from_t1_bank_0_to_t1_iter1__empty_n = from_t1_bank_0_to_t1_iter1_if_empty_n;
  assign from_t1_bank_0_to_t1_iter1__full_n = from_t1_bank_0_to_t1_iter1_if_full_n;
  assign from_t1_bank_0_to_t1_iter1_if_read = from_t1_bank_0_to_t1_iter1__read;
  assign from_t1_bank_0_to_t1_iter1_if_read_ce = 1'b1;
  assign from_t1_bank_0_to_t1_iter1_if_write = from_t1_bank_0_to_t1_iter1__write;
  assign from_t1_bank_0_to_t1_iter1_if_write_ce = 1'b1;
  assign from_t1_bank_0_to_t1_iter1_reset = ~ ap_rst_n;
  assign from_t1_iter100_to_t1_iter101_clk = ap_clk;
  assign from_t1_iter100_to_t1_iter101_if_din = from_t1_iter100_to_t1_iter101__din;
  assign from_t1_iter100_to_t1_iter101__dout = from_t1_iter100_to_t1_iter101_if_dout;
  assign from_t1_iter100_to_t1_iter101__empty_n = from_t1_iter100_to_t1_iter101_if_empty_n;
  assign from_t1_iter100_to_t1_iter101__full_n = from_t1_iter100_to_t1_iter101_if_full_n;
  assign from_t1_iter100_to_t1_iter101_if_read = from_t1_iter100_to_t1_iter101__read;
  assign from_t1_iter100_to_t1_iter101_if_read_ce = 1'b1;
  assign from_t1_iter100_to_t1_iter101_if_write = from_t1_iter100_to_t1_iter101__write;
  assign from_t1_iter100_to_t1_iter101_if_write_ce = 1'b1;
  assign from_t1_iter100_to_t1_iter101_reset = ~ ap_rst_n;
  assign from_t1_iter101_to_t1_iter102_clk = ap_clk;
  assign from_t1_iter101_to_t1_iter102_if_din = from_t1_iter101_to_t1_iter102__din;
  assign from_t1_iter101_to_t1_iter102__dout = from_t1_iter101_to_t1_iter102_if_dout;
  assign from_t1_iter101_to_t1_iter102__empty_n = from_t1_iter101_to_t1_iter102_if_empty_n;
  assign from_t1_iter101_to_t1_iter102__full_n = from_t1_iter101_to_t1_iter102_if_full_n;
  assign from_t1_iter101_to_t1_iter102_if_read = from_t1_iter101_to_t1_iter102__read;
  assign from_t1_iter101_to_t1_iter102_if_read_ce = 1'b1;
  assign from_t1_iter101_to_t1_iter102_if_write = from_t1_iter101_to_t1_iter102__write;
  assign from_t1_iter101_to_t1_iter102_if_write_ce = 1'b1;
  assign from_t1_iter101_to_t1_iter102_reset = ~ ap_rst_n;
  assign from_t1_iter102_to_t1_iter103_clk = ap_clk;
  assign from_t1_iter102_to_t1_iter103_if_din = from_t1_iter102_to_t1_iter103__din;
  assign from_t1_iter102_to_t1_iter103__dout = from_t1_iter102_to_t1_iter103_if_dout;
  assign from_t1_iter102_to_t1_iter103__empty_n = from_t1_iter102_to_t1_iter103_if_empty_n;
  assign from_t1_iter102_to_t1_iter103__full_n = from_t1_iter102_to_t1_iter103_if_full_n;
  assign from_t1_iter102_to_t1_iter103_if_read = from_t1_iter102_to_t1_iter103__read;
  assign from_t1_iter102_to_t1_iter103_if_read_ce = 1'b1;
  assign from_t1_iter102_to_t1_iter103_if_write = from_t1_iter102_to_t1_iter103__write;
  assign from_t1_iter102_to_t1_iter103_if_write_ce = 1'b1;
  assign from_t1_iter102_to_t1_iter103_reset = ~ ap_rst_n;
  assign from_t1_iter103_to_t1_iter104_clk = ap_clk;
  assign from_t1_iter103_to_t1_iter104_if_din = from_t1_iter103_to_t1_iter104__din;
  assign from_t1_iter103_to_t1_iter104__dout = from_t1_iter103_to_t1_iter104_if_dout;
  assign from_t1_iter103_to_t1_iter104__empty_n = from_t1_iter103_to_t1_iter104_if_empty_n;
  assign from_t1_iter103_to_t1_iter104__full_n = from_t1_iter103_to_t1_iter104_if_full_n;
  assign from_t1_iter103_to_t1_iter104_if_read = from_t1_iter103_to_t1_iter104__read;
  assign from_t1_iter103_to_t1_iter104_if_read_ce = 1'b1;
  assign from_t1_iter103_to_t1_iter104_if_write = from_t1_iter103_to_t1_iter104__write;
  assign from_t1_iter103_to_t1_iter104_if_write_ce = 1'b1;
  assign from_t1_iter103_to_t1_iter104_reset = ~ ap_rst_n;
  assign from_t1_iter104_to_t1_iter105_clk = ap_clk;
  assign from_t1_iter104_to_t1_iter105_if_din = from_t1_iter104_to_t1_iter105__din;
  assign from_t1_iter104_to_t1_iter105__dout = from_t1_iter104_to_t1_iter105_if_dout;
  assign from_t1_iter104_to_t1_iter105__empty_n = from_t1_iter104_to_t1_iter105_if_empty_n;
  assign from_t1_iter104_to_t1_iter105__full_n = from_t1_iter104_to_t1_iter105_if_full_n;
  assign from_t1_iter104_to_t1_iter105_if_read = from_t1_iter104_to_t1_iter105__read;
  assign from_t1_iter104_to_t1_iter105_if_read_ce = 1'b1;
  assign from_t1_iter104_to_t1_iter105_if_write = from_t1_iter104_to_t1_iter105__write;
  assign from_t1_iter104_to_t1_iter105_if_write_ce = 1'b1;
  assign from_t1_iter104_to_t1_iter105_reset = ~ ap_rst_n;
  assign from_t1_iter105_to_t1_iter106_clk = ap_clk;
  assign from_t1_iter105_to_t1_iter106_if_din = from_t1_iter105_to_t1_iter106__din;
  assign from_t1_iter105_to_t1_iter106__dout = from_t1_iter105_to_t1_iter106_if_dout;
  assign from_t1_iter105_to_t1_iter106__empty_n = from_t1_iter105_to_t1_iter106_if_empty_n;
  assign from_t1_iter105_to_t1_iter106__full_n = from_t1_iter105_to_t1_iter106_if_full_n;
  assign from_t1_iter105_to_t1_iter106_if_read = from_t1_iter105_to_t1_iter106__read;
  assign from_t1_iter105_to_t1_iter106_if_read_ce = 1'b1;
  assign from_t1_iter105_to_t1_iter106_if_write = from_t1_iter105_to_t1_iter106__write;
  assign from_t1_iter105_to_t1_iter106_if_write_ce = 1'b1;
  assign from_t1_iter105_to_t1_iter106_reset = ~ ap_rst_n;
  assign from_t1_iter106_to_t1_iter107_clk = ap_clk;
  assign from_t1_iter106_to_t1_iter107_if_din = from_t1_iter106_to_t1_iter107__din;
  assign from_t1_iter106_to_t1_iter107__dout = from_t1_iter106_to_t1_iter107_if_dout;
  assign from_t1_iter106_to_t1_iter107__empty_n = from_t1_iter106_to_t1_iter107_if_empty_n;
  assign from_t1_iter106_to_t1_iter107__full_n = from_t1_iter106_to_t1_iter107_if_full_n;
  assign from_t1_iter106_to_t1_iter107_if_read = from_t1_iter106_to_t1_iter107__read;
  assign from_t1_iter106_to_t1_iter107_if_read_ce = 1'b1;
  assign from_t1_iter106_to_t1_iter107_if_write = from_t1_iter106_to_t1_iter107__write;
  assign from_t1_iter106_to_t1_iter107_if_write_ce = 1'b1;
  assign from_t1_iter106_to_t1_iter107_reset = ~ ap_rst_n;
  assign from_t1_iter107_to_t1_iter108_clk = ap_clk;
  assign from_t1_iter107_to_t1_iter108_if_din = from_t1_iter107_to_t1_iter108__din;
  assign from_t1_iter107_to_t1_iter108__dout = from_t1_iter107_to_t1_iter108_if_dout;
  assign from_t1_iter107_to_t1_iter108__empty_n = from_t1_iter107_to_t1_iter108_if_empty_n;
  assign from_t1_iter107_to_t1_iter108__full_n = from_t1_iter107_to_t1_iter108_if_full_n;
  assign from_t1_iter107_to_t1_iter108_if_read = from_t1_iter107_to_t1_iter108__read;
  assign from_t1_iter107_to_t1_iter108_if_read_ce = 1'b1;
  assign from_t1_iter107_to_t1_iter108_if_write = from_t1_iter107_to_t1_iter108__write;
  assign from_t1_iter107_to_t1_iter108_if_write_ce = 1'b1;
  assign from_t1_iter107_to_t1_iter108_reset = ~ ap_rst_n;
  assign from_t1_iter108_to_t0_clk = ap_clk;
  assign from_t1_iter108_to_t0_if_din = from_t1_iter108_to_t0__din;
  assign from_t1_iter108_to_t0__dout = from_t1_iter108_to_t0_if_dout;
  assign from_t1_iter108_to_t0__empty_n = from_t1_iter108_to_t0_if_empty_n;
  assign from_t1_iter108_to_t0__full_n = from_t1_iter108_to_t0_if_full_n;
  assign from_t1_iter108_to_t0_if_read = from_t1_iter108_to_t0__read;
  assign from_t1_iter108_to_t0_if_read_ce = 1'b1;
  assign from_t1_iter108_to_t0_if_write = from_t1_iter108_to_t0__write;
  assign from_t1_iter108_to_t0_if_write_ce = 1'b1;
  assign from_t1_iter108_to_t0_reset = ~ ap_rst_n;
  assign from_t1_iter10_to_t1_iter11_clk = ap_clk;
  assign from_t1_iter10_to_t1_iter11_if_din = from_t1_iter10_to_t1_iter11__din;
  assign from_t1_iter10_to_t1_iter11__dout = from_t1_iter10_to_t1_iter11_if_dout;
  assign from_t1_iter10_to_t1_iter11__empty_n = from_t1_iter10_to_t1_iter11_if_empty_n;
  assign from_t1_iter10_to_t1_iter11__full_n = from_t1_iter10_to_t1_iter11_if_full_n;
  assign from_t1_iter10_to_t1_iter11_if_read = from_t1_iter10_to_t1_iter11__read;
  assign from_t1_iter10_to_t1_iter11_if_read_ce = 1'b1;
  assign from_t1_iter10_to_t1_iter11_if_write = from_t1_iter10_to_t1_iter11__write;
  assign from_t1_iter10_to_t1_iter11_if_write_ce = 1'b1;
  assign from_t1_iter10_to_t1_iter11_reset = ~ ap_rst_n;
  assign from_t1_iter11_to_t1_iter12_clk = ap_clk;
  assign from_t1_iter11_to_t1_iter12_if_din = from_t1_iter11_to_t1_iter12__din;
  assign from_t1_iter11_to_t1_iter12__dout = from_t1_iter11_to_t1_iter12_if_dout;
  assign from_t1_iter11_to_t1_iter12__empty_n = from_t1_iter11_to_t1_iter12_if_empty_n;
  assign from_t1_iter11_to_t1_iter12__full_n = from_t1_iter11_to_t1_iter12_if_full_n;
  assign from_t1_iter11_to_t1_iter12_if_read = from_t1_iter11_to_t1_iter12__read;
  assign from_t1_iter11_to_t1_iter12_if_read_ce = 1'b1;
  assign from_t1_iter11_to_t1_iter12_if_write = from_t1_iter11_to_t1_iter12__write;
  assign from_t1_iter11_to_t1_iter12_if_write_ce = 1'b1;
  assign from_t1_iter11_to_t1_iter12_reset = ~ ap_rst_n;
  assign from_t1_iter12_to_t1_iter13_clk = ap_clk;
  assign from_t1_iter12_to_t1_iter13_if_din = from_t1_iter12_to_t1_iter13__din;
  assign from_t1_iter12_to_t1_iter13__dout = from_t1_iter12_to_t1_iter13_if_dout;
  assign from_t1_iter12_to_t1_iter13__empty_n = from_t1_iter12_to_t1_iter13_if_empty_n;
  assign from_t1_iter12_to_t1_iter13__full_n = from_t1_iter12_to_t1_iter13_if_full_n;
  assign from_t1_iter12_to_t1_iter13_if_read = from_t1_iter12_to_t1_iter13__read;
  assign from_t1_iter12_to_t1_iter13_if_read_ce = 1'b1;
  assign from_t1_iter12_to_t1_iter13_if_write = from_t1_iter12_to_t1_iter13__write;
  assign from_t1_iter12_to_t1_iter13_if_write_ce = 1'b1;
  assign from_t1_iter12_to_t1_iter13_reset = ~ ap_rst_n;
  assign from_t1_iter13_to_t1_iter14_clk = ap_clk;
  assign from_t1_iter13_to_t1_iter14_if_din = from_t1_iter13_to_t1_iter14__din;
  assign from_t1_iter13_to_t1_iter14__dout = from_t1_iter13_to_t1_iter14_if_dout;
  assign from_t1_iter13_to_t1_iter14__empty_n = from_t1_iter13_to_t1_iter14_if_empty_n;
  assign from_t1_iter13_to_t1_iter14__full_n = from_t1_iter13_to_t1_iter14_if_full_n;
  assign from_t1_iter13_to_t1_iter14_if_read = from_t1_iter13_to_t1_iter14__read;
  assign from_t1_iter13_to_t1_iter14_if_read_ce = 1'b1;
  assign from_t1_iter13_to_t1_iter14_if_write = from_t1_iter13_to_t1_iter14__write;
  assign from_t1_iter13_to_t1_iter14_if_write_ce = 1'b1;
  assign from_t1_iter13_to_t1_iter14_reset = ~ ap_rst_n;
  assign from_t1_iter14_to_t1_iter15_clk = ap_clk;
  assign from_t1_iter14_to_t1_iter15_if_din = from_t1_iter14_to_t1_iter15__din;
  assign from_t1_iter14_to_t1_iter15__dout = from_t1_iter14_to_t1_iter15_if_dout;
  assign from_t1_iter14_to_t1_iter15__empty_n = from_t1_iter14_to_t1_iter15_if_empty_n;
  assign from_t1_iter14_to_t1_iter15__full_n = from_t1_iter14_to_t1_iter15_if_full_n;
  assign from_t1_iter14_to_t1_iter15_if_read = from_t1_iter14_to_t1_iter15__read;
  assign from_t1_iter14_to_t1_iter15_if_read_ce = 1'b1;
  assign from_t1_iter14_to_t1_iter15_if_write = from_t1_iter14_to_t1_iter15__write;
  assign from_t1_iter14_to_t1_iter15_if_write_ce = 1'b1;
  assign from_t1_iter14_to_t1_iter15_reset = ~ ap_rst_n;
  assign from_t1_iter15_to_t1_iter16_clk = ap_clk;
  assign from_t1_iter15_to_t1_iter16_if_din = from_t1_iter15_to_t1_iter16__din;
  assign from_t1_iter15_to_t1_iter16__dout = from_t1_iter15_to_t1_iter16_if_dout;
  assign from_t1_iter15_to_t1_iter16__empty_n = from_t1_iter15_to_t1_iter16_if_empty_n;
  assign from_t1_iter15_to_t1_iter16__full_n = from_t1_iter15_to_t1_iter16_if_full_n;
  assign from_t1_iter15_to_t1_iter16_if_read = from_t1_iter15_to_t1_iter16__read;
  assign from_t1_iter15_to_t1_iter16_if_read_ce = 1'b1;
  assign from_t1_iter15_to_t1_iter16_if_write = from_t1_iter15_to_t1_iter16__write;
  assign from_t1_iter15_to_t1_iter16_if_write_ce = 1'b1;
  assign from_t1_iter15_to_t1_iter16_reset = ~ ap_rst_n;
  assign from_t1_iter16_to_t1_iter17_clk = ap_clk;
  assign from_t1_iter16_to_t1_iter17_if_din = from_t1_iter16_to_t1_iter17__din;
  assign from_t1_iter16_to_t1_iter17__dout = from_t1_iter16_to_t1_iter17_if_dout;
  assign from_t1_iter16_to_t1_iter17__empty_n = from_t1_iter16_to_t1_iter17_if_empty_n;
  assign from_t1_iter16_to_t1_iter17__full_n = from_t1_iter16_to_t1_iter17_if_full_n;
  assign from_t1_iter16_to_t1_iter17_if_read = from_t1_iter16_to_t1_iter17__read;
  assign from_t1_iter16_to_t1_iter17_if_read_ce = 1'b1;
  assign from_t1_iter16_to_t1_iter17_if_write = from_t1_iter16_to_t1_iter17__write;
  assign from_t1_iter16_to_t1_iter17_if_write_ce = 1'b1;
  assign from_t1_iter16_to_t1_iter17_reset = ~ ap_rst_n;
  assign from_t1_iter17_to_t1_iter18_clk = ap_clk;
  assign from_t1_iter17_to_t1_iter18_if_din = from_t1_iter17_to_t1_iter18__din;
  assign from_t1_iter17_to_t1_iter18__dout = from_t1_iter17_to_t1_iter18_if_dout;
  assign from_t1_iter17_to_t1_iter18__empty_n = from_t1_iter17_to_t1_iter18_if_empty_n;
  assign from_t1_iter17_to_t1_iter18__full_n = from_t1_iter17_to_t1_iter18_if_full_n;
  assign from_t1_iter17_to_t1_iter18_if_read = from_t1_iter17_to_t1_iter18__read;
  assign from_t1_iter17_to_t1_iter18_if_read_ce = 1'b1;
  assign from_t1_iter17_to_t1_iter18_if_write = from_t1_iter17_to_t1_iter18__write;
  assign from_t1_iter17_to_t1_iter18_if_write_ce = 1'b1;
  assign from_t1_iter17_to_t1_iter18_reset = ~ ap_rst_n;
  assign from_t1_iter18_to_t1_iter19_clk = ap_clk;
  assign from_t1_iter18_to_t1_iter19_if_din = from_t1_iter18_to_t1_iter19__din;
  assign from_t1_iter18_to_t1_iter19__dout = from_t1_iter18_to_t1_iter19_if_dout;
  assign from_t1_iter18_to_t1_iter19__empty_n = from_t1_iter18_to_t1_iter19_if_empty_n;
  assign from_t1_iter18_to_t1_iter19__full_n = from_t1_iter18_to_t1_iter19_if_full_n;
  assign from_t1_iter18_to_t1_iter19_if_read = from_t1_iter18_to_t1_iter19__read;
  assign from_t1_iter18_to_t1_iter19_if_read_ce = 1'b1;
  assign from_t1_iter18_to_t1_iter19_if_write = from_t1_iter18_to_t1_iter19__write;
  assign from_t1_iter18_to_t1_iter19_if_write_ce = 1'b1;
  assign from_t1_iter18_to_t1_iter19_reset = ~ ap_rst_n;
  assign from_t1_iter19_to_t1_iter20_clk = ap_clk;
  assign from_t1_iter19_to_t1_iter20_if_din = from_t1_iter19_to_t1_iter20__din;
  assign from_t1_iter19_to_t1_iter20__dout = from_t1_iter19_to_t1_iter20_if_dout;
  assign from_t1_iter19_to_t1_iter20__empty_n = from_t1_iter19_to_t1_iter20_if_empty_n;
  assign from_t1_iter19_to_t1_iter20__full_n = from_t1_iter19_to_t1_iter20_if_full_n;
  assign from_t1_iter19_to_t1_iter20_if_read = from_t1_iter19_to_t1_iter20__read;
  assign from_t1_iter19_to_t1_iter20_if_read_ce = 1'b1;
  assign from_t1_iter19_to_t1_iter20_if_write = from_t1_iter19_to_t1_iter20__write;
  assign from_t1_iter19_to_t1_iter20_if_write_ce = 1'b1;
  assign from_t1_iter19_to_t1_iter20_reset = ~ ap_rst_n;
  assign from_t1_iter1_to_t1_iter2_clk = ap_clk;
  assign from_t1_iter1_to_t1_iter2_if_din = from_t1_iter1_to_t1_iter2__din;
  assign from_t1_iter1_to_t1_iter2__dout = from_t1_iter1_to_t1_iter2_if_dout;
  assign from_t1_iter1_to_t1_iter2__empty_n = from_t1_iter1_to_t1_iter2_if_empty_n;
  assign from_t1_iter1_to_t1_iter2__full_n = from_t1_iter1_to_t1_iter2_if_full_n;
  assign from_t1_iter1_to_t1_iter2_if_read = from_t1_iter1_to_t1_iter2__read;
  assign from_t1_iter1_to_t1_iter2_if_read_ce = 1'b1;
  assign from_t1_iter1_to_t1_iter2_if_write = from_t1_iter1_to_t1_iter2__write;
  assign from_t1_iter1_to_t1_iter2_if_write_ce = 1'b1;
  assign from_t1_iter1_to_t1_iter2_reset = ~ ap_rst_n;
  assign from_t1_iter20_to_t1_iter21_clk = ap_clk;
  assign from_t1_iter20_to_t1_iter21_if_din = from_t1_iter20_to_t1_iter21__din;
  assign from_t1_iter20_to_t1_iter21__dout = from_t1_iter20_to_t1_iter21_if_dout;
  assign from_t1_iter20_to_t1_iter21__empty_n = from_t1_iter20_to_t1_iter21_if_empty_n;
  assign from_t1_iter20_to_t1_iter21__full_n = from_t1_iter20_to_t1_iter21_if_full_n;
  assign from_t1_iter20_to_t1_iter21_if_read = from_t1_iter20_to_t1_iter21__read;
  assign from_t1_iter20_to_t1_iter21_if_read_ce = 1'b1;
  assign from_t1_iter20_to_t1_iter21_if_write = from_t1_iter20_to_t1_iter21__write;
  assign from_t1_iter20_to_t1_iter21_if_write_ce = 1'b1;
  assign from_t1_iter20_to_t1_iter21_reset = ~ ap_rst_n;
  assign from_t1_iter21_to_t1_iter22_clk = ap_clk;
  assign from_t1_iter21_to_t1_iter22_if_din = from_t1_iter21_to_t1_iter22__din;
  assign from_t1_iter21_to_t1_iter22__dout = from_t1_iter21_to_t1_iter22_if_dout;
  assign from_t1_iter21_to_t1_iter22__empty_n = from_t1_iter21_to_t1_iter22_if_empty_n;
  assign from_t1_iter21_to_t1_iter22__full_n = from_t1_iter21_to_t1_iter22_if_full_n;
  assign from_t1_iter21_to_t1_iter22_if_read = from_t1_iter21_to_t1_iter22__read;
  assign from_t1_iter21_to_t1_iter22_if_read_ce = 1'b1;
  assign from_t1_iter21_to_t1_iter22_if_write = from_t1_iter21_to_t1_iter22__write;
  assign from_t1_iter21_to_t1_iter22_if_write_ce = 1'b1;
  assign from_t1_iter21_to_t1_iter22_reset = ~ ap_rst_n;
  assign from_t1_iter22_to_t1_iter23_clk = ap_clk;
  assign from_t1_iter22_to_t1_iter23_if_din = from_t1_iter22_to_t1_iter23__din;
  assign from_t1_iter22_to_t1_iter23__dout = from_t1_iter22_to_t1_iter23_if_dout;
  assign from_t1_iter22_to_t1_iter23__empty_n = from_t1_iter22_to_t1_iter23_if_empty_n;
  assign from_t1_iter22_to_t1_iter23__full_n = from_t1_iter22_to_t1_iter23_if_full_n;
  assign from_t1_iter22_to_t1_iter23_if_read = from_t1_iter22_to_t1_iter23__read;
  assign from_t1_iter22_to_t1_iter23_if_read_ce = 1'b1;
  assign from_t1_iter22_to_t1_iter23_if_write = from_t1_iter22_to_t1_iter23__write;
  assign from_t1_iter22_to_t1_iter23_if_write_ce = 1'b1;
  assign from_t1_iter22_to_t1_iter23_reset = ~ ap_rst_n;
  assign from_t1_iter23_to_t1_iter24_clk = ap_clk;
  assign from_t1_iter23_to_t1_iter24_if_din = from_t1_iter23_to_t1_iter24__din;
  assign from_t1_iter23_to_t1_iter24__dout = from_t1_iter23_to_t1_iter24_if_dout;
  assign from_t1_iter23_to_t1_iter24__empty_n = from_t1_iter23_to_t1_iter24_if_empty_n;
  assign from_t1_iter23_to_t1_iter24__full_n = from_t1_iter23_to_t1_iter24_if_full_n;
  assign from_t1_iter23_to_t1_iter24_if_read = from_t1_iter23_to_t1_iter24__read;
  assign from_t1_iter23_to_t1_iter24_if_read_ce = 1'b1;
  assign from_t1_iter23_to_t1_iter24_if_write = from_t1_iter23_to_t1_iter24__write;
  assign from_t1_iter23_to_t1_iter24_if_write_ce = 1'b1;
  assign from_t1_iter23_to_t1_iter24_reset = ~ ap_rst_n;
  assign from_t1_iter24_to_t1_iter25_clk = ap_clk;
  assign from_t1_iter24_to_t1_iter25_if_din = from_t1_iter24_to_t1_iter25__din;
  assign from_t1_iter24_to_t1_iter25__dout = from_t1_iter24_to_t1_iter25_if_dout;
  assign from_t1_iter24_to_t1_iter25__empty_n = from_t1_iter24_to_t1_iter25_if_empty_n;
  assign from_t1_iter24_to_t1_iter25__full_n = from_t1_iter24_to_t1_iter25_if_full_n;
  assign from_t1_iter24_to_t1_iter25_if_read = from_t1_iter24_to_t1_iter25__read;
  assign from_t1_iter24_to_t1_iter25_if_read_ce = 1'b1;
  assign from_t1_iter24_to_t1_iter25_if_write = from_t1_iter24_to_t1_iter25__write;
  assign from_t1_iter24_to_t1_iter25_if_write_ce = 1'b1;
  assign from_t1_iter24_to_t1_iter25_reset = ~ ap_rst_n;
  assign from_t1_iter25_to_t1_iter26_clk = ap_clk;
  assign from_t1_iter25_to_t1_iter26_if_din = from_t1_iter25_to_t1_iter26__din;
  assign from_t1_iter25_to_t1_iter26__dout = from_t1_iter25_to_t1_iter26_if_dout;
  assign from_t1_iter25_to_t1_iter26__empty_n = from_t1_iter25_to_t1_iter26_if_empty_n;
  assign from_t1_iter25_to_t1_iter26__full_n = from_t1_iter25_to_t1_iter26_if_full_n;
  assign from_t1_iter25_to_t1_iter26_if_read = from_t1_iter25_to_t1_iter26__read;
  assign from_t1_iter25_to_t1_iter26_if_read_ce = 1'b1;
  assign from_t1_iter25_to_t1_iter26_if_write = from_t1_iter25_to_t1_iter26__write;
  assign from_t1_iter25_to_t1_iter26_if_write_ce = 1'b1;
  assign from_t1_iter25_to_t1_iter26_reset = ~ ap_rst_n;
  assign from_t1_iter26_to_t1_iter27_clk = ap_clk;
  assign from_t1_iter26_to_t1_iter27_if_din = from_t1_iter26_to_t1_iter27__din;
  assign from_t1_iter26_to_t1_iter27__dout = from_t1_iter26_to_t1_iter27_if_dout;
  assign from_t1_iter26_to_t1_iter27__empty_n = from_t1_iter26_to_t1_iter27_if_empty_n;
  assign from_t1_iter26_to_t1_iter27__full_n = from_t1_iter26_to_t1_iter27_if_full_n;
  assign from_t1_iter26_to_t1_iter27_if_read = from_t1_iter26_to_t1_iter27__read;
  assign from_t1_iter26_to_t1_iter27_if_read_ce = 1'b1;
  assign from_t1_iter26_to_t1_iter27_if_write = from_t1_iter26_to_t1_iter27__write;
  assign from_t1_iter26_to_t1_iter27_if_write_ce = 1'b1;
  assign from_t1_iter26_to_t1_iter27_reset = ~ ap_rst_n;
  assign from_t1_iter27_to_t1_iter28_clk = ap_clk;
  assign from_t1_iter27_to_t1_iter28_if_din = from_t1_iter27_to_t1_iter28__din;
  assign from_t1_iter27_to_t1_iter28__dout = from_t1_iter27_to_t1_iter28_if_dout;
  assign from_t1_iter27_to_t1_iter28__empty_n = from_t1_iter27_to_t1_iter28_if_empty_n;
  assign from_t1_iter27_to_t1_iter28__full_n = from_t1_iter27_to_t1_iter28_if_full_n;
  assign from_t1_iter27_to_t1_iter28_if_read = from_t1_iter27_to_t1_iter28__read;
  assign from_t1_iter27_to_t1_iter28_if_read_ce = 1'b1;
  assign from_t1_iter27_to_t1_iter28_if_write = from_t1_iter27_to_t1_iter28__write;
  assign from_t1_iter27_to_t1_iter28_if_write_ce = 1'b1;
  assign from_t1_iter27_to_t1_iter28_reset = ~ ap_rst_n;
  assign from_t1_iter28_to_t1_iter29_clk = ap_clk;
  assign from_t1_iter28_to_t1_iter29_if_din = from_t1_iter28_to_t1_iter29__din;
  assign from_t1_iter28_to_t1_iter29__dout = from_t1_iter28_to_t1_iter29_if_dout;
  assign from_t1_iter28_to_t1_iter29__empty_n = from_t1_iter28_to_t1_iter29_if_empty_n;
  assign from_t1_iter28_to_t1_iter29__full_n = from_t1_iter28_to_t1_iter29_if_full_n;
  assign from_t1_iter28_to_t1_iter29_if_read = from_t1_iter28_to_t1_iter29__read;
  assign from_t1_iter28_to_t1_iter29_if_read_ce = 1'b1;
  assign from_t1_iter28_to_t1_iter29_if_write = from_t1_iter28_to_t1_iter29__write;
  assign from_t1_iter28_to_t1_iter29_if_write_ce = 1'b1;
  assign from_t1_iter28_to_t1_iter29_reset = ~ ap_rst_n;
  assign from_t1_iter29_to_t1_iter30_clk = ap_clk;
  assign from_t1_iter29_to_t1_iter30_if_din = from_t1_iter29_to_t1_iter30__din;
  assign from_t1_iter29_to_t1_iter30__dout = from_t1_iter29_to_t1_iter30_if_dout;
  assign from_t1_iter29_to_t1_iter30__empty_n = from_t1_iter29_to_t1_iter30_if_empty_n;
  assign from_t1_iter29_to_t1_iter30__full_n = from_t1_iter29_to_t1_iter30_if_full_n;
  assign from_t1_iter29_to_t1_iter30_if_read = from_t1_iter29_to_t1_iter30__read;
  assign from_t1_iter29_to_t1_iter30_if_read_ce = 1'b1;
  assign from_t1_iter29_to_t1_iter30_if_write = from_t1_iter29_to_t1_iter30__write;
  assign from_t1_iter29_to_t1_iter30_if_write_ce = 1'b1;
  assign from_t1_iter29_to_t1_iter30_reset = ~ ap_rst_n;
  assign from_t1_iter2_to_t1_iter3_clk = ap_clk;
  assign from_t1_iter2_to_t1_iter3_if_din = from_t1_iter2_to_t1_iter3__din;
  assign from_t1_iter2_to_t1_iter3__dout = from_t1_iter2_to_t1_iter3_if_dout;
  assign from_t1_iter2_to_t1_iter3__empty_n = from_t1_iter2_to_t1_iter3_if_empty_n;
  assign from_t1_iter2_to_t1_iter3__full_n = from_t1_iter2_to_t1_iter3_if_full_n;
  assign from_t1_iter2_to_t1_iter3_if_read = from_t1_iter2_to_t1_iter3__read;
  assign from_t1_iter2_to_t1_iter3_if_read_ce = 1'b1;
  assign from_t1_iter2_to_t1_iter3_if_write = from_t1_iter2_to_t1_iter3__write;
  assign from_t1_iter2_to_t1_iter3_if_write_ce = 1'b1;
  assign from_t1_iter2_to_t1_iter3_reset = ~ ap_rst_n;
  assign from_t1_iter30_to_t1_iter31_clk = ap_clk;
  assign from_t1_iter30_to_t1_iter31_if_din = from_t1_iter30_to_t1_iter31__din;
  assign from_t1_iter30_to_t1_iter31__dout = from_t1_iter30_to_t1_iter31_if_dout;
  assign from_t1_iter30_to_t1_iter31__empty_n = from_t1_iter30_to_t1_iter31_if_empty_n;
  assign from_t1_iter30_to_t1_iter31__full_n = from_t1_iter30_to_t1_iter31_if_full_n;
  assign from_t1_iter30_to_t1_iter31_if_read = from_t1_iter30_to_t1_iter31__read;
  assign from_t1_iter30_to_t1_iter31_if_read_ce = 1'b1;
  assign from_t1_iter30_to_t1_iter31_if_write = from_t1_iter30_to_t1_iter31__write;
  assign from_t1_iter30_to_t1_iter31_if_write_ce = 1'b1;
  assign from_t1_iter30_to_t1_iter31_reset = ~ ap_rst_n;
  assign from_t1_iter31_to_t1_iter32_clk = ap_clk;
  assign from_t1_iter31_to_t1_iter32_if_din = from_t1_iter31_to_t1_iter32__din;
  assign from_t1_iter31_to_t1_iter32__dout = from_t1_iter31_to_t1_iter32_if_dout;
  assign from_t1_iter31_to_t1_iter32__empty_n = from_t1_iter31_to_t1_iter32_if_empty_n;
  assign from_t1_iter31_to_t1_iter32__full_n = from_t1_iter31_to_t1_iter32_if_full_n;
  assign from_t1_iter31_to_t1_iter32_if_read = from_t1_iter31_to_t1_iter32__read;
  assign from_t1_iter31_to_t1_iter32_if_read_ce = 1'b1;
  assign from_t1_iter31_to_t1_iter32_if_write = from_t1_iter31_to_t1_iter32__write;
  assign from_t1_iter31_to_t1_iter32_if_write_ce = 1'b1;
  assign from_t1_iter31_to_t1_iter32_reset = ~ ap_rst_n;
  assign from_t1_iter32_to_t1_iter33_clk = ap_clk;
  assign from_t1_iter32_to_t1_iter33_if_din = from_t1_iter32_to_t1_iter33__din;
  assign from_t1_iter32_to_t1_iter33__dout = from_t1_iter32_to_t1_iter33_if_dout;
  assign from_t1_iter32_to_t1_iter33__empty_n = from_t1_iter32_to_t1_iter33_if_empty_n;
  assign from_t1_iter32_to_t1_iter33__full_n = from_t1_iter32_to_t1_iter33_if_full_n;
  assign from_t1_iter32_to_t1_iter33_if_read = from_t1_iter32_to_t1_iter33__read;
  assign from_t1_iter32_to_t1_iter33_if_read_ce = 1'b1;
  assign from_t1_iter32_to_t1_iter33_if_write = from_t1_iter32_to_t1_iter33__write;
  assign from_t1_iter32_to_t1_iter33_if_write_ce = 1'b1;
  assign from_t1_iter32_to_t1_iter33_reset = ~ ap_rst_n;
  assign from_t1_iter33_to_t1_iter34_clk = ap_clk;
  assign from_t1_iter33_to_t1_iter34_if_din = from_t1_iter33_to_t1_iter34__din;
  assign from_t1_iter33_to_t1_iter34__dout = from_t1_iter33_to_t1_iter34_if_dout;
  assign from_t1_iter33_to_t1_iter34__empty_n = from_t1_iter33_to_t1_iter34_if_empty_n;
  assign from_t1_iter33_to_t1_iter34__full_n = from_t1_iter33_to_t1_iter34_if_full_n;
  assign from_t1_iter33_to_t1_iter34_if_read = from_t1_iter33_to_t1_iter34__read;
  assign from_t1_iter33_to_t1_iter34_if_read_ce = 1'b1;
  assign from_t1_iter33_to_t1_iter34_if_write = from_t1_iter33_to_t1_iter34__write;
  assign from_t1_iter33_to_t1_iter34_if_write_ce = 1'b1;
  assign from_t1_iter33_to_t1_iter34_reset = ~ ap_rst_n;
  assign from_t1_iter34_to_t1_iter35_clk = ap_clk;
  assign from_t1_iter34_to_t1_iter35_if_din = from_t1_iter34_to_t1_iter35__din;
  assign from_t1_iter34_to_t1_iter35__dout = from_t1_iter34_to_t1_iter35_if_dout;
  assign from_t1_iter34_to_t1_iter35__empty_n = from_t1_iter34_to_t1_iter35_if_empty_n;
  assign from_t1_iter34_to_t1_iter35__full_n = from_t1_iter34_to_t1_iter35_if_full_n;
  assign from_t1_iter34_to_t1_iter35_if_read = from_t1_iter34_to_t1_iter35__read;
  assign from_t1_iter34_to_t1_iter35_if_read_ce = 1'b1;
  assign from_t1_iter34_to_t1_iter35_if_write = from_t1_iter34_to_t1_iter35__write;
  assign from_t1_iter34_to_t1_iter35_if_write_ce = 1'b1;
  assign from_t1_iter34_to_t1_iter35_reset = ~ ap_rst_n;
  assign from_t1_iter35_to_t1_iter36_clk = ap_clk;
  assign from_t1_iter35_to_t1_iter36_if_din = from_t1_iter35_to_t1_iter36__din;
  assign from_t1_iter35_to_t1_iter36__dout = from_t1_iter35_to_t1_iter36_if_dout;
  assign from_t1_iter35_to_t1_iter36__empty_n = from_t1_iter35_to_t1_iter36_if_empty_n;
  assign from_t1_iter35_to_t1_iter36__full_n = from_t1_iter35_to_t1_iter36_if_full_n;
  assign from_t1_iter35_to_t1_iter36_if_read = from_t1_iter35_to_t1_iter36__read;
  assign from_t1_iter35_to_t1_iter36_if_read_ce = 1'b1;
  assign from_t1_iter35_to_t1_iter36_if_write = from_t1_iter35_to_t1_iter36__write;
  assign from_t1_iter35_to_t1_iter36_if_write_ce = 1'b1;
  assign from_t1_iter35_to_t1_iter36_reset = ~ ap_rst_n;
  assign from_t1_iter36_to_t1_iter37_clk = ap_clk;
  assign from_t1_iter36_to_t1_iter37_if_din = from_t1_iter36_to_t1_iter37__din;
  assign from_t1_iter36_to_t1_iter37__dout = from_t1_iter36_to_t1_iter37_if_dout;
  assign from_t1_iter36_to_t1_iter37__empty_n = from_t1_iter36_to_t1_iter37_if_empty_n;
  assign from_t1_iter36_to_t1_iter37__full_n = from_t1_iter36_to_t1_iter37_if_full_n;
  assign from_t1_iter36_to_t1_iter37_if_read = from_t1_iter36_to_t1_iter37__read;
  assign from_t1_iter36_to_t1_iter37_if_read_ce = 1'b1;
  assign from_t1_iter36_to_t1_iter37_if_write = from_t1_iter36_to_t1_iter37__write;
  assign from_t1_iter36_to_t1_iter37_if_write_ce = 1'b1;
  assign from_t1_iter36_to_t1_iter37_reset = ~ ap_rst_n;
  assign from_t1_iter37_to_t1_iter38_clk = ap_clk;
  assign from_t1_iter37_to_t1_iter38_if_din = from_t1_iter37_to_t1_iter38__din;
  assign from_t1_iter37_to_t1_iter38__dout = from_t1_iter37_to_t1_iter38_if_dout;
  assign from_t1_iter37_to_t1_iter38__empty_n = from_t1_iter37_to_t1_iter38_if_empty_n;
  assign from_t1_iter37_to_t1_iter38__full_n = from_t1_iter37_to_t1_iter38_if_full_n;
  assign from_t1_iter37_to_t1_iter38_if_read = from_t1_iter37_to_t1_iter38__read;
  assign from_t1_iter37_to_t1_iter38_if_read_ce = 1'b1;
  assign from_t1_iter37_to_t1_iter38_if_write = from_t1_iter37_to_t1_iter38__write;
  assign from_t1_iter37_to_t1_iter38_if_write_ce = 1'b1;
  assign from_t1_iter37_to_t1_iter38_reset = ~ ap_rst_n;
  assign from_t1_iter38_to_t1_iter39_clk = ap_clk;
  assign from_t1_iter38_to_t1_iter39_if_din = from_t1_iter38_to_t1_iter39__din;
  assign from_t1_iter38_to_t1_iter39__dout = from_t1_iter38_to_t1_iter39_if_dout;
  assign from_t1_iter38_to_t1_iter39__empty_n = from_t1_iter38_to_t1_iter39_if_empty_n;
  assign from_t1_iter38_to_t1_iter39__full_n = from_t1_iter38_to_t1_iter39_if_full_n;
  assign from_t1_iter38_to_t1_iter39_if_read = from_t1_iter38_to_t1_iter39__read;
  assign from_t1_iter38_to_t1_iter39_if_read_ce = 1'b1;
  assign from_t1_iter38_to_t1_iter39_if_write = from_t1_iter38_to_t1_iter39__write;
  assign from_t1_iter38_to_t1_iter39_if_write_ce = 1'b1;
  assign from_t1_iter38_to_t1_iter39_reset = ~ ap_rst_n;
  assign from_t1_iter39_to_t1_iter40_clk = ap_clk;
  assign from_t1_iter39_to_t1_iter40_if_din = from_t1_iter39_to_t1_iter40__din;
  assign from_t1_iter39_to_t1_iter40__dout = from_t1_iter39_to_t1_iter40_if_dout;
  assign from_t1_iter39_to_t1_iter40__empty_n = from_t1_iter39_to_t1_iter40_if_empty_n;
  assign from_t1_iter39_to_t1_iter40__full_n = from_t1_iter39_to_t1_iter40_if_full_n;
  assign from_t1_iter39_to_t1_iter40_if_read = from_t1_iter39_to_t1_iter40__read;
  assign from_t1_iter39_to_t1_iter40_if_read_ce = 1'b1;
  assign from_t1_iter39_to_t1_iter40_if_write = from_t1_iter39_to_t1_iter40__write;
  assign from_t1_iter39_to_t1_iter40_if_write_ce = 1'b1;
  assign from_t1_iter39_to_t1_iter40_reset = ~ ap_rst_n;
  assign from_t1_iter3_to_t1_iter4_clk = ap_clk;
  assign from_t1_iter3_to_t1_iter4_if_din = from_t1_iter3_to_t1_iter4__din;
  assign from_t1_iter3_to_t1_iter4__dout = from_t1_iter3_to_t1_iter4_if_dout;
  assign from_t1_iter3_to_t1_iter4__empty_n = from_t1_iter3_to_t1_iter4_if_empty_n;
  assign from_t1_iter3_to_t1_iter4__full_n = from_t1_iter3_to_t1_iter4_if_full_n;
  assign from_t1_iter3_to_t1_iter4_if_read = from_t1_iter3_to_t1_iter4__read;
  assign from_t1_iter3_to_t1_iter4_if_read_ce = 1'b1;
  assign from_t1_iter3_to_t1_iter4_if_write = from_t1_iter3_to_t1_iter4__write;
  assign from_t1_iter3_to_t1_iter4_if_write_ce = 1'b1;
  assign from_t1_iter3_to_t1_iter4_reset = ~ ap_rst_n;
  assign from_t1_iter40_to_t1_iter41_clk = ap_clk;
  assign from_t1_iter40_to_t1_iter41_if_din = from_t1_iter40_to_t1_iter41__din;
  assign from_t1_iter40_to_t1_iter41__dout = from_t1_iter40_to_t1_iter41_if_dout;
  assign from_t1_iter40_to_t1_iter41__empty_n = from_t1_iter40_to_t1_iter41_if_empty_n;
  assign from_t1_iter40_to_t1_iter41__full_n = from_t1_iter40_to_t1_iter41_if_full_n;
  assign from_t1_iter40_to_t1_iter41_if_read = from_t1_iter40_to_t1_iter41__read;
  assign from_t1_iter40_to_t1_iter41_if_read_ce = 1'b1;
  assign from_t1_iter40_to_t1_iter41_if_write = from_t1_iter40_to_t1_iter41__write;
  assign from_t1_iter40_to_t1_iter41_if_write_ce = 1'b1;
  assign from_t1_iter40_to_t1_iter41_reset = ~ ap_rst_n;
  assign from_t1_iter41_to_t1_iter42_clk = ap_clk;
  assign from_t1_iter41_to_t1_iter42_if_din = from_t1_iter41_to_t1_iter42__din;
  assign from_t1_iter41_to_t1_iter42__dout = from_t1_iter41_to_t1_iter42_if_dout;
  assign from_t1_iter41_to_t1_iter42__empty_n = from_t1_iter41_to_t1_iter42_if_empty_n;
  assign from_t1_iter41_to_t1_iter42__full_n = from_t1_iter41_to_t1_iter42_if_full_n;
  assign from_t1_iter41_to_t1_iter42_if_read = from_t1_iter41_to_t1_iter42__read;
  assign from_t1_iter41_to_t1_iter42_if_read_ce = 1'b1;
  assign from_t1_iter41_to_t1_iter42_if_write = from_t1_iter41_to_t1_iter42__write;
  assign from_t1_iter41_to_t1_iter42_if_write_ce = 1'b1;
  assign from_t1_iter41_to_t1_iter42_reset = ~ ap_rst_n;
  assign from_t1_iter42_to_t1_iter43_clk = ap_clk;
  assign from_t1_iter42_to_t1_iter43_if_din = from_t1_iter42_to_t1_iter43__din;
  assign from_t1_iter42_to_t1_iter43__dout = from_t1_iter42_to_t1_iter43_if_dout;
  assign from_t1_iter42_to_t1_iter43__empty_n = from_t1_iter42_to_t1_iter43_if_empty_n;
  assign from_t1_iter42_to_t1_iter43__full_n = from_t1_iter42_to_t1_iter43_if_full_n;
  assign from_t1_iter42_to_t1_iter43_if_read = from_t1_iter42_to_t1_iter43__read;
  assign from_t1_iter42_to_t1_iter43_if_read_ce = 1'b1;
  assign from_t1_iter42_to_t1_iter43_if_write = from_t1_iter42_to_t1_iter43__write;
  assign from_t1_iter42_to_t1_iter43_if_write_ce = 1'b1;
  assign from_t1_iter42_to_t1_iter43_reset = ~ ap_rst_n;
  assign from_t1_iter43_to_t1_iter44_clk = ap_clk;
  assign from_t1_iter43_to_t1_iter44_if_din = from_t1_iter43_to_t1_iter44__din;
  assign from_t1_iter43_to_t1_iter44__dout = from_t1_iter43_to_t1_iter44_if_dout;
  assign from_t1_iter43_to_t1_iter44__empty_n = from_t1_iter43_to_t1_iter44_if_empty_n;
  assign from_t1_iter43_to_t1_iter44__full_n = from_t1_iter43_to_t1_iter44_if_full_n;
  assign from_t1_iter43_to_t1_iter44_if_read = from_t1_iter43_to_t1_iter44__read;
  assign from_t1_iter43_to_t1_iter44_if_read_ce = 1'b1;
  assign from_t1_iter43_to_t1_iter44_if_write = from_t1_iter43_to_t1_iter44__write;
  assign from_t1_iter43_to_t1_iter44_if_write_ce = 1'b1;
  assign from_t1_iter43_to_t1_iter44_reset = ~ ap_rst_n;
  assign from_t1_iter44_to_t1_iter45_clk = ap_clk;
  assign from_t1_iter44_to_t1_iter45_if_din = from_t1_iter44_to_t1_iter45__din;
  assign from_t1_iter44_to_t1_iter45__dout = from_t1_iter44_to_t1_iter45_if_dout;
  assign from_t1_iter44_to_t1_iter45__empty_n = from_t1_iter44_to_t1_iter45_if_empty_n;
  assign from_t1_iter44_to_t1_iter45__full_n = from_t1_iter44_to_t1_iter45_if_full_n;
  assign from_t1_iter44_to_t1_iter45_if_read = from_t1_iter44_to_t1_iter45__read;
  assign from_t1_iter44_to_t1_iter45_if_read_ce = 1'b1;
  assign from_t1_iter44_to_t1_iter45_if_write = from_t1_iter44_to_t1_iter45__write;
  assign from_t1_iter44_to_t1_iter45_if_write_ce = 1'b1;
  assign from_t1_iter44_to_t1_iter45_reset = ~ ap_rst_n;
  assign from_t1_iter45_to_t1_iter46_clk = ap_clk;
  assign from_t1_iter45_to_t1_iter46_if_din = from_t1_iter45_to_t1_iter46__din;
  assign from_t1_iter45_to_t1_iter46__dout = from_t1_iter45_to_t1_iter46_if_dout;
  assign from_t1_iter45_to_t1_iter46__empty_n = from_t1_iter45_to_t1_iter46_if_empty_n;
  assign from_t1_iter45_to_t1_iter46__full_n = from_t1_iter45_to_t1_iter46_if_full_n;
  assign from_t1_iter45_to_t1_iter46_if_read = from_t1_iter45_to_t1_iter46__read;
  assign from_t1_iter45_to_t1_iter46_if_read_ce = 1'b1;
  assign from_t1_iter45_to_t1_iter46_if_write = from_t1_iter45_to_t1_iter46__write;
  assign from_t1_iter45_to_t1_iter46_if_write_ce = 1'b1;
  assign from_t1_iter45_to_t1_iter46_reset = ~ ap_rst_n;
  assign from_t1_iter46_to_t1_iter47_clk = ap_clk;
  assign from_t1_iter46_to_t1_iter47_if_din = from_t1_iter46_to_t1_iter47__din;
  assign from_t1_iter46_to_t1_iter47__dout = from_t1_iter46_to_t1_iter47_if_dout;
  assign from_t1_iter46_to_t1_iter47__empty_n = from_t1_iter46_to_t1_iter47_if_empty_n;
  assign from_t1_iter46_to_t1_iter47__full_n = from_t1_iter46_to_t1_iter47_if_full_n;
  assign from_t1_iter46_to_t1_iter47_if_read = from_t1_iter46_to_t1_iter47__read;
  assign from_t1_iter46_to_t1_iter47_if_read_ce = 1'b1;
  assign from_t1_iter46_to_t1_iter47_if_write = from_t1_iter46_to_t1_iter47__write;
  assign from_t1_iter46_to_t1_iter47_if_write_ce = 1'b1;
  assign from_t1_iter46_to_t1_iter47_reset = ~ ap_rst_n;
  assign from_t1_iter47_to_t1_iter48_clk = ap_clk;
  assign from_t1_iter47_to_t1_iter48_if_din = from_t1_iter47_to_t1_iter48__din;
  assign from_t1_iter47_to_t1_iter48__dout = from_t1_iter47_to_t1_iter48_if_dout;
  assign from_t1_iter47_to_t1_iter48__empty_n = from_t1_iter47_to_t1_iter48_if_empty_n;
  assign from_t1_iter47_to_t1_iter48__full_n = from_t1_iter47_to_t1_iter48_if_full_n;
  assign from_t1_iter47_to_t1_iter48_if_read = from_t1_iter47_to_t1_iter48__read;
  assign from_t1_iter47_to_t1_iter48_if_read_ce = 1'b1;
  assign from_t1_iter47_to_t1_iter48_if_write = from_t1_iter47_to_t1_iter48__write;
  assign from_t1_iter47_to_t1_iter48_if_write_ce = 1'b1;
  assign from_t1_iter47_to_t1_iter48_reset = ~ ap_rst_n;
  assign from_t1_iter48_to_t1_iter49_clk = ap_clk;
  assign from_t1_iter48_to_t1_iter49_if_din = from_t1_iter48_to_t1_iter49__din;
  assign from_t1_iter48_to_t1_iter49__dout = from_t1_iter48_to_t1_iter49_if_dout;
  assign from_t1_iter48_to_t1_iter49__empty_n = from_t1_iter48_to_t1_iter49_if_empty_n;
  assign from_t1_iter48_to_t1_iter49__full_n = from_t1_iter48_to_t1_iter49_if_full_n;
  assign from_t1_iter48_to_t1_iter49_if_read = from_t1_iter48_to_t1_iter49__read;
  assign from_t1_iter48_to_t1_iter49_if_read_ce = 1'b1;
  assign from_t1_iter48_to_t1_iter49_if_write = from_t1_iter48_to_t1_iter49__write;
  assign from_t1_iter48_to_t1_iter49_if_write_ce = 1'b1;
  assign from_t1_iter48_to_t1_iter49_reset = ~ ap_rst_n;
  assign from_t1_iter49_to_t1_iter50_clk = ap_clk;
  assign from_t1_iter49_to_t1_iter50_if_din = from_t1_iter49_to_t1_iter50__din;
  assign from_t1_iter49_to_t1_iter50__dout = from_t1_iter49_to_t1_iter50_if_dout;
  assign from_t1_iter49_to_t1_iter50__empty_n = from_t1_iter49_to_t1_iter50_if_empty_n;
  assign from_t1_iter49_to_t1_iter50__full_n = from_t1_iter49_to_t1_iter50_if_full_n;
  assign from_t1_iter49_to_t1_iter50_if_read = from_t1_iter49_to_t1_iter50__read;
  assign from_t1_iter49_to_t1_iter50_if_read_ce = 1'b1;
  assign from_t1_iter49_to_t1_iter50_if_write = from_t1_iter49_to_t1_iter50__write;
  assign from_t1_iter49_to_t1_iter50_if_write_ce = 1'b1;
  assign from_t1_iter49_to_t1_iter50_reset = ~ ap_rst_n;
  assign from_t1_iter4_to_t1_iter5_clk = ap_clk;
  assign from_t1_iter4_to_t1_iter5_if_din = from_t1_iter4_to_t1_iter5__din;
  assign from_t1_iter4_to_t1_iter5__dout = from_t1_iter4_to_t1_iter5_if_dout;
  assign from_t1_iter4_to_t1_iter5__empty_n = from_t1_iter4_to_t1_iter5_if_empty_n;
  assign from_t1_iter4_to_t1_iter5__full_n = from_t1_iter4_to_t1_iter5_if_full_n;
  assign from_t1_iter4_to_t1_iter5_if_read = from_t1_iter4_to_t1_iter5__read;
  assign from_t1_iter4_to_t1_iter5_if_read_ce = 1'b1;
  assign from_t1_iter4_to_t1_iter5_if_write = from_t1_iter4_to_t1_iter5__write;
  assign from_t1_iter4_to_t1_iter5_if_write_ce = 1'b1;
  assign from_t1_iter4_to_t1_iter5_reset = ~ ap_rst_n;
  assign from_t1_iter50_to_t1_iter51_clk = ap_clk;
  assign from_t1_iter50_to_t1_iter51_if_din = from_t1_iter50_to_t1_iter51__din;
  assign from_t1_iter50_to_t1_iter51__dout = from_t1_iter50_to_t1_iter51_if_dout;
  assign from_t1_iter50_to_t1_iter51__empty_n = from_t1_iter50_to_t1_iter51_if_empty_n;
  assign from_t1_iter50_to_t1_iter51__full_n = from_t1_iter50_to_t1_iter51_if_full_n;
  assign from_t1_iter50_to_t1_iter51_if_read = from_t1_iter50_to_t1_iter51__read;
  assign from_t1_iter50_to_t1_iter51_if_read_ce = 1'b1;
  assign from_t1_iter50_to_t1_iter51_if_write = from_t1_iter50_to_t1_iter51__write;
  assign from_t1_iter50_to_t1_iter51_if_write_ce = 1'b1;
  assign from_t1_iter50_to_t1_iter51_reset = ~ ap_rst_n;
  assign from_t1_iter51_to_t1_iter52_clk = ap_clk;
  assign from_t1_iter51_to_t1_iter52_if_din = from_t1_iter51_to_t1_iter52__din;
  assign from_t1_iter51_to_t1_iter52__dout = from_t1_iter51_to_t1_iter52_if_dout;
  assign from_t1_iter51_to_t1_iter52__empty_n = from_t1_iter51_to_t1_iter52_if_empty_n;
  assign from_t1_iter51_to_t1_iter52__full_n = from_t1_iter51_to_t1_iter52_if_full_n;
  assign from_t1_iter51_to_t1_iter52_if_read = from_t1_iter51_to_t1_iter52__read;
  assign from_t1_iter51_to_t1_iter52_if_read_ce = 1'b1;
  assign from_t1_iter51_to_t1_iter52_if_write = from_t1_iter51_to_t1_iter52__write;
  assign from_t1_iter51_to_t1_iter52_if_write_ce = 1'b1;
  assign from_t1_iter51_to_t1_iter52_reset = ~ ap_rst_n;
  assign from_t1_iter52_to_t1_iter53_clk = ap_clk;
  assign from_t1_iter52_to_t1_iter53_if_din = from_t1_iter52_to_t1_iter53__din;
  assign from_t1_iter52_to_t1_iter53__dout = from_t1_iter52_to_t1_iter53_if_dout;
  assign from_t1_iter52_to_t1_iter53__empty_n = from_t1_iter52_to_t1_iter53_if_empty_n;
  assign from_t1_iter52_to_t1_iter53__full_n = from_t1_iter52_to_t1_iter53_if_full_n;
  assign from_t1_iter52_to_t1_iter53_if_read = from_t1_iter52_to_t1_iter53__read;
  assign from_t1_iter52_to_t1_iter53_if_read_ce = 1'b1;
  assign from_t1_iter52_to_t1_iter53_if_write = from_t1_iter52_to_t1_iter53__write;
  assign from_t1_iter52_to_t1_iter53_if_write_ce = 1'b1;
  assign from_t1_iter52_to_t1_iter53_reset = ~ ap_rst_n;
  assign from_t1_iter53_to_t1_iter54_clk = ap_clk;
  assign from_t1_iter53_to_t1_iter54_if_din = from_t1_iter53_to_t1_iter54__din;
  assign from_t1_iter53_to_t1_iter54__dout = from_t1_iter53_to_t1_iter54_if_dout;
  assign from_t1_iter53_to_t1_iter54__empty_n = from_t1_iter53_to_t1_iter54_if_empty_n;
  assign from_t1_iter53_to_t1_iter54__full_n = from_t1_iter53_to_t1_iter54_if_full_n;
  assign from_t1_iter53_to_t1_iter54_if_read = from_t1_iter53_to_t1_iter54__read;
  assign from_t1_iter53_to_t1_iter54_if_read_ce = 1'b1;
  assign from_t1_iter53_to_t1_iter54_if_write = from_t1_iter53_to_t1_iter54__write;
  assign from_t1_iter53_to_t1_iter54_if_write_ce = 1'b1;
  assign from_t1_iter53_to_t1_iter54_reset = ~ ap_rst_n;
  assign from_t1_iter54_to_t1_iter55_clk = ap_clk;
  assign from_t1_iter54_to_t1_iter55_if_din = from_t1_iter54_to_t1_iter55__din;
  assign from_t1_iter54_to_t1_iter55__dout = from_t1_iter54_to_t1_iter55_if_dout;
  assign from_t1_iter54_to_t1_iter55__empty_n = from_t1_iter54_to_t1_iter55_if_empty_n;
  assign from_t1_iter54_to_t1_iter55__full_n = from_t1_iter54_to_t1_iter55_if_full_n;
  assign from_t1_iter54_to_t1_iter55_if_read = from_t1_iter54_to_t1_iter55__read;
  assign from_t1_iter54_to_t1_iter55_if_read_ce = 1'b1;
  assign from_t1_iter54_to_t1_iter55_if_write = from_t1_iter54_to_t1_iter55__write;
  assign from_t1_iter54_to_t1_iter55_if_write_ce = 1'b1;
  assign from_t1_iter54_to_t1_iter55_reset = ~ ap_rst_n;
  assign from_t1_iter55_to_t1_iter56_clk = ap_clk;
  assign from_t1_iter55_to_t1_iter56_if_din = from_t1_iter55_to_t1_iter56__din;
  assign from_t1_iter55_to_t1_iter56__dout = from_t1_iter55_to_t1_iter56_if_dout;
  assign from_t1_iter55_to_t1_iter56__empty_n = from_t1_iter55_to_t1_iter56_if_empty_n;
  assign from_t1_iter55_to_t1_iter56__full_n = from_t1_iter55_to_t1_iter56_if_full_n;
  assign from_t1_iter55_to_t1_iter56_if_read = from_t1_iter55_to_t1_iter56__read;
  assign from_t1_iter55_to_t1_iter56_if_read_ce = 1'b1;
  assign from_t1_iter55_to_t1_iter56_if_write = from_t1_iter55_to_t1_iter56__write;
  assign from_t1_iter55_to_t1_iter56_if_write_ce = 1'b1;
  assign from_t1_iter55_to_t1_iter56_reset = ~ ap_rst_n;
  assign from_t1_iter56_to_t1_iter57_clk = ap_clk;
  assign from_t1_iter56_to_t1_iter57_if_din = from_t1_iter56_to_t1_iter57__din;
  assign from_t1_iter56_to_t1_iter57__dout = from_t1_iter56_to_t1_iter57_if_dout;
  assign from_t1_iter56_to_t1_iter57__empty_n = from_t1_iter56_to_t1_iter57_if_empty_n;
  assign from_t1_iter56_to_t1_iter57__full_n = from_t1_iter56_to_t1_iter57_if_full_n;
  assign from_t1_iter56_to_t1_iter57_if_read = from_t1_iter56_to_t1_iter57__read;
  assign from_t1_iter56_to_t1_iter57_if_read_ce = 1'b1;
  assign from_t1_iter56_to_t1_iter57_if_write = from_t1_iter56_to_t1_iter57__write;
  assign from_t1_iter56_to_t1_iter57_if_write_ce = 1'b1;
  assign from_t1_iter56_to_t1_iter57_reset = ~ ap_rst_n;
  assign from_t1_iter57_to_t1_iter58_clk = ap_clk;
  assign from_t1_iter57_to_t1_iter58_if_din = from_t1_iter57_to_t1_iter58__din;
  assign from_t1_iter57_to_t1_iter58__dout = from_t1_iter57_to_t1_iter58_if_dout;
  assign from_t1_iter57_to_t1_iter58__empty_n = from_t1_iter57_to_t1_iter58_if_empty_n;
  assign from_t1_iter57_to_t1_iter58__full_n = from_t1_iter57_to_t1_iter58_if_full_n;
  assign from_t1_iter57_to_t1_iter58_if_read = from_t1_iter57_to_t1_iter58__read;
  assign from_t1_iter57_to_t1_iter58_if_read_ce = 1'b1;
  assign from_t1_iter57_to_t1_iter58_if_write = from_t1_iter57_to_t1_iter58__write;
  assign from_t1_iter57_to_t1_iter58_if_write_ce = 1'b1;
  assign from_t1_iter57_to_t1_iter58_reset = ~ ap_rst_n;
  assign from_t1_iter58_to_t1_iter59_clk = ap_clk;
  assign from_t1_iter58_to_t1_iter59_if_din = from_t1_iter58_to_t1_iter59__din;
  assign from_t1_iter58_to_t1_iter59__dout = from_t1_iter58_to_t1_iter59_if_dout;
  assign from_t1_iter58_to_t1_iter59__empty_n = from_t1_iter58_to_t1_iter59_if_empty_n;
  assign from_t1_iter58_to_t1_iter59__full_n = from_t1_iter58_to_t1_iter59_if_full_n;
  assign from_t1_iter58_to_t1_iter59_if_read = from_t1_iter58_to_t1_iter59__read;
  assign from_t1_iter58_to_t1_iter59_if_read_ce = 1'b1;
  assign from_t1_iter58_to_t1_iter59_if_write = from_t1_iter58_to_t1_iter59__write;
  assign from_t1_iter58_to_t1_iter59_if_write_ce = 1'b1;
  assign from_t1_iter58_to_t1_iter59_reset = ~ ap_rst_n;
  assign from_t1_iter59_to_t1_iter60_clk = ap_clk;
  assign from_t1_iter59_to_t1_iter60_if_din = from_t1_iter59_to_t1_iter60__din;
  assign from_t1_iter59_to_t1_iter60__dout = from_t1_iter59_to_t1_iter60_if_dout;
  assign from_t1_iter59_to_t1_iter60__empty_n = from_t1_iter59_to_t1_iter60_if_empty_n;
  assign from_t1_iter59_to_t1_iter60__full_n = from_t1_iter59_to_t1_iter60_if_full_n;
  assign from_t1_iter59_to_t1_iter60_if_read = from_t1_iter59_to_t1_iter60__read;
  assign from_t1_iter59_to_t1_iter60_if_read_ce = 1'b1;
  assign from_t1_iter59_to_t1_iter60_if_write = from_t1_iter59_to_t1_iter60__write;
  assign from_t1_iter59_to_t1_iter60_if_write_ce = 1'b1;
  assign from_t1_iter59_to_t1_iter60_reset = ~ ap_rst_n;
  assign from_t1_iter5_to_t1_iter6_clk = ap_clk;
  assign from_t1_iter5_to_t1_iter6_if_din = from_t1_iter5_to_t1_iter6__din;
  assign from_t1_iter5_to_t1_iter6__dout = from_t1_iter5_to_t1_iter6_if_dout;
  assign from_t1_iter5_to_t1_iter6__empty_n = from_t1_iter5_to_t1_iter6_if_empty_n;
  assign from_t1_iter5_to_t1_iter6__full_n = from_t1_iter5_to_t1_iter6_if_full_n;
  assign from_t1_iter5_to_t1_iter6_if_read = from_t1_iter5_to_t1_iter6__read;
  assign from_t1_iter5_to_t1_iter6_if_read_ce = 1'b1;
  assign from_t1_iter5_to_t1_iter6_if_write = from_t1_iter5_to_t1_iter6__write;
  assign from_t1_iter5_to_t1_iter6_if_write_ce = 1'b1;
  assign from_t1_iter5_to_t1_iter6_reset = ~ ap_rst_n;
  assign from_t1_iter60_to_t1_iter61_clk = ap_clk;
  assign from_t1_iter60_to_t1_iter61_if_din = from_t1_iter60_to_t1_iter61__din;
  assign from_t1_iter60_to_t1_iter61__dout = from_t1_iter60_to_t1_iter61_if_dout;
  assign from_t1_iter60_to_t1_iter61__empty_n = from_t1_iter60_to_t1_iter61_if_empty_n;
  assign from_t1_iter60_to_t1_iter61__full_n = from_t1_iter60_to_t1_iter61_if_full_n;
  assign from_t1_iter60_to_t1_iter61_if_read = from_t1_iter60_to_t1_iter61__read;
  assign from_t1_iter60_to_t1_iter61_if_read_ce = 1'b1;
  assign from_t1_iter60_to_t1_iter61_if_write = from_t1_iter60_to_t1_iter61__write;
  assign from_t1_iter60_to_t1_iter61_if_write_ce = 1'b1;
  assign from_t1_iter60_to_t1_iter61_reset = ~ ap_rst_n;
  assign from_t1_iter61_to_t1_iter62_clk = ap_clk;
  assign from_t1_iter61_to_t1_iter62_if_din = from_t1_iter61_to_t1_iter62__din;
  assign from_t1_iter61_to_t1_iter62__dout = from_t1_iter61_to_t1_iter62_if_dout;
  assign from_t1_iter61_to_t1_iter62__empty_n = from_t1_iter61_to_t1_iter62_if_empty_n;
  assign from_t1_iter61_to_t1_iter62__full_n = from_t1_iter61_to_t1_iter62_if_full_n;
  assign from_t1_iter61_to_t1_iter62_if_read = from_t1_iter61_to_t1_iter62__read;
  assign from_t1_iter61_to_t1_iter62_if_read_ce = 1'b1;
  assign from_t1_iter61_to_t1_iter62_if_write = from_t1_iter61_to_t1_iter62__write;
  assign from_t1_iter61_to_t1_iter62_if_write_ce = 1'b1;
  assign from_t1_iter61_to_t1_iter62_reset = ~ ap_rst_n;
  assign from_t1_iter62_to_t1_iter63_clk = ap_clk;
  assign from_t1_iter62_to_t1_iter63_if_din = from_t1_iter62_to_t1_iter63__din;
  assign from_t1_iter62_to_t1_iter63__dout = from_t1_iter62_to_t1_iter63_if_dout;
  assign from_t1_iter62_to_t1_iter63__empty_n = from_t1_iter62_to_t1_iter63_if_empty_n;
  assign from_t1_iter62_to_t1_iter63__full_n = from_t1_iter62_to_t1_iter63_if_full_n;
  assign from_t1_iter62_to_t1_iter63_if_read = from_t1_iter62_to_t1_iter63__read;
  assign from_t1_iter62_to_t1_iter63_if_read_ce = 1'b1;
  assign from_t1_iter62_to_t1_iter63_if_write = from_t1_iter62_to_t1_iter63__write;
  assign from_t1_iter62_to_t1_iter63_if_write_ce = 1'b1;
  assign from_t1_iter62_to_t1_iter63_reset = ~ ap_rst_n;
  assign from_t1_iter63_to_t1_iter64_clk = ap_clk;
  assign from_t1_iter63_to_t1_iter64_if_din = from_t1_iter63_to_t1_iter64__din;
  assign from_t1_iter63_to_t1_iter64__dout = from_t1_iter63_to_t1_iter64_if_dout;
  assign from_t1_iter63_to_t1_iter64__empty_n = from_t1_iter63_to_t1_iter64_if_empty_n;
  assign from_t1_iter63_to_t1_iter64__full_n = from_t1_iter63_to_t1_iter64_if_full_n;
  assign from_t1_iter63_to_t1_iter64_if_read = from_t1_iter63_to_t1_iter64__read;
  assign from_t1_iter63_to_t1_iter64_if_read_ce = 1'b1;
  assign from_t1_iter63_to_t1_iter64_if_write = from_t1_iter63_to_t1_iter64__write;
  assign from_t1_iter63_to_t1_iter64_if_write_ce = 1'b1;
  assign from_t1_iter63_to_t1_iter64_reset = ~ ap_rst_n;
  assign from_t1_iter64_to_t1_iter65_clk = ap_clk;
  assign from_t1_iter64_to_t1_iter65_if_din = from_t1_iter64_to_t1_iter65__din;
  assign from_t1_iter64_to_t1_iter65__dout = from_t1_iter64_to_t1_iter65_if_dout;
  assign from_t1_iter64_to_t1_iter65__empty_n = from_t1_iter64_to_t1_iter65_if_empty_n;
  assign from_t1_iter64_to_t1_iter65__full_n = from_t1_iter64_to_t1_iter65_if_full_n;
  assign from_t1_iter64_to_t1_iter65_if_read = from_t1_iter64_to_t1_iter65__read;
  assign from_t1_iter64_to_t1_iter65_if_read_ce = 1'b1;
  assign from_t1_iter64_to_t1_iter65_if_write = from_t1_iter64_to_t1_iter65__write;
  assign from_t1_iter64_to_t1_iter65_if_write_ce = 1'b1;
  assign from_t1_iter64_to_t1_iter65_reset = ~ ap_rst_n;
  assign from_t1_iter65_to_t1_iter66_clk = ap_clk;
  assign from_t1_iter65_to_t1_iter66_if_din = from_t1_iter65_to_t1_iter66__din;
  assign from_t1_iter65_to_t1_iter66__dout = from_t1_iter65_to_t1_iter66_if_dout;
  assign from_t1_iter65_to_t1_iter66__empty_n = from_t1_iter65_to_t1_iter66_if_empty_n;
  assign from_t1_iter65_to_t1_iter66__full_n = from_t1_iter65_to_t1_iter66_if_full_n;
  assign from_t1_iter65_to_t1_iter66_if_read = from_t1_iter65_to_t1_iter66__read;
  assign from_t1_iter65_to_t1_iter66_if_read_ce = 1'b1;
  assign from_t1_iter65_to_t1_iter66_if_write = from_t1_iter65_to_t1_iter66__write;
  assign from_t1_iter65_to_t1_iter66_if_write_ce = 1'b1;
  assign from_t1_iter65_to_t1_iter66_reset = ~ ap_rst_n;
  assign from_t1_iter66_to_t1_iter67_clk = ap_clk;
  assign from_t1_iter66_to_t1_iter67_if_din = from_t1_iter66_to_t1_iter67__din;
  assign from_t1_iter66_to_t1_iter67__dout = from_t1_iter66_to_t1_iter67_if_dout;
  assign from_t1_iter66_to_t1_iter67__empty_n = from_t1_iter66_to_t1_iter67_if_empty_n;
  assign from_t1_iter66_to_t1_iter67__full_n = from_t1_iter66_to_t1_iter67_if_full_n;
  assign from_t1_iter66_to_t1_iter67_if_read = from_t1_iter66_to_t1_iter67__read;
  assign from_t1_iter66_to_t1_iter67_if_read_ce = 1'b1;
  assign from_t1_iter66_to_t1_iter67_if_write = from_t1_iter66_to_t1_iter67__write;
  assign from_t1_iter66_to_t1_iter67_if_write_ce = 1'b1;
  assign from_t1_iter66_to_t1_iter67_reset = ~ ap_rst_n;
  assign from_t1_iter67_to_t1_iter68_clk = ap_clk;
  assign from_t1_iter67_to_t1_iter68_if_din = from_t1_iter67_to_t1_iter68__din;
  assign from_t1_iter67_to_t1_iter68__dout = from_t1_iter67_to_t1_iter68_if_dout;
  assign from_t1_iter67_to_t1_iter68__empty_n = from_t1_iter67_to_t1_iter68_if_empty_n;
  assign from_t1_iter67_to_t1_iter68__full_n = from_t1_iter67_to_t1_iter68_if_full_n;
  assign from_t1_iter67_to_t1_iter68_if_read = from_t1_iter67_to_t1_iter68__read;
  assign from_t1_iter67_to_t1_iter68_if_read_ce = 1'b1;
  assign from_t1_iter67_to_t1_iter68_if_write = from_t1_iter67_to_t1_iter68__write;
  assign from_t1_iter67_to_t1_iter68_if_write_ce = 1'b1;
  assign from_t1_iter67_to_t1_iter68_reset = ~ ap_rst_n;
  assign from_t1_iter68_to_t1_iter69_clk = ap_clk;
  assign from_t1_iter68_to_t1_iter69_if_din = from_t1_iter68_to_t1_iter69__din;
  assign from_t1_iter68_to_t1_iter69__dout = from_t1_iter68_to_t1_iter69_if_dout;
  assign from_t1_iter68_to_t1_iter69__empty_n = from_t1_iter68_to_t1_iter69_if_empty_n;
  assign from_t1_iter68_to_t1_iter69__full_n = from_t1_iter68_to_t1_iter69_if_full_n;
  assign from_t1_iter68_to_t1_iter69_if_read = from_t1_iter68_to_t1_iter69__read;
  assign from_t1_iter68_to_t1_iter69_if_read_ce = 1'b1;
  assign from_t1_iter68_to_t1_iter69_if_write = from_t1_iter68_to_t1_iter69__write;
  assign from_t1_iter68_to_t1_iter69_if_write_ce = 1'b1;
  assign from_t1_iter68_to_t1_iter69_reset = ~ ap_rst_n;
  assign from_t1_iter69_to_t1_iter70_clk = ap_clk;
  assign from_t1_iter69_to_t1_iter70_if_din = from_t1_iter69_to_t1_iter70__din;
  assign from_t1_iter69_to_t1_iter70__dout = from_t1_iter69_to_t1_iter70_if_dout;
  assign from_t1_iter69_to_t1_iter70__empty_n = from_t1_iter69_to_t1_iter70_if_empty_n;
  assign from_t1_iter69_to_t1_iter70__full_n = from_t1_iter69_to_t1_iter70_if_full_n;
  assign from_t1_iter69_to_t1_iter70_if_read = from_t1_iter69_to_t1_iter70__read;
  assign from_t1_iter69_to_t1_iter70_if_read_ce = 1'b1;
  assign from_t1_iter69_to_t1_iter70_if_write = from_t1_iter69_to_t1_iter70__write;
  assign from_t1_iter69_to_t1_iter70_if_write_ce = 1'b1;
  assign from_t1_iter69_to_t1_iter70_reset = ~ ap_rst_n;
  assign from_t1_iter6_to_t1_iter7_clk = ap_clk;
  assign from_t1_iter6_to_t1_iter7_if_din = from_t1_iter6_to_t1_iter7__din;
  assign from_t1_iter6_to_t1_iter7__dout = from_t1_iter6_to_t1_iter7_if_dout;
  assign from_t1_iter6_to_t1_iter7__empty_n = from_t1_iter6_to_t1_iter7_if_empty_n;
  assign from_t1_iter6_to_t1_iter7__full_n = from_t1_iter6_to_t1_iter7_if_full_n;
  assign from_t1_iter6_to_t1_iter7_if_read = from_t1_iter6_to_t1_iter7__read;
  assign from_t1_iter6_to_t1_iter7_if_read_ce = 1'b1;
  assign from_t1_iter6_to_t1_iter7_if_write = from_t1_iter6_to_t1_iter7__write;
  assign from_t1_iter6_to_t1_iter7_if_write_ce = 1'b1;
  assign from_t1_iter6_to_t1_iter7_reset = ~ ap_rst_n;
  assign from_t1_iter70_to_t1_iter71_clk = ap_clk;
  assign from_t1_iter70_to_t1_iter71_if_din = from_t1_iter70_to_t1_iter71__din;
  assign from_t1_iter70_to_t1_iter71__dout = from_t1_iter70_to_t1_iter71_if_dout;
  assign from_t1_iter70_to_t1_iter71__empty_n = from_t1_iter70_to_t1_iter71_if_empty_n;
  assign from_t1_iter70_to_t1_iter71__full_n = from_t1_iter70_to_t1_iter71_if_full_n;
  assign from_t1_iter70_to_t1_iter71_if_read = from_t1_iter70_to_t1_iter71__read;
  assign from_t1_iter70_to_t1_iter71_if_read_ce = 1'b1;
  assign from_t1_iter70_to_t1_iter71_if_write = from_t1_iter70_to_t1_iter71__write;
  assign from_t1_iter70_to_t1_iter71_if_write_ce = 1'b1;
  assign from_t1_iter70_to_t1_iter71_reset = ~ ap_rst_n;
  assign from_t1_iter71_to_t1_iter72_clk = ap_clk;
  assign from_t1_iter71_to_t1_iter72_if_din = from_t1_iter71_to_t1_iter72__din;
  assign from_t1_iter71_to_t1_iter72__dout = from_t1_iter71_to_t1_iter72_if_dout;
  assign from_t1_iter71_to_t1_iter72__empty_n = from_t1_iter71_to_t1_iter72_if_empty_n;
  assign from_t1_iter71_to_t1_iter72__full_n = from_t1_iter71_to_t1_iter72_if_full_n;
  assign from_t1_iter71_to_t1_iter72_if_read = from_t1_iter71_to_t1_iter72__read;
  assign from_t1_iter71_to_t1_iter72_if_read_ce = 1'b1;
  assign from_t1_iter71_to_t1_iter72_if_write = from_t1_iter71_to_t1_iter72__write;
  assign from_t1_iter71_to_t1_iter72_if_write_ce = 1'b1;
  assign from_t1_iter71_to_t1_iter72_reset = ~ ap_rst_n;
  assign from_t1_iter72_to_t1_iter73_clk = ap_clk;
  assign from_t1_iter72_to_t1_iter73_if_din = from_t1_iter72_to_t1_iter73__din;
  assign from_t1_iter72_to_t1_iter73__dout = from_t1_iter72_to_t1_iter73_if_dout;
  assign from_t1_iter72_to_t1_iter73__empty_n = from_t1_iter72_to_t1_iter73_if_empty_n;
  assign from_t1_iter72_to_t1_iter73__full_n = from_t1_iter72_to_t1_iter73_if_full_n;
  assign from_t1_iter72_to_t1_iter73_if_read = from_t1_iter72_to_t1_iter73__read;
  assign from_t1_iter72_to_t1_iter73_if_read_ce = 1'b1;
  assign from_t1_iter72_to_t1_iter73_if_write = from_t1_iter72_to_t1_iter73__write;
  assign from_t1_iter72_to_t1_iter73_if_write_ce = 1'b1;
  assign from_t1_iter72_to_t1_iter73_reset = ~ ap_rst_n;
  assign from_t1_iter73_to_t1_iter74_clk = ap_clk;
  assign from_t1_iter73_to_t1_iter74_if_din = from_t1_iter73_to_t1_iter74__din;
  assign from_t1_iter73_to_t1_iter74__dout = from_t1_iter73_to_t1_iter74_if_dout;
  assign from_t1_iter73_to_t1_iter74__empty_n = from_t1_iter73_to_t1_iter74_if_empty_n;
  assign from_t1_iter73_to_t1_iter74__full_n = from_t1_iter73_to_t1_iter74_if_full_n;
  assign from_t1_iter73_to_t1_iter74_if_read = from_t1_iter73_to_t1_iter74__read;
  assign from_t1_iter73_to_t1_iter74_if_read_ce = 1'b1;
  assign from_t1_iter73_to_t1_iter74_if_write = from_t1_iter73_to_t1_iter74__write;
  assign from_t1_iter73_to_t1_iter74_if_write_ce = 1'b1;
  assign from_t1_iter73_to_t1_iter74_reset = ~ ap_rst_n;
  assign from_t1_iter74_to_t1_iter75_clk = ap_clk;
  assign from_t1_iter74_to_t1_iter75_if_din = from_t1_iter74_to_t1_iter75__din;
  assign from_t1_iter74_to_t1_iter75__dout = from_t1_iter74_to_t1_iter75_if_dout;
  assign from_t1_iter74_to_t1_iter75__empty_n = from_t1_iter74_to_t1_iter75_if_empty_n;
  assign from_t1_iter74_to_t1_iter75__full_n = from_t1_iter74_to_t1_iter75_if_full_n;
  assign from_t1_iter74_to_t1_iter75_if_read = from_t1_iter74_to_t1_iter75__read;
  assign from_t1_iter74_to_t1_iter75_if_read_ce = 1'b1;
  assign from_t1_iter74_to_t1_iter75_if_write = from_t1_iter74_to_t1_iter75__write;
  assign from_t1_iter74_to_t1_iter75_if_write_ce = 1'b1;
  assign from_t1_iter74_to_t1_iter75_reset = ~ ap_rst_n;
  assign from_t1_iter75_to_t1_iter76_clk = ap_clk;
  assign from_t1_iter75_to_t1_iter76_if_din = from_t1_iter75_to_t1_iter76__din;
  assign from_t1_iter75_to_t1_iter76__dout = from_t1_iter75_to_t1_iter76_if_dout;
  assign from_t1_iter75_to_t1_iter76__empty_n = from_t1_iter75_to_t1_iter76_if_empty_n;
  assign from_t1_iter75_to_t1_iter76__full_n = from_t1_iter75_to_t1_iter76_if_full_n;
  assign from_t1_iter75_to_t1_iter76_if_read = from_t1_iter75_to_t1_iter76__read;
  assign from_t1_iter75_to_t1_iter76_if_read_ce = 1'b1;
  assign from_t1_iter75_to_t1_iter76_if_write = from_t1_iter75_to_t1_iter76__write;
  assign from_t1_iter75_to_t1_iter76_if_write_ce = 1'b1;
  assign from_t1_iter75_to_t1_iter76_reset = ~ ap_rst_n;
  assign from_t1_iter76_to_t1_iter77_clk = ap_clk;
  assign from_t1_iter76_to_t1_iter77_if_din = from_t1_iter76_to_t1_iter77__din;
  assign from_t1_iter76_to_t1_iter77__dout = from_t1_iter76_to_t1_iter77_if_dout;
  assign from_t1_iter76_to_t1_iter77__empty_n = from_t1_iter76_to_t1_iter77_if_empty_n;
  assign from_t1_iter76_to_t1_iter77__full_n = from_t1_iter76_to_t1_iter77_if_full_n;
  assign from_t1_iter76_to_t1_iter77_if_read = from_t1_iter76_to_t1_iter77__read;
  assign from_t1_iter76_to_t1_iter77_if_read_ce = 1'b1;
  assign from_t1_iter76_to_t1_iter77_if_write = from_t1_iter76_to_t1_iter77__write;
  assign from_t1_iter76_to_t1_iter77_if_write_ce = 1'b1;
  assign from_t1_iter76_to_t1_iter77_reset = ~ ap_rst_n;
  assign from_t1_iter77_to_t1_iter78_clk = ap_clk;
  assign from_t1_iter77_to_t1_iter78_if_din = from_t1_iter77_to_t1_iter78__din;
  assign from_t1_iter77_to_t1_iter78__dout = from_t1_iter77_to_t1_iter78_if_dout;
  assign from_t1_iter77_to_t1_iter78__empty_n = from_t1_iter77_to_t1_iter78_if_empty_n;
  assign from_t1_iter77_to_t1_iter78__full_n = from_t1_iter77_to_t1_iter78_if_full_n;
  assign from_t1_iter77_to_t1_iter78_if_read = from_t1_iter77_to_t1_iter78__read;
  assign from_t1_iter77_to_t1_iter78_if_read_ce = 1'b1;
  assign from_t1_iter77_to_t1_iter78_if_write = from_t1_iter77_to_t1_iter78__write;
  assign from_t1_iter77_to_t1_iter78_if_write_ce = 1'b1;
  assign from_t1_iter77_to_t1_iter78_reset = ~ ap_rst_n;
  assign from_t1_iter78_to_t1_iter79_clk = ap_clk;
  assign from_t1_iter78_to_t1_iter79_if_din = from_t1_iter78_to_t1_iter79__din;
  assign from_t1_iter78_to_t1_iter79__dout = from_t1_iter78_to_t1_iter79_if_dout;
  assign from_t1_iter78_to_t1_iter79__empty_n = from_t1_iter78_to_t1_iter79_if_empty_n;
  assign from_t1_iter78_to_t1_iter79__full_n = from_t1_iter78_to_t1_iter79_if_full_n;
  assign from_t1_iter78_to_t1_iter79_if_read = from_t1_iter78_to_t1_iter79__read;
  assign from_t1_iter78_to_t1_iter79_if_read_ce = 1'b1;
  assign from_t1_iter78_to_t1_iter79_if_write = from_t1_iter78_to_t1_iter79__write;
  assign from_t1_iter78_to_t1_iter79_if_write_ce = 1'b1;
  assign from_t1_iter78_to_t1_iter79_reset = ~ ap_rst_n;
  assign from_t1_iter79_to_t1_iter80_clk = ap_clk;
  assign from_t1_iter79_to_t1_iter80_if_din = from_t1_iter79_to_t1_iter80__din;
  assign from_t1_iter79_to_t1_iter80__dout = from_t1_iter79_to_t1_iter80_if_dout;
  assign from_t1_iter79_to_t1_iter80__empty_n = from_t1_iter79_to_t1_iter80_if_empty_n;
  assign from_t1_iter79_to_t1_iter80__full_n = from_t1_iter79_to_t1_iter80_if_full_n;
  assign from_t1_iter79_to_t1_iter80_if_read = from_t1_iter79_to_t1_iter80__read;
  assign from_t1_iter79_to_t1_iter80_if_read_ce = 1'b1;
  assign from_t1_iter79_to_t1_iter80_if_write = from_t1_iter79_to_t1_iter80__write;
  assign from_t1_iter79_to_t1_iter80_if_write_ce = 1'b1;
  assign from_t1_iter79_to_t1_iter80_reset = ~ ap_rst_n;
  assign from_t1_iter7_to_t1_iter8_clk = ap_clk;
  assign from_t1_iter7_to_t1_iter8_if_din = from_t1_iter7_to_t1_iter8__din;
  assign from_t1_iter7_to_t1_iter8__dout = from_t1_iter7_to_t1_iter8_if_dout;
  assign from_t1_iter7_to_t1_iter8__empty_n = from_t1_iter7_to_t1_iter8_if_empty_n;
  assign from_t1_iter7_to_t1_iter8__full_n = from_t1_iter7_to_t1_iter8_if_full_n;
  assign from_t1_iter7_to_t1_iter8_if_read = from_t1_iter7_to_t1_iter8__read;
  assign from_t1_iter7_to_t1_iter8_if_read_ce = 1'b1;
  assign from_t1_iter7_to_t1_iter8_if_write = from_t1_iter7_to_t1_iter8__write;
  assign from_t1_iter7_to_t1_iter8_if_write_ce = 1'b1;
  assign from_t1_iter7_to_t1_iter8_reset = ~ ap_rst_n;
  assign from_t1_iter80_to_t1_iter81_clk = ap_clk;
  assign from_t1_iter80_to_t1_iter81_if_din = from_t1_iter80_to_t1_iter81__din;
  assign from_t1_iter80_to_t1_iter81__dout = from_t1_iter80_to_t1_iter81_if_dout;
  assign from_t1_iter80_to_t1_iter81__empty_n = from_t1_iter80_to_t1_iter81_if_empty_n;
  assign from_t1_iter80_to_t1_iter81__full_n = from_t1_iter80_to_t1_iter81_if_full_n;
  assign from_t1_iter80_to_t1_iter81_if_read = from_t1_iter80_to_t1_iter81__read;
  assign from_t1_iter80_to_t1_iter81_if_read_ce = 1'b1;
  assign from_t1_iter80_to_t1_iter81_if_write = from_t1_iter80_to_t1_iter81__write;
  assign from_t1_iter80_to_t1_iter81_if_write_ce = 1'b1;
  assign from_t1_iter80_to_t1_iter81_reset = ~ ap_rst_n;
  assign from_t1_iter81_to_t1_iter82_clk = ap_clk;
  assign from_t1_iter81_to_t1_iter82_if_din = from_t1_iter81_to_t1_iter82__din;
  assign from_t1_iter81_to_t1_iter82__dout = from_t1_iter81_to_t1_iter82_if_dout;
  assign from_t1_iter81_to_t1_iter82__empty_n = from_t1_iter81_to_t1_iter82_if_empty_n;
  assign from_t1_iter81_to_t1_iter82__full_n = from_t1_iter81_to_t1_iter82_if_full_n;
  assign from_t1_iter81_to_t1_iter82_if_read = from_t1_iter81_to_t1_iter82__read;
  assign from_t1_iter81_to_t1_iter82_if_read_ce = 1'b1;
  assign from_t1_iter81_to_t1_iter82_if_write = from_t1_iter81_to_t1_iter82__write;
  assign from_t1_iter81_to_t1_iter82_if_write_ce = 1'b1;
  assign from_t1_iter81_to_t1_iter82_reset = ~ ap_rst_n;
  assign from_t1_iter82_to_t1_iter83_clk = ap_clk;
  assign from_t1_iter82_to_t1_iter83_if_din = from_t1_iter82_to_t1_iter83__din;
  assign from_t1_iter82_to_t1_iter83__dout = from_t1_iter82_to_t1_iter83_if_dout;
  assign from_t1_iter82_to_t1_iter83__empty_n = from_t1_iter82_to_t1_iter83_if_empty_n;
  assign from_t1_iter82_to_t1_iter83__full_n = from_t1_iter82_to_t1_iter83_if_full_n;
  assign from_t1_iter82_to_t1_iter83_if_read = from_t1_iter82_to_t1_iter83__read;
  assign from_t1_iter82_to_t1_iter83_if_read_ce = 1'b1;
  assign from_t1_iter82_to_t1_iter83_if_write = from_t1_iter82_to_t1_iter83__write;
  assign from_t1_iter82_to_t1_iter83_if_write_ce = 1'b1;
  assign from_t1_iter82_to_t1_iter83_reset = ~ ap_rst_n;
  assign from_t1_iter83_to_t1_iter84_clk = ap_clk;
  assign from_t1_iter83_to_t1_iter84_if_din = from_t1_iter83_to_t1_iter84__din;
  assign from_t1_iter83_to_t1_iter84__dout = from_t1_iter83_to_t1_iter84_if_dout;
  assign from_t1_iter83_to_t1_iter84__empty_n = from_t1_iter83_to_t1_iter84_if_empty_n;
  assign from_t1_iter83_to_t1_iter84__full_n = from_t1_iter83_to_t1_iter84_if_full_n;
  assign from_t1_iter83_to_t1_iter84_if_read = from_t1_iter83_to_t1_iter84__read;
  assign from_t1_iter83_to_t1_iter84_if_read_ce = 1'b1;
  assign from_t1_iter83_to_t1_iter84_if_write = from_t1_iter83_to_t1_iter84__write;
  assign from_t1_iter83_to_t1_iter84_if_write_ce = 1'b1;
  assign from_t1_iter83_to_t1_iter84_reset = ~ ap_rst_n;
  assign from_t1_iter84_to_t1_iter85_clk = ap_clk;
  assign from_t1_iter84_to_t1_iter85_if_din = from_t1_iter84_to_t1_iter85__din;
  assign from_t1_iter84_to_t1_iter85__dout = from_t1_iter84_to_t1_iter85_if_dout;
  assign from_t1_iter84_to_t1_iter85__empty_n = from_t1_iter84_to_t1_iter85_if_empty_n;
  assign from_t1_iter84_to_t1_iter85__full_n = from_t1_iter84_to_t1_iter85_if_full_n;
  assign from_t1_iter84_to_t1_iter85_if_read = from_t1_iter84_to_t1_iter85__read;
  assign from_t1_iter84_to_t1_iter85_if_read_ce = 1'b1;
  assign from_t1_iter84_to_t1_iter85_if_write = from_t1_iter84_to_t1_iter85__write;
  assign from_t1_iter84_to_t1_iter85_if_write_ce = 1'b1;
  assign from_t1_iter84_to_t1_iter85_reset = ~ ap_rst_n;
  assign from_t1_iter85_to_t1_iter86_clk = ap_clk;
  assign from_t1_iter85_to_t1_iter86_if_din = from_t1_iter85_to_t1_iter86__din;
  assign from_t1_iter85_to_t1_iter86__dout = from_t1_iter85_to_t1_iter86_if_dout;
  assign from_t1_iter85_to_t1_iter86__empty_n = from_t1_iter85_to_t1_iter86_if_empty_n;
  assign from_t1_iter85_to_t1_iter86__full_n = from_t1_iter85_to_t1_iter86_if_full_n;
  assign from_t1_iter85_to_t1_iter86_if_read = from_t1_iter85_to_t1_iter86__read;
  assign from_t1_iter85_to_t1_iter86_if_read_ce = 1'b1;
  assign from_t1_iter85_to_t1_iter86_if_write = from_t1_iter85_to_t1_iter86__write;
  assign from_t1_iter85_to_t1_iter86_if_write_ce = 1'b1;
  assign from_t1_iter85_to_t1_iter86_reset = ~ ap_rst_n;
  assign from_t1_iter86_to_t1_iter87_clk = ap_clk;
  assign from_t1_iter86_to_t1_iter87_if_din = from_t1_iter86_to_t1_iter87__din;
  assign from_t1_iter86_to_t1_iter87__dout = from_t1_iter86_to_t1_iter87_if_dout;
  assign from_t1_iter86_to_t1_iter87__empty_n = from_t1_iter86_to_t1_iter87_if_empty_n;
  assign from_t1_iter86_to_t1_iter87__full_n = from_t1_iter86_to_t1_iter87_if_full_n;
  assign from_t1_iter86_to_t1_iter87_if_read = from_t1_iter86_to_t1_iter87__read;
  assign from_t1_iter86_to_t1_iter87_if_read_ce = 1'b1;
  assign from_t1_iter86_to_t1_iter87_if_write = from_t1_iter86_to_t1_iter87__write;
  assign from_t1_iter86_to_t1_iter87_if_write_ce = 1'b1;
  assign from_t1_iter86_to_t1_iter87_reset = ~ ap_rst_n;
  assign from_t1_iter87_to_t1_iter88_clk = ap_clk;
  assign from_t1_iter87_to_t1_iter88_if_din = from_t1_iter87_to_t1_iter88__din;
  assign from_t1_iter87_to_t1_iter88__dout = from_t1_iter87_to_t1_iter88_if_dout;
  assign from_t1_iter87_to_t1_iter88__empty_n = from_t1_iter87_to_t1_iter88_if_empty_n;
  assign from_t1_iter87_to_t1_iter88__full_n = from_t1_iter87_to_t1_iter88_if_full_n;
  assign from_t1_iter87_to_t1_iter88_if_read = from_t1_iter87_to_t1_iter88__read;
  assign from_t1_iter87_to_t1_iter88_if_read_ce = 1'b1;
  assign from_t1_iter87_to_t1_iter88_if_write = from_t1_iter87_to_t1_iter88__write;
  assign from_t1_iter87_to_t1_iter88_if_write_ce = 1'b1;
  assign from_t1_iter87_to_t1_iter88_reset = ~ ap_rst_n;
  assign from_t1_iter88_to_t1_iter89_clk = ap_clk;
  assign from_t1_iter88_to_t1_iter89_if_din = from_t1_iter88_to_t1_iter89__din;
  assign from_t1_iter88_to_t1_iter89__dout = from_t1_iter88_to_t1_iter89_if_dout;
  assign from_t1_iter88_to_t1_iter89__empty_n = from_t1_iter88_to_t1_iter89_if_empty_n;
  assign from_t1_iter88_to_t1_iter89__full_n = from_t1_iter88_to_t1_iter89_if_full_n;
  assign from_t1_iter88_to_t1_iter89_if_read = from_t1_iter88_to_t1_iter89__read;
  assign from_t1_iter88_to_t1_iter89_if_read_ce = 1'b1;
  assign from_t1_iter88_to_t1_iter89_if_write = from_t1_iter88_to_t1_iter89__write;
  assign from_t1_iter88_to_t1_iter89_if_write_ce = 1'b1;
  assign from_t1_iter88_to_t1_iter89_reset = ~ ap_rst_n;
  assign from_t1_iter89_to_t1_iter90_clk = ap_clk;
  assign from_t1_iter89_to_t1_iter90_if_din = from_t1_iter89_to_t1_iter90__din;
  assign from_t1_iter89_to_t1_iter90__dout = from_t1_iter89_to_t1_iter90_if_dout;
  assign from_t1_iter89_to_t1_iter90__empty_n = from_t1_iter89_to_t1_iter90_if_empty_n;
  assign from_t1_iter89_to_t1_iter90__full_n = from_t1_iter89_to_t1_iter90_if_full_n;
  assign from_t1_iter89_to_t1_iter90_if_read = from_t1_iter89_to_t1_iter90__read;
  assign from_t1_iter89_to_t1_iter90_if_read_ce = 1'b1;
  assign from_t1_iter89_to_t1_iter90_if_write = from_t1_iter89_to_t1_iter90__write;
  assign from_t1_iter89_to_t1_iter90_if_write_ce = 1'b1;
  assign from_t1_iter89_to_t1_iter90_reset = ~ ap_rst_n;
  assign from_t1_iter8_to_t1_iter9_clk = ap_clk;
  assign from_t1_iter8_to_t1_iter9_if_din = from_t1_iter8_to_t1_iter9__din;
  assign from_t1_iter8_to_t1_iter9__dout = from_t1_iter8_to_t1_iter9_if_dout;
  assign from_t1_iter8_to_t1_iter9__empty_n = from_t1_iter8_to_t1_iter9_if_empty_n;
  assign from_t1_iter8_to_t1_iter9__full_n = from_t1_iter8_to_t1_iter9_if_full_n;
  assign from_t1_iter8_to_t1_iter9_if_read = from_t1_iter8_to_t1_iter9__read;
  assign from_t1_iter8_to_t1_iter9_if_read_ce = 1'b1;
  assign from_t1_iter8_to_t1_iter9_if_write = from_t1_iter8_to_t1_iter9__write;
  assign from_t1_iter8_to_t1_iter9_if_write_ce = 1'b1;
  assign from_t1_iter8_to_t1_iter9_reset = ~ ap_rst_n;
  assign from_t1_iter90_to_t1_iter91_clk = ap_clk;
  assign from_t1_iter90_to_t1_iter91_if_din = from_t1_iter90_to_t1_iter91__din;
  assign from_t1_iter90_to_t1_iter91__dout = from_t1_iter90_to_t1_iter91_if_dout;
  assign from_t1_iter90_to_t1_iter91__empty_n = from_t1_iter90_to_t1_iter91_if_empty_n;
  assign from_t1_iter90_to_t1_iter91__full_n = from_t1_iter90_to_t1_iter91_if_full_n;
  assign from_t1_iter90_to_t1_iter91_if_read = from_t1_iter90_to_t1_iter91__read;
  assign from_t1_iter90_to_t1_iter91_if_read_ce = 1'b1;
  assign from_t1_iter90_to_t1_iter91_if_write = from_t1_iter90_to_t1_iter91__write;
  assign from_t1_iter90_to_t1_iter91_if_write_ce = 1'b1;
  assign from_t1_iter90_to_t1_iter91_reset = ~ ap_rst_n;
  assign from_t1_iter91_to_t1_iter92_clk = ap_clk;
  assign from_t1_iter91_to_t1_iter92_if_din = from_t1_iter91_to_t1_iter92__din;
  assign from_t1_iter91_to_t1_iter92__dout = from_t1_iter91_to_t1_iter92_if_dout;
  assign from_t1_iter91_to_t1_iter92__empty_n = from_t1_iter91_to_t1_iter92_if_empty_n;
  assign from_t1_iter91_to_t1_iter92__full_n = from_t1_iter91_to_t1_iter92_if_full_n;
  assign from_t1_iter91_to_t1_iter92_if_read = from_t1_iter91_to_t1_iter92__read;
  assign from_t1_iter91_to_t1_iter92_if_read_ce = 1'b1;
  assign from_t1_iter91_to_t1_iter92_if_write = from_t1_iter91_to_t1_iter92__write;
  assign from_t1_iter91_to_t1_iter92_if_write_ce = 1'b1;
  assign from_t1_iter91_to_t1_iter92_reset = ~ ap_rst_n;
  assign from_t1_iter92_to_t1_iter93_clk = ap_clk;
  assign from_t1_iter92_to_t1_iter93_if_din = from_t1_iter92_to_t1_iter93__din;
  assign from_t1_iter92_to_t1_iter93__dout = from_t1_iter92_to_t1_iter93_if_dout;
  assign from_t1_iter92_to_t1_iter93__empty_n = from_t1_iter92_to_t1_iter93_if_empty_n;
  assign from_t1_iter92_to_t1_iter93__full_n = from_t1_iter92_to_t1_iter93_if_full_n;
  assign from_t1_iter92_to_t1_iter93_if_read = from_t1_iter92_to_t1_iter93__read;
  assign from_t1_iter92_to_t1_iter93_if_read_ce = 1'b1;
  assign from_t1_iter92_to_t1_iter93_if_write = from_t1_iter92_to_t1_iter93__write;
  assign from_t1_iter92_to_t1_iter93_if_write_ce = 1'b1;
  assign from_t1_iter92_to_t1_iter93_reset = ~ ap_rst_n;
  assign from_t1_iter93_to_t1_iter94_clk = ap_clk;
  assign from_t1_iter93_to_t1_iter94_if_din = from_t1_iter93_to_t1_iter94__din;
  assign from_t1_iter93_to_t1_iter94__dout = from_t1_iter93_to_t1_iter94_if_dout;
  assign from_t1_iter93_to_t1_iter94__empty_n = from_t1_iter93_to_t1_iter94_if_empty_n;
  assign from_t1_iter93_to_t1_iter94__full_n = from_t1_iter93_to_t1_iter94_if_full_n;
  assign from_t1_iter93_to_t1_iter94_if_read = from_t1_iter93_to_t1_iter94__read;
  assign from_t1_iter93_to_t1_iter94_if_read_ce = 1'b1;
  assign from_t1_iter93_to_t1_iter94_if_write = from_t1_iter93_to_t1_iter94__write;
  assign from_t1_iter93_to_t1_iter94_if_write_ce = 1'b1;
  assign from_t1_iter93_to_t1_iter94_reset = ~ ap_rst_n;
  assign from_t1_iter94_to_t1_iter95_clk = ap_clk;
  assign from_t1_iter94_to_t1_iter95_if_din = from_t1_iter94_to_t1_iter95__din;
  assign from_t1_iter94_to_t1_iter95__dout = from_t1_iter94_to_t1_iter95_if_dout;
  assign from_t1_iter94_to_t1_iter95__empty_n = from_t1_iter94_to_t1_iter95_if_empty_n;
  assign from_t1_iter94_to_t1_iter95__full_n = from_t1_iter94_to_t1_iter95_if_full_n;
  assign from_t1_iter94_to_t1_iter95_if_read = from_t1_iter94_to_t1_iter95__read;
  assign from_t1_iter94_to_t1_iter95_if_read_ce = 1'b1;
  assign from_t1_iter94_to_t1_iter95_if_write = from_t1_iter94_to_t1_iter95__write;
  assign from_t1_iter94_to_t1_iter95_if_write_ce = 1'b1;
  assign from_t1_iter94_to_t1_iter95_reset = ~ ap_rst_n;
  assign from_t1_iter95_to_t1_iter96_clk = ap_clk;
  assign from_t1_iter95_to_t1_iter96_if_din = from_t1_iter95_to_t1_iter96__din;
  assign from_t1_iter95_to_t1_iter96__dout = from_t1_iter95_to_t1_iter96_if_dout;
  assign from_t1_iter95_to_t1_iter96__empty_n = from_t1_iter95_to_t1_iter96_if_empty_n;
  assign from_t1_iter95_to_t1_iter96__full_n = from_t1_iter95_to_t1_iter96_if_full_n;
  assign from_t1_iter95_to_t1_iter96_if_read = from_t1_iter95_to_t1_iter96__read;
  assign from_t1_iter95_to_t1_iter96_if_read_ce = 1'b1;
  assign from_t1_iter95_to_t1_iter96_if_write = from_t1_iter95_to_t1_iter96__write;
  assign from_t1_iter95_to_t1_iter96_if_write_ce = 1'b1;
  assign from_t1_iter95_to_t1_iter96_reset = ~ ap_rst_n;
  assign from_t1_iter96_to_t1_iter97_clk = ap_clk;
  assign from_t1_iter96_to_t1_iter97_if_din = from_t1_iter96_to_t1_iter97__din;
  assign from_t1_iter96_to_t1_iter97__dout = from_t1_iter96_to_t1_iter97_if_dout;
  assign from_t1_iter96_to_t1_iter97__empty_n = from_t1_iter96_to_t1_iter97_if_empty_n;
  assign from_t1_iter96_to_t1_iter97__full_n = from_t1_iter96_to_t1_iter97_if_full_n;
  assign from_t1_iter96_to_t1_iter97_if_read = from_t1_iter96_to_t1_iter97__read;
  assign from_t1_iter96_to_t1_iter97_if_read_ce = 1'b1;
  assign from_t1_iter96_to_t1_iter97_if_write = from_t1_iter96_to_t1_iter97__write;
  assign from_t1_iter96_to_t1_iter97_if_write_ce = 1'b1;
  assign from_t1_iter96_to_t1_iter97_reset = ~ ap_rst_n;
  assign from_t1_iter97_to_t1_iter98_clk = ap_clk;
  assign from_t1_iter97_to_t1_iter98_if_din = from_t1_iter97_to_t1_iter98__din;
  assign from_t1_iter97_to_t1_iter98__dout = from_t1_iter97_to_t1_iter98_if_dout;
  assign from_t1_iter97_to_t1_iter98__empty_n = from_t1_iter97_to_t1_iter98_if_empty_n;
  assign from_t1_iter97_to_t1_iter98__full_n = from_t1_iter97_to_t1_iter98_if_full_n;
  assign from_t1_iter97_to_t1_iter98_if_read = from_t1_iter97_to_t1_iter98__read;
  assign from_t1_iter97_to_t1_iter98_if_read_ce = 1'b1;
  assign from_t1_iter97_to_t1_iter98_if_write = from_t1_iter97_to_t1_iter98__write;
  assign from_t1_iter97_to_t1_iter98_if_write_ce = 1'b1;
  assign from_t1_iter97_to_t1_iter98_reset = ~ ap_rst_n;
  assign from_t1_iter98_to_t1_iter99_clk = ap_clk;
  assign from_t1_iter98_to_t1_iter99_if_din = from_t1_iter98_to_t1_iter99__din;
  assign from_t1_iter98_to_t1_iter99__dout = from_t1_iter98_to_t1_iter99_if_dout;
  assign from_t1_iter98_to_t1_iter99__empty_n = from_t1_iter98_to_t1_iter99_if_empty_n;
  assign from_t1_iter98_to_t1_iter99__full_n = from_t1_iter98_to_t1_iter99_if_full_n;
  assign from_t1_iter98_to_t1_iter99_if_read = from_t1_iter98_to_t1_iter99__read;
  assign from_t1_iter98_to_t1_iter99_if_read_ce = 1'b1;
  assign from_t1_iter98_to_t1_iter99_if_write = from_t1_iter98_to_t1_iter99__write;
  assign from_t1_iter98_to_t1_iter99_if_write_ce = 1'b1;
  assign from_t1_iter98_to_t1_iter99_reset = ~ ap_rst_n;
  assign from_t1_iter99_to_t1_iter100_clk = ap_clk;
  assign from_t1_iter99_to_t1_iter100_if_din = from_t1_iter99_to_t1_iter100__din;
  assign from_t1_iter99_to_t1_iter100__dout = from_t1_iter99_to_t1_iter100_if_dout;
  assign from_t1_iter99_to_t1_iter100__empty_n = from_t1_iter99_to_t1_iter100_if_empty_n;
  assign from_t1_iter99_to_t1_iter100__full_n = from_t1_iter99_to_t1_iter100_if_full_n;
  assign from_t1_iter99_to_t1_iter100_if_read = from_t1_iter99_to_t1_iter100__read;
  assign from_t1_iter99_to_t1_iter100_if_read_ce = 1'b1;
  assign from_t1_iter99_to_t1_iter100_if_write = from_t1_iter99_to_t1_iter100__write;
  assign from_t1_iter99_to_t1_iter100_if_write_ce = 1'b1;
  assign from_t1_iter99_to_t1_iter100_reset = ~ ap_rst_n;
  assign from_t1_iter9_to_t1_iter10_clk = ap_clk;
  assign from_t1_iter9_to_t1_iter10_if_din = from_t1_iter9_to_t1_iter10__din;
  assign from_t1_iter9_to_t1_iter10__dout = from_t1_iter9_to_t1_iter10_if_dout;
  assign from_t1_iter9_to_t1_iter10__empty_n = from_t1_iter9_to_t1_iter10_if_empty_n;
  assign from_t1_iter9_to_t1_iter10__full_n = from_t1_iter9_to_t1_iter10_if_full_n;
  assign from_t1_iter9_to_t1_iter10_if_read = from_t1_iter9_to_t1_iter10__read;
  assign from_t1_iter9_to_t1_iter10_if_read_ce = 1'b1;
  assign from_t1_iter9_to_t1_iter10_if_write = from_t1_iter9_to_t1_iter10__write;
  assign from_t1_iter9_to_t1_iter10_if_write_ce = 1'b1;
  assign from_t1_iter9_to_t1_iter10_reset = ~ ap_rst_n;
  assign BurstRead_floatx16_0_ap_clk = ap_clk;
  assign BurstRead_floatx16_0__ap_done = BurstRead_floatx16_0_ap_done;
  assign BurstRead_floatx16_0__ap_idle = BurstRead_floatx16_0_ap_idle;
  assign BurstRead_floatx16_0__ap_ready = BurstRead_floatx16_0_ap_ready;
  assign BurstRead_floatx16_0_ap_rst_n = ap_rst_n;
  assign BurstRead_floatx16_0_ap_start = BurstRead_floatx16_0__ap_start;
  assign bank_0_t1_buf__din = BurstRead_floatx16_0_dest_din;
  assign BurstRead_floatx16_0_dest_full_n = bank_0_t1_buf__full_n;
  assign bank_0_t1_buf__write = BurstRead_floatx16_0_dest_write;
  assign BurstRead_floatx16_0_n = BurstRead_floatx16_0___coalesced_data_num__q0;
  assign BurstRead_floatx16_0_src_read_addr_offset = BurstRead_floatx16_0___bank_0_t1__q0;
  assign bank_0_t1_read_addr__din = BurstRead_floatx16_0_src_read_addr_s_din;
  assign BurstRead_floatx16_0_src_read_addr_s_full_n = bank_0_t1_read_addr__full_n;
  assign bank_0_t1_read_addr__write = BurstRead_floatx16_0_src_read_addr_s_write;
  assign BurstRead_floatx16_0_src_read_data_peek_dout = { 1'b0 , bank_0_t1_read_data__dout };
  assign BurstRead_floatx16_0_src_read_data_peek_empty_n = bank_0_t1_read_data__empty_n;
  assign BurstRead_floatx16_0_src_read_data_s_dout = { 1'b0 , bank_0_t1_read_data__dout };
  assign BurstRead_floatx16_0_src_read_data_s_empty_n = bank_0_t1_read_data__empty_n;
  assign bank_0_t1_read_data__read = BurstRead_floatx16_0_src_read_data_s_read;
  assign BurstRead_floatx16_0_src_write_addr_offset = BurstRead_floatx16_0___bank_0_t1__q0;
  assign bank_0_t1_write_addr__din = BurstRead_floatx16_0_src_write_addr_s_din;
  assign BurstRead_floatx16_0_src_write_addr_s_full_n = bank_0_t1_write_addr__full_n;
  assign bank_0_t1_write_addr__write = BurstRead_floatx16_0_src_write_addr_s_write;
  assign bank_0_t1_write_data__din = BurstRead_floatx16_0_src_write_data_din;
  assign BurstRead_floatx16_0_src_write_data_full_n = bank_0_t1_write_data__full_n;
  assign bank_0_t1_write_data__write = BurstRead_floatx16_0_src_write_data_write;
  assign BurstRead_floatx16_0_src_write_resp_peek_dout = { 1'b0 , bank_0_t1_write_resp__dout };
  assign BurstRead_floatx16_0_src_write_resp_peek_empty_n = bank_0_t1_write_resp__empty_n;
  assign BurstRead_floatx16_0_src_write_resp_s_dout = { 1'b0 , bank_0_t1_write_resp__dout };
  assign BurstRead_floatx16_0_src_write_resp_s_empty_n = bank_0_t1_write_resp__empty_n;
  assign bank_0_t1_write_resp__read = BurstRead_floatx16_0_src_write_resp_s_read;
  assign BurstWrite_floatx16_0_ap_clk = ap_clk;
  assign BurstWrite_floatx16_0__ap_done = BurstWrite_floatx16_0_ap_done;
  assign BurstWrite_floatx16_0__ap_idle = BurstWrite_floatx16_0_ap_idle;
  assign BurstWrite_floatx16_0__ap_ready = BurstWrite_floatx16_0_ap_ready;
  assign BurstWrite_floatx16_0_ap_rst_n = ap_rst_n;
  assign BurstWrite_floatx16_0_ap_start = BurstWrite_floatx16_0__ap_start;
  assign BurstWrite_floatx16_0_dest_read_addr_offset = BurstWrite_floatx16_0___bank_1_t0__q0;
  assign bank_1_t0_read_addr__din = BurstWrite_floatx16_0_dest_read_addr_s_din;
  assign BurstWrite_floatx16_0_dest_read_addr_s_full_n = bank_1_t0_read_addr__full_n;
  assign bank_1_t0_read_addr__write = BurstWrite_floatx16_0_dest_read_addr_s_write;
  assign BurstWrite_floatx16_0_dest_read_data_peek_dout = { 1'b0 , bank_1_t0_read_data__dout };
  assign BurstWrite_floatx16_0_dest_read_data_peek_empty_n = bank_1_t0_read_data__empty_n;
  assign BurstWrite_floatx16_0_dest_read_data_s_dout = { 1'b0 , bank_1_t0_read_data__dout };
  assign BurstWrite_floatx16_0_dest_read_data_s_empty_n = bank_1_t0_read_data__empty_n;
  assign bank_1_t0_read_data__read = BurstWrite_floatx16_0_dest_read_data_s_read;
  assign BurstWrite_floatx16_0_dest_write_addr_offset = BurstWrite_floatx16_0___bank_1_t0__q0;
  assign bank_1_t0_write_addr__din = BurstWrite_floatx16_0_dest_write_addr_s_din;
  assign BurstWrite_floatx16_0_dest_write_addr_s_full_n = bank_1_t0_write_addr__full_n;
  assign bank_1_t0_write_addr__write = BurstWrite_floatx16_0_dest_write_addr_s_write;
  assign bank_1_t0_write_data__din = BurstWrite_floatx16_0_dest_write_data_din;
  assign BurstWrite_floatx16_0_dest_write_data_full_n = bank_1_t0_write_data__full_n;
  assign bank_1_t0_write_data__write = BurstWrite_floatx16_0_dest_write_data_write;
  assign BurstWrite_floatx16_0_dest_write_resp_peek_dout = { 1'b0 , bank_1_t0_write_resp__dout };
  assign BurstWrite_floatx16_0_dest_write_resp_peek_empty_n = bank_1_t0_write_resp__empty_n;
  assign BurstWrite_floatx16_0_dest_write_resp_s_dout = { 1'b0 , bank_1_t0_write_resp__dout };
  assign BurstWrite_floatx16_0_dest_write_resp_s_empty_n = bank_1_t0_write_resp__empty_n;
  assign bank_1_t0_write_resp__read = BurstWrite_floatx16_0_dest_write_resp_s_read;
  assign BurstWrite_floatx16_0_n = BurstWrite_floatx16_0___coalesced_data_num__q0;
  assign BurstWrite_floatx16_0_src_peek_dout = bank_1_t0_buf__dout;
  assign BurstWrite_floatx16_0_src_peek_empty_n = bank_1_t0_buf__empty_n;
  assign BurstWrite_floatx16_0_src_s_dout = bank_1_t0_buf__dout;
  assign BurstWrite_floatx16_0_src_s_empty_n = bank_1_t0_buf__empty_n;
  assign bank_1_t0_buf__read = BurstWrite_floatx16_0_src_s_read;
  assign Module0Func_0_ap_clk = ap_clk;
  assign Module0Func_0_ap_rst_n = ap_rst_n;
  assign Module0Func_0_ap_start = Module0Func_0__ap_start;
  assign Module0Func_0_dram_t1_bank_0_fifo_peek_dout = bank_0_t1_buf__dout;
  assign Module0Func_0_dram_t1_bank_0_fifo_peek_empty_n = bank_0_t1_buf__empty_n;
  assign Module0Func_0_dram_t1_bank_0_fifo_s_dout = bank_0_t1_buf__dout;
  assign Module0Func_0_dram_t1_bank_0_fifo_s_empty_n = bank_0_t1_buf__empty_n;
  assign bank_0_t1_buf__read = Module0Func_0_dram_t1_bank_0_fifo_s_read;
  assign from_t1_bank_0_to_t1_iter1__din = Module0Func_0_fifo_st_0_din;
  assign Module0Func_0_fifo_st_0_full_n = from_t1_bank_0_to_t1_iter1__full_n;
  assign from_t1_bank_0_to_t1_iter1__write = Module0Func_0_fifo_st_0_write;
  assign Module1Func_0_ap_clk = ap_clk;
  assign Module1Func_0_ap_rst_n = ap_rst_n;
  assign Module1Func_0_ap_start = Module1Func_0__ap_start;
  assign Module1Func_0_fifo_ld_0_peek_dout = from_t1_bank_0_to_t1_iter1__dout;
  assign Module1Func_0_fifo_ld_0_peek_empty_n = from_t1_bank_0_to_t1_iter1__empty_n;
  assign Module1Func_0_fifo_ld_0_s_dout = from_t1_bank_0_to_t1_iter1__dout;
  assign Module1Func_0_fifo_ld_0_s_empty_n = from_t1_bank_0_to_t1_iter1__empty_n;
  assign from_t1_bank_0_to_t1_iter1__read = Module1Func_0_fifo_ld_0_s_read;
  assign from_t1_iter1_to_t1_iter2__din = Module1Func_0_fifo_st_0_din;
  assign Module1Func_0_fifo_st_0_full_n = from_t1_iter1_to_t1_iter2__full_n;
  assign from_t1_iter1_to_t1_iter2__write = Module1Func_0_fifo_st_0_write;
  assign Module2Func_0_ap_clk = ap_clk;
  assign Module2Func_0_ap_rst_n = ap_rst_n;
  assign Module2Func_0_ap_start = Module2Func_0__ap_start;
  assign Module2Func_0_fifo_ld_0_peek_dout = from_t1_iter1_to_t1_iter2__dout;
  assign Module2Func_0_fifo_ld_0_peek_empty_n = from_t1_iter1_to_t1_iter2__empty_n;
  assign Module2Func_0_fifo_ld_0_s_dout = from_t1_iter1_to_t1_iter2__dout;
  assign Module2Func_0_fifo_ld_0_s_empty_n = from_t1_iter1_to_t1_iter2__empty_n;
  assign from_t1_iter1_to_t1_iter2__read = Module2Func_0_fifo_ld_0_s_read;
  assign from_t1_iter2_to_t1_iter3__din = Module2Func_0_fifo_st_0_din;
  assign Module2Func_0_fifo_st_0_full_n = from_t1_iter2_to_t1_iter3__full_n;
  assign from_t1_iter2_to_t1_iter3__write = Module2Func_0_fifo_st_0_write;
  assign Module2Func_1_ap_clk = ap_clk;
  assign Module2Func_1_ap_rst_n = ap_rst_n;
  assign Module2Func_1_ap_start = Module2Func_1__ap_start;
  assign Module2Func_1_fifo_ld_0_peek_dout = from_t1_iter2_to_t1_iter3__dout;
  assign Module2Func_1_fifo_ld_0_peek_empty_n = from_t1_iter2_to_t1_iter3__empty_n;
  assign Module2Func_1_fifo_ld_0_s_dout = from_t1_iter2_to_t1_iter3__dout;
  assign Module2Func_1_fifo_ld_0_s_empty_n = from_t1_iter2_to_t1_iter3__empty_n;
  assign from_t1_iter2_to_t1_iter3__read = Module2Func_1_fifo_ld_0_s_read;
  assign from_t1_iter3_to_t1_iter4__din = Module2Func_1_fifo_st_0_din;
  assign Module2Func_1_fifo_st_0_full_n = from_t1_iter3_to_t1_iter4__full_n;
  assign from_t1_iter3_to_t1_iter4__write = Module2Func_1_fifo_st_0_write;
  assign Module2Func_2_ap_clk = ap_clk;
  assign Module2Func_2_ap_rst_n = ap_rst_n;
  assign Module2Func_2_ap_start = Module2Func_2__ap_start;
  assign Module2Func_2_fifo_ld_0_peek_dout = from_t1_iter3_to_t1_iter4__dout;
  assign Module2Func_2_fifo_ld_0_peek_empty_n = from_t1_iter3_to_t1_iter4__empty_n;
  assign Module2Func_2_fifo_ld_0_s_dout = from_t1_iter3_to_t1_iter4__dout;
  assign Module2Func_2_fifo_ld_0_s_empty_n = from_t1_iter3_to_t1_iter4__empty_n;
  assign from_t1_iter3_to_t1_iter4__read = Module2Func_2_fifo_ld_0_s_read;
  assign from_t1_iter4_to_t1_iter5__din = Module2Func_2_fifo_st_0_din;
  assign Module2Func_2_fifo_st_0_full_n = from_t1_iter4_to_t1_iter5__full_n;
  assign from_t1_iter4_to_t1_iter5__write = Module2Func_2_fifo_st_0_write;
  assign Module2Func_3_ap_clk = ap_clk;
  assign Module2Func_3_ap_rst_n = ap_rst_n;
  assign Module2Func_3_ap_start = Module2Func_3__ap_start;
  assign Module2Func_3_fifo_ld_0_peek_dout = from_t1_iter4_to_t1_iter5__dout;
  assign Module2Func_3_fifo_ld_0_peek_empty_n = from_t1_iter4_to_t1_iter5__empty_n;
  assign Module2Func_3_fifo_ld_0_s_dout = from_t1_iter4_to_t1_iter5__dout;
  assign Module2Func_3_fifo_ld_0_s_empty_n = from_t1_iter4_to_t1_iter5__empty_n;
  assign from_t1_iter4_to_t1_iter5__read = Module2Func_3_fifo_ld_0_s_read;
  assign from_t1_iter5_to_t1_iter6__din = Module2Func_3_fifo_st_0_din;
  assign Module2Func_3_fifo_st_0_full_n = from_t1_iter5_to_t1_iter6__full_n;
  assign from_t1_iter5_to_t1_iter6__write = Module2Func_3_fifo_st_0_write;
  assign Module2Func_4_ap_clk = ap_clk;
  assign Module2Func_4_ap_rst_n = ap_rst_n;
  assign Module2Func_4_ap_start = Module2Func_4__ap_start;
  assign Module2Func_4_fifo_ld_0_peek_dout = from_t1_iter5_to_t1_iter6__dout;
  assign Module2Func_4_fifo_ld_0_peek_empty_n = from_t1_iter5_to_t1_iter6__empty_n;
  assign Module2Func_4_fifo_ld_0_s_dout = from_t1_iter5_to_t1_iter6__dout;
  assign Module2Func_4_fifo_ld_0_s_empty_n = from_t1_iter5_to_t1_iter6__empty_n;
  assign from_t1_iter5_to_t1_iter6__read = Module2Func_4_fifo_ld_0_s_read;
  assign from_t1_iter6_to_t1_iter7__din = Module2Func_4_fifo_st_0_din;
  assign Module2Func_4_fifo_st_0_full_n = from_t1_iter6_to_t1_iter7__full_n;
  assign from_t1_iter6_to_t1_iter7__write = Module2Func_4_fifo_st_0_write;
  assign Module2Func_5_ap_clk = ap_clk;
  assign Module2Func_5_ap_rst_n = ap_rst_n;
  assign Module2Func_5_ap_start = Module2Func_5__ap_start;
  assign Module2Func_5_fifo_ld_0_peek_dout = from_t1_iter6_to_t1_iter7__dout;
  assign Module2Func_5_fifo_ld_0_peek_empty_n = from_t1_iter6_to_t1_iter7__empty_n;
  assign Module2Func_5_fifo_ld_0_s_dout = from_t1_iter6_to_t1_iter7__dout;
  assign Module2Func_5_fifo_ld_0_s_empty_n = from_t1_iter6_to_t1_iter7__empty_n;
  assign from_t1_iter6_to_t1_iter7__read = Module2Func_5_fifo_ld_0_s_read;
  assign from_t1_iter7_to_t1_iter8__din = Module2Func_5_fifo_st_0_din;
  assign Module2Func_5_fifo_st_0_full_n = from_t1_iter7_to_t1_iter8__full_n;
  assign from_t1_iter7_to_t1_iter8__write = Module2Func_5_fifo_st_0_write;
  assign Module2Func_6_ap_clk = ap_clk;
  assign Module2Func_6_ap_rst_n = ap_rst_n;
  assign Module2Func_6_ap_start = Module2Func_6__ap_start;
  assign Module2Func_6_fifo_ld_0_peek_dout = from_t1_iter7_to_t1_iter8__dout;
  assign Module2Func_6_fifo_ld_0_peek_empty_n = from_t1_iter7_to_t1_iter8__empty_n;
  assign Module2Func_6_fifo_ld_0_s_dout = from_t1_iter7_to_t1_iter8__dout;
  assign Module2Func_6_fifo_ld_0_s_empty_n = from_t1_iter7_to_t1_iter8__empty_n;
  assign from_t1_iter7_to_t1_iter8__read = Module2Func_6_fifo_ld_0_s_read;
  assign from_t1_iter8_to_t1_iter9__din = Module2Func_6_fifo_st_0_din;
  assign Module2Func_6_fifo_st_0_full_n = from_t1_iter8_to_t1_iter9__full_n;
  assign from_t1_iter8_to_t1_iter9__write = Module2Func_6_fifo_st_0_write;
  assign Module2Func_7_ap_clk = ap_clk;
  assign Module2Func_7_ap_rst_n = ap_rst_n;
  assign Module2Func_7_ap_start = Module2Func_7__ap_start;
  assign Module2Func_7_fifo_ld_0_peek_dout = from_t1_iter8_to_t1_iter9__dout;
  assign Module2Func_7_fifo_ld_0_peek_empty_n = from_t1_iter8_to_t1_iter9__empty_n;
  assign Module2Func_7_fifo_ld_0_s_dout = from_t1_iter8_to_t1_iter9__dout;
  assign Module2Func_7_fifo_ld_0_s_empty_n = from_t1_iter8_to_t1_iter9__empty_n;
  assign from_t1_iter8_to_t1_iter9__read = Module2Func_7_fifo_ld_0_s_read;
  assign from_t1_iter9_to_t1_iter10__din = Module2Func_7_fifo_st_0_din;
  assign Module2Func_7_fifo_st_0_full_n = from_t1_iter9_to_t1_iter10__full_n;
  assign from_t1_iter9_to_t1_iter10__write = Module2Func_7_fifo_st_0_write;
  assign Module2Func_8_ap_clk = ap_clk;
  assign Module2Func_8_ap_rst_n = ap_rst_n;
  assign Module2Func_8_ap_start = Module2Func_8__ap_start;
  assign Module2Func_8_fifo_ld_0_peek_dout = from_t1_iter9_to_t1_iter10__dout;
  assign Module2Func_8_fifo_ld_0_peek_empty_n = from_t1_iter9_to_t1_iter10__empty_n;
  assign Module2Func_8_fifo_ld_0_s_dout = from_t1_iter9_to_t1_iter10__dout;
  assign Module2Func_8_fifo_ld_0_s_empty_n = from_t1_iter9_to_t1_iter10__empty_n;
  assign from_t1_iter9_to_t1_iter10__read = Module2Func_8_fifo_ld_0_s_read;
  assign from_t1_iter10_to_t1_iter11__din = Module2Func_8_fifo_st_0_din;
  assign Module2Func_8_fifo_st_0_full_n = from_t1_iter10_to_t1_iter11__full_n;
  assign from_t1_iter10_to_t1_iter11__write = Module2Func_8_fifo_st_0_write;
  assign Module2Func_9_ap_clk = ap_clk;
  assign Module2Func_9_ap_rst_n = ap_rst_n;
  assign Module2Func_9_ap_start = Module2Func_9__ap_start;
  assign Module2Func_9_fifo_ld_0_peek_dout = from_t1_iter10_to_t1_iter11__dout;
  assign Module2Func_9_fifo_ld_0_peek_empty_n = from_t1_iter10_to_t1_iter11__empty_n;
  assign Module2Func_9_fifo_ld_0_s_dout = from_t1_iter10_to_t1_iter11__dout;
  assign Module2Func_9_fifo_ld_0_s_empty_n = from_t1_iter10_to_t1_iter11__empty_n;
  assign from_t1_iter10_to_t1_iter11__read = Module2Func_9_fifo_ld_0_s_read;
  assign from_t1_iter11_to_t1_iter12__din = Module2Func_9_fifo_st_0_din;
  assign Module2Func_9_fifo_st_0_full_n = from_t1_iter11_to_t1_iter12__full_n;
  assign from_t1_iter11_to_t1_iter12__write = Module2Func_9_fifo_st_0_write;
  assign Module2Func_10_ap_clk = ap_clk;
  assign Module2Func_10_ap_rst_n = ap_rst_n;
  assign Module2Func_10_ap_start = Module2Func_10__ap_start;
  assign Module2Func_10_fifo_ld_0_peek_dout = from_t1_iter11_to_t1_iter12__dout;
  assign Module2Func_10_fifo_ld_0_peek_empty_n = from_t1_iter11_to_t1_iter12__empty_n;
  assign Module2Func_10_fifo_ld_0_s_dout = from_t1_iter11_to_t1_iter12__dout;
  assign Module2Func_10_fifo_ld_0_s_empty_n = from_t1_iter11_to_t1_iter12__empty_n;
  assign from_t1_iter11_to_t1_iter12__read = Module2Func_10_fifo_ld_0_s_read;
  assign from_t1_iter12_to_t1_iter13__din = Module2Func_10_fifo_st_0_din;
  assign Module2Func_10_fifo_st_0_full_n = from_t1_iter12_to_t1_iter13__full_n;
  assign from_t1_iter12_to_t1_iter13__write = Module2Func_10_fifo_st_0_write;
  assign Module2Func_11_ap_clk = ap_clk;
  assign Module2Func_11_ap_rst_n = ap_rst_n;
  assign Module2Func_11_ap_start = Module2Func_11__ap_start;
  assign Module2Func_11_fifo_ld_0_peek_dout = from_t1_iter12_to_t1_iter13__dout;
  assign Module2Func_11_fifo_ld_0_peek_empty_n = from_t1_iter12_to_t1_iter13__empty_n;
  assign Module2Func_11_fifo_ld_0_s_dout = from_t1_iter12_to_t1_iter13__dout;
  assign Module2Func_11_fifo_ld_0_s_empty_n = from_t1_iter12_to_t1_iter13__empty_n;
  assign from_t1_iter12_to_t1_iter13__read = Module2Func_11_fifo_ld_0_s_read;
  assign from_t1_iter13_to_t1_iter14__din = Module2Func_11_fifo_st_0_din;
  assign Module2Func_11_fifo_st_0_full_n = from_t1_iter13_to_t1_iter14__full_n;
  assign from_t1_iter13_to_t1_iter14__write = Module2Func_11_fifo_st_0_write;
  assign Module2Func_12_ap_clk = ap_clk;
  assign Module2Func_12_ap_rst_n = ap_rst_n;
  assign Module2Func_12_ap_start = Module2Func_12__ap_start;
  assign Module2Func_12_fifo_ld_0_peek_dout = from_t1_iter13_to_t1_iter14__dout;
  assign Module2Func_12_fifo_ld_0_peek_empty_n = from_t1_iter13_to_t1_iter14__empty_n;
  assign Module2Func_12_fifo_ld_0_s_dout = from_t1_iter13_to_t1_iter14__dout;
  assign Module2Func_12_fifo_ld_0_s_empty_n = from_t1_iter13_to_t1_iter14__empty_n;
  assign from_t1_iter13_to_t1_iter14__read = Module2Func_12_fifo_ld_0_s_read;
  assign from_t1_iter14_to_t1_iter15__din = Module2Func_12_fifo_st_0_din;
  assign Module2Func_12_fifo_st_0_full_n = from_t1_iter14_to_t1_iter15__full_n;
  assign from_t1_iter14_to_t1_iter15__write = Module2Func_12_fifo_st_0_write;
  assign Module2Func_13_ap_clk = ap_clk;
  assign Module2Func_13_ap_rst_n = ap_rst_n;
  assign Module2Func_13_ap_start = Module2Func_13__ap_start;
  assign Module2Func_13_fifo_ld_0_peek_dout = from_t1_iter14_to_t1_iter15__dout;
  assign Module2Func_13_fifo_ld_0_peek_empty_n = from_t1_iter14_to_t1_iter15__empty_n;
  assign Module2Func_13_fifo_ld_0_s_dout = from_t1_iter14_to_t1_iter15__dout;
  assign Module2Func_13_fifo_ld_0_s_empty_n = from_t1_iter14_to_t1_iter15__empty_n;
  assign from_t1_iter14_to_t1_iter15__read = Module2Func_13_fifo_ld_0_s_read;
  assign from_t1_iter15_to_t1_iter16__din = Module2Func_13_fifo_st_0_din;
  assign Module2Func_13_fifo_st_0_full_n = from_t1_iter15_to_t1_iter16__full_n;
  assign from_t1_iter15_to_t1_iter16__write = Module2Func_13_fifo_st_0_write;
  assign Module2Func_14_ap_clk = ap_clk;
  assign Module2Func_14_ap_rst_n = ap_rst_n;
  assign Module2Func_14_ap_start = Module2Func_14__ap_start;
  assign Module2Func_14_fifo_ld_0_peek_dout = from_t1_iter15_to_t1_iter16__dout;
  assign Module2Func_14_fifo_ld_0_peek_empty_n = from_t1_iter15_to_t1_iter16__empty_n;
  assign Module2Func_14_fifo_ld_0_s_dout = from_t1_iter15_to_t1_iter16__dout;
  assign Module2Func_14_fifo_ld_0_s_empty_n = from_t1_iter15_to_t1_iter16__empty_n;
  assign from_t1_iter15_to_t1_iter16__read = Module2Func_14_fifo_ld_0_s_read;
  assign from_t1_iter16_to_t1_iter17__din = Module2Func_14_fifo_st_0_din;
  assign Module2Func_14_fifo_st_0_full_n = from_t1_iter16_to_t1_iter17__full_n;
  assign from_t1_iter16_to_t1_iter17__write = Module2Func_14_fifo_st_0_write;
  assign Module2Func_15_ap_clk = ap_clk;
  assign Module2Func_15_ap_rst_n = ap_rst_n;
  assign Module2Func_15_ap_start = Module2Func_15__ap_start;
  assign Module2Func_15_fifo_ld_0_peek_dout = from_t1_iter16_to_t1_iter17__dout;
  assign Module2Func_15_fifo_ld_0_peek_empty_n = from_t1_iter16_to_t1_iter17__empty_n;
  assign Module2Func_15_fifo_ld_0_s_dout = from_t1_iter16_to_t1_iter17__dout;
  assign Module2Func_15_fifo_ld_0_s_empty_n = from_t1_iter16_to_t1_iter17__empty_n;
  assign from_t1_iter16_to_t1_iter17__read = Module2Func_15_fifo_ld_0_s_read;
  assign from_t1_iter17_to_t1_iter18__din = Module2Func_15_fifo_st_0_din;
  assign Module2Func_15_fifo_st_0_full_n = from_t1_iter17_to_t1_iter18__full_n;
  assign from_t1_iter17_to_t1_iter18__write = Module2Func_15_fifo_st_0_write;
  assign Module2Func_16_ap_clk = ap_clk;
  assign Module2Func_16_ap_rst_n = ap_rst_n;
  assign Module2Func_16_ap_start = Module2Func_16__ap_start;
  assign Module2Func_16_fifo_ld_0_peek_dout = from_t1_iter17_to_t1_iter18__dout;
  assign Module2Func_16_fifo_ld_0_peek_empty_n = from_t1_iter17_to_t1_iter18__empty_n;
  assign Module2Func_16_fifo_ld_0_s_dout = from_t1_iter17_to_t1_iter18__dout;
  assign Module2Func_16_fifo_ld_0_s_empty_n = from_t1_iter17_to_t1_iter18__empty_n;
  assign from_t1_iter17_to_t1_iter18__read = Module2Func_16_fifo_ld_0_s_read;
  assign from_t1_iter18_to_t1_iter19__din = Module2Func_16_fifo_st_0_din;
  assign Module2Func_16_fifo_st_0_full_n = from_t1_iter18_to_t1_iter19__full_n;
  assign from_t1_iter18_to_t1_iter19__write = Module2Func_16_fifo_st_0_write;
  assign Module2Func_17_ap_clk = ap_clk;
  assign Module2Func_17_ap_rst_n = ap_rst_n;
  assign Module2Func_17_ap_start = Module2Func_17__ap_start;
  assign Module2Func_17_fifo_ld_0_peek_dout = from_t1_iter18_to_t1_iter19__dout;
  assign Module2Func_17_fifo_ld_0_peek_empty_n = from_t1_iter18_to_t1_iter19__empty_n;
  assign Module2Func_17_fifo_ld_0_s_dout = from_t1_iter18_to_t1_iter19__dout;
  assign Module2Func_17_fifo_ld_0_s_empty_n = from_t1_iter18_to_t1_iter19__empty_n;
  assign from_t1_iter18_to_t1_iter19__read = Module2Func_17_fifo_ld_0_s_read;
  assign from_t1_iter19_to_t1_iter20__din = Module2Func_17_fifo_st_0_din;
  assign Module2Func_17_fifo_st_0_full_n = from_t1_iter19_to_t1_iter20__full_n;
  assign from_t1_iter19_to_t1_iter20__write = Module2Func_17_fifo_st_0_write;
  assign Module2Func_18_ap_clk = ap_clk;
  assign Module2Func_18_ap_rst_n = ap_rst_n;
  assign Module2Func_18_ap_start = Module2Func_18__ap_start;
  assign Module2Func_18_fifo_ld_0_peek_dout = from_t1_iter19_to_t1_iter20__dout;
  assign Module2Func_18_fifo_ld_0_peek_empty_n = from_t1_iter19_to_t1_iter20__empty_n;
  assign Module2Func_18_fifo_ld_0_s_dout = from_t1_iter19_to_t1_iter20__dout;
  assign Module2Func_18_fifo_ld_0_s_empty_n = from_t1_iter19_to_t1_iter20__empty_n;
  assign from_t1_iter19_to_t1_iter20__read = Module2Func_18_fifo_ld_0_s_read;
  assign from_t1_iter20_to_t1_iter21__din = Module2Func_18_fifo_st_0_din;
  assign Module2Func_18_fifo_st_0_full_n = from_t1_iter20_to_t1_iter21__full_n;
  assign from_t1_iter20_to_t1_iter21__write = Module2Func_18_fifo_st_0_write;
  assign Module2Func_19_ap_clk = ap_clk;
  assign Module2Func_19_ap_rst_n = ap_rst_n;
  assign Module2Func_19_ap_start = Module2Func_19__ap_start;
  assign Module2Func_19_fifo_ld_0_peek_dout = from_t1_iter20_to_t1_iter21__dout;
  assign Module2Func_19_fifo_ld_0_peek_empty_n = from_t1_iter20_to_t1_iter21__empty_n;
  assign Module2Func_19_fifo_ld_0_s_dout = from_t1_iter20_to_t1_iter21__dout;
  assign Module2Func_19_fifo_ld_0_s_empty_n = from_t1_iter20_to_t1_iter21__empty_n;
  assign from_t1_iter20_to_t1_iter21__read = Module2Func_19_fifo_ld_0_s_read;
  assign from_t1_iter21_to_t1_iter22__din = Module2Func_19_fifo_st_0_din;
  assign Module2Func_19_fifo_st_0_full_n = from_t1_iter21_to_t1_iter22__full_n;
  assign from_t1_iter21_to_t1_iter22__write = Module2Func_19_fifo_st_0_write;
  assign Module2Func_20_ap_clk = ap_clk;
  assign Module2Func_20_ap_rst_n = ap_rst_n;
  assign Module2Func_20_ap_start = Module2Func_20__ap_start;
  assign Module2Func_20_fifo_ld_0_peek_dout = from_t1_iter21_to_t1_iter22__dout;
  assign Module2Func_20_fifo_ld_0_peek_empty_n = from_t1_iter21_to_t1_iter22__empty_n;
  assign Module2Func_20_fifo_ld_0_s_dout = from_t1_iter21_to_t1_iter22__dout;
  assign Module2Func_20_fifo_ld_0_s_empty_n = from_t1_iter21_to_t1_iter22__empty_n;
  assign from_t1_iter21_to_t1_iter22__read = Module2Func_20_fifo_ld_0_s_read;
  assign from_t1_iter22_to_t1_iter23__din = Module2Func_20_fifo_st_0_din;
  assign Module2Func_20_fifo_st_0_full_n = from_t1_iter22_to_t1_iter23__full_n;
  assign from_t1_iter22_to_t1_iter23__write = Module2Func_20_fifo_st_0_write;
  assign Module2Func_21_ap_clk = ap_clk;
  assign Module2Func_21_ap_rst_n = ap_rst_n;
  assign Module2Func_21_ap_start = Module2Func_21__ap_start;
  assign Module2Func_21_fifo_ld_0_peek_dout = from_t1_iter22_to_t1_iter23__dout;
  assign Module2Func_21_fifo_ld_0_peek_empty_n = from_t1_iter22_to_t1_iter23__empty_n;
  assign Module2Func_21_fifo_ld_0_s_dout = from_t1_iter22_to_t1_iter23__dout;
  assign Module2Func_21_fifo_ld_0_s_empty_n = from_t1_iter22_to_t1_iter23__empty_n;
  assign from_t1_iter22_to_t1_iter23__read = Module2Func_21_fifo_ld_0_s_read;
  assign from_t1_iter23_to_t1_iter24__din = Module2Func_21_fifo_st_0_din;
  assign Module2Func_21_fifo_st_0_full_n = from_t1_iter23_to_t1_iter24__full_n;
  assign from_t1_iter23_to_t1_iter24__write = Module2Func_21_fifo_st_0_write;
  assign Module2Func_22_ap_clk = ap_clk;
  assign Module2Func_22_ap_rst_n = ap_rst_n;
  assign Module2Func_22_ap_start = Module2Func_22__ap_start;
  assign Module2Func_22_fifo_ld_0_peek_dout = from_t1_iter23_to_t1_iter24__dout;
  assign Module2Func_22_fifo_ld_0_peek_empty_n = from_t1_iter23_to_t1_iter24__empty_n;
  assign Module2Func_22_fifo_ld_0_s_dout = from_t1_iter23_to_t1_iter24__dout;
  assign Module2Func_22_fifo_ld_0_s_empty_n = from_t1_iter23_to_t1_iter24__empty_n;
  assign from_t1_iter23_to_t1_iter24__read = Module2Func_22_fifo_ld_0_s_read;
  assign from_t1_iter24_to_t1_iter25__din = Module2Func_22_fifo_st_0_din;
  assign Module2Func_22_fifo_st_0_full_n = from_t1_iter24_to_t1_iter25__full_n;
  assign from_t1_iter24_to_t1_iter25__write = Module2Func_22_fifo_st_0_write;
  assign Module2Func_23_ap_clk = ap_clk;
  assign Module2Func_23_ap_rst_n = ap_rst_n;
  assign Module2Func_23_ap_start = Module2Func_23__ap_start;
  assign Module2Func_23_fifo_ld_0_peek_dout = from_t1_iter24_to_t1_iter25__dout;
  assign Module2Func_23_fifo_ld_0_peek_empty_n = from_t1_iter24_to_t1_iter25__empty_n;
  assign Module2Func_23_fifo_ld_0_s_dout = from_t1_iter24_to_t1_iter25__dout;
  assign Module2Func_23_fifo_ld_0_s_empty_n = from_t1_iter24_to_t1_iter25__empty_n;
  assign from_t1_iter24_to_t1_iter25__read = Module2Func_23_fifo_ld_0_s_read;
  assign from_t1_iter25_to_t1_iter26__din = Module2Func_23_fifo_st_0_din;
  assign Module2Func_23_fifo_st_0_full_n = from_t1_iter25_to_t1_iter26__full_n;
  assign from_t1_iter25_to_t1_iter26__write = Module2Func_23_fifo_st_0_write;
  assign Module2Func_24_ap_clk = ap_clk;
  assign Module2Func_24_ap_rst_n = ap_rst_n;
  assign Module2Func_24_ap_start = Module2Func_24__ap_start;
  assign Module2Func_24_fifo_ld_0_peek_dout = from_t1_iter25_to_t1_iter26__dout;
  assign Module2Func_24_fifo_ld_0_peek_empty_n = from_t1_iter25_to_t1_iter26__empty_n;
  assign Module2Func_24_fifo_ld_0_s_dout = from_t1_iter25_to_t1_iter26__dout;
  assign Module2Func_24_fifo_ld_0_s_empty_n = from_t1_iter25_to_t1_iter26__empty_n;
  assign from_t1_iter25_to_t1_iter26__read = Module2Func_24_fifo_ld_0_s_read;
  assign from_t1_iter26_to_t1_iter27__din = Module2Func_24_fifo_st_0_din;
  assign Module2Func_24_fifo_st_0_full_n = from_t1_iter26_to_t1_iter27__full_n;
  assign from_t1_iter26_to_t1_iter27__write = Module2Func_24_fifo_st_0_write;
  assign Module2Func_25_ap_clk = ap_clk;
  assign Module2Func_25_ap_rst_n = ap_rst_n;
  assign Module2Func_25_ap_start = Module2Func_25__ap_start;
  assign Module2Func_25_fifo_ld_0_peek_dout = from_t1_iter26_to_t1_iter27__dout;
  assign Module2Func_25_fifo_ld_0_peek_empty_n = from_t1_iter26_to_t1_iter27__empty_n;
  assign Module2Func_25_fifo_ld_0_s_dout = from_t1_iter26_to_t1_iter27__dout;
  assign Module2Func_25_fifo_ld_0_s_empty_n = from_t1_iter26_to_t1_iter27__empty_n;
  assign from_t1_iter26_to_t1_iter27__read = Module2Func_25_fifo_ld_0_s_read;
  assign from_t1_iter27_to_t1_iter28__din = Module2Func_25_fifo_st_0_din;
  assign Module2Func_25_fifo_st_0_full_n = from_t1_iter27_to_t1_iter28__full_n;
  assign from_t1_iter27_to_t1_iter28__write = Module2Func_25_fifo_st_0_write;
  assign Module2Func_26_ap_clk = ap_clk;
  assign Module2Func_26_ap_rst_n = ap_rst_n;
  assign Module2Func_26_ap_start = Module2Func_26__ap_start;
  assign Module2Func_26_fifo_ld_0_peek_dout = from_t1_iter27_to_t1_iter28__dout;
  assign Module2Func_26_fifo_ld_0_peek_empty_n = from_t1_iter27_to_t1_iter28__empty_n;
  assign Module2Func_26_fifo_ld_0_s_dout = from_t1_iter27_to_t1_iter28__dout;
  assign Module2Func_26_fifo_ld_0_s_empty_n = from_t1_iter27_to_t1_iter28__empty_n;
  assign from_t1_iter27_to_t1_iter28__read = Module2Func_26_fifo_ld_0_s_read;
  assign from_t1_iter28_to_t1_iter29__din = Module2Func_26_fifo_st_0_din;
  assign Module2Func_26_fifo_st_0_full_n = from_t1_iter28_to_t1_iter29__full_n;
  assign from_t1_iter28_to_t1_iter29__write = Module2Func_26_fifo_st_0_write;
  assign Module2Func_27_ap_clk = ap_clk;
  assign Module2Func_27_ap_rst_n = ap_rst_n;
  assign Module2Func_27_ap_start = Module2Func_27__ap_start;
  assign Module2Func_27_fifo_ld_0_peek_dout = from_t1_iter28_to_t1_iter29__dout;
  assign Module2Func_27_fifo_ld_0_peek_empty_n = from_t1_iter28_to_t1_iter29__empty_n;
  assign Module2Func_27_fifo_ld_0_s_dout = from_t1_iter28_to_t1_iter29__dout;
  assign Module2Func_27_fifo_ld_0_s_empty_n = from_t1_iter28_to_t1_iter29__empty_n;
  assign from_t1_iter28_to_t1_iter29__read = Module2Func_27_fifo_ld_0_s_read;
  assign from_t1_iter29_to_t1_iter30__din = Module2Func_27_fifo_st_0_din;
  assign Module2Func_27_fifo_st_0_full_n = from_t1_iter29_to_t1_iter30__full_n;
  assign from_t1_iter29_to_t1_iter30__write = Module2Func_27_fifo_st_0_write;
  assign Module2Func_28_ap_clk = ap_clk;
  assign Module2Func_28_ap_rst_n = ap_rst_n;
  assign Module2Func_28_ap_start = Module2Func_28__ap_start;
  assign Module2Func_28_fifo_ld_0_peek_dout = from_t1_iter29_to_t1_iter30__dout;
  assign Module2Func_28_fifo_ld_0_peek_empty_n = from_t1_iter29_to_t1_iter30__empty_n;
  assign Module2Func_28_fifo_ld_0_s_dout = from_t1_iter29_to_t1_iter30__dout;
  assign Module2Func_28_fifo_ld_0_s_empty_n = from_t1_iter29_to_t1_iter30__empty_n;
  assign from_t1_iter29_to_t1_iter30__read = Module2Func_28_fifo_ld_0_s_read;
  assign from_t1_iter30_to_t1_iter31__din = Module2Func_28_fifo_st_0_din;
  assign Module2Func_28_fifo_st_0_full_n = from_t1_iter30_to_t1_iter31__full_n;
  assign from_t1_iter30_to_t1_iter31__write = Module2Func_28_fifo_st_0_write;
  assign Module2Func_29_ap_clk = ap_clk;
  assign Module2Func_29_ap_rst_n = ap_rst_n;
  assign Module2Func_29_ap_start = Module2Func_29__ap_start;
  assign Module2Func_29_fifo_ld_0_peek_dout = from_t1_iter30_to_t1_iter31__dout;
  assign Module2Func_29_fifo_ld_0_peek_empty_n = from_t1_iter30_to_t1_iter31__empty_n;
  assign Module2Func_29_fifo_ld_0_s_dout = from_t1_iter30_to_t1_iter31__dout;
  assign Module2Func_29_fifo_ld_0_s_empty_n = from_t1_iter30_to_t1_iter31__empty_n;
  assign from_t1_iter30_to_t1_iter31__read = Module2Func_29_fifo_ld_0_s_read;
  assign from_t1_iter31_to_t1_iter32__din = Module2Func_29_fifo_st_0_din;
  assign Module2Func_29_fifo_st_0_full_n = from_t1_iter31_to_t1_iter32__full_n;
  assign from_t1_iter31_to_t1_iter32__write = Module2Func_29_fifo_st_0_write;
  assign Module2Func_30_ap_clk = ap_clk;
  assign Module2Func_30_ap_rst_n = ap_rst_n;
  assign Module2Func_30_ap_start = Module2Func_30__ap_start;
  assign Module2Func_30_fifo_ld_0_peek_dout = from_t1_iter31_to_t1_iter32__dout;
  assign Module2Func_30_fifo_ld_0_peek_empty_n = from_t1_iter31_to_t1_iter32__empty_n;
  assign Module2Func_30_fifo_ld_0_s_dout = from_t1_iter31_to_t1_iter32__dout;
  assign Module2Func_30_fifo_ld_0_s_empty_n = from_t1_iter31_to_t1_iter32__empty_n;
  assign from_t1_iter31_to_t1_iter32__read = Module2Func_30_fifo_ld_0_s_read;
  assign from_t1_iter32_to_t1_iter33__din = Module2Func_30_fifo_st_0_din;
  assign Module2Func_30_fifo_st_0_full_n = from_t1_iter32_to_t1_iter33__full_n;
  assign from_t1_iter32_to_t1_iter33__write = Module2Func_30_fifo_st_0_write;
  assign Module2Func_31_ap_clk = ap_clk;
  assign Module2Func_31_ap_rst_n = ap_rst_n;
  assign Module2Func_31_ap_start = Module2Func_31__ap_start;
  assign Module2Func_31_fifo_ld_0_peek_dout = from_t1_iter32_to_t1_iter33__dout;
  assign Module2Func_31_fifo_ld_0_peek_empty_n = from_t1_iter32_to_t1_iter33__empty_n;
  assign Module2Func_31_fifo_ld_0_s_dout = from_t1_iter32_to_t1_iter33__dout;
  assign Module2Func_31_fifo_ld_0_s_empty_n = from_t1_iter32_to_t1_iter33__empty_n;
  assign from_t1_iter32_to_t1_iter33__read = Module2Func_31_fifo_ld_0_s_read;
  assign from_t1_iter33_to_t1_iter34__din = Module2Func_31_fifo_st_0_din;
  assign Module2Func_31_fifo_st_0_full_n = from_t1_iter33_to_t1_iter34__full_n;
  assign from_t1_iter33_to_t1_iter34__write = Module2Func_31_fifo_st_0_write;
  assign Module2Func_32_ap_clk = ap_clk;
  assign Module2Func_32_ap_rst_n = ap_rst_n;
  assign Module2Func_32_ap_start = Module2Func_32__ap_start;
  assign Module2Func_32_fifo_ld_0_peek_dout = from_t1_iter33_to_t1_iter34__dout;
  assign Module2Func_32_fifo_ld_0_peek_empty_n = from_t1_iter33_to_t1_iter34__empty_n;
  assign Module2Func_32_fifo_ld_0_s_dout = from_t1_iter33_to_t1_iter34__dout;
  assign Module2Func_32_fifo_ld_0_s_empty_n = from_t1_iter33_to_t1_iter34__empty_n;
  assign from_t1_iter33_to_t1_iter34__read = Module2Func_32_fifo_ld_0_s_read;
  assign from_t1_iter34_to_t1_iter35__din = Module2Func_32_fifo_st_0_din;
  assign Module2Func_32_fifo_st_0_full_n = from_t1_iter34_to_t1_iter35__full_n;
  assign from_t1_iter34_to_t1_iter35__write = Module2Func_32_fifo_st_0_write;
  assign Module2Func_33_ap_clk = ap_clk;
  assign Module2Func_33_ap_rst_n = ap_rst_n;
  assign Module2Func_33_ap_start = Module2Func_33__ap_start;
  assign Module2Func_33_fifo_ld_0_peek_dout = from_t1_iter34_to_t1_iter35__dout;
  assign Module2Func_33_fifo_ld_0_peek_empty_n = from_t1_iter34_to_t1_iter35__empty_n;
  assign Module2Func_33_fifo_ld_0_s_dout = from_t1_iter34_to_t1_iter35__dout;
  assign Module2Func_33_fifo_ld_0_s_empty_n = from_t1_iter34_to_t1_iter35__empty_n;
  assign from_t1_iter34_to_t1_iter35__read = Module2Func_33_fifo_ld_0_s_read;
  assign from_t1_iter35_to_t1_iter36__din = Module2Func_33_fifo_st_0_din;
  assign Module2Func_33_fifo_st_0_full_n = from_t1_iter35_to_t1_iter36__full_n;
  assign from_t1_iter35_to_t1_iter36__write = Module2Func_33_fifo_st_0_write;
  assign Module2Func_34_ap_clk = ap_clk;
  assign Module2Func_34_ap_rst_n = ap_rst_n;
  assign Module2Func_34_ap_start = Module2Func_34__ap_start;
  assign Module2Func_34_fifo_ld_0_peek_dout = from_t1_iter35_to_t1_iter36__dout;
  assign Module2Func_34_fifo_ld_0_peek_empty_n = from_t1_iter35_to_t1_iter36__empty_n;
  assign Module2Func_34_fifo_ld_0_s_dout = from_t1_iter35_to_t1_iter36__dout;
  assign Module2Func_34_fifo_ld_0_s_empty_n = from_t1_iter35_to_t1_iter36__empty_n;
  assign from_t1_iter35_to_t1_iter36__read = Module2Func_34_fifo_ld_0_s_read;
  assign from_t1_iter36_to_t1_iter37__din = Module2Func_34_fifo_st_0_din;
  assign Module2Func_34_fifo_st_0_full_n = from_t1_iter36_to_t1_iter37__full_n;
  assign from_t1_iter36_to_t1_iter37__write = Module2Func_34_fifo_st_0_write;
  assign Module2Func_35_ap_clk = ap_clk;
  assign Module2Func_35_ap_rst_n = ap_rst_n;
  assign Module2Func_35_ap_start = Module2Func_35__ap_start;
  assign Module2Func_35_fifo_ld_0_peek_dout = from_t1_iter36_to_t1_iter37__dout;
  assign Module2Func_35_fifo_ld_0_peek_empty_n = from_t1_iter36_to_t1_iter37__empty_n;
  assign Module2Func_35_fifo_ld_0_s_dout = from_t1_iter36_to_t1_iter37__dout;
  assign Module2Func_35_fifo_ld_0_s_empty_n = from_t1_iter36_to_t1_iter37__empty_n;
  assign from_t1_iter36_to_t1_iter37__read = Module2Func_35_fifo_ld_0_s_read;
  assign from_t1_iter37_to_t1_iter38__din = Module2Func_35_fifo_st_0_din;
  assign Module2Func_35_fifo_st_0_full_n = from_t1_iter37_to_t1_iter38__full_n;
  assign from_t1_iter37_to_t1_iter38__write = Module2Func_35_fifo_st_0_write;
  assign Module2Func_36_ap_clk = ap_clk;
  assign Module2Func_36_ap_rst_n = ap_rst_n;
  assign Module2Func_36_ap_start = Module2Func_36__ap_start;
  assign Module2Func_36_fifo_ld_0_peek_dout = from_t1_iter37_to_t1_iter38__dout;
  assign Module2Func_36_fifo_ld_0_peek_empty_n = from_t1_iter37_to_t1_iter38__empty_n;
  assign Module2Func_36_fifo_ld_0_s_dout = from_t1_iter37_to_t1_iter38__dout;
  assign Module2Func_36_fifo_ld_0_s_empty_n = from_t1_iter37_to_t1_iter38__empty_n;
  assign from_t1_iter37_to_t1_iter38__read = Module2Func_36_fifo_ld_0_s_read;
  assign from_t1_iter38_to_t1_iter39__din = Module2Func_36_fifo_st_0_din;
  assign Module2Func_36_fifo_st_0_full_n = from_t1_iter38_to_t1_iter39__full_n;
  assign from_t1_iter38_to_t1_iter39__write = Module2Func_36_fifo_st_0_write;
  assign Module2Func_37_ap_clk = ap_clk;
  assign Module2Func_37_ap_rst_n = ap_rst_n;
  assign Module2Func_37_ap_start = Module2Func_37__ap_start;
  assign Module2Func_37_fifo_ld_0_peek_dout = from_t1_iter38_to_t1_iter39__dout;
  assign Module2Func_37_fifo_ld_0_peek_empty_n = from_t1_iter38_to_t1_iter39__empty_n;
  assign Module2Func_37_fifo_ld_0_s_dout = from_t1_iter38_to_t1_iter39__dout;
  assign Module2Func_37_fifo_ld_0_s_empty_n = from_t1_iter38_to_t1_iter39__empty_n;
  assign from_t1_iter38_to_t1_iter39__read = Module2Func_37_fifo_ld_0_s_read;
  assign from_t1_iter39_to_t1_iter40__din = Module2Func_37_fifo_st_0_din;
  assign Module2Func_37_fifo_st_0_full_n = from_t1_iter39_to_t1_iter40__full_n;
  assign from_t1_iter39_to_t1_iter40__write = Module2Func_37_fifo_st_0_write;
  assign Module2Func_38_ap_clk = ap_clk;
  assign Module2Func_38_ap_rst_n = ap_rst_n;
  assign Module2Func_38_ap_start = Module2Func_38__ap_start;
  assign Module2Func_38_fifo_ld_0_peek_dout = from_t1_iter39_to_t1_iter40__dout;
  assign Module2Func_38_fifo_ld_0_peek_empty_n = from_t1_iter39_to_t1_iter40__empty_n;
  assign Module2Func_38_fifo_ld_0_s_dout = from_t1_iter39_to_t1_iter40__dout;
  assign Module2Func_38_fifo_ld_0_s_empty_n = from_t1_iter39_to_t1_iter40__empty_n;
  assign from_t1_iter39_to_t1_iter40__read = Module2Func_38_fifo_ld_0_s_read;
  assign from_t1_iter40_to_t1_iter41__din = Module2Func_38_fifo_st_0_din;
  assign Module2Func_38_fifo_st_0_full_n = from_t1_iter40_to_t1_iter41__full_n;
  assign from_t1_iter40_to_t1_iter41__write = Module2Func_38_fifo_st_0_write;
  assign Module2Func_39_ap_clk = ap_clk;
  assign Module2Func_39_ap_rst_n = ap_rst_n;
  assign Module2Func_39_ap_start = Module2Func_39__ap_start;
  assign Module2Func_39_fifo_ld_0_peek_dout = from_t1_iter40_to_t1_iter41__dout;
  assign Module2Func_39_fifo_ld_0_peek_empty_n = from_t1_iter40_to_t1_iter41__empty_n;
  assign Module2Func_39_fifo_ld_0_s_dout = from_t1_iter40_to_t1_iter41__dout;
  assign Module2Func_39_fifo_ld_0_s_empty_n = from_t1_iter40_to_t1_iter41__empty_n;
  assign from_t1_iter40_to_t1_iter41__read = Module2Func_39_fifo_ld_0_s_read;
  assign from_t1_iter41_to_t1_iter42__din = Module2Func_39_fifo_st_0_din;
  assign Module2Func_39_fifo_st_0_full_n = from_t1_iter41_to_t1_iter42__full_n;
  assign from_t1_iter41_to_t1_iter42__write = Module2Func_39_fifo_st_0_write;
  assign Module2Func_40_ap_clk = ap_clk;
  assign Module2Func_40_ap_rst_n = ap_rst_n;
  assign Module2Func_40_ap_start = Module2Func_40__ap_start;
  assign Module2Func_40_fifo_ld_0_peek_dout = from_t1_iter41_to_t1_iter42__dout;
  assign Module2Func_40_fifo_ld_0_peek_empty_n = from_t1_iter41_to_t1_iter42__empty_n;
  assign Module2Func_40_fifo_ld_0_s_dout = from_t1_iter41_to_t1_iter42__dout;
  assign Module2Func_40_fifo_ld_0_s_empty_n = from_t1_iter41_to_t1_iter42__empty_n;
  assign from_t1_iter41_to_t1_iter42__read = Module2Func_40_fifo_ld_0_s_read;
  assign from_t1_iter42_to_t1_iter43__din = Module2Func_40_fifo_st_0_din;
  assign Module2Func_40_fifo_st_0_full_n = from_t1_iter42_to_t1_iter43__full_n;
  assign from_t1_iter42_to_t1_iter43__write = Module2Func_40_fifo_st_0_write;
  assign Module2Func_41_ap_clk = ap_clk;
  assign Module2Func_41_ap_rst_n = ap_rst_n;
  assign Module2Func_41_ap_start = Module2Func_41__ap_start;
  assign Module2Func_41_fifo_ld_0_peek_dout = from_t1_iter42_to_t1_iter43__dout;
  assign Module2Func_41_fifo_ld_0_peek_empty_n = from_t1_iter42_to_t1_iter43__empty_n;
  assign Module2Func_41_fifo_ld_0_s_dout = from_t1_iter42_to_t1_iter43__dout;
  assign Module2Func_41_fifo_ld_0_s_empty_n = from_t1_iter42_to_t1_iter43__empty_n;
  assign from_t1_iter42_to_t1_iter43__read = Module2Func_41_fifo_ld_0_s_read;
  assign from_t1_iter43_to_t1_iter44__din = Module2Func_41_fifo_st_0_din;
  assign Module2Func_41_fifo_st_0_full_n = from_t1_iter43_to_t1_iter44__full_n;
  assign from_t1_iter43_to_t1_iter44__write = Module2Func_41_fifo_st_0_write;
  assign Module2Func_42_ap_clk = ap_clk;
  assign Module2Func_42_ap_rst_n = ap_rst_n;
  assign Module2Func_42_ap_start = Module2Func_42__ap_start;
  assign Module2Func_42_fifo_ld_0_peek_dout = from_t1_iter43_to_t1_iter44__dout;
  assign Module2Func_42_fifo_ld_0_peek_empty_n = from_t1_iter43_to_t1_iter44__empty_n;
  assign Module2Func_42_fifo_ld_0_s_dout = from_t1_iter43_to_t1_iter44__dout;
  assign Module2Func_42_fifo_ld_0_s_empty_n = from_t1_iter43_to_t1_iter44__empty_n;
  assign from_t1_iter43_to_t1_iter44__read = Module2Func_42_fifo_ld_0_s_read;
  assign from_t1_iter44_to_t1_iter45__din = Module2Func_42_fifo_st_0_din;
  assign Module2Func_42_fifo_st_0_full_n = from_t1_iter44_to_t1_iter45__full_n;
  assign from_t1_iter44_to_t1_iter45__write = Module2Func_42_fifo_st_0_write;
  assign Module2Func_43_ap_clk = ap_clk;
  assign Module2Func_43_ap_rst_n = ap_rst_n;
  assign Module2Func_43_ap_start = Module2Func_43__ap_start;
  assign Module2Func_43_fifo_ld_0_peek_dout = from_t1_iter44_to_t1_iter45__dout;
  assign Module2Func_43_fifo_ld_0_peek_empty_n = from_t1_iter44_to_t1_iter45__empty_n;
  assign Module2Func_43_fifo_ld_0_s_dout = from_t1_iter44_to_t1_iter45__dout;
  assign Module2Func_43_fifo_ld_0_s_empty_n = from_t1_iter44_to_t1_iter45__empty_n;
  assign from_t1_iter44_to_t1_iter45__read = Module2Func_43_fifo_ld_0_s_read;
  assign from_t1_iter45_to_t1_iter46__din = Module2Func_43_fifo_st_0_din;
  assign Module2Func_43_fifo_st_0_full_n = from_t1_iter45_to_t1_iter46__full_n;
  assign from_t1_iter45_to_t1_iter46__write = Module2Func_43_fifo_st_0_write;
  assign Module2Func_44_ap_clk = ap_clk;
  assign Module2Func_44_ap_rst_n = ap_rst_n;
  assign Module2Func_44_ap_start = Module2Func_44__ap_start;
  assign Module2Func_44_fifo_ld_0_peek_dout = from_t1_iter45_to_t1_iter46__dout;
  assign Module2Func_44_fifo_ld_0_peek_empty_n = from_t1_iter45_to_t1_iter46__empty_n;
  assign Module2Func_44_fifo_ld_0_s_dout = from_t1_iter45_to_t1_iter46__dout;
  assign Module2Func_44_fifo_ld_0_s_empty_n = from_t1_iter45_to_t1_iter46__empty_n;
  assign from_t1_iter45_to_t1_iter46__read = Module2Func_44_fifo_ld_0_s_read;
  assign from_t1_iter46_to_t1_iter47__din = Module2Func_44_fifo_st_0_din;
  assign Module2Func_44_fifo_st_0_full_n = from_t1_iter46_to_t1_iter47__full_n;
  assign from_t1_iter46_to_t1_iter47__write = Module2Func_44_fifo_st_0_write;
  assign Module2Func_45_ap_clk = ap_clk;
  assign Module2Func_45_ap_rst_n = ap_rst_n;
  assign Module2Func_45_ap_start = Module2Func_45__ap_start;
  assign Module2Func_45_fifo_ld_0_peek_dout = from_t1_iter46_to_t1_iter47__dout;
  assign Module2Func_45_fifo_ld_0_peek_empty_n = from_t1_iter46_to_t1_iter47__empty_n;
  assign Module2Func_45_fifo_ld_0_s_dout = from_t1_iter46_to_t1_iter47__dout;
  assign Module2Func_45_fifo_ld_0_s_empty_n = from_t1_iter46_to_t1_iter47__empty_n;
  assign from_t1_iter46_to_t1_iter47__read = Module2Func_45_fifo_ld_0_s_read;
  assign from_t1_iter47_to_t1_iter48__din = Module2Func_45_fifo_st_0_din;
  assign Module2Func_45_fifo_st_0_full_n = from_t1_iter47_to_t1_iter48__full_n;
  assign from_t1_iter47_to_t1_iter48__write = Module2Func_45_fifo_st_0_write;
  assign Module2Func_46_ap_clk = ap_clk;
  assign Module2Func_46_ap_rst_n = ap_rst_n;
  assign Module2Func_46_ap_start = Module2Func_46__ap_start;
  assign Module2Func_46_fifo_ld_0_peek_dout = from_t1_iter47_to_t1_iter48__dout;
  assign Module2Func_46_fifo_ld_0_peek_empty_n = from_t1_iter47_to_t1_iter48__empty_n;
  assign Module2Func_46_fifo_ld_0_s_dout = from_t1_iter47_to_t1_iter48__dout;
  assign Module2Func_46_fifo_ld_0_s_empty_n = from_t1_iter47_to_t1_iter48__empty_n;
  assign from_t1_iter47_to_t1_iter48__read = Module2Func_46_fifo_ld_0_s_read;
  assign from_t1_iter48_to_t1_iter49__din = Module2Func_46_fifo_st_0_din;
  assign Module2Func_46_fifo_st_0_full_n = from_t1_iter48_to_t1_iter49__full_n;
  assign from_t1_iter48_to_t1_iter49__write = Module2Func_46_fifo_st_0_write;
  assign Module2Func_47_ap_clk = ap_clk;
  assign Module2Func_47_ap_rst_n = ap_rst_n;
  assign Module2Func_47_ap_start = Module2Func_47__ap_start;
  assign Module2Func_47_fifo_ld_0_peek_dout = from_t1_iter48_to_t1_iter49__dout;
  assign Module2Func_47_fifo_ld_0_peek_empty_n = from_t1_iter48_to_t1_iter49__empty_n;
  assign Module2Func_47_fifo_ld_0_s_dout = from_t1_iter48_to_t1_iter49__dout;
  assign Module2Func_47_fifo_ld_0_s_empty_n = from_t1_iter48_to_t1_iter49__empty_n;
  assign from_t1_iter48_to_t1_iter49__read = Module2Func_47_fifo_ld_0_s_read;
  assign from_t1_iter49_to_t1_iter50__din = Module2Func_47_fifo_st_0_din;
  assign Module2Func_47_fifo_st_0_full_n = from_t1_iter49_to_t1_iter50__full_n;
  assign from_t1_iter49_to_t1_iter50__write = Module2Func_47_fifo_st_0_write;
  assign Module2Func_48_ap_clk = ap_clk;
  assign Module2Func_48_ap_rst_n = ap_rst_n;
  assign Module2Func_48_ap_start = Module2Func_48__ap_start;
  assign Module2Func_48_fifo_ld_0_peek_dout = from_t1_iter49_to_t1_iter50__dout;
  assign Module2Func_48_fifo_ld_0_peek_empty_n = from_t1_iter49_to_t1_iter50__empty_n;
  assign Module2Func_48_fifo_ld_0_s_dout = from_t1_iter49_to_t1_iter50__dout;
  assign Module2Func_48_fifo_ld_0_s_empty_n = from_t1_iter49_to_t1_iter50__empty_n;
  assign from_t1_iter49_to_t1_iter50__read = Module2Func_48_fifo_ld_0_s_read;
  assign from_t1_iter50_to_t1_iter51__din = Module2Func_48_fifo_st_0_din;
  assign Module2Func_48_fifo_st_0_full_n = from_t1_iter50_to_t1_iter51__full_n;
  assign from_t1_iter50_to_t1_iter51__write = Module2Func_48_fifo_st_0_write;
  assign Module2Func_49_ap_clk = ap_clk;
  assign Module2Func_49_ap_rst_n = ap_rst_n;
  assign Module2Func_49_ap_start = Module2Func_49__ap_start;
  assign Module2Func_49_fifo_ld_0_peek_dout = from_t1_iter50_to_t1_iter51__dout;
  assign Module2Func_49_fifo_ld_0_peek_empty_n = from_t1_iter50_to_t1_iter51__empty_n;
  assign Module2Func_49_fifo_ld_0_s_dout = from_t1_iter50_to_t1_iter51__dout;
  assign Module2Func_49_fifo_ld_0_s_empty_n = from_t1_iter50_to_t1_iter51__empty_n;
  assign from_t1_iter50_to_t1_iter51__read = Module2Func_49_fifo_ld_0_s_read;
  assign from_t1_iter51_to_t1_iter52__din = Module2Func_49_fifo_st_0_din;
  assign Module2Func_49_fifo_st_0_full_n = from_t1_iter51_to_t1_iter52__full_n;
  assign from_t1_iter51_to_t1_iter52__write = Module2Func_49_fifo_st_0_write;
  assign Module2Func_50_ap_clk = ap_clk;
  assign Module2Func_50_ap_rst_n = ap_rst_n;
  assign Module2Func_50_ap_start = Module2Func_50__ap_start;
  assign Module2Func_50_fifo_ld_0_peek_dout = from_t1_iter51_to_t1_iter52__dout;
  assign Module2Func_50_fifo_ld_0_peek_empty_n = from_t1_iter51_to_t1_iter52__empty_n;
  assign Module2Func_50_fifo_ld_0_s_dout = from_t1_iter51_to_t1_iter52__dout;
  assign Module2Func_50_fifo_ld_0_s_empty_n = from_t1_iter51_to_t1_iter52__empty_n;
  assign from_t1_iter51_to_t1_iter52__read = Module2Func_50_fifo_ld_0_s_read;
  assign from_t1_iter52_to_t1_iter53__din = Module2Func_50_fifo_st_0_din;
  assign Module2Func_50_fifo_st_0_full_n = from_t1_iter52_to_t1_iter53__full_n;
  assign from_t1_iter52_to_t1_iter53__write = Module2Func_50_fifo_st_0_write;
  assign Module2Func_51_ap_clk = ap_clk;
  assign Module2Func_51_ap_rst_n = ap_rst_n;
  assign Module2Func_51_ap_start = Module2Func_51__ap_start;
  assign Module2Func_51_fifo_ld_0_peek_dout = from_t1_iter52_to_t1_iter53__dout;
  assign Module2Func_51_fifo_ld_0_peek_empty_n = from_t1_iter52_to_t1_iter53__empty_n;
  assign Module2Func_51_fifo_ld_0_s_dout = from_t1_iter52_to_t1_iter53__dout;
  assign Module2Func_51_fifo_ld_0_s_empty_n = from_t1_iter52_to_t1_iter53__empty_n;
  assign from_t1_iter52_to_t1_iter53__read = Module2Func_51_fifo_ld_0_s_read;
  assign from_t1_iter53_to_t1_iter54__din = Module2Func_51_fifo_st_0_din;
  assign Module2Func_51_fifo_st_0_full_n = from_t1_iter53_to_t1_iter54__full_n;
  assign from_t1_iter53_to_t1_iter54__write = Module2Func_51_fifo_st_0_write;
  assign Module2Func_52_ap_clk = ap_clk;
  assign Module2Func_52_ap_rst_n = ap_rst_n;
  assign Module2Func_52_ap_start = Module2Func_52__ap_start;
  assign Module2Func_52_fifo_ld_0_peek_dout = from_t1_iter53_to_t1_iter54__dout;
  assign Module2Func_52_fifo_ld_0_peek_empty_n = from_t1_iter53_to_t1_iter54__empty_n;
  assign Module2Func_52_fifo_ld_0_s_dout = from_t1_iter53_to_t1_iter54__dout;
  assign Module2Func_52_fifo_ld_0_s_empty_n = from_t1_iter53_to_t1_iter54__empty_n;
  assign from_t1_iter53_to_t1_iter54__read = Module2Func_52_fifo_ld_0_s_read;
  assign from_t1_iter54_to_t1_iter55__din = Module2Func_52_fifo_st_0_din;
  assign Module2Func_52_fifo_st_0_full_n = from_t1_iter54_to_t1_iter55__full_n;
  assign from_t1_iter54_to_t1_iter55__write = Module2Func_52_fifo_st_0_write;
  assign Module2Func_53_ap_clk = ap_clk;
  assign Module2Func_53_ap_rst_n = ap_rst_n;
  assign Module2Func_53_ap_start = Module2Func_53__ap_start;
  assign Module2Func_53_fifo_ld_0_peek_dout = from_t1_iter54_to_t1_iter55__dout;
  assign Module2Func_53_fifo_ld_0_peek_empty_n = from_t1_iter54_to_t1_iter55__empty_n;
  assign Module2Func_53_fifo_ld_0_s_dout = from_t1_iter54_to_t1_iter55__dout;
  assign Module2Func_53_fifo_ld_0_s_empty_n = from_t1_iter54_to_t1_iter55__empty_n;
  assign from_t1_iter54_to_t1_iter55__read = Module2Func_53_fifo_ld_0_s_read;
  assign from_t1_iter55_to_t1_iter56__din = Module2Func_53_fifo_st_0_din;
  assign Module2Func_53_fifo_st_0_full_n = from_t1_iter55_to_t1_iter56__full_n;
  assign from_t1_iter55_to_t1_iter56__write = Module2Func_53_fifo_st_0_write;
  assign Module2Func_54_ap_clk = ap_clk;
  assign Module2Func_54_ap_rst_n = ap_rst_n;
  assign Module2Func_54_ap_start = Module2Func_54__ap_start;
  assign Module2Func_54_fifo_ld_0_peek_dout = from_t1_iter55_to_t1_iter56__dout;
  assign Module2Func_54_fifo_ld_0_peek_empty_n = from_t1_iter55_to_t1_iter56__empty_n;
  assign Module2Func_54_fifo_ld_0_s_dout = from_t1_iter55_to_t1_iter56__dout;
  assign Module2Func_54_fifo_ld_0_s_empty_n = from_t1_iter55_to_t1_iter56__empty_n;
  assign from_t1_iter55_to_t1_iter56__read = Module2Func_54_fifo_ld_0_s_read;
  assign from_t1_iter56_to_t1_iter57__din = Module2Func_54_fifo_st_0_din;
  assign Module2Func_54_fifo_st_0_full_n = from_t1_iter56_to_t1_iter57__full_n;
  assign from_t1_iter56_to_t1_iter57__write = Module2Func_54_fifo_st_0_write;
  assign Module2Func_55_ap_clk = ap_clk;
  assign Module2Func_55_ap_rst_n = ap_rst_n;
  assign Module2Func_55_ap_start = Module2Func_55__ap_start;
  assign Module2Func_55_fifo_ld_0_peek_dout = from_t1_iter56_to_t1_iter57__dout;
  assign Module2Func_55_fifo_ld_0_peek_empty_n = from_t1_iter56_to_t1_iter57__empty_n;
  assign Module2Func_55_fifo_ld_0_s_dout = from_t1_iter56_to_t1_iter57__dout;
  assign Module2Func_55_fifo_ld_0_s_empty_n = from_t1_iter56_to_t1_iter57__empty_n;
  assign from_t1_iter56_to_t1_iter57__read = Module2Func_55_fifo_ld_0_s_read;
  assign from_t1_iter57_to_t1_iter58__din = Module2Func_55_fifo_st_0_din;
  assign Module2Func_55_fifo_st_0_full_n = from_t1_iter57_to_t1_iter58__full_n;
  assign from_t1_iter57_to_t1_iter58__write = Module2Func_55_fifo_st_0_write;
  assign Module2Func_56_ap_clk = ap_clk;
  assign Module2Func_56_ap_rst_n = ap_rst_n;
  assign Module2Func_56_ap_start = Module2Func_56__ap_start;
  assign Module2Func_56_fifo_ld_0_peek_dout = from_t1_iter57_to_t1_iter58__dout;
  assign Module2Func_56_fifo_ld_0_peek_empty_n = from_t1_iter57_to_t1_iter58__empty_n;
  assign Module2Func_56_fifo_ld_0_s_dout = from_t1_iter57_to_t1_iter58__dout;
  assign Module2Func_56_fifo_ld_0_s_empty_n = from_t1_iter57_to_t1_iter58__empty_n;
  assign from_t1_iter57_to_t1_iter58__read = Module2Func_56_fifo_ld_0_s_read;
  assign from_t1_iter58_to_t1_iter59__din = Module2Func_56_fifo_st_0_din;
  assign Module2Func_56_fifo_st_0_full_n = from_t1_iter58_to_t1_iter59__full_n;
  assign from_t1_iter58_to_t1_iter59__write = Module2Func_56_fifo_st_0_write;
  assign Module2Func_57_ap_clk = ap_clk;
  assign Module2Func_57_ap_rst_n = ap_rst_n;
  assign Module2Func_57_ap_start = Module2Func_57__ap_start;
  assign Module2Func_57_fifo_ld_0_peek_dout = from_t1_iter58_to_t1_iter59__dout;
  assign Module2Func_57_fifo_ld_0_peek_empty_n = from_t1_iter58_to_t1_iter59__empty_n;
  assign Module2Func_57_fifo_ld_0_s_dout = from_t1_iter58_to_t1_iter59__dout;
  assign Module2Func_57_fifo_ld_0_s_empty_n = from_t1_iter58_to_t1_iter59__empty_n;
  assign from_t1_iter58_to_t1_iter59__read = Module2Func_57_fifo_ld_0_s_read;
  assign from_t1_iter59_to_t1_iter60__din = Module2Func_57_fifo_st_0_din;
  assign Module2Func_57_fifo_st_0_full_n = from_t1_iter59_to_t1_iter60__full_n;
  assign from_t1_iter59_to_t1_iter60__write = Module2Func_57_fifo_st_0_write;
  assign Module2Func_58_ap_clk = ap_clk;
  assign Module2Func_58_ap_rst_n = ap_rst_n;
  assign Module2Func_58_ap_start = Module2Func_58__ap_start;
  assign Module2Func_58_fifo_ld_0_peek_dout = from_t1_iter59_to_t1_iter60__dout;
  assign Module2Func_58_fifo_ld_0_peek_empty_n = from_t1_iter59_to_t1_iter60__empty_n;
  assign Module2Func_58_fifo_ld_0_s_dout = from_t1_iter59_to_t1_iter60__dout;
  assign Module2Func_58_fifo_ld_0_s_empty_n = from_t1_iter59_to_t1_iter60__empty_n;
  assign from_t1_iter59_to_t1_iter60__read = Module2Func_58_fifo_ld_0_s_read;
  assign from_t1_iter60_to_t1_iter61__din = Module2Func_58_fifo_st_0_din;
  assign Module2Func_58_fifo_st_0_full_n = from_t1_iter60_to_t1_iter61__full_n;
  assign from_t1_iter60_to_t1_iter61__write = Module2Func_58_fifo_st_0_write;
  assign Module2Func_59_ap_clk = ap_clk;
  assign Module2Func_59_ap_rst_n = ap_rst_n;
  assign Module2Func_59_ap_start = Module2Func_59__ap_start;
  assign Module2Func_59_fifo_ld_0_peek_dout = from_t1_iter60_to_t1_iter61__dout;
  assign Module2Func_59_fifo_ld_0_peek_empty_n = from_t1_iter60_to_t1_iter61__empty_n;
  assign Module2Func_59_fifo_ld_0_s_dout = from_t1_iter60_to_t1_iter61__dout;
  assign Module2Func_59_fifo_ld_0_s_empty_n = from_t1_iter60_to_t1_iter61__empty_n;
  assign from_t1_iter60_to_t1_iter61__read = Module2Func_59_fifo_ld_0_s_read;
  assign from_t1_iter61_to_t1_iter62__din = Module2Func_59_fifo_st_0_din;
  assign Module2Func_59_fifo_st_0_full_n = from_t1_iter61_to_t1_iter62__full_n;
  assign from_t1_iter61_to_t1_iter62__write = Module2Func_59_fifo_st_0_write;
  assign Module2Func_60_ap_clk = ap_clk;
  assign Module2Func_60_ap_rst_n = ap_rst_n;
  assign Module2Func_60_ap_start = Module2Func_60__ap_start;
  assign Module2Func_60_fifo_ld_0_peek_dout = from_t1_iter61_to_t1_iter62__dout;
  assign Module2Func_60_fifo_ld_0_peek_empty_n = from_t1_iter61_to_t1_iter62__empty_n;
  assign Module2Func_60_fifo_ld_0_s_dout = from_t1_iter61_to_t1_iter62__dout;
  assign Module2Func_60_fifo_ld_0_s_empty_n = from_t1_iter61_to_t1_iter62__empty_n;
  assign from_t1_iter61_to_t1_iter62__read = Module2Func_60_fifo_ld_0_s_read;
  assign from_t1_iter62_to_t1_iter63__din = Module2Func_60_fifo_st_0_din;
  assign Module2Func_60_fifo_st_0_full_n = from_t1_iter62_to_t1_iter63__full_n;
  assign from_t1_iter62_to_t1_iter63__write = Module2Func_60_fifo_st_0_write;
  assign Module2Func_61_ap_clk = ap_clk;
  assign Module2Func_61_ap_rst_n = ap_rst_n;
  assign Module2Func_61_ap_start = Module2Func_61__ap_start;
  assign Module2Func_61_fifo_ld_0_peek_dout = from_t1_iter62_to_t1_iter63__dout;
  assign Module2Func_61_fifo_ld_0_peek_empty_n = from_t1_iter62_to_t1_iter63__empty_n;
  assign Module2Func_61_fifo_ld_0_s_dout = from_t1_iter62_to_t1_iter63__dout;
  assign Module2Func_61_fifo_ld_0_s_empty_n = from_t1_iter62_to_t1_iter63__empty_n;
  assign from_t1_iter62_to_t1_iter63__read = Module2Func_61_fifo_ld_0_s_read;
  assign from_t1_iter63_to_t1_iter64__din = Module2Func_61_fifo_st_0_din;
  assign Module2Func_61_fifo_st_0_full_n = from_t1_iter63_to_t1_iter64__full_n;
  assign from_t1_iter63_to_t1_iter64__write = Module2Func_61_fifo_st_0_write;
  assign Module2Func_62_ap_clk = ap_clk;
  assign Module2Func_62_ap_rst_n = ap_rst_n;
  assign Module2Func_62_ap_start = Module2Func_62__ap_start;
  assign Module2Func_62_fifo_ld_0_peek_dout = from_t1_iter63_to_t1_iter64__dout;
  assign Module2Func_62_fifo_ld_0_peek_empty_n = from_t1_iter63_to_t1_iter64__empty_n;
  assign Module2Func_62_fifo_ld_0_s_dout = from_t1_iter63_to_t1_iter64__dout;
  assign Module2Func_62_fifo_ld_0_s_empty_n = from_t1_iter63_to_t1_iter64__empty_n;
  assign from_t1_iter63_to_t1_iter64__read = Module2Func_62_fifo_ld_0_s_read;
  assign from_t1_iter64_to_t1_iter65__din = Module2Func_62_fifo_st_0_din;
  assign Module2Func_62_fifo_st_0_full_n = from_t1_iter64_to_t1_iter65__full_n;
  assign from_t1_iter64_to_t1_iter65__write = Module2Func_62_fifo_st_0_write;
  assign Module2Func_63_ap_clk = ap_clk;
  assign Module2Func_63_ap_rst_n = ap_rst_n;
  assign Module2Func_63_ap_start = Module2Func_63__ap_start;
  assign Module2Func_63_fifo_ld_0_peek_dout = from_t1_iter64_to_t1_iter65__dout;
  assign Module2Func_63_fifo_ld_0_peek_empty_n = from_t1_iter64_to_t1_iter65__empty_n;
  assign Module2Func_63_fifo_ld_0_s_dout = from_t1_iter64_to_t1_iter65__dout;
  assign Module2Func_63_fifo_ld_0_s_empty_n = from_t1_iter64_to_t1_iter65__empty_n;
  assign from_t1_iter64_to_t1_iter65__read = Module2Func_63_fifo_ld_0_s_read;
  assign from_t1_iter65_to_t1_iter66__din = Module2Func_63_fifo_st_0_din;
  assign Module2Func_63_fifo_st_0_full_n = from_t1_iter65_to_t1_iter66__full_n;
  assign from_t1_iter65_to_t1_iter66__write = Module2Func_63_fifo_st_0_write;
  assign Module2Func_64_ap_clk = ap_clk;
  assign Module2Func_64_ap_rst_n = ap_rst_n;
  assign Module2Func_64_ap_start = Module2Func_64__ap_start;
  assign Module2Func_64_fifo_ld_0_peek_dout = from_t1_iter65_to_t1_iter66__dout;
  assign Module2Func_64_fifo_ld_0_peek_empty_n = from_t1_iter65_to_t1_iter66__empty_n;
  assign Module2Func_64_fifo_ld_0_s_dout = from_t1_iter65_to_t1_iter66__dout;
  assign Module2Func_64_fifo_ld_0_s_empty_n = from_t1_iter65_to_t1_iter66__empty_n;
  assign from_t1_iter65_to_t1_iter66__read = Module2Func_64_fifo_ld_0_s_read;
  assign from_t1_iter66_to_t1_iter67__din = Module2Func_64_fifo_st_0_din;
  assign Module2Func_64_fifo_st_0_full_n = from_t1_iter66_to_t1_iter67__full_n;
  assign from_t1_iter66_to_t1_iter67__write = Module2Func_64_fifo_st_0_write;
  assign Module2Func_65_ap_clk = ap_clk;
  assign Module2Func_65_ap_rst_n = ap_rst_n;
  assign Module2Func_65_ap_start = Module2Func_65__ap_start;
  assign Module2Func_65_fifo_ld_0_peek_dout = from_t1_iter66_to_t1_iter67__dout;
  assign Module2Func_65_fifo_ld_0_peek_empty_n = from_t1_iter66_to_t1_iter67__empty_n;
  assign Module2Func_65_fifo_ld_0_s_dout = from_t1_iter66_to_t1_iter67__dout;
  assign Module2Func_65_fifo_ld_0_s_empty_n = from_t1_iter66_to_t1_iter67__empty_n;
  assign from_t1_iter66_to_t1_iter67__read = Module2Func_65_fifo_ld_0_s_read;
  assign from_t1_iter67_to_t1_iter68__din = Module2Func_65_fifo_st_0_din;
  assign Module2Func_65_fifo_st_0_full_n = from_t1_iter67_to_t1_iter68__full_n;
  assign from_t1_iter67_to_t1_iter68__write = Module2Func_65_fifo_st_0_write;
  assign Module2Func_66_ap_clk = ap_clk;
  assign Module2Func_66_ap_rst_n = ap_rst_n;
  assign Module2Func_66_ap_start = Module2Func_66__ap_start;
  assign Module2Func_66_fifo_ld_0_peek_dout = from_t1_iter67_to_t1_iter68__dout;
  assign Module2Func_66_fifo_ld_0_peek_empty_n = from_t1_iter67_to_t1_iter68__empty_n;
  assign Module2Func_66_fifo_ld_0_s_dout = from_t1_iter67_to_t1_iter68__dout;
  assign Module2Func_66_fifo_ld_0_s_empty_n = from_t1_iter67_to_t1_iter68__empty_n;
  assign from_t1_iter67_to_t1_iter68__read = Module2Func_66_fifo_ld_0_s_read;
  assign from_t1_iter68_to_t1_iter69__din = Module2Func_66_fifo_st_0_din;
  assign Module2Func_66_fifo_st_0_full_n = from_t1_iter68_to_t1_iter69__full_n;
  assign from_t1_iter68_to_t1_iter69__write = Module2Func_66_fifo_st_0_write;
  assign Module2Func_67_ap_clk = ap_clk;
  assign Module2Func_67_ap_rst_n = ap_rst_n;
  assign Module2Func_67_ap_start = Module2Func_67__ap_start;
  assign Module2Func_67_fifo_ld_0_peek_dout = from_t1_iter68_to_t1_iter69__dout;
  assign Module2Func_67_fifo_ld_0_peek_empty_n = from_t1_iter68_to_t1_iter69__empty_n;
  assign Module2Func_67_fifo_ld_0_s_dout = from_t1_iter68_to_t1_iter69__dout;
  assign Module2Func_67_fifo_ld_0_s_empty_n = from_t1_iter68_to_t1_iter69__empty_n;
  assign from_t1_iter68_to_t1_iter69__read = Module2Func_67_fifo_ld_0_s_read;
  assign from_t1_iter69_to_t1_iter70__din = Module2Func_67_fifo_st_0_din;
  assign Module2Func_67_fifo_st_0_full_n = from_t1_iter69_to_t1_iter70__full_n;
  assign from_t1_iter69_to_t1_iter70__write = Module2Func_67_fifo_st_0_write;
  assign Module2Func_68_ap_clk = ap_clk;
  assign Module2Func_68_ap_rst_n = ap_rst_n;
  assign Module2Func_68_ap_start = Module2Func_68__ap_start;
  assign Module2Func_68_fifo_ld_0_peek_dout = from_t1_iter69_to_t1_iter70__dout;
  assign Module2Func_68_fifo_ld_0_peek_empty_n = from_t1_iter69_to_t1_iter70__empty_n;
  assign Module2Func_68_fifo_ld_0_s_dout = from_t1_iter69_to_t1_iter70__dout;
  assign Module2Func_68_fifo_ld_0_s_empty_n = from_t1_iter69_to_t1_iter70__empty_n;
  assign from_t1_iter69_to_t1_iter70__read = Module2Func_68_fifo_ld_0_s_read;
  assign from_t1_iter70_to_t1_iter71__din = Module2Func_68_fifo_st_0_din;
  assign Module2Func_68_fifo_st_0_full_n = from_t1_iter70_to_t1_iter71__full_n;
  assign from_t1_iter70_to_t1_iter71__write = Module2Func_68_fifo_st_0_write;
  assign Module2Func_69_ap_clk = ap_clk;
  assign Module2Func_69_ap_rst_n = ap_rst_n;
  assign Module2Func_69_ap_start = Module2Func_69__ap_start;
  assign Module2Func_69_fifo_ld_0_peek_dout = from_t1_iter70_to_t1_iter71__dout;
  assign Module2Func_69_fifo_ld_0_peek_empty_n = from_t1_iter70_to_t1_iter71__empty_n;
  assign Module2Func_69_fifo_ld_0_s_dout = from_t1_iter70_to_t1_iter71__dout;
  assign Module2Func_69_fifo_ld_0_s_empty_n = from_t1_iter70_to_t1_iter71__empty_n;
  assign from_t1_iter70_to_t1_iter71__read = Module2Func_69_fifo_ld_0_s_read;
  assign from_t1_iter71_to_t1_iter72__din = Module2Func_69_fifo_st_0_din;
  assign Module2Func_69_fifo_st_0_full_n = from_t1_iter71_to_t1_iter72__full_n;
  assign from_t1_iter71_to_t1_iter72__write = Module2Func_69_fifo_st_0_write;
  assign Module2Func_70_ap_clk = ap_clk;
  assign Module2Func_70_ap_rst_n = ap_rst_n;
  assign Module2Func_70_ap_start = Module2Func_70__ap_start;
  assign Module2Func_70_fifo_ld_0_peek_dout = from_t1_iter71_to_t1_iter72__dout;
  assign Module2Func_70_fifo_ld_0_peek_empty_n = from_t1_iter71_to_t1_iter72__empty_n;
  assign Module2Func_70_fifo_ld_0_s_dout = from_t1_iter71_to_t1_iter72__dout;
  assign Module2Func_70_fifo_ld_0_s_empty_n = from_t1_iter71_to_t1_iter72__empty_n;
  assign from_t1_iter71_to_t1_iter72__read = Module2Func_70_fifo_ld_0_s_read;
  assign from_t1_iter72_to_t1_iter73__din = Module2Func_70_fifo_st_0_din;
  assign Module2Func_70_fifo_st_0_full_n = from_t1_iter72_to_t1_iter73__full_n;
  assign from_t1_iter72_to_t1_iter73__write = Module2Func_70_fifo_st_0_write;
  assign Module2Func_71_ap_clk = ap_clk;
  assign Module2Func_71_ap_rst_n = ap_rst_n;
  assign Module2Func_71_ap_start = Module2Func_71__ap_start;
  assign Module2Func_71_fifo_ld_0_peek_dout = from_t1_iter72_to_t1_iter73__dout;
  assign Module2Func_71_fifo_ld_0_peek_empty_n = from_t1_iter72_to_t1_iter73__empty_n;
  assign Module2Func_71_fifo_ld_0_s_dout = from_t1_iter72_to_t1_iter73__dout;
  assign Module2Func_71_fifo_ld_0_s_empty_n = from_t1_iter72_to_t1_iter73__empty_n;
  assign from_t1_iter72_to_t1_iter73__read = Module2Func_71_fifo_ld_0_s_read;
  assign from_t1_iter73_to_t1_iter74__din = Module2Func_71_fifo_st_0_din;
  assign Module2Func_71_fifo_st_0_full_n = from_t1_iter73_to_t1_iter74__full_n;
  assign from_t1_iter73_to_t1_iter74__write = Module2Func_71_fifo_st_0_write;
  assign Module2Func_72_ap_clk = ap_clk;
  assign Module2Func_72_ap_rst_n = ap_rst_n;
  assign Module2Func_72_ap_start = Module2Func_72__ap_start;
  assign Module2Func_72_fifo_ld_0_peek_dout = from_t1_iter73_to_t1_iter74__dout;
  assign Module2Func_72_fifo_ld_0_peek_empty_n = from_t1_iter73_to_t1_iter74__empty_n;
  assign Module2Func_72_fifo_ld_0_s_dout = from_t1_iter73_to_t1_iter74__dout;
  assign Module2Func_72_fifo_ld_0_s_empty_n = from_t1_iter73_to_t1_iter74__empty_n;
  assign from_t1_iter73_to_t1_iter74__read = Module2Func_72_fifo_ld_0_s_read;
  assign from_t1_iter74_to_t1_iter75__din = Module2Func_72_fifo_st_0_din;
  assign Module2Func_72_fifo_st_0_full_n = from_t1_iter74_to_t1_iter75__full_n;
  assign from_t1_iter74_to_t1_iter75__write = Module2Func_72_fifo_st_0_write;
  assign Module2Func_73_ap_clk = ap_clk;
  assign Module2Func_73_ap_rst_n = ap_rst_n;
  assign Module2Func_73_ap_start = Module2Func_73__ap_start;
  assign Module2Func_73_fifo_ld_0_peek_dout = from_t1_iter74_to_t1_iter75__dout;
  assign Module2Func_73_fifo_ld_0_peek_empty_n = from_t1_iter74_to_t1_iter75__empty_n;
  assign Module2Func_73_fifo_ld_0_s_dout = from_t1_iter74_to_t1_iter75__dout;
  assign Module2Func_73_fifo_ld_0_s_empty_n = from_t1_iter74_to_t1_iter75__empty_n;
  assign from_t1_iter74_to_t1_iter75__read = Module2Func_73_fifo_ld_0_s_read;
  assign from_t1_iter75_to_t1_iter76__din = Module2Func_73_fifo_st_0_din;
  assign Module2Func_73_fifo_st_0_full_n = from_t1_iter75_to_t1_iter76__full_n;
  assign from_t1_iter75_to_t1_iter76__write = Module2Func_73_fifo_st_0_write;
  assign Module2Func_74_ap_clk = ap_clk;
  assign Module2Func_74_ap_rst_n = ap_rst_n;
  assign Module2Func_74_ap_start = Module2Func_74__ap_start;
  assign Module2Func_74_fifo_ld_0_peek_dout = from_t1_iter75_to_t1_iter76__dout;
  assign Module2Func_74_fifo_ld_0_peek_empty_n = from_t1_iter75_to_t1_iter76__empty_n;
  assign Module2Func_74_fifo_ld_0_s_dout = from_t1_iter75_to_t1_iter76__dout;
  assign Module2Func_74_fifo_ld_0_s_empty_n = from_t1_iter75_to_t1_iter76__empty_n;
  assign from_t1_iter75_to_t1_iter76__read = Module2Func_74_fifo_ld_0_s_read;
  assign from_t1_iter76_to_t1_iter77__din = Module2Func_74_fifo_st_0_din;
  assign Module2Func_74_fifo_st_0_full_n = from_t1_iter76_to_t1_iter77__full_n;
  assign from_t1_iter76_to_t1_iter77__write = Module2Func_74_fifo_st_0_write;
  assign Module2Func_75_ap_clk = ap_clk;
  assign Module2Func_75_ap_rst_n = ap_rst_n;
  assign Module2Func_75_ap_start = Module2Func_75__ap_start;
  assign Module2Func_75_fifo_ld_0_peek_dout = from_t1_iter76_to_t1_iter77__dout;
  assign Module2Func_75_fifo_ld_0_peek_empty_n = from_t1_iter76_to_t1_iter77__empty_n;
  assign Module2Func_75_fifo_ld_0_s_dout = from_t1_iter76_to_t1_iter77__dout;
  assign Module2Func_75_fifo_ld_0_s_empty_n = from_t1_iter76_to_t1_iter77__empty_n;
  assign from_t1_iter76_to_t1_iter77__read = Module2Func_75_fifo_ld_0_s_read;
  assign from_t1_iter77_to_t1_iter78__din = Module2Func_75_fifo_st_0_din;
  assign Module2Func_75_fifo_st_0_full_n = from_t1_iter77_to_t1_iter78__full_n;
  assign from_t1_iter77_to_t1_iter78__write = Module2Func_75_fifo_st_0_write;
  assign Module2Func_76_ap_clk = ap_clk;
  assign Module2Func_76_ap_rst_n = ap_rst_n;
  assign Module2Func_76_ap_start = Module2Func_76__ap_start;
  assign Module2Func_76_fifo_ld_0_peek_dout = from_t1_iter77_to_t1_iter78__dout;
  assign Module2Func_76_fifo_ld_0_peek_empty_n = from_t1_iter77_to_t1_iter78__empty_n;
  assign Module2Func_76_fifo_ld_0_s_dout = from_t1_iter77_to_t1_iter78__dout;
  assign Module2Func_76_fifo_ld_0_s_empty_n = from_t1_iter77_to_t1_iter78__empty_n;
  assign from_t1_iter77_to_t1_iter78__read = Module2Func_76_fifo_ld_0_s_read;
  assign from_t1_iter78_to_t1_iter79__din = Module2Func_76_fifo_st_0_din;
  assign Module2Func_76_fifo_st_0_full_n = from_t1_iter78_to_t1_iter79__full_n;
  assign from_t1_iter78_to_t1_iter79__write = Module2Func_76_fifo_st_0_write;
  assign Module2Func_77_ap_clk = ap_clk;
  assign Module2Func_77_ap_rst_n = ap_rst_n;
  assign Module2Func_77_ap_start = Module2Func_77__ap_start;
  assign Module2Func_77_fifo_ld_0_peek_dout = from_t1_iter78_to_t1_iter79__dout;
  assign Module2Func_77_fifo_ld_0_peek_empty_n = from_t1_iter78_to_t1_iter79__empty_n;
  assign Module2Func_77_fifo_ld_0_s_dout = from_t1_iter78_to_t1_iter79__dout;
  assign Module2Func_77_fifo_ld_0_s_empty_n = from_t1_iter78_to_t1_iter79__empty_n;
  assign from_t1_iter78_to_t1_iter79__read = Module2Func_77_fifo_ld_0_s_read;
  assign from_t1_iter79_to_t1_iter80__din = Module2Func_77_fifo_st_0_din;
  assign Module2Func_77_fifo_st_0_full_n = from_t1_iter79_to_t1_iter80__full_n;
  assign from_t1_iter79_to_t1_iter80__write = Module2Func_77_fifo_st_0_write;
  assign Module2Func_78_ap_clk = ap_clk;
  assign Module2Func_78_ap_rst_n = ap_rst_n;
  assign Module2Func_78_ap_start = Module2Func_78__ap_start;
  assign Module2Func_78_fifo_ld_0_peek_dout = from_t1_iter79_to_t1_iter80__dout;
  assign Module2Func_78_fifo_ld_0_peek_empty_n = from_t1_iter79_to_t1_iter80__empty_n;
  assign Module2Func_78_fifo_ld_0_s_dout = from_t1_iter79_to_t1_iter80__dout;
  assign Module2Func_78_fifo_ld_0_s_empty_n = from_t1_iter79_to_t1_iter80__empty_n;
  assign from_t1_iter79_to_t1_iter80__read = Module2Func_78_fifo_ld_0_s_read;
  assign from_t1_iter80_to_t1_iter81__din = Module2Func_78_fifo_st_0_din;
  assign Module2Func_78_fifo_st_0_full_n = from_t1_iter80_to_t1_iter81__full_n;
  assign from_t1_iter80_to_t1_iter81__write = Module2Func_78_fifo_st_0_write;
  assign Module2Func_79_ap_clk = ap_clk;
  assign Module2Func_79_ap_rst_n = ap_rst_n;
  assign Module2Func_79_ap_start = Module2Func_79__ap_start;
  assign Module2Func_79_fifo_ld_0_peek_dout = from_t1_iter80_to_t1_iter81__dout;
  assign Module2Func_79_fifo_ld_0_peek_empty_n = from_t1_iter80_to_t1_iter81__empty_n;
  assign Module2Func_79_fifo_ld_0_s_dout = from_t1_iter80_to_t1_iter81__dout;
  assign Module2Func_79_fifo_ld_0_s_empty_n = from_t1_iter80_to_t1_iter81__empty_n;
  assign from_t1_iter80_to_t1_iter81__read = Module2Func_79_fifo_ld_0_s_read;
  assign from_t1_iter81_to_t1_iter82__din = Module2Func_79_fifo_st_0_din;
  assign Module2Func_79_fifo_st_0_full_n = from_t1_iter81_to_t1_iter82__full_n;
  assign from_t1_iter81_to_t1_iter82__write = Module2Func_79_fifo_st_0_write;
  assign Module2Func_80_ap_clk = ap_clk;
  assign Module2Func_80_ap_rst_n = ap_rst_n;
  assign Module2Func_80_ap_start = Module2Func_80__ap_start;
  assign Module2Func_80_fifo_ld_0_peek_dout = from_t1_iter81_to_t1_iter82__dout;
  assign Module2Func_80_fifo_ld_0_peek_empty_n = from_t1_iter81_to_t1_iter82__empty_n;
  assign Module2Func_80_fifo_ld_0_s_dout = from_t1_iter81_to_t1_iter82__dout;
  assign Module2Func_80_fifo_ld_0_s_empty_n = from_t1_iter81_to_t1_iter82__empty_n;
  assign from_t1_iter81_to_t1_iter82__read = Module2Func_80_fifo_ld_0_s_read;
  assign from_t1_iter82_to_t1_iter83__din = Module2Func_80_fifo_st_0_din;
  assign Module2Func_80_fifo_st_0_full_n = from_t1_iter82_to_t1_iter83__full_n;
  assign from_t1_iter82_to_t1_iter83__write = Module2Func_80_fifo_st_0_write;
  assign Module2Func_81_ap_clk = ap_clk;
  assign Module2Func_81_ap_rst_n = ap_rst_n;
  assign Module2Func_81_ap_start = Module2Func_81__ap_start;
  assign Module2Func_81_fifo_ld_0_peek_dout = from_t1_iter82_to_t1_iter83__dout;
  assign Module2Func_81_fifo_ld_0_peek_empty_n = from_t1_iter82_to_t1_iter83__empty_n;
  assign Module2Func_81_fifo_ld_0_s_dout = from_t1_iter82_to_t1_iter83__dout;
  assign Module2Func_81_fifo_ld_0_s_empty_n = from_t1_iter82_to_t1_iter83__empty_n;
  assign from_t1_iter82_to_t1_iter83__read = Module2Func_81_fifo_ld_0_s_read;
  assign from_t1_iter83_to_t1_iter84__din = Module2Func_81_fifo_st_0_din;
  assign Module2Func_81_fifo_st_0_full_n = from_t1_iter83_to_t1_iter84__full_n;
  assign from_t1_iter83_to_t1_iter84__write = Module2Func_81_fifo_st_0_write;
  assign Module2Func_82_ap_clk = ap_clk;
  assign Module2Func_82_ap_rst_n = ap_rst_n;
  assign Module2Func_82_ap_start = Module2Func_82__ap_start;
  assign Module2Func_82_fifo_ld_0_peek_dout = from_t1_iter83_to_t1_iter84__dout;
  assign Module2Func_82_fifo_ld_0_peek_empty_n = from_t1_iter83_to_t1_iter84__empty_n;
  assign Module2Func_82_fifo_ld_0_s_dout = from_t1_iter83_to_t1_iter84__dout;
  assign Module2Func_82_fifo_ld_0_s_empty_n = from_t1_iter83_to_t1_iter84__empty_n;
  assign from_t1_iter83_to_t1_iter84__read = Module2Func_82_fifo_ld_0_s_read;
  assign from_t1_iter84_to_t1_iter85__din = Module2Func_82_fifo_st_0_din;
  assign Module2Func_82_fifo_st_0_full_n = from_t1_iter84_to_t1_iter85__full_n;
  assign from_t1_iter84_to_t1_iter85__write = Module2Func_82_fifo_st_0_write;
  assign Module2Func_83_ap_clk = ap_clk;
  assign Module2Func_83_ap_rst_n = ap_rst_n;
  assign Module2Func_83_ap_start = Module2Func_83__ap_start;
  assign Module2Func_83_fifo_ld_0_peek_dout = from_t1_iter84_to_t1_iter85__dout;
  assign Module2Func_83_fifo_ld_0_peek_empty_n = from_t1_iter84_to_t1_iter85__empty_n;
  assign Module2Func_83_fifo_ld_0_s_dout = from_t1_iter84_to_t1_iter85__dout;
  assign Module2Func_83_fifo_ld_0_s_empty_n = from_t1_iter84_to_t1_iter85__empty_n;
  assign from_t1_iter84_to_t1_iter85__read = Module2Func_83_fifo_ld_0_s_read;
  assign from_t1_iter85_to_t1_iter86__din = Module2Func_83_fifo_st_0_din;
  assign Module2Func_83_fifo_st_0_full_n = from_t1_iter85_to_t1_iter86__full_n;
  assign from_t1_iter85_to_t1_iter86__write = Module2Func_83_fifo_st_0_write;
  assign Module2Func_84_ap_clk = ap_clk;
  assign Module2Func_84_ap_rst_n = ap_rst_n;
  assign Module2Func_84_ap_start = Module2Func_84__ap_start;
  assign Module2Func_84_fifo_ld_0_peek_dout = from_t1_iter85_to_t1_iter86__dout;
  assign Module2Func_84_fifo_ld_0_peek_empty_n = from_t1_iter85_to_t1_iter86__empty_n;
  assign Module2Func_84_fifo_ld_0_s_dout = from_t1_iter85_to_t1_iter86__dout;
  assign Module2Func_84_fifo_ld_0_s_empty_n = from_t1_iter85_to_t1_iter86__empty_n;
  assign from_t1_iter85_to_t1_iter86__read = Module2Func_84_fifo_ld_0_s_read;
  assign from_t1_iter86_to_t1_iter87__din = Module2Func_84_fifo_st_0_din;
  assign Module2Func_84_fifo_st_0_full_n = from_t1_iter86_to_t1_iter87__full_n;
  assign from_t1_iter86_to_t1_iter87__write = Module2Func_84_fifo_st_0_write;
  assign Module2Func_85_ap_clk = ap_clk;
  assign Module2Func_85_ap_rst_n = ap_rst_n;
  assign Module2Func_85_ap_start = Module2Func_85__ap_start;
  assign Module2Func_85_fifo_ld_0_peek_dout = from_t1_iter86_to_t1_iter87__dout;
  assign Module2Func_85_fifo_ld_0_peek_empty_n = from_t1_iter86_to_t1_iter87__empty_n;
  assign Module2Func_85_fifo_ld_0_s_dout = from_t1_iter86_to_t1_iter87__dout;
  assign Module2Func_85_fifo_ld_0_s_empty_n = from_t1_iter86_to_t1_iter87__empty_n;
  assign from_t1_iter86_to_t1_iter87__read = Module2Func_85_fifo_ld_0_s_read;
  assign from_t1_iter87_to_t1_iter88__din = Module2Func_85_fifo_st_0_din;
  assign Module2Func_85_fifo_st_0_full_n = from_t1_iter87_to_t1_iter88__full_n;
  assign from_t1_iter87_to_t1_iter88__write = Module2Func_85_fifo_st_0_write;
  assign Module2Func_86_ap_clk = ap_clk;
  assign Module2Func_86_ap_rst_n = ap_rst_n;
  assign Module2Func_86_ap_start = Module2Func_86__ap_start;
  assign Module2Func_86_fifo_ld_0_peek_dout = from_t1_iter87_to_t1_iter88__dout;
  assign Module2Func_86_fifo_ld_0_peek_empty_n = from_t1_iter87_to_t1_iter88__empty_n;
  assign Module2Func_86_fifo_ld_0_s_dout = from_t1_iter87_to_t1_iter88__dout;
  assign Module2Func_86_fifo_ld_0_s_empty_n = from_t1_iter87_to_t1_iter88__empty_n;
  assign from_t1_iter87_to_t1_iter88__read = Module2Func_86_fifo_ld_0_s_read;
  assign from_t1_iter88_to_t1_iter89__din = Module2Func_86_fifo_st_0_din;
  assign Module2Func_86_fifo_st_0_full_n = from_t1_iter88_to_t1_iter89__full_n;
  assign from_t1_iter88_to_t1_iter89__write = Module2Func_86_fifo_st_0_write;
  assign Module2Func_87_ap_clk = ap_clk;
  assign Module2Func_87_ap_rst_n = ap_rst_n;
  assign Module2Func_87_ap_start = Module2Func_87__ap_start;
  assign Module2Func_87_fifo_ld_0_peek_dout = from_t1_iter88_to_t1_iter89__dout;
  assign Module2Func_87_fifo_ld_0_peek_empty_n = from_t1_iter88_to_t1_iter89__empty_n;
  assign Module2Func_87_fifo_ld_0_s_dout = from_t1_iter88_to_t1_iter89__dout;
  assign Module2Func_87_fifo_ld_0_s_empty_n = from_t1_iter88_to_t1_iter89__empty_n;
  assign from_t1_iter88_to_t1_iter89__read = Module2Func_87_fifo_ld_0_s_read;
  assign from_t1_iter89_to_t1_iter90__din = Module2Func_87_fifo_st_0_din;
  assign Module2Func_87_fifo_st_0_full_n = from_t1_iter89_to_t1_iter90__full_n;
  assign from_t1_iter89_to_t1_iter90__write = Module2Func_87_fifo_st_0_write;
  assign Module2Func_88_ap_clk = ap_clk;
  assign Module2Func_88_ap_rst_n = ap_rst_n;
  assign Module2Func_88_ap_start = Module2Func_88__ap_start;
  assign Module2Func_88_fifo_ld_0_peek_dout = from_t1_iter89_to_t1_iter90__dout;
  assign Module2Func_88_fifo_ld_0_peek_empty_n = from_t1_iter89_to_t1_iter90__empty_n;
  assign Module2Func_88_fifo_ld_0_s_dout = from_t1_iter89_to_t1_iter90__dout;
  assign Module2Func_88_fifo_ld_0_s_empty_n = from_t1_iter89_to_t1_iter90__empty_n;
  assign from_t1_iter89_to_t1_iter90__read = Module2Func_88_fifo_ld_0_s_read;
  assign from_t1_iter90_to_t1_iter91__din = Module2Func_88_fifo_st_0_din;
  assign Module2Func_88_fifo_st_0_full_n = from_t1_iter90_to_t1_iter91__full_n;
  assign from_t1_iter90_to_t1_iter91__write = Module2Func_88_fifo_st_0_write;
  assign Module2Func_89_ap_clk = ap_clk;
  assign Module2Func_89_ap_rst_n = ap_rst_n;
  assign Module2Func_89_ap_start = Module2Func_89__ap_start;
  assign Module2Func_89_fifo_ld_0_peek_dout = from_t1_iter90_to_t1_iter91__dout;
  assign Module2Func_89_fifo_ld_0_peek_empty_n = from_t1_iter90_to_t1_iter91__empty_n;
  assign Module2Func_89_fifo_ld_0_s_dout = from_t1_iter90_to_t1_iter91__dout;
  assign Module2Func_89_fifo_ld_0_s_empty_n = from_t1_iter90_to_t1_iter91__empty_n;
  assign from_t1_iter90_to_t1_iter91__read = Module2Func_89_fifo_ld_0_s_read;
  assign from_t1_iter91_to_t1_iter92__din = Module2Func_89_fifo_st_0_din;
  assign Module2Func_89_fifo_st_0_full_n = from_t1_iter91_to_t1_iter92__full_n;
  assign from_t1_iter91_to_t1_iter92__write = Module2Func_89_fifo_st_0_write;
  assign Module2Func_90_ap_clk = ap_clk;
  assign Module2Func_90_ap_rst_n = ap_rst_n;
  assign Module2Func_90_ap_start = Module2Func_90__ap_start;
  assign Module2Func_90_fifo_ld_0_peek_dout = from_t1_iter91_to_t1_iter92__dout;
  assign Module2Func_90_fifo_ld_0_peek_empty_n = from_t1_iter91_to_t1_iter92__empty_n;
  assign Module2Func_90_fifo_ld_0_s_dout = from_t1_iter91_to_t1_iter92__dout;
  assign Module2Func_90_fifo_ld_0_s_empty_n = from_t1_iter91_to_t1_iter92__empty_n;
  assign from_t1_iter91_to_t1_iter92__read = Module2Func_90_fifo_ld_0_s_read;
  assign from_t1_iter92_to_t1_iter93__din = Module2Func_90_fifo_st_0_din;
  assign Module2Func_90_fifo_st_0_full_n = from_t1_iter92_to_t1_iter93__full_n;
  assign from_t1_iter92_to_t1_iter93__write = Module2Func_90_fifo_st_0_write;
  assign Module2Func_91_ap_clk = ap_clk;
  assign Module2Func_91_ap_rst_n = ap_rst_n;
  assign Module2Func_91_ap_start = Module2Func_91__ap_start;
  assign Module2Func_91_fifo_ld_0_peek_dout = from_t1_iter92_to_t1_iter93__dout;
  assign Module2Func_91_fifo_ld_0_peek_empty_n = from_t1_iter92_to_t1_iter93__empty_n;
  assign Module2Func_91_fifo_ld_0_s_dout = from_t1_iter92_to_t1_iter93__dout;
  assign Module2Func_91_fifo_ld_0_s_empty_n = from_t1_iter92_to_t1_iter93__empty_n;
  assign from_t1_iter92_to_t1_iter93__read = Module2Func_91_fifo_ld_0_s_read;
  assign from_t1_iter93_to_t1_iter94__din = Module2Func_91_fifo_st_0_din;
  assign Module2Func_91_fifo_st_0_full_n = from_t1_iter93_to_t1_iter94__full_n;
  assign from_t1_iter93_to_t1_iter94__write = Module2Func_91_fifo_st_0_write;
  assign Module2Func_92_ap_clk = ap_clk;
  assign Module2Func_92_ap_rst_n = ap_rst_n;
  assign Module2Func_92_ap_start = Module2Func_92__ap_start;
  assign Module2Func_92_fifo_ld_0_peek_dout = from_t1_iter93_to_t1_iter94__dout;
  assign Module2Func_92_fifo_ld_0_peek_empty_n = from_t1_iter93_to_t1_iter94__empty_n;
  assign Module2Func_92_fifo_ld_0_s_dout = from_t1_iter93_to_t1_iter94__dout;
  assign Module2Func_92_fifo_ld_0_s_empty_n = from_t1_iter93_to_t1_iter94__empty_n;
  assign from_t1_iter93_to_t1_iter94__read = Module2Func_92_fifo_ld_0_s_read;
  assign from_t1_iter94_to_t1_iter95__din = Module2Func_92_fifo_st_0_din;
  assign Module2Func_92_fifo_st_0_full_n = from_t1_iter94_to_t1_iter95__full_n;
  assign from_t1_iter94_to_t1_iter95__write = Module2Func_92_fifo_st_0_write;
  assign Module2Func_93_ap_clk = ap_clk;
  assign Module2Func_93_ap_rst_n = ap_rst_n;
  assign Module2Func_93_ap_start = Module2Func_93__ap_start;
  assign Module2Func_93_fifo_ld_0_peek_dout = from_t1_iter94_to_t1_iter95__dout;
  assign Module2Func_93_fifo_ld_0_peek_empty_n = from_t1_iter94_to_t1_iter95__empty_n;
  assign Module2Func_93_fifo_ld_0_s_dout = from_t1_iter94_to_t1_iter95__dout;
  assign Module2Func_93_fifo_ld_0_s_empty_n = from_t1_iter94_to_t1_iter95__empty_n;
  assign from_t1_iter94_to_t1_iter95__read = Module2Func_93_fifo_ld_0_s_read;
  assign from_t1_iter95_to_t1_iter96__din = Module2Func_93_fifo_st_0_din;
  assign Module2Func_93_fifo_st_0_full_n = from_t1_iter95_to_t1_iter96__full_n;
  assign from_t1_iter95_to_t1_iter96__write = Module2Func_93_fifo_st_0_write;
  assign Module2Func_94_ap_clk = ap_clk;
  assign Module2Func_94_ap_rst_n = ap_rst_n;
  assign Module2Func_94_ap_start = Module2Func_94__ap_start;
  assign Module2Func_94_fifo_ld_0_peek_dout = from_t1_iter95_to_t1_iter96__dout;
  assign Module2Func_94_fifo_ld_0_peek_empty_n = from_t1_iter95_to_t1_iter96__empty_n;
  assign Module2Func_94_fifo_ld_0_s_dout = from_t1_iter95_to_t1_iter96__dout;
  assign Module2Func_94_fifo_ld_0_s_empty_n = from_t1_iter95_to_t1_iter96__empty_n;
  assign from_t1_iter95_to_t1_iter96__read = Module2Func_94_fifo_ld_0_s_read;
  assign from_t1_iter96_to_t1_iter97__din = Module2Func_94_fifo_st_0_din;
  assign Module2Func_94_fifo_st_0_full_n = from_t1_iter96_to_t1_iter97__full_n;
  assign from_t1_iter96_to_t1_iter97__write = Module2Func_94_fifo_st_0_write;
  assign Module2Func_95_ap_clk = ap_clk;
  assign Module2Func_95_ap_rst_n = ap_rst_n;
  assign Module2Func_95_ap_start = Module2Func_95__ap_start;
  assign Module2Func_95_fifo_ld_0_peek_dout = from_t1_iter96_to_t1_iter97__dout;
  assign Module2Func_95_fifo_ld_0_peek_empty_n = from_t1_iter96_to_t1_iter97__empty_n;
  assign Module2Func_95_fifo_ld_0_s_dout = from_t1_iter96_to_t1_iter97__dout;
  assign Module2Func_95_fifo_ld_0_s_empty_n = from_t1_iter96_to_t1_iter97__empty_n;
  assign from_t1_iter96_to_t1_iter97__read = Module2Func_95_fifo_ld_0_s_read;
  assign from_t1_iter97_to_t1_iter98__din = Module2Func_95_fifo_st_0_din;
  assign Module2Func_95_fifo_st_0_full_n = from_t1_iter97_to_t1_iter98__full_n;
  assign from_t1_iter97_to_t1_iter98__write = Module2Func_95_fifo_st_0_write;
  assign Module2Func_96_ap_clk = ap_clk;
  assign Module2Func_96_ap_rst_n = ap_rst_n;
  assign Module2Func_96_ap_start = Module2Func_96__ap_start;
  assign Module2Func_96_fifo_ld_0_peek_dout = from_t1_iter97_to_t1_iter98__dout;
  assign Module2Func_96_fifo_ld_0_peek_empty_n = from_t1_iter97_to_t1_iter98__empty_n;
  assign Module2Func_96_fifo_ld_0_s_dout = from_t1_iter97_to_t1_iter98__dout;
  assign Module2Func_96_fifo_ld_0_s_empty_n = from_t1_iter97_to_t1_iter98__empty_n;
  assign from_t1_iter97_to_t1_iter98__read = Module2Func_96_fifo_ld_0_s_read;
  assign from_t1_iter98_to_t1_iter99__din = Module2Func_96_fifo_st_0_din;
  assign Module2Func_96_fifo_st_0_full_n = from_t1_iter98_to_t1_iter99__full_n;
  assign from_t1_iter98_to_t1_iter99__write = Module2Func_96_fifo_st_0_write;
  assign Module2Func_97_ap_clk = ap_clk;
  assign Module2Func_97_ap_rst_n = ap_rst_n;
  assign Module2Func_97_ap_start = Module2Func_97__ap_start;
  assign Module2Func_97_fifo_ld_0_peek_dout = from_t1_iter98_to_t1_iter99__dout;
  assign Module2Func_97_fifo_ld_0_peek_empty_n = from_t1_iter98_to_t1_iter99__empty_n;
  assign Module2Func_97_fifo_ld_0_s_dout = from_t1_iter98_to_t1_iter99__dout;
  assign Module2Func_97_fifo_ld_0_s_empty_n = from_t1_iter98_to_t1_iter99__empty_n;
  assign from_t1_iter98_to_t1_iter99__read = Module2Func_97_fifo_ld_0_s_read;
  assign from_t1_iter99_to_t1_iter100__din = Module2Func_97_fifo_st_0_din;
  assign Module2Func_97_fifo_st_0_full_n = from_t1_iter99_to_t1_iter100__full_n;
  assign from_t1_iter99_to_t1_iter100__write = Module2Func_97_fifo_st_0_write;
  assign Module2Func_98_ap_clk = ap_clk;
  assign Module2Func_98_ap_rst_n = ap_rst_n;
  assign Module2Func_98_ap_start = Module2Func_98__ap_start;
  assign Module2Func_98_fifo_ld_0_peek_dout = from_t1_iter99_to_t1_iter100__dout;
  assign Module2Func_98_fifo_ld_0_peek_empty_n = from_t1_iter99_to_t1_iter100__empty_n;
  assign Module2Func_98_fifo_ld_0_s_dout = from_t1_iter99_to_t1_iter100__dout;
  assign Module2Func_98_fifo_ld_0_s_empty_n = from_t1_iter99_to_t1_iter100__empty_n;
  assign from_t1_iter99_to_t1_iter100__read = Module2Func_98_fifo_ld_0_s_read;
  assign from_t1_iter100_to_t1_iter101__din = Module2Func_98_fifo_st_0_din;
  assign Module2Func_98_fifo_st_0_full_n = from_t1_iter100_to_t1_iter101__full_n;
  assign from_t1_iter100_to_t1_iter101__write = Module2Func_98_fifo_st_0_write;
  assign Module2Func_99_ap_clk = ap_clk;
  assign Module2Func_99_ap_rst_n = ap_rst_n;
  assign Module2Func_99_ap_start = Module2Func_99__ap_start;
  assign Module2Func_99_fifo_ld_0_peek_dout = from_t1_iter100_to_t1_iter101__dout;
  assign Module2Func_99_fifo_ld_0_peek_empty_n = from_t1_iter100_to_t1_iter101__empty_n;
  assign Module2Func_99_fifo_ld_0_s_dout = from_t1_iter100_to_t1_iter101__dout;
  assign Module2Func_99_fifo_ld_0_s_empty_n = from_t1_iter100_to_t1_iter101__empty_n;
  assign from_t1_iter100_to_t1_iter101__read = Module2Func_99_fifo_ld_0_s_read;
  assign from_t1_iter101_to_t1_iter102__din = Module2Func_99_fifo_st_0_din;
  assign Module2Func_99_fifo_st_0_full_n = from_t1_iter101_to_t1_iter102__full_n;
  assign from_t1_iter101_to_t1_iter102__write = Module2Func_99_fifo_st_0_write;
  assign Module2Func_100_ap_clk = ap_clk;
  assign Module2Func_100_ap_rst_n = ap_rst_n;
  assign Module2Func_100_ap_start = Module2Func_100__ap_start;
  assign Module2Func_100_fifo_ld_0_peek_dout = from_t1_iter101_to_t1_iter102__dout;
  assign Module2Func_100_fifo_ld_0_peek_empty_n = from_t1_iter101_to_t1_iter102__empty_n;
  assign Module2Func_100_fifo_ld_0_s_dout = from_t1_iter101_to_t1_iter102__dout;
  assign Module2Func_100_fifo_ld_0_s_empty_n = from_t1_iter101_to_t1_iter102__empty_n;
  assign from_t1_iter101_to_t1_iter102__read = Module2Func_100_fifo_ld_0_s_read;
  assign from_t1_iter102_to_t1_iter103__din = Module2Func_100_fifo_st_0_din;
  assign Module2Func_100_fifo_st_0_full_n = from_t1_iter102_to_t1_iter103__full_n;
  assign from_t1_iter102_to_t1_iter103__write = Module2Func_100_fifo_st_0_write;
  assign Module2Func_101_ap_clk = ap_clk;
  assign Module2Func_101_ap_rst_n = ap_rst_n;
  assign Module2Func_101_ap_start = Module2Func_101__ap_start;
  assign Module2Func_101_fifo_ld_0_peek_dout = from_t1_iter102_to_t1_iter103__dout;
  assign Module2Func_101_fifo_ld_0_peek_empty_n = from_t1_iter102_to_t1_iter103__empty_n;
  assign Module2Func_101_fifo_ld_0_s_dout = from_t1_iter102_to_t1_iter103__dout;
  assign Module2Func_101_fifo_ld_0_s_empty_n = from_t1_iter102_to_t1_iter103__empty_n;
  assign from_t1_iter102_to_t1_iter103__read = Module2Func_101_fifo_ld_0_s_read;
  assign from_t1_iter103_to_t1_iter104__din = Module2Func_101_fifo_st_0_din;
  assign Module2Func_101_fifo_st_0_full_n = from_t1_iter103_to_t1_iter104__full_n;
  assign from_t1_iter103_to_t1_iter104__write = Module2Func_101_fifo_st_0_write;
  assign Module2Func_102_ap_clk = ap_clk;
  assign Module2Func_102_ap_rst_n = ap_rst_n;
  assign Module2Func_102_ap_start = Module2Func_102__ap_start;
  assign Module2Func_102_fifo_ld_0_peek_dout = from_t1_iter103_to_t1_iter104__dout;
  assign Module2Func_102_fifo_ld_0_peek_empty_n = from_t1_iter103_to_t1_iter104__empty_n;
  assign Module2Func_102_fifo_ld_0_s_dout = from_t1_iter103_to_t1_iter104__dout;
  assign Module2Func_102_fifo_ld_0_s_empty_n = from_t1_iter103_to_t1_iter104__empty_n;
  assign from_t1_iter103_to_t1_iter104__read = Module2Func_102_fifo_ld_0_s_read;
  assign from_t1_iter104_to_t1_iter105__din = Module2Func_102_fifo_st_0_din;
  assign Module2Func_102_fifo_st_0_full_n = from_t1_iter104_to_t1_iter105__full_n;
  assign from_t1_iter104_to_t1_iter105__write = Module2Func_102_fifo_st_0_write;
  assign Module2Func_103_ap_clk = ap_clk;
  assign Module2Func_103_ap_rst_n = ap_rst_n;
  assign Module2Func_103_ap_start = Module2Func_103__ap_start;
  assign Module2Func_103_fifo_ld_0_peek_dout = from_t1_iter104_to_t1_iter105__dout;
  assign Module2Func_103_fifo_ld_0_peek_empty_n = from_t1_iter104_to_t1_iter105__empty_n;
  assign Module2Func_103_fifo_ld_0_s_dout = from_t1_iter104_to_t1_iter105__dout;
  assign Module2Func_103_fifo_ld_0_s_empty_n = from_t1_iter104_to_t1_iter105__empty_n;
  assign from_t1_iter104_to_t1_iter105__read = Module2Func_103_fifo_ld_0_s_read;
  assign from_t1_iter105_to_t1_iter106__din = Module2Func_103_fifo_st_0_din;
  assign Module2Func_103_fifo_st_0_full_n = from_t1_iter105_to_t1_iter106__full_n;
  assign from_t1_iter105_to_t1_iter106__write = Module2Func_103_fifo_st_0_write;
  assign Module2Func_104_ap_clk = ap_clk;
  assign Module2Func_104_ap_rst_n = ap_rst_n;
  assign Module2Func_104_ap_start = Module2Func_104__ap_start;
  assign Module2Func_104_fifo_ld_0_peek_dout = from_t1_iter105_to_t1_iter106__dout;
  assign Module2Func_104_fifo_ld_0_peek_empty_n = from_t1_iter105_to_t1_iter106__empty_n;
  assign Module2Func_104_fifo_ld_0_s_dout = from_t1_iter105_to_t1_iter106__dout;
  assign Module2Func_104_fifo_ld_0_s_empty_n = from_t1_iter105_to_t1_iter106__empty_n;
  assign from_t1_iter105_to_t1_iter106__read = Module2Func_104_fifo_ld_0_s_read;
  assign from_t1_iter106_to_t1_iter107__din = Module2Func_104_fifo_st_0_din;
  assign Module2Func_104_fifo_st_0_full_n = from_t1_iter106_to_t1_iter107__full_n;
  assign from_t1_iter106_to_t1_iter107__write = Module2Func_104_fifo_st_0_write;
  assign Module2Func_105_ap_clk = ap_clk;
  assign Module2Func_105_ap_rst_n = ap_rst_n;
  assign Module2Func_105_ap_start = Module2Func_105__ap_start;
  assign Module2Func_105_fifo_ld_0_peek_dout = from_t1_iter106_to_t1_iter107__dout;
  assign Module2Func_105_fifo_ld_0_peek_empty_n = from_t1_iter106_to_t1_iter107__empty_n;
  assign Module2Func_105_fifo_ld_0_s_dout = from_t1_iter106_to_t1_iter107__dout;
  assign Module2Func_105_fifo_ld_0_s_empty_n = from_t1_iter106_to_t1_iter107__empty_n;
  assign from_t1_iter106_to_t1_iter107__read = Module2Func_105_fifo_ld_0_s_read;
  assign from_t1_iter107_to_t1_iter108__din = Module2Func_105_fifo_st_0_din;
  assign Module2Func_105_fifo_st_0_full_n = from_t1_iter107_to_t1_iter108__full_n;
  assign from_t1_iter107_to_t1_iter108__write = Module2Func_105_fifo_st_0_write;
  assign Module2Func_106_ap_clk = ap_clk;
  assign Module2Func_106_ap_rst_n = ap_rst_n;
  assign Module2Func_106_ap_start = Module2Func_106__ap_start;
  assign Module2Func_106_fifo_ld_0_peek_dout = from_t1_iter107_to_t1_iter108__dout;
  assign Module2Func_106_fifo_ld_0_peek_empty_n = from_t1_iter107_to_t1_iter108__empty_n;
  assign Module2Func_106_fifo_ld_0_s_dout = from_t1_iter107_to_t1_iter108__dout;
  assign Module2Func_106_fifo_ld_0_s_empty_n = from_t1_iter107_to_t1_iter108__empty_n;
  assign from_t1_iter107_to_t1_iter108__read = Module2Func_106_fifo_ld_0_s_read;
  assign from_t1_iter108_to_t0__din = Module2Func_106_fifo_st_0_din;
  assign Module2Func_106_fifo_st_0_full_n = from_t1_iter108_to_t0__full_n;
  assign from_t1_iter108_to_t0__write = Module2Func_106_fifo_st_0_write;
  assign Module2Func_107_ap_clk = ap_clk;
  assign Module2Func_107_ap_rst_n = ap_rst_n;
  assign Module2Func_107_ap_start = Module2Func_107__ap_start;
  assign Module2Func_107_fifo_ld_0_peek_dout = from_t1_iter108_to_t0__dout;
  assign Module2Func_107_fifo_ld_0_peek_empty_n = from_t1_iter108_to_t0__empty_n;
  assign Module2Func_107_fifo_ld_0_s_dout = from_t1_iter108_to_t0__dout;
  assign Module2Func_107_fifo_ld_0_s_empty_n = from_t1_iter108_to_t0__empty_n;
  assign from_t1_iter108_to_t0__read = Module2Func_107_fifo_ld_0_s_read;
  assign from_t0_to_t0_bank_1__din = Module2Func_107_fifo_st_0_din;
  assign Module2Func_107_fifo_st_0_full_n = from_t0_to_t0_bank_1__full_n;
  assign from_t0_to_t0_bank_1__write = Module2Func_107_fifo_st_0_write;
  assign Module3Func_0_ap_clk = ap_clk;
  assign Module3Func_0_ap_rst_n = ap_rst_n;
  assign Module3Func_0_ap_start = Module3Func_0__ap_start;
  assign bank_1_t0_buf__din = Module3Func_0_dram_t0_bank_1_fifo_din;
  assign Module3Func_0_dram_t0_bank_1_fifo_full_n = bank_1_t0_buf__full_n;
  assign bank_1_t0_buf__write = Module3Func_0_dram_t0_bank_1_fifo_write;
  assign Module3Func_0_fifo_ld_0_peek_dout = from_t0_to_t0_bank_1__dout;
  assign Module3Func_0_fifo_ld_0_peek_empty_n = from_t0_to_t0_bank_1__empty_n;
  assign Module3Func_0_fifo_ld_0_s_dout = from_t0_to_t0_bank_1__dout;
  assign Module3Func_0_fifo_ld_0_s_empty_n = from_t0_to_t0_bank_1__empty_n;
  assign from_t0_to_t0_bank_1__read = Module3Func_0_fifo_ld_0_s_read;
  assign bank_0_t1__m_axi_clk = ap_clk;
  assign m_axi_bank_0_t1_ARADDR = bank_0_t1__m_axi_m_axi_ARADDR;
  assign m_axi_bank_0_t1_ARBURST = bank_0_t1__m_axi_m_axi_ARBURST;
  assign m_axi_bank_0_t1_ARCACHE = bank_0_t1__m_axi_m_axi_ARCACHE;
  assign m_axi_bank_0_t1_ARID = bank_0_t1__m_axi_m_axi_ARID;
  assign m_axi_bank_0_t1_ARLEN = bank_0_t1__m_axi_m_axi_ARLEN;
  assign m_axi_bank_0_t1_ARLOCK = bank_0_t1__m_axi_m_axi_ARLOCK;
  assign m_axi_bank_0_t1_ARPROT = bank_0_t1__m_axi_m_axi_ARPROT;
  assign m_axi_bank_0_t1_ARQOS = bank_0_t1__m_axi_m_axi_ARQOS;
  assign bank_0_t1__m_axi_m_axi_ARREADY = m_axi_bank_0_t1_ARREADY;
  assign m_axi_bank_0_t1_ARSIZE = bank_0_t1__m_axi_m_axi_ARSIZE;
  assign m_axi_bank_0_t1_ARVALID = bank_0_t1__m_axi_m_axi_ARVALID;
  assign m_axi_bank_0_t1_AWADDR = bank_0_t1__m_axi_m_axi_AWADDR;
  assign m_axi_bank_0_t1_AWBURST = bank_0_t1__m_axi_m_axi_AWBURST;
  assign m_axi_bank_0_t1_AWCACHE = bank_0_t1__m_axi_m_axi_AWCACHE;
  assign m_axi_bank_0_t1_AWID = bank_0_t1__m_axi_m_axi_AWID;
  assign m_axi_bank_0_t1_AWLEN = bank_0_t1__m_axi_m_axi_AWLEN;
  assign m_axi_bank_0_t1_AWLOCK = bank_0_t1__m_axi_m_axi_AWLOCK;
  assign m_axi_bank_0_t1_AWPROT = bank_0_t1__m_axi_m_axi_AWPROT;
  assign m_axi_bank_0_t1_AWQOS = bank_0_t1__m_axi_m_axi_AWQOS;
  assign bank_0_t1__m_axi_m_axi_AWREADY = m_axi_bank_0_t1_AWREADY;
  assign m_axi_bank_0_t1_AWSIZE = bank_0_t1__m_axi_m_axi_AWSIZE;
  assign m_axi_bank_0_t1_AWVALID = bank_0_t1__m_axi_m_axi_AWVALID;
  assign bank_0_t1__m_axi_m_axi_BID = m_axi_bank_0_t1_BID;
  assign m_axi_bank_0_t1_BREADY = bank_0_t1__m_axi_m_axi_BREADY;
  assign bank_0_t1__m_axi_m_axi_BRESP = m_axi_bank_0_t1_BRESP;
  assign bank_0_t1__m_axi_m_axi_BVALID = m_axi_bank_0_t1_BVALID;
  assign bank_0_t1__m_axi_m_axi_RDATA = m_axi_bank_0_t1_RDATA;
  assign bank_0_t1__m_axi_m_axi_RID = m_axi_bank_0_t1_RID;
  assign bank_0_t1__m_axi_m_axi_RLAST = m_axi_bank_0_t1_RLAST;
  assign m_axi_bank_0_t1_RREADY = bank_0_t1__m_axi_m_axi_RREADY;
  assign bank_0_t1__m_axi_m_axi_RRESP = m_axi_bank_0_t1_RRESP;
  assign bank_0_t1__m_axi_m_axi_RVALID = m_axi_bank_0_t1_RVALID;
  assign m_axi_bank_0_t1_WDATA = bank_0_t1__m_axi_m_axi_WDATA;
  assign m_axi_bank_0_t1_WLAST = bank_0_t1__m_axi_m_axi_WLAST;
  assign bank_0_t1__m_axi_m_axi_WREADY = m_axi_bank_0_t1_WREADY;
  assign m_axi_bank_0_t1_WSTRB = bank_0_t1__m_axi_m_axi_WSTRB;
  assign m_axi_bank_0_t1_WVALID = bank_0_t1__m_axi_m_axi_WVALID;
  assign bank_0_t1__m_axi_read_addr_din = bank_0_t1_read_addr__din;
  assign bank_0_t1_read_addr__full_n = bank_0_t1__m_axi_read_addr_full_n;
  assign bank_0_t1__m_axi_read_addr_write = bank_0_t1_read_addr__write;
  assign bank_0_t1_read_data__dout = bank_0_t1__m_axi_read_data_dout;
  assign bank_0_t1_read_data__empty_n = bank_0_t1__m_axi_read_data_empty_n;
  assign bank_0_t1__m_axi_read_data_read = bank_0_t1_read_data__read;
  assign bank_0_t1__m_axi_rst = ~ ap_rst_n;
  assign bank_0_t1__m_axi_write_addr_din = bank_0_t1_write_addr__din;
  assign bank_0_t1_write_addr__full_n = bank_0_t1__m_axi_write_addr_full_n;
  assign bank_0_t1__m_axi_write_addr_write = bank_0_t1_write_addr__write;
  assign bank_0_t1__m_axi_write_data_din = bank_0_t1_write_data__din;
  assign bank_0_t1_write_data__full_n = bank_0_t1__m_axi_write_data_full_n;
  assign bank_0_t1__m_axi_write_data_write = bank_0_t1_write_data__write;
  assign bank_0_t1_write_resp__dout = bank_0_t1__m_axi_write_resp_dout;
  assign bank_0_t1_write_resp__empty_n = bank_0_t1__m_axi_write_resp_empty_n;
  assign bank_0_t1__m_axi_write_resp_read = bank_0_t1_write_resp__read;
  assign bank_1_t0__m_axi_clk = ap_clk;
  assign m_axi_bank_1_t0_ARADDR = bank_1_t0__m_axi_m_axi_ARADDR;
  assign m_axi_bank_1_t0_ARBURST = bank_1_t0__m_axi_m_axi_ARBURST;
  assign m_axi_bank_1_t0_ARCACHE = bank_1_t0__m_axi_m_axi_ARCACHE;
  assign m_axi_bank_1_t0_ARID = bank_1_t0__m_axi_m_axi_ARID;
  assign m_axi_bank_1_t0_ARLEN = bank_1_t0__m_axi_m_axi_ARLEN;
  assign m_axi_bank_1_t0_ARLOCK = bank_1_t0__m_axi_m_axi_ARLOCK;
  assign m_axi_bank_1_t0_ARPROT = bank_1_t0__m_axi_m_axi_ARPROT;
  assign m_axi_bank_1_t0_ARQOS = bank_1_t0__m_axi_m_axi_ARQOS;
  assign bank_1_t0__m_axi_m_axi_ARREADY = m_axi_bank_1_t0_ARREADY;
  assign m_axi_bank_1_t0_ARSIZE = bank_1_t0__m_axi_m_axi_ARSIZE;
  assign m_axi_bank_1_t0_ARVALID = bank_1_t0__m_axi_m_axi_ARVALID;
  assign m_axi_bank_1_t0_AWADDR = bank_1_t0__m_axi_m_axi_AWADDR;
  assign m_axi_bank_1_t0_AWBURST = bank_1_t0__m_axi_m_axi_AWBURST;
  assign m_axi_bank_1_t0_AWCACHE = bank_1_t0__m_axi_m_axi_AWCACHE;
  assign m_axi_bank_1_t0_AWID = bank_1_t0__m_axi_m_axi_AWID;
  assign m_axi_bank_1_t0_AWLEN = bank_1_t0__m_axi_m_axi_AWLEN;
  assign m_axi_bank_1_t0_AWLOCK = bank_1_t0__m_axi_m_axi_AWLOCK;
  assign m_axi_bank_1_t0_AWPROT = bank_1_t0__m_axi_m_axi_AWPROT;
  assign m_axi_bank_1_t0_AWQOS = bank_1_t0__m_axi_m_axi_AWQOS;
  assign bank_1_t0__m_axi_m_axi_AWREADY = m_axi_bank_1_t0_AWREADY;
  assign m_axi_bank_1_t0_AWSIZE = bank_1_t0__m_axi_m_axi_AWSIZE;
  assign m_axi_bank_1_t0_AWVALID = bank_1_t0__m_axi_m_axi_AWVALID;
  assign bank_1_t0__m_axi_m_axi_BID = m_axi_bank_1_t0_BID;
  assign m_axi_bank_1_t0_BREADY = bank_1_t0__m_axi_m_axi_BREADY;
  assign bank_1_t0__m_axi_m_axi_BRESP = m_axi_bank_1_t0_BRESP;
  assign bank_1_t0__m_axi_m_axi_BVALID = m_axi_bank_1_t0_BVALID;
  assign bank_1_t0__m_axi_m_axi_RDATA = m_axi_bank_1_t0_RDATA;
  assign bank_1_t0__m_axi_m_axi_RID = m_axi_bank_1_t0_RID;
  assign bank_1_t0__m_axi_m_axi_RLAST = m_axi_bank_1_t0_RLAST;
  assign m_axi_bank_1_t0_RREADY = bank_1_t0__m_axi_m_axi_RREADY;
  assign bank_1_t0__m_axi_m_axi_RRESP = m_axi_bank_1_t0_RRESP;
  assign bank_1_t0__m_axi_m_axi_RVALID = m_axi_bank_1_t0_RVALID;
  assign m_axi_bank_1_t0_WDATA = bank_1_t0__m_axi_m_axi_WDATA;
  assign m_axi_bank_1_t0_WLAST = bank_1_t0__m_axi_m_axi_WLAST;
  assign bank_1_t0__m_axi_m_axi_WREADY = m_axi_bank_1_t0_WREADY;
  assign m_axi_bank_1_t0_WSTRB = bank_1_t0__m_axi_m_axi_WSTRB;
  assign m_axi_bank_1_t0_WVALID = bank_1_t0__m_axi_m_axi_WVALID;
  assign bank_1_t0__m_axi_read_addr_din = bank_1_t0_read_addr__din;
  assign bank_1_t0_read_addr__full_n = bank_1_t0__m_axi_read_addr_full_n;
  assign bank_1_t0__m_axi_read_addr_write = bank_1_t0_read_addr__write;
  assign bank_1_t0_read_data__dout = bank_1_t0__m_axi_read_data_dout;
  assign bank_1_t0_read_data__empty_n = bank_1_t0__m_axi_read_data_empty_n;
  assign bank_1_t0__m_axi_read_data_read = bank_1_t0_read_data__read;
  assign bank_1_t0__m_axi_rst = ~ ap_rst_n;
  assign bank_1_t0__m_axi_write_addr_din = bank_1_t0_write_addr__din;
  assign bank_1_t0_write_addr__full_n = bank_1_t0__m_axi_write_addr_full_n;
  assign bank_1_t0__m_axi_write_addr_write = bank_1_t0_write_addr__write;
  assign bank_1_t0__m_axi_write_data_din = bank_1_t0_write_data__din;
  assign bank_1_t0_write_data__full_n = bank_1_t0__m_axi_write_data_full_n;
  assign bank_1_t0__m_axi_write_data_write = bank_1_t0_write_data__write;
  assign bank_1_t0_write_resp__dout = bank_1_t0__m_axi_write_resp_dout;
  assign bank_1_t0_write_resp__empty_n = bank_1_t0__m_axi_write_resp_empty_n;
  assign bank_1_t0__m_axi_write_resp_read = bank_1_t0_write_resp__read;
  assign BurstRead_floatx16_0___bank_0_t1__q0 = __tapa_fsm_unit_BurstRead_floatx16_0___bank_0_t1__q0;
  assign BurstRead_floatx16_0___coalesced_data_num__q0 = __tapa_fsm_unit_BurstRead_floatx16_0___coalesced_data_num__q0;
  assign __tapa_fsm_unit_BurstRead_floatx16_0__ap_done = BurstRead_floatx16_0__ap_done;
  assign __tapa_fsm_unit_BurstRead_floatx16_0__ap_idle = BurstRead_floatx16_0__ap_idle;
  assign __tapa_fsm_unit_BurstRead_floatx16_0__ap_ready = BurstRead_floatx16_0__ap_ready;
  assign BurstRead_floatx16_0__ap_start = __tapa_fsm_unit_BurstRead_floatx16_0__ap_start;
  assign BurstWrite_floatx16_0___bank_1_t0__q0 = __tapa_fsm_unit_BurstWrite_floatx16_0___bank_1_t0__q0;
  assign BurstWrite_floatx16_0___coalesced_data_num__q0 = __tapa_fsm_unit_BurstWrite_floatx16_0___coalesced_data_num__q0;
  assign __tapa_fsm_unit_BurstWrite_floatx16_0__ap_done = BurstWrite_floatx16_0__ap_done;
  assign __tapa_fsm_unit_BurstWrite_floatx16_0__ap_idle = BurstWrite_floatx16_0__ap_idle;
  assign __tapa_fsm_unit_BurstWrite_floatx16_0__ap_ready = BurstWrite_floatx16_0__ap_ready;
  assign BurstWrite_floatx16_0__ap_start = __tapa_fsm_unit_BurstWrite_floatx16_0__ap_start;
  assign Module0Func_0__ap_start = __tapa_fsm_unit_Module0Func_0__ap_start;
  assign Module1Func_0__ap_start = __tapa_fsm_unit_Module1Func_0__ap_start;
  assign Module2Func_0__ap_start = __tapa_fsm_unit_Module2Func_0__ap_start;
  assign Module2Func_100__ap_start = __tapa_fsm_unit_Module2Func_100__ap_start;
  assign Module2Func_101__ap_start = __tapa_fsm_unit_Module2Func_101__ap_start;
  assign Module2Func_102__ap_start = __tapa_fsm_unit_Module2Func_102__ap_start;
  assign Module2Func_103__ap_start = __tapa_fsm_unit_Module2Func_103__ap_start;
  assign Module2Func_104__ap_start = __tapa_fsm_unit_Module2Func_104__ap_start;
  assign Module2Func_105__ap_start = __tapa_fsm_unit_Module2Func_105__ap_start;
  assign Module2Func_106__ap_start = __tapa_fsm_unit_Module2Func_106__ap_start;
  assign Module2Func_107__ap_start = __tapa_fsm_unit_Module2Func_107__ap_start;
  assign Module2Func_10__ap_start = __tapa_fsm_unit_Module2Func_10__ap_start;
  assign Module2Func_11__ap_start = __tapa_fsm_unit_Module2Func_11__ap_start;
  assign Module2Func_12__ap_start = __tapa_fsm_unit_Module2Func_12__ap_start;
  assign Module2Func_13__ap_start = __tapa_fsm_unit_Module2Func_13__ap_start;
  assign Module2Func_14__ap_start = __tapa_fsm_unit_Module2Func_14__ap_start;
  assign Module2Func_15__ap_start = __tapa_fsm_unit_Module2Func_15__ap_start;
  assign Module2Func_16__ap_start = __tapa_fsm_unit_Module2Func_16__ap_start;
  assign Module2Func_17__ap_start = __tapa_fsm_unit_Module2Func_17__ap_start;
  assign Module2Func_18__ap_start = __tapa_fsm_unit_Module2Func_18__ap_start;
  assign Module2Func_19__ap_start = __tapa_fsm_unit_Module2Func_19__ap_start;
  assign Module2Func_1__ap_start = __tapa_fsm_unit_Module2Func_1__ap_start;
  assign Module2Func_20__ap_start = __tapa_fsm_unit_Module2Func_20__ap_start;
  assign Module2Func_21__ap_start = __tapa_fsm_unit_Module2Func_21__ap_start;
  assign Module2Func_22__ap_start = __tapa_fsm_unit_Module2Func_22__ap_start;
  assign Module2Func_23__ap_start = __tapa_fsm_unit_Module2Func_23__ap_start;
  assign Module2Func_24__ap_start = __tapa_fsm_unit_Module2Func_24__ap_start;
  assign Module2Func_25__ap_start = __tapa_fsm_unit_Module2Func_25__ap_start;
  assign Module2Func_26__ap_start = __tapa_fsm_unit_Module2Func_26__ap_start;
  assign Module2Func_27__ap_start = __tapa_fsm_unit_Module2Func_27__ap_start;
  assign Module2Func_28__ap_start = __tapa_fsm_unit_Module2Func_28__ap_start;
  assign Module2Func_29__ap_start = __tapa_fsm_unit_Module2Func_29__ap_start;
  assign Module2Func_2__ap_start = __tapa_fsm_unit_Module2Func_2__ap_start;
  assign Module2Func_30__ap_start = __tapa_fsm_unit_Module2Func_30__ap_start;
  assign Module2Func_31__ap_start = __tapa_fsm_unit_Module2Func_31__ap_start;
  assign Module2Func_32__ap_start = __tapa_fsm_unit_Module2Func_32__ap_start;
  assign Module2Func_33__ap_start = __tapa_fsm_unit_Module2Func_33__ap_start;
  assign Module2Func_34__ap_start = __tapa_fsm_unit_Module2Func_34__ap_start;
  assign Module2Func_35__ap_start = __tapa_fsm_unit_Module2Func_35__ap_start;
  assign Module2Func_36__ap_start = __tapa_fsm_unit_Module2Func_36__ap_start;
  assign Module2Func_37__ap_start = __tapa_fsm_unit_Module2Func_37__ap_start;
  assign Module2Func_38__ap_start = __tapa_fsm_unit_Module2Func_38__ap_start;
  assign Module2Func_39__ap_start = __tapa_fsm_unit_Module2Func_39__ap_start;
  assign Module2Func_3__ap_start = __tapa_fsm_unit_Module2Func_3__ap_start;
  assign Module2Func_40__ap_start = __tapa_fsm_unit_Module2Func_40__ap_start;
  assign Module2Func_41__ap_start = __tapa_fsm_unit_Module2Func_41__ap_start;
  assign Module2Func_42__ap_start = __tapa_fsm_unit_Module2Func_42__ap_start;
  assign Module2Func_43__ap_start = __tapa_fsm_unit_Module2Func_43__ap_start;
  assign Module2Func_44__ap_start = __tapa_fsm_unit_Module2Func_44__ap_start;
  assign Module2Func_45__ap_start = __tapa_fsm_unit_Module2Func_45__ap_start;
  assign Module2Func_46__ap_start = __tapa_fsm_unit_Module2Func_46__ap_start;
  assign Module2Func_47__ap_start = __tapa_fsm_unit_Module2Func_47__ap_start;
  assign Module2Func_48__ap_start = __tapa_fsm_unit_Module2Func_48__ap_start;
  assign Module2Func_49__ap_start = __tapa_fsm_unit_Module2Func_49__ap_start;
  assign Module2Func_4__ap_start = __tapa_fsm_unit_Module2Func_4__ap_start;
  assign Module2Func_50__ap_start = __tapa_fsm_unit_Module2Func_50__ap_start;
  assign Module2Func_51__ap_start = __tapa_fsm_unit_Module2Func_51__ap_start;
  assign Module2Func_52__ap_start = __tapa_fsm_unit_Module2Func_52__ap_start;
  assign Module2Func_53__ap_start = __tapa_fsm_unit_Module2Func_53__ap_start;
  assign Module2Func_54__ap_start = __tapa_fsm_unit_Module2Func_54__ap_start;
  assign Module2Func_55__ap_start = __tapa_fsm_unit_Module2Func_55__ap_start;
  assign Module2Func_56__ap_start = __tapa_fsm_unit_Module2Func_56__ap_start;
  assign Module2Func_57__ap_start = __tapa_fsm_unit_Module2Func_57__ap_start;
  assign Module2Func_58__ap_start = __tapa_fsm_unit_Module2Func_58__ap_start;
  assign Module2Func_59__ap_start = __tapa_fsm_unit_Module2Func_59__ap_start;
  assign Module2Func_5__ap_start = __tapa_fsm_unit_Module2Func_5__ap_start;
  assign Module2Func_60__ap_start = __tapa_fsm_unit_Module2Func_60__ap_start;
  assign Module2Func_61__ap_start = __tapa_fsm_unit_Module2Func_61__ap_start;
  assign Module2Func_62__ap_start = __tapa_fsm_unit_Module2Func_62__ap_start;
  assign Module2Func_63__ap_start = __tapa_fsm_unit_Module2Func_63__ap_start;
  assign Module2Func_64__ap_start = __tapa_fsm_unit_Module2Func_64__ap_start;
  assign Module2Func_65__ap_start = __tapa_fsm_unit_Module2Func_65__ap_start;
  assign Module2Func_66__ap_start = __tapa_fsm_unit_Module2Func_66__ap_start;
  assign Module2Func_67__ap_start = __tapa_fsm_unit_Module2Func_67__ap_start;
  assign Module2Func_68__ap_start = __tapa_fsm_unit_Module2Func_68__ap_start;
  assign Module2Func_69__ap_start = __tapa_fsm_unit_Module2Func_69__ap_start;
  assign Module2Func_6__ap_start = __tapa_fsm_unit_Module2Func_6__ap_start;
  assign Module2Func_70__ap_start = __tapa_fsm_unit_Module2Func_70__ap_start;
  assign Module2Func_71__ap_start = __tapa_fsm_unit_Module2Func_71__ap_start;
  assign Module2Func_72__ap_start = __tapa_fsm_unit_Module2Func_72__ap_start;
  assign Module2Func_73__ap_start = __tapa_fsm_unit_Module2Func_73__ap_start;
  assign Module2Func_74__ap_start = __tapa_fsm_unit_Module2Func_74__ap_start;
  assign Module2Func_75__ap_start = __tapa_fsm_unit_Module2Func_75__ap_start;
  assign Module2Func_76__ap_start = __tapa_fsm_unit_Module2Func_76__ap_start;
  assign Module2Func_77__ap_start = __tapa_fsm_unit_Module2Func_77__ap_start;
  assign Module2Func_78__ap_start = __tapa_fsm_unit_Module2Func_78__ap_start;
  assign Module2Func_79__ap_start = __tapa_fsm_unit_Module2Func_79__ap_start;
  assign Module2Func_7__ap_start = __tapa_fsm_unit_Module2Func_7__ap_start;
  assign Module2Func_80__ap_start = __tapa_fsm_unit_Module2Func_80__ap_start;
  assign Module2Func_81__ap_start = __tapa_fsm_unit_Module2Func_81__ap_start;
  assign Module2Func_82__ap_start = __tapa_fsm_unit_Module2Func_82__ap_start;
  assign Module2Func_83__ap_start = __tapa_fsm_unit_Module2Func_83__ap_start;
  assign Module2Func_84__ap_start = __tapa_fsm_unit_Module2Func_84__ap_start;
  assign Module2Func_85__ap_start = __tapa_fsm_unit_Module2Func_85__ap_start;
  assign Module2Func_86__ap_start = __tapa_fsm_unit_Module2Func_86__ap_start;
  assign Module2Func_87__ap_start = __tapa_fsm_unit_Module2Func_87__ap_start;
  assign Module2Func_88__ap_start = __tapa_fsm_unit_Module2Func_88__ap_start;
  assign Module2Func_89__ap_start = __tapa_fsm_unit_Module2Func_89__ap_start;
  assign Module2Func_8__ap_start = __tapa_fsm_unit_Module2Func_8__ap_start;
  assign Module2Func_90__ap_start = __tapa_fsm_unit_Module2Func_90__ap_start;
  assign Module2Func_91__ap_start = __tapa_fsm_unit_Module2Func_91__ap_start;
  assign Module2Func_92__ap_start = __tapa_fsm_unit_Module2Func_92__ap_start;
  assign Module2Func_93__ap_start = __tapa_fsm_unit_Module2Func_93__ap_start;
  assign Module2Func_94__ap_start = __tapa_fsm_unit_Module2Func_94__ap_start;
  assign Module2Func_95__ap_start = __tapa_fsm_unit_Module2Func_95__ap_start;
  assign Module2Func_96__ap_start = __tapa_fsm_unit_Module2Func_96__ap_start;
  assign Module2Func_97__ap_start = __tapa_fsm_unit_Module2Func_97__ap_start;
  assign Module2Func_98__ap_start = __tapa_fsm_unit_Module2Func_98__ap_start;
  assign Module2Func_99__ap_start = __tapa_fsm_unit_Module2Func_99__ap_start;
  assign Module2Func_9__ap_start = __tapa_fsm_unit_Module2Func_9__ap_start;
  assign Module3Func_0__ap_start = __tapa_fsm_unit_Module3Func_0__ap_start;
  assign __tapa_fsm_unit_ap_clk = ap_clk;
  assign ap_done = __tapa_fsm_unit_ap_done;
  assign ap_idle = __tapa_fsm_unit_ap_idle;
  assign ap_ready = __tapa_fsm_unit_ap_ready;
  assign __tapa_fsm_unit_ap_rst_n = ap_rst_n;
  assign __tapa_fsm_unit_ap_start = ap_start;
  assign __tapa_fsm_unit_bank_0_t1 = bank_0_t1;
  assign __tapa_fsm_unit_bank_1_t0 = bank_1_t0;
  assign __tapa_fsm_unit_coalesced_data_num = coalesced_data_num;
endmodule