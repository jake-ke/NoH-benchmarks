`timescale 1 ns / 1 ps 

(* CORE_GENERATION_INFO = "Knn_Knn,hls_ip_2023_2_2,{HLS_INPUT_TYPE=cxx,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=0,HLS_INPUT_PART=xcvh1582-vsva3697-2MP-e-S,HLS_INPUT_CLOCK=3.330000,HLS_INPUT_ARCH=others,HLS_SYN_CLOCK=1.000000,HLS_SYN_LAT=0,HLS_SYN_TPT=none,HLS_SYN_MEM=0,HLS_SYN_DSP=0,HLS_SYN_FF=2066,HLS_SYN_LUT=3752,HLS_VERSION=2023_2_2}" *)


module Knn
(
  s_axi_control_AWVALID,
  s_axi_control_AWREADY,
  s_axi_control_AWADDR,
  s_axi_control_WVALID,
  s_axi_control_WREADY,
  s_axi_control_WDATA,
  s_axi_control_WSTRB,
  s_axi_control_ARVALID,
  s_axi_control_ARREADY,
  s_axi_control_ARADDR,
  s_axi_control_RVALID,
  s_axi_control_RREADY,
  s_axi_control_RDATA,
  s_axi_control_RRESP,
  s_axi_control_BVALID,
  s_axi_control_BREADY,
  s_axi_control_BRESP,
  ap_clk,
  ap_rst_n,
  interrupt,
  m_axi_L3_out_dist_ARADDR,
  m_axi_L3_out_dist_ARBURST,
  m_axi_L3_out_dist_ARCACHE,
  m_axi_L3_out_dist_ARID,
  m_axi_L3_out_dist_ARLEN,
  m_axi_L3_out_dist_ARLOCK,
  m_axi_L3_out_dist_ARPROT,
  m_axi_L3_out_dist_ARQOS,
  m_axi_L3_out_dist_ARREADY,
  m_axi_L3_out_dist_ARSIZE,
  m_axi_L3_out_dist_ARVALID,
  m_axi_L3_out_dist_AWADDR,
  m_axi_L3_out_dist_AWBURST,
  m_axi_L3_out_dist_AWCACHE,
  m_axi_L3_out_dist_AWID,
  m_axi_L3_out_dist_AWLEN,
  m_axi_L3_out_dist_AWLOCK,
  m_axi_L3_out_dist_AWPROT,
  m_axi_L3_out_dist_AWQOS,
  m_axi_L3_out_dist_AWREADY,
  m_axi_L3_out_dist_AWSIZE,
  m_axi_L3_out_dist_AWVALID,
  m_axi_L3_out_dist_BID,
  m_axi_L3_out_dist_BREADY,
  m_axi_L3_out_dist_BRESP,
  m_axi_L3_out_dist_BVALID,
  m_axi_L3_out_dist_RDATA,
  m_axi_L3_out_dist_RID,
  m_axi_L3_out_dist_RLAST,
  m_axi_L3_out_dist_RREADY,
  m_axi_L3_out_dist_RRESP,
  m_axi_L3_out_dist_RVALID,
  m_axi_L3_out_dist_WDATA,
  m_axi_L3_out_dist_WLAST,
  m_axi_L3_out_dist_WREADY,
  m_axi_L3_out_dist_WSTRB,
  m_axi_L3_out_dist_WVALID,
  m_axi_L3_out_id_ARADDR,
  m_axi_L3_out_id_ARBURST,
  m_axi_L3_out_id_ARCACHE,
  m_axi_L3_out_id_ARID,
  m_axi_L3_out_id_ARLEN,
  m_axi_L3_out_id_ARLOCK,
  m_axi_L3_out_id_ARPROT,
  m_axi_L3_out_id_ARQOS,
  m_axi_L3_out_id_ARREADY,
  m_axi_L3_out_id_ARSIZE,
  m_axi_L3_out_id_ARVALID,
  m_axi_L3_out_id_AWADDR,
  m_axi_L3_out_id_AWBURST,
  m_axi_L3_out_id_AWCACHE,
  m_axi_L3_out_id_AWID,
  m_axi_L3_out_id_AWLEN,
  m_axi_L3_out_id_AWLOCK,
  m_axi_L3_out_id_AWPROT,
  m_axi_L3_out_id_AWQOS,
  m_axi_L3_out_id_AWREADY,
  m_axi_L3_out_id_AWSIZE,
  m_axi_L3_out_id_AWVALID,
  m_axi_L3_out_id_BID,
  m_axi_L3_out_id_BREADY,
  m_axi_L3_out_id_BRESP,
  m_axi_L3_out_id_BVALID,
  m_axi_L3_out_id_RDATA,
  m_axi_L3_out_id_RID,
  m_axi_L3_out_id_RLAST,
  m_axi_L3_out_id_RREADY,
  m_axi_L3_out_id_RRESP,
  m_axi_L3_out_id_RVALID,
  m_axi_L3_out_id_WDATA,
  m_axi_L3_out_id_WLAST,
  m_axi_L3_out_id_WREADY,
  m_axi_L3_out_id_WSTRB,
  m_axi_L3_out_id_WVALID,
  m_axi_in_0_ARADDR,
  m_axi_in_0_ARBURST,
  m_axi_in_0_ARCACHE,
  m_axi_in_0_ARID,
  m_axi_in_0_ARLEN,
  m_axi_in_0_ARLOCK,
  m_axi_in_0_ARPROT,
  m_axi_in_0_ARQOS,
  m_axi_in_0_ARREADY,
  m_axi_in_0_ARSIZE,
  m_axi_in_0_ARVALID,
  m_axi_in_0_AWADDR,
  m_axi_in_0_AWBURST,
  m_axi_in_0_AWCACHE,
  m_axi_in_0_AWID,
  m_axi_in_0_AWLEN,
  m_axi_in_0_AWLOCK,
  m_axi_in_0_AWPROT,
  m_axi_in_0_AWQOS,
  m_axi_in_0_AWREADY,
  m_axi_in_0_AWSIZE,
  m_axi_in_0_AWVALID,
  m_axi_in_0_BID,
  m_axi_in_0_BREADY,
  m_axi_in_0_BRESP,
  m_axi_in_0_BVALID,
  m_axi_in_0_RDATA,
  m_axi_in_0_RID,
  m_axi_in_0_RLAST,
  m_axi_in_0_RREADY,
  m_axi_in_0_RRESP,
  m_axi_in_0_RVALID,
  m_axi_in_0_WDATA,
  m_axi_in_0_WLAST,
  m_axi_in_0_WREADY,
  m_axi_in_0_WSTRB,
  m_axi_in_0_WVALID,
  m_axi_in_1_ARADDR,
  m_axi_in_1_ARBURST,
  m_axi_in_1_ARCACHE,
  m_axi_in_1_ARID,
  m_axi_in_1_ARLEN,
  m_axi_in_1_ARLOCK,
  m_axi_in_1_ARPROT,
  m_axi_in_1_ARQOS,
  m_axi_in_1_ARREADY,
  m_axi_in_1_ARSIZE,
  m_axi_in_1_ARVALID,
  m_axi_in_1_AWADDR,
  m_axi_in_1_AWBURST,
  m_axi_in_1_AWCACHE,
  m_axi_in_1_AWID,
  m_axi_in_1_AWLEN,
  m_axi_in_1_AWLOCK,
  m_axi_in_1_AWPROT,
  m_axi_in_1_AWQOS,
  m_axi_in_1_AWREADY,
  m_axi_in_1_AWSIZE,
  m_axi_in_1_AWVALID,
  m_axi_in_1_BID,
  m_axi_in_1_BREADY,
  m_axi_in_1_BRESP,
  m_axi_in_1_BVALID,
  m_axi_in_1_RDATA,
  m_axi_in_1_RID,
  m_axi_in_1_RLAST,
  m_axi_in_1_RREADY,
  m_axi_in_1_RRESP,
  m_axi_in_1_RVALID,
  m_axi_in_1_WDATA,
  m_axi_in_1_WLAST,
  m_axi_in_1_WREADY,
  m_axi_in_1_WSTRB,
  m_axi_in_1_WVALID,
  m_axi_in_10_ARADDR,
  m_axi_in_10_ARBURST,
  m_axi_in_10_ARCACHE,
  m_axi_in_10_ARID,
  m_axi_in_10_ARLEN,
  m_axi_in_10_ARLOCK,
  m_axi_in_10_ARPROT,
  m_axi_in_10_ARQOS,
  m_axi_in_10_ARREADY,
  m_axi_in_10_ARSIZE,
  m_axi_in_10_ARVALID,
  m_axi_in_10_AWADDR,
  m_axi_in_10_AWBURST,
  m_axi_in_10_AWCACHE,
  m_axi_in_10_AWID,
  m_axi_in_10_AWLEN,
  m_axi_in_10_AWLOCK,
  m_axi_in_10_AWPROT,
  m_axi_in_10_AWQOS,
  m_axi_in_10_AWREADY,
  m_axi_in_10_AWSIZE,
  m_axi_in_10_AWVALID,
  m_axi_in_10_BID,
  m_axi_in_10_BREADY,
  m_axi_in_10_BRESP,
  m_axi_in_10_BVALID,
  m_axi_in_10_RDATA,
  m_axi_in_10_RID,
  m_axi_in_10_RLAST,
  m_axi_in_10_RREADY,
  m_axi_in_10_RRESP,
  m_axi_in_10_RVALID,
  m_axi_in_10_WDATA,
  m_axi_in_10_WLAST,
  m_axi_in_10_WREADY,
  m_axi_in_10_WSTRB,
  m_axi_in_10_WVALID,
  m_axi_in_11_ARADDR,
  m_axi_in_11_ARBURST,
  m_axi_in_11_ARCACHE,
  m_axi_in_11_ARID,
  m_axi_in_11_ARLEN,
  m_axi_in_11_ARLOCK,
  m_axi_in_11_ARPROT,
  m_axi_in_11_ARQOS,
  m_axi_in_11_ARREADY,
  m_axi_in_11_ARSIZE,
  m_axi_in_11_ARVALID,
  m_axi_in_11_AWADDR,
  m_axi_in_11_AWBURST,
  m_axi_in_11_AWCACHE,
  m_axi_in_11_AWID,
  m_axi_in_11_AWLEN,
  m_axi_in_11_AWLOCK,
  m_axi_in_11_AWPROT,
  m_axi_in_11_AWQOS,
  m_axi_in_11_AWREADY,
  m_axi_in_11_AWSIZE,
  m_axi_in_11_AWVALID,
  m_axi_in_11_BID,
  m_axi_in_11_BREADY,
  m_axi_in_11_BRESP,
  m_axi_in_11_BVALID,
  m_axi_in_11_RDATA,
  m_axi_in_11_RID,
  m_axi_in_11_RLAST,
  m_axi_in_11_RREADY,
  m_axi_in_11_RRESP,
  m_axi_in_11_RVALID,
  m_axi_in_11_WDATA,
  m_axi_in_11_WLAST,
  m_axi_in_11_WREADY,
  m_axi_in_11_WSTRB,
  m_axi_in_11_WVALID,
  m_axi_in_12_ARADDR,
  m_axi_in_12_ARBURST,
  m_axi_in_12_ARCACHE,
  m_axi_in_12_ARID,
  m_axi_in_12_ARLEN,
  m_axi_in_12_ARLOCK,
  m_axi_in_12_ARPROT,
  m_axi_in_12_ARQOS,
  m_axi_in_12_ARREADY,
  m_axi_in_12_ARSIZE,
  m_axi_in_12_ARVALID,
  m_axi_in_12_AWADDR,
  m_axi_in_12_AWBURST,
  m_axi_in_12_AWCACHE,
  m_axi_in_12_AWID,
  m_axi_in_12_AWLEN,
  m_axi_in_12_AWLOCK,
  m_axi_in_12_AWPROT,
  m_axi_in_12_AWQOS,
  m_axi_in_12_AWREADY,
  m_axi_in_12_AWSIZE,
  m_axi_in_12_AWVALID,
  m_axi_in_12_BID,
  m_axi_in_12_BREADY,
  m_axi_in_12_BRESP,
  m_axi_in_12_BVALID,
  m_axi_in_12_RDATA,
  m_axi_in_12_RID,
  m_axi_in_12_RLAST,
  m_axi_in_12_RREADY,
  m_axi_in_12_RRESP,
  m_axi_in_12_RVALID,
  m_axi_in_12_WDATA,
  m_axi_in_12_WLAST,
  m_axi_in_12_WREADY,
  m_axi_in_12_WSTRB,
  m_axi_in_12_WVALID,
  m_axi_in_13_ARADDR,
  m_axi_in_13_ARBURST,
  m_axi_in_13_ARCACHE,
  m_axi_in_13_ARID,
  m_axi_in_13_ARLEN,
  m_axi_in_13_ARLOCK,
  m_axi_in_13_ARPROT,
  m_axi_in_13_ARQOS,
  m_axi_in_13_ARREADY,
  m_axi_in_13_ARSIZE,
  m_axi_in_13_ARVALID,
  m_axi_in_13_AWADDR,
  m_axi_in_13_AWBURST,
  m_axi_in_13_AWCACHE,
  m_axi_in_13_AWID,
  m_axi_in_13_AWLEN,
  m_axi_in_13_AWLOCK,
  m_axi_in_13_AWPROT,
  m_axi_in_13_AWQOS,
  m_axi_in_13_AWREADY,
  m_axi_in_13_AWSIZE,
  m_axi_in_13_AWVALID,
  m_axi_in_13_BID,
  m_axi_in_13_BREADY,
  m_axi_in_13_BRESP,
  m_axi_in_13_BVALID,
  m_axi_in_13_RDATA,
  m_axi_in_13_RID,
  m_axi_in_13_RLAST,
  m_axi_in_13_RREADY,
  m_axi_in_13_RRESP,
  m_axi_in_13_RVALID,
  m_axi_in_13_WDATA,
  m_axi_in_13_WLAST,
  m_axi_in_13_WREADY,
  m_axi_in_13_WSTRB,
  m_axi_in_13_WVALID,
  m_axi_in_14_ARADDR,
  m_axi_in_14_ARBURST,
  m_axi_in_14_ARCACHE,
  m_axi_in_14_ARID,
  m_axi_in_14_ARLEN,
  m_axi_in_14_ARLOCK,
  m_axi_in_14_ARPROT,
  m_axi_in_14_ARQOS,
  m_axi_in_14_ARREADY,
  m_axi_in_14_ARSIZE,
  m_axi_in_14_ARVALID,
  m_axi_in_14_AWADDR,
  m_axi_in_14_AWBURST,
  m_axi_in_14_AWCACHE,
  m_axi_in_14_AWID,
  m_axi_in_14_AWLEN,
  m_axi_in_14_AWLOCK,
  m_axi_in_14_AWPROT,
  m_axi_in_14_AWQOS,
  m_axi_in_14_AWREADY,
  m_axi_in_14_AWSIZE,
  m_axi_in_14_AWVALID,
  m_axi_in_14_BID,
  m_axi_in_14_BREADY,
  m_axi_in_14_BRESP,
  m_axi_in_14_BVALID,
  m_axi_in_14_RDATA,
  m_axi_in_14_RID,
  m_axi_in_14_RLAST,
  m_axi_in_14_RREADY,
  m_axi_in_14_RRESP,
  m_axi_in_14_RVALID,
  m_axi_in_14_WDATA,
  m_axi_in_14_WLAST,
  m_axi_in_14_WREADY,
  m_axi_in_14_WSTRB,
  m_axi_in_14_WVALID,
  m_axi_in_15_ARADDR,
  m_axi_in_15_ARBURST,
  m_axi_in_15_ARCACHE,
  m_axi_in_15_ARID,
  m_axi_in_15_ARLEN,
  m_axi_in_15_ARLOCK,
  m_axi_in_15_ARPROT,
  m_axi_in_15_ARQOS,
  m_axi_in_15_ARREADY,
  m_axi_in_15_ARSIZE,
  m_axi_in_15_ARVALID,
  m_axi_in_15_AWADDR,
  m_axi_in_15_AWBURST,
  m_axi_in_15_AWCACHE,
  m_axi_in_15_AWID,
  m_axi_in_15_AWLEN,
  m_axi_in_15_AWLOCK,
  m_axi_in_15_AWPROT,
  m_axi_in_15_AWQOS,
  m_axi_in_15_AWREADY,
  m_axi_in_15_AWSIZE,
  m_axi_in_15_AWVALID,
  m_axi_in_15_BID,
  m_axi_in_15_BREADY,
  m_axi_in_15_BRESP,
  m_axi_in_15_BVALID,
  m_axi_in_15_RDATA,
  m_axi_in_15_RID,
  m_axi_in_15_RLAST,
  m_axi_in_15_RREADY,
  m_axi_in_15_RRESP,
  m_axi_in_15_RVALID,
  m_axi_in_15_WDATA,
  m_axi_in_15_WLAST,
  m_axi_in_15_WREADY,
  m_axi_in_15_WSTRB,
  m_axi_in_15_WVALID,
  m_axi_in_16_ARADDR,
  m_axi_in_16_ARBURST,
  m_axi_in_16_ARCACHE,
  m_axi_in_16_ARID,
  m_axi_in_16_ARLEN,
  m_axi_in_16_ARLOCK,
  m_axi_in_16_ARPROT,
  m_axi_in_16_ARQOS,
  m_axi_in_16_ARREADY,
  m_axi_in_16_ARSIZE,
  m_axi_in_16_ARVALID,
  m_axi_in_16_AWADDR,
  m_axi_in_16_AWBURST,
  m_axi_in_16_AWCACHE,
  m_axi_in_16_AWID,
  m_axi_in_16_AWLEN,
  m_axi_in_16_AWLOCK,
  m_axi_in_16_AWPROT,
  m_axi_in_16_AWQOS,
  m_axi_in_16_AWREADY,
  m_axi_in_16_AWSIZE,
  m_axi_in_16_AWVALID,
  m_axi_in_16_BID,
  m_axi_in_16_BREADY,
  m_axi_in_16_BRESP,
  m_axi_in_16_BVALID,
  m_axi_in_16_RDATA,
  m_axi_in_16_RID,
  m_axi_in_16_RLAST,
  m_axi_in_16_RREADY,
  m_axi_in_16_RRESP,
  m_axi_in_16_RVALID,
  m_axi_in_16_WDATA,
  m_axi_in_16_WLAST,
  m_axi_in_16_WREADY,
  m_axi_in_16_WSTRB,
  m_axi_in_16_WVALID,
  m_axi_in_17_ARADDR,
  m_axi_in_17_ARBURST,
  m_axi_in_17_ARCACHE,
  m_axi_in_17_ARID,
  m_axi_in_17_ARLEN,
  m_axi_in_17_ARLOCK,
  m_axi_in_17_ARPROT,
  m_axi_in_17_ARQOS,
  m_axi_in_17_ARREADY,
  m_axi_in_17_ARSIZE,
  m_axi_in_17_ARVALID,
  m_axi_in_17_AWADDR,
  m_axi_in_17_AWBURST,
  m_axi_in_17_AWCACHE,
  m_axi_in_17_AWID,
  m_axi_in_17_AWLEN,
  m_axi_in_17_AWLOCK,
  m_axi_in_17_AWPROT,
  m_axi_in_17_AWQOS,
  m_axi_in_17_AWREADY,
  m_axi_in_17_AWSIZE,
  m_axi_in_17_AWVALID,
  m_axi_in_17_BID,
  m_axi_in_17_BREADY,
  m_axi_in_17_BRESP,
  m_axi_in_17_BVALID,
  m_axi_in_17_RDATA,
  m_axi_in_17_RID,
  m_axi_in_17_RLAST,
  m_axi_in_17_RREADY,
  m_axi_in_17_RRESP,
  m_axi_in_17_RVALID,
  m_axi_in_17_WDATA,
  m_axi_in_17_WLAST,
  m_axi_in_17_WREADY,
  m_axi_in_17_WSTRB,
  m_axi_in_17_WVALID,
  m_axi_in_18_ARADDR,
  m_axi_in_18_ARBURST,
  m_axi_in_18_ARCACHE,
  m_axi_in_18_ARID,
  m_axi_in_18_ARLEN,
  m_axi_in_18_ARLOCK,
  m_axi_in_18_ARPROT,
  m_axi_in_18_ARQOS,
  m_axi_in_18_ARREADY,
  m_axi_in_18_ARSIZE,
  m_axi_in_18_ARVALID,
  m_axi_in_18_AWADDR,
  m_axi_in_18_AWBURST,
  m_axi_in_18_AWCACHE,
  m_axi_in_18_AWID,
  m_axi_in_18_AWLEN,
  m_axi_in_18_AWLOCK,
  m_axi_in_18_AWPROT,
  m_axi_in_18_AWQOS,
  m_axi_in_18_AWREADY,
  m_axi_in_18_AWSIZE,
  m_axi_in_18_AWVALID,
  m_axi_in_18_BID,
  m_axi_in_18_BREADY,
  m_axi_in_18_BRESP,
  m_axi_in_18_BVALID,
  m_axi_in_18_RDATA,
  m_axi_in_18_RID,
  m_axi_in_18_RLAST,
  m_axi_in_18_RREADY,
  m_axi_in_18_RRESP,
  m_axi_in_18_RVALID,
  m_axi_in_18_WDATA,
  m_axi_in_18_WLAST,
  m_axi_in_18_WREADY,
  m_axi_in_18_WSTRB,
  m_axi_in_18_WVALID,
  m_axi_in_19_ARADDR,
  m_axi_in_19_ARBURST,
  m_axi_in_19_ARCACHE,
  m_axi_in_19_ARID,
  m_axi_in_19_ARLEN,
  m_axi_in_19_ARLOCK,
  m_axi_in_19_ARPROT,
  m_axi_in_19_ARQOS,
  m_axi_in_19_ARREADY,
  m_axi_in_19_ARSIZE,
  m_axi_in_19_ARVALID,
  m_axi_in_19_AWADDR,
  m_axi_in_19_AWBURST,
  m_axi_in_19_AWCACHE,
  m_axi_in_19_AWID,
  m_axi_in_19_AWLEN,
  m_axi_in_19_AWLOCK,
  m_axi_in_19_AWPROT,
  m_axi_in_19_AWQOS,
  m_axi_in_19_AWREADY,
  m_axi_in_19_AWSIZE,
  m_axi_in_19_AWVALID,
  m_axi_in_19_BID,
  m_axi_in_19_BREADY,
  m_axi_in_19_BRESP,
  m_axi_in_19_BVALID,
  m_axi_in_19_RDATA,
  m_axi_in_19_RID,
  m_axi_in_19_RLAST,
  m_axi_in_19_RREADY,
  m_axi_in_19_RRESP,
  m_axi_in_19_RVALID,
  m_axi_in_19_WDATA,
  m_axi_in_19_WLAST,
  m_axi_in_19_WREADY,
  m_axi_in_19_WSTRB,
  m_axi_in_19_WVALID,
  m_axi_in_2_ARADDR,
  m_axi_in_2_ARBURST,
  m_axi_in_2_ARCACHE,
  m_axi_in_2_ARID,
  m_axi_in_2_ARLEN,
  m_axi_in_2_ARLOCK,
  m_axi_in_2_ARPROT,
  m_axi_in_2_ARQOS,
  m_axi_in_2_ARREADY,
  m_axi_in_2_ARSIZE,
  m_axi_in_2_ARVALID,
  m_axi_in_2_AWADDR,
  m_axi_in_2_AWBURST,
  m_axi_in_2_AWCACHE,
  m_axi_in_2_AWID,
  m_axi_in_2_AWLEN,
  m_axi_in_2_AWLOCK,
  m_axi_in_2_AWPROT,
  m_axi_in_2_AWQOS,
  m_axi_in_2_AWREADY,
  m_axi_in_2_AWSIZE,
  m_axi_in_2_AWVALID,
  m_axi_in_2_BID,
  m_axi_in_2_BREADY,
  m_axi_in_2_BRESP,
  m_axi_in_2_BVALID,
  m_axi_in_2_RDATA,
  m_axi_in_2_RID,
  m_axi_in_2_RLAST,
  m_axi_in_2_RREADY,
  m_axi_in_2_RRESP,
  m_axi_in_2_RVALID,
  m_axi_in_2_WDATA,
  m_axi_in_2_WLAST,
  m_axi_in_2_WREADY,
  m_axi_in_2_WSTRB,
  m_axi_in_2_WVALID,
  m_axi_in_20_ARADDR,
  m_axi_in_20_ARBURST,
  m_axi_in_20_ARCACHE,
  m_axi_in_20_ARID,
  m_axi_in_20_ARLEN,
  m_axi_in_20_ARLOCK,
  m_axi_in_20_ARPROT,
  m_axi_in_20_ARQOS,
  m_axi_in_20_ARREADY,
  m_axi_in_20_ARSIZE,
  m_axi_in_20_ARVALID,
  m_axi_in_20_AWADDR,
  m_axi_in_20_AWBURST,
  m_axi_in_20_AWCACHE,
  m_axi_in_20_AWID,
  m_axi_in_20_AWLEN,
  m_axi_in_20_AWLOCK,
  m_axi_in_20_AWPROT,
  m_axi_in_20_AWQOS,
  m_axi_in_20_AWREADY,
  m_axi_in_20_AWSIZE,
  m_axi_in_20_AWVALID,
  m_axi_in_20_BID,
  m_axi_in_20_BREADY,
  m_axi_in_20_BRESP,
  m_axi_in_20_BVALID,
  m_axi_in_20_RDATA,
  m_axi_in_20_RID,
  m_axi_in_20_RLAST,
  m_axi_in_20_RREADY,
  m_axi_in_20_RRESP,
  m_axi_in_20_RVALID,
  m_axi_in_20_WDATA,
  m_axi_in_20_WLAST,
  m_axi_in_20_WREADY,
  m_axi_in_20_WSTRB,
  m_axi_in_20_WVALID,
  m_axi_in_21_ARADDR,
  m_axi_in_21_ARBURST,
  m_axi_in_21_ARCACHE,
  m_axi_in_21_ARID,
  m_axi_in_21_ARLEN,
  m_axi_in_21_ARLOCK,
  m_axi_in_21_ARPROT,
  m_axi_in_21_ARQOS,
  m_axi_in_21_ARREADY,
  m_axi_in_21_ARSIZE,
  m_axi_in_21_ARVALID,
  m_axi_in_21_AWADDR,
  m_axi_in_21_AWBURST,
  m_axi_in_21_AWCACHE,
  m_axi_in_21_AWID,
  m_axi_in_21_AWLEN,
  m_axi_in_21_AWLOCK,
  m_axi_in_21_AWPROT,
  m_axi_in_21_AWQOS,
  m_axi_in_21_AWREADY,
  m_axi_in_21_AWSIZE,
  m_axi_in_21_AWVALID,
  m_axi_in_21_BID,
  m_axi_in_21_BREADY,
  m_axi_in_21_BRESP,
  m_axi_in_21_BVALID,
  m_axi_in_21_RDATA,
  m_axi_in_21_RID,
  m_axi_in_21_RLAST,
  m_axi_in_21_RREADY,
  m_axi_in_21_RRESP,
  m_axi_in_21_RVALID,
  m_axi_in_21_WDATA,
  m_axi_in_21_WLAST,
  m_axi_in_21_WREADY,
  m_axi_in_21_WSTRB,
  m_axi_in_21_WVALID,
  m_axi_in_22_ARADDR,
  m_axi_in_22_ARBURST,
  m_axi_in_22_ARCACHE,
  m_axi_in_22_ARID,
  m_axi_in_22_ARLEN,
  m_axi_in_22_ARLOCK,
  m_axi_in_22_ARPROT,
  m_axi_in_22_ARQOS,
  m_axi_in_22_ARREADY,
  m_axi_in_22_ARSIZE,
  m_axi_in_22_ARVALID,
  m_axi_in_22_AWADDR,
  m_axi_in_22_AWBURST,
  m_axi_in_22_AWCACHE,
  m_axi_in_22_AWID,
  m_axi_in_22_AWLEN,
  m_axi_in_22_AWLOCK,
  m_axi_in_22_AWPROT,
  m_axi_in_22_AWQOS,
  m_axi_in_22_AWREADY,
  m_axi_in_22_AWSIZE,
  m_axi_in_22_AWVALID,
  m_axi_in_22_BID,
  m_axi_in_22_BREADY,
  m_axi_in_22_BRESP,
  m_axi_in_22_BVALID,
  m_axi_in_22_RDATA,
  m_axi_in_22_RID,
  m_axi_in_22_RLAST,
  m_axi_in_22_RREADY,
  m_axi_in_22_RRESP,
  m_axi_in_22_RVALID,
  m_axi_in_22_WDATA,
  m_axi_in_22_WLAST,
  m_axi_in_22_WREADY,
  m_axi_in_22_WSTRB,
  m_axi_in_22_WVALID,
  m_axi_in_23_ARADDR,
  m_axi_in_23_ARBURST,
  m_axi_in_23_ARCACHE,
  m_axi_in_23_ARID,
  m_axi_in_23_ARLEN,
  m_axi_in_23_ARLOCK,
  m_axi_in_23_ARPROT,
  m_axi_in_23_ARQOS,
  m_axi_in_23_ARREADY,
  m_axi_in_23_ARSIZE,
  m_axi_in_23_ARVALID,
  m_axi_in_23_AWADDR,
  m_axi_in_23_AWBURST,
  m_axi_in_23_AWCACHE,
  m_axi_in_23_AWID,
  m_axi_in_23_AWLEN,
  m_axi_in_23_AWLOCK,
  m_axi_in_23_AWPROT,
  m_axi_in_23_AWQOS,
  m_axi_in_23_AWREADY,
  m_axi_in_23_AWSIZE,
  m_axi_in_23_AWVALID,
  m_axi_in_23_BID,
  m_axi_in_23_BREADY,
  m_axi_in_23_BRESP,
  m_axi_in_23_BVALID,
  m_axi_in_23_RDATA,
  m_axi_in_23_RID,
  m_axi_in_23_RLAST,
  m_axi_in_23_RREADY,
  m_axi_in_23_RRESP,
  m_axi_in_23_RVALID,
  m_axi_in_23_WDATA,
  m_axi_in_23_WLAST,
  m_axi_in_23_WREADY,
  m_axi_in_23_WSTRB,
  m_axi_in_23_WVALID,
  m_axi_in_24_ARADDR,
  m_axi_in_24_ARBURST,
  m_axi_in_24_ARCACHE,
  m_axi_in_24_ARID,
  m_axi_in_24_ARLEN,
  m_axi_in_24_ARLOCK,
  m_axi_in_24_ARPROT,
  m_axi_in_24_ARQOS,
  m_axi_in_24_ARREADY,
  m_axi_in_24_ARSIZE,
  m_axi_in_24_ARVALID,
  m_axi_in_24_AWADDR,
  m_axi_in_24_AWBURST,
  m_axi_in_24_AWCACHE,
  m_axi_in_24_AWID,
  m_axi_in_24_AWLEN,
  m_axi_in_24_AWLOCK,
  m_axi_in_24_AWPROT,
  m_axi_in_24_AWQOS,
  m_axi_in_24_AWREADY,
  m_axi_in_24_AWSIZE,
  m_axi_in_24_AWVALID,
  m_axi_in_24_BID,
  m_axi_in_24_BREADY,
  m_axi_in_24_BRESP,
  m_axi_in_24_BVALID,
  m_axi_in_24_RDATA,
  m_axi_in_24_RID,
  m_axi_in_24_RLAST,
  m_axi_in_24_RREADY,
  m_axi_in_24_RRESP,
  m_axi_in_24_RVALID,
  m_axi_in_24_WDATA,
  m_axi_in_24_WLAST,
  m_axi_in_24_WREADY,
  m_axi_in_24_WSTRB,
  m_axi_in_24_WVALID,
  m_axi_in_25_ARADDR,
  m_axi_in_25_ARBURST,
  m_axi_in_25_ARCACHE,
  m_axi_in_25_ARID,
  m_axi_in_25_ARLEN,
  m_axi_in_25_ARLOCK,
  m_axi_in_25_ARPROT,
  m_axi_in_25_ARQOS,
  m_axi_in_25_ARREADY,
  m_axi_in_25_ARSIZE,
  m_axi_in_25_ARVALID,
  m_axi_in_25_AWADDR,
  m_axi_in_25_AWBURST,
  m_axi_in_25_AWCACHE,
  m_axi_in_25_AWID,
  m_axi_in_25_AWLEN,
  m_axi_in_25_AWLOCK,
  m_axi_in_25_AWPROT,
  m_axi_in_25_AWQOS,
  m_axi_in_25_AWREADY,
  m_axi_in_25_AWSIZE,
  m_axi_in_25_AWVALID,
  m_axi_in_25_BID,
  m_axi_in_25_BREADY,
  m_axi_in_25_BRESP,
  m_axi_in_25_BVALID,
  m_axi_in_25_RDATA,
  m_axi_in_25_RID,
  m_axi_in_25_RLAST,
  m_axi_in_25_RREADY,
  m_axi_in_25_RRESP,
  m_axi_in_25_RVALID,
  m_axi_in_25_WDATA,
  m_axi_in_25_WLAST,
  m_axi_in_25_WREADY,
  m_axi_in_25_WSTRB,
  m_axi_in_25_WVALID,
  m_axi_in_26_ARADDR,
  m_axi_in_26_ARBURST,
  m_axi_in_26_ARCACHE,
  m_axi_in_26_ARID,
  m_axi_in_26_ARLEN,
  m_axi_in_26_ARLOCK,
  m_axi_in_26_ARPROT,
  m_axi_in_26_ARQOS,
  m_axi_in_26_ARREADY,
  m_axi_in_26_ARSIZE,
  m_axi_in_26_ARVALID,
  m_axi_in_26_AWADDR,
  m_axi_in_26_AWBURST,
  m_axi_in_26_AWCACHE,
  m_axi_in_26_AWID,
  m_axi_in_26_AWLEN,
  m_axi_in_26_AWLOCK,
  m_axi_in_26_AWPROT,
  m_axi_in_26_AWQOS,
  m_axi_in_26_AWREADY,
  m_axi_in_26_AWSIZE,
  m_axi_in_26_AWVALID,
  m_axi_in_26_BID,
  m_axi_in_26_BREADY,
  m_axi_in_26_BRESP,
  m_axi_in_26_BVALID,
  m_axi_in_26_RDATA,
  m_axi_in_26_RID,
  m_axi_in_26_RLAST,
  m_axi_in_26_RREADY,
  m_axi_in_26_RRESP,
  m_axi_in_26_RVALID,
  m_axi_in_26_WDATA,
  m_axi_in_26_WLAST,
  m_axi_in_26_WREADY,
  m_axi_in_26_WSTRB,
  m_axi_in_26_WVALID,
  m_axi_in_3_ARADDR,
  m_axi_in_3_ARBURST,
  m_axi_in_3_ARCACHE,
  m_axi_in_3_ARID,
  m_axi_in_3_ARLEN,
  m_axi_in_3_ARLOCK,
  m_axi_in_3_ARPROT,
  m_axi_in_3_ARQOS,
  m_axi_in_3_ARREADY,
  m_axi_in_3_ARSIZE,
  m_axi_in_3_ARVALID,
  m_axi_in_3_AWADDR,
  m_axi_in_3_AWBURST,
  m_axi_in_3_AWCACHE,
  m_axi_in_3_AWID,
  m_axi_in_3_AWLEN,
  m_axi_in_3_AWLOCK,
  m_axi_in_3_AWPROT,
  m_axi_in_3_AWQOS,
  m_axi_in_3_AWREADY,
  m_axi_in_3_AWSIZE,
  m_axi_in_3_AWVALID,
  m_axi_in_3_BID,
  m_axi_in_3_BREADY,
  m_axi_in_3_BRESP,
  m_axi_in_3_BVALID,
  m_axi_in_3_RDATA,
  m_axi_in_3_RID,
  m_axi_in_3_RLAST,
  m_axi_in_3_RREADY,
  m_axi_in_3_RRESP,
  m_axi_in_3_RVALID,
  m_axi_in_3_WDATA,
  m_axi_in_3_WLAST,
  m_axi_in_3_WREADY,
  m_axi_in_3_WSTRB,
  m_axi_in_3_WVALID,
  m_axi_in_4_ARADDR,
  m_axi_in_4_ARBURST,
  m_axi_in_4_ARCACHE,
  m_axi_in_4_ARID,
  m_axi_in_4_ARLEN,
  m_axi_in_4_ARLOCK,
  m_axi_in_4_ARPROT,
  m_axi_in_4_ARQOS,
  m_axi_in_4_ARREADY,
  m_axi_in_4_ARSIZE,
  m_axi_in_4_ARVALID,
  m_axi_in_4_AWADDR,
  m_axi_in_4_AWBURST,
  m_axi_in_4_AWCACHE,
  m_axi_in_4_AWID,
  m_axi_in_4_AWLEN,
  m_axi_in_4_AWLOCK,
  m_axi_in_4_AWPROT,
  m_axi_in_4_AWQOS,
  m_axi_in_4_AWREADY,
  m_axi_in_4_AWSIZE,
  m_axi_in_4_AWVALID,
  m_axi_in_4_BID,
  m_axi_in_4_BREADY,
  m_axi_in_4_BRESP,
  m_axi_in_4_BVALID,
  m_axi_in_4_RDATA,
  m_axi_in_4_RID,
  m_axi_in_4_RLAST,
  m_axi_in_4_RREADY,
  m_axi_in_4_RRESP,
  m_axi_in_4_RVALID,
  m_axi_in_4_WDATA,
  m_axi_in_4_WLAST,
  m_axi_in_4_WREADY,
  m_axi_in_4_WSTRB,
  m_axi_in_4_WVALID,
  m_axi_in_5_ARADDR,
  m_axi_in_5_ARBURST,
  m_axi_in_5_ARCACHE,
  m_axi_in_5_ARID,
  m_axi_in_5_ARLEN,
  m_axi_in_5_ARLOCK,
  m_axi_in_5_ARPROT,
  m_axi_in_5_ARQOS,
  m_axi_in_5_ARREADY,
  m_axi_in_5_ARSIZE,
  m_axi_in_5_ARVALID,
  m_axi_in_5_AWADDR,
  m_axi_in_5_AWBURST,
  m_axi_in_5_AWCACHE,
  m_axi_in_5_AWID,
  m_axi_in_5_AWLEN,
  m_axi_in_5_AWLOCK,
  m_axi_in_5_AWPROT,
  m_axi_in_5_AWQOS,
  m_axi_in_5_AWREADY,
  m_axi_in_5_AWSIZE,
  m_axi_in_5_AWVALID,
  m_axi_in_5_BID,
  m_axi_in_5_BREADY,
  m_axi_in_5_BRESP,
  m_axi_in_5_BVALID,
  m_axi_in_5_RDATA,
  m_axi_in_5_RID,
  m_axi_in_5_RLAST,
  m_axi_in_5_RREADY,
  m_axi_in_5_RRESP,
  m_axi_in_5_RVALID,
  m_axi_in_5_WDATA,
  m_axi_in_5_WLAST,
  m_axi_in_5_WREADY,
  m_axi_in_5_WSTRB,
  m_axi_in_5_WVALID,
  m_axi_in_6_ARADDR,
  m_axi_in_6_ARBURST,
  m_axi_in_6_ARCACHE,
  m_axi_in_6_ARID,
  m_axi_in_6_ARLEN,
  m_axi_in_6_ARLOCK,
  m_axi_in_6_ARPROT,
  m_axi_in_6_ARQOS,
  m_axi_in_6_ARREADY,
  m_axi_in_6_ARSIZE,
  m_axi_in_6_ARVALID,
  m_axi_in_6_AWADDR,
  m_axi_in_6_AWBURST,
  m_axi_in_6_AWCACHE,
  m_axi_in_6_AWID,
  m_axi_in_6_AWLEN,
  m_axi_in_6_AWLOCK,
  m_axi_in_6_AWPROT,
  m_axi_in_6_AWQOS,
  m_axi_in_6_AWREADY,
  m_axi_in_6_AWSIZE,
  m_axi_in_6_AWVALID,
  m_axi_in_6_BID,
  m_axi_in_6_BREADY,
  m_axi_in_6_BRESP,
  m_axi_in_6_BVALID,
  m_axi_in_6_RDATA,
  m_axi_in_6_RID,
  m_axi_in_6_RLAST,
  m_axi_in_6_RREADY,
  m_axi_in_6_RRESP,
  m_axi_in_6_RVALID,
  m_axi_in_6_WDATA,
  m_axi_in_6_WLAST,
  m_axi_in_6_WREADY,
  m_axi_in_6_WSTRB,
  m_axi_in_6_WVALID,
  m_axi_in_7_ARADDR,
  m_axi_in_7_ARBURST,
  m_axi_in_7_ARCACHE,
  m_axi_in_7_ARID,
  m_axi_in_7_ARLEN,
  m_axi_in_7_ARLOCK,
  m_axi_in_7_ARPROT,
  m_axi_in_7_ARQOS,
  m_axi_in_7_ARREADY,
  m_axi_in_7_ARSIZE,
  m_axi_in_7_ARVALID,
  m_axi_in_7_AWADDR,
  m_axi_in_7_AWBURST,
  m_axi_in_7_AWCACHE,
  m_axi_in_7_AWID,
  m_axi_in_7_AWLEN,
  m_axi_in_7_AWLOCK,
  m_axi_in_7_AWPROT,
  m_axi_in_7_AWQOS,
  m_axi_in_7_AWREADY,
  m_axi_in_7_AWSIZE,
  m_axi_in_7_AWVALID,
  m_axi_in_7_BID,
  m_axi_in_7_BREADY,
  m_axi_in_7_BRESP,
  m_axi_in_7_BVALID,
  m_axi_in_7_RDATA,
  m_axi_in_7_RID,
  m_axi_in_7_RLAST,
  m_axi_in_7_RREADY,
  m_axi_in_7_RRESP,
  m_axi_in_7_RVALID,
  m_axi_in_7_WDATA,
  m_axi_in_7_WLAST,
  m_axi_in_7_WREADY,
  m_axi_in_7_WSTRB,
  m_axi_in_7_WVALID,
  m_axi_in_8_ARADDR,
  m_axi_in_8_ARBURST,
  m_axi_in_8_ARCACHE,
  m_axi_in_8_ARID,
  m_axi_in_8_ARLEN,
  m_axi_in_8_ARLOCK,
  m_axi_in_8_ARPROT,
  m_axi_in_8_ARQOS,
  m_axi_in_8_ARREADY,
  m_axi_in_8_ARSIZE,
  m_axi_in_8_ARVALID,
  m_axi_in_8_AWADDR,
  m_axi_in_8_AWBURST,
  m_axi_in_8_AWCACHE,
  m_axi_in_8_AWID,
  m_axi_in_8_AWLEN,
  m_axi_in_8_AWLOCK,
  m_axi_in_8_AWPROT,
  m_axi_in_8_AWQOS,
  m_axi_in_8_AWREADY,
  m_axi_in_8_AWSIZE,
  m_axi_in_8_AWVALID,
  m_axi_in_8_BID,
  m_axi_in_8_BREADY,
  m_axi_in_8_BRESP,
  m_axi_in_8_BVALID,
  m_axi_in_8_RDATA,
  m_axi_in_8_RID,
  m_axi_in_8_RLAST,
  m_axi_in_8_RREADY,
  m_axi_in_8_RRESP,
  m_axi_in_8_RVALID,
  m_axi_in_8_WDATA,
  m_axi_in_8_WLAST,
  m_axi_in_8_WREADY,
  m_axi_in_8_WSTRB,
  m_axi_in_8_WVALID,
  m_axi_in_9_ARADDR,
  m_axi_in_9_ARBURST,
  m_axi_in_9_ARCACHE,
  m_axi_in_9_ARID,
  m_axi_in_9_ARLEN,
  m_axi_in_9_ARLOCK,
  m_axi_in_9_ARPROT,
  m_axi_in_9_ARQOS,
  m_axi_in_9_ARREADY,
  m_axi_in_9_ARSIZE,
  m_axi_in_9_ARVALID,
  m_axi_in_9_AWADDR,
  m_axi_in_9_AWBURST,
  m_axi_in_9_AWCACHE,
  m_axi_in_9_AWID,
  m_axi_in_9_AWLEN,
  m_axi_in_9_AWLOCK,
  m_axi_in_9_AWPROT,
  m_axi_in_9_AWQOS,
  m_axi_in_9_AWREADY,
  m_axi_in_9_AWSIZE,
  m_axi_in_9_AWVALID,
  m_axi_in_9_BID,
  m_axi_in_9_BREADY,
  m_axi_in_9_BRESP,
  m_axi_in_9_BVALID,
  m_axi_in_9_RDATA,
  m_axi_in_9_RID,
  m_axi_in_9_RLAST,
  m_axi_in_9_RREADY,
  m_axi_in_9_RRESP,
  m_axi_in_9_RVALID,
  m_axi_in_9_WDATA,
  m_axi_in_9_WLAST,
  m_axi_in_9_WREADY,
  m_axi_in_9_WSTRB,
  m_axi_in_9_WVALID
);

  parameter C_S_AXI_CONTROL_DATA_WIDTH = 32;
  parameter C_S_AXI_CONTROL_ADDR_WIDTH = 9;
  parameter C_S_AXI_DATA_WIDTH = 32;
  parameter C_S_AXI_CONTROL_WSTRB_WIDTH = 32 / 8;
  parameter C_S_AXI_WSTRB_WIDTH = 32 / 8;
  (* RS_HS = "s_axi_control_AW.valid" *)input s_axi_control_AWVALID;
  (* RS_HS = "s_axi_control_AW.ready" *)output s_axi_control_AWREADY;
  (* RS_HS = "s_axi_control_AW.data" *)input [C_S_AXI_CONTROL_ADDR_WIDTH-1:0] s_axi_control_AWADDR;
  (* RS_HS = "s_axi_control_W.valid" *)input s_axi_control_WVALID;
  (* RS_HS = "s_axi_control_W.ready" *)output s_axi_control_WREADY;
  (* RS_HS = "s_axi_control_W.data" *)input [C_S_AXI_CONTROL_DATA_WIDTH-1:0] s_axi_control_WDATA;
  (* RS_HS = "s_axi_control_W.data" *)input [C_S_AXI_CONTROL_WSTRB_WIDTH-1:0] s_axi_control_WSTRB;
  (* RS_HS = "s_axi_control_AR.valid" *)input s_axi_control_ARVALID;
  (* RS_HS = "s_axi_control_AR.ready" *)output s_axi_control_ARREADY;
  (* RS_HS = "s_axi_control_AR.data" *)input [C_S_AXI_CONTROL_ADDR_WIDTH-1:0] s_axi_control_ARADDR;
  (* RS_HS = "s_axi_control_R.valid" *)output s_axi_control_RVALID;
  (* RS_HS = "s_axi_control_R.ready" *)input s_axi_control_RREADY;
  (* RS_HS = "s_axi_control_R.data" *)output [C_S_AXI_CONTROL_DATA_WIDTH-1:0] s_axi_control_RDATA;
  (* RS_HS = "s_axi_control_R.data" *)output [1:0] s_axi_control_RRESP;
  (* RS_HS = "s_axi_control_B.valid" *)output s_axi_control_BVALID;
  (* RS_HS = "s_axi_control_B.ready" *)input s_axi_control_BREADY;
  (* RS_HS = "s_axi_control_B.data" *)output [1:0] s_axi_control_BRESP;
  (* RS_CLK *)input ap_clk;
  (* RS_RST = "ff" *)input ap_rst_n;
  (* RS_FF = "interrupt" *)output interrupt;
  (* RS_HS = "m_axi_L3_out_dist_AR.data" *)output [63:0] m_axi_L3_out_dist_ARADDR;
  (* RS_HS = "m_axi_L3_out_dist_AR.data" *)output [1:0] m_axi_L3_out_dist_ARBURST;
  (* RS_HS = "m_axi_L3_out_dist_AR.data" *)output [3:0] m_axi_L3_out_dist_ARCACHE;
  (* RS_HS = "m_axi_L3_out_dist_AR.data" *)output [0:0] m_axi_L3_out_dist_ARID;
  (* RS_HS = "m_axi_L3_out_dist_AR.data" *)output [7:0] m_axi_L3_out_dist_ARLEN;
  (* RS_HS = "m_axi_L3_out_dist_AR.data" *)output m_axi_L3_out_dist_ARLOCK;
  (* RS_HS = "m_axi_L3_out_dist_AR.data" *)output [2:0] m_axi_L3_out_dist_ARPROT;
  (* RS_HS = "m_axi_L3_out_dist_AR.data" *)output [3:0] m_axi_L3_out_dist_ARQOS;
  (* RS_HS = "m_axi_L3_out_dist_AR.ready" *)input m_axi_L3_out_dist_ARREADY;
  (* RS_HS = "m_axi_L3_out_dist_AR.data" *)output [2:0] m_axi_L3_out_dist_ARSIZE;
  (* RS_HS = "m_axi_L3_out_dist_AR.valid" *)output m_axi_L3_out_dist_ARVALID;
  (* RS_HS = "m_axi_L3_out_dist_AW.data" *)output [63:0] m_axi_L3_out_dist_AWADDR;
  (* RS_HS = "m_axi_L3_out_dist_AW.data" *)output [1:0] m_axi_L3_out_dist_AWBURST;
  (* RS_HS = "m_axi_L3_out_dist_AW.data" *)output [3:0] m_axi_L3_out_dist_AWCACHE;
  (* RS_HS = "m_axi_L3_out_dist_AW.data" *)output [0:0] m_axi_L3_out_dist_AWID;
  (* RS_HS = "m_axi_L3_out_dist_AW.data" *)output [7:0] m_axi_L3_out_dist_AWLEN;
  (* RS_HS = "m_axi_L3_out_dist_AW.data" *)output m_axi_L3_out_dist_AWLOCK;
  (* RS_HS = "m_axi_L3_out_dist_AW.data" *)output [2:0] m_axi_L3_out_dist_AWPROT;
  (* RS_HS = "m_axi_L3_out_dist_AW.data" *)output [3:0] m_axi_L3_out_dist_AWQOS;
  (* RS_HS = "m_axi_L3_out_dist_AW.ready" *)input m_axi_L3_out_dist_AWREADY;
  (* RS_HS = "m_axi_L3_out_dist_AW.data" *)output [2:0] m_axi_L3_out_dist_AWSIZE;
  (* RS_HS = "m_axi_L3_out_dist_AW.valid" *)output m_axi_L3_out_dist_AWVALID;
  (* RS_HS = "m_axi_L3_out_dist_B.data" *)input [0:0] m_axi_L3_out_dist_BID;
  (* RS_HS = "m_axi_L3_out_dist_B.ready" *)output m_axi_L3_out_dist_BREADY;
  (* RS_HS = "m_axi_L3_out_dist_B.data" *)input [1:0] m_axi_L3_out_dist_BRESP;
  (* RS_HS = "m_axi_L3_out_dist_B.valid" *)input m_axi_L3_out_dist_BVALID;
  (* RS_HS = "m_axi_L3_out_dist_R.data" *)input [31:0] m_axi_L3_out_dist_RDATA;
  (* RS_HS = "m_axi_L3_out_dist_R.data" *)input [0:0] m_axi_L3_out_dist_RID;
  (* RS_HS = "m_axi_L3_out_dist_R.data" *)input m_axi_L3_out_dist_RLAST;
  (* RS_HS = "m_axi_L3_out_dist_R.ready" *)output m_axi_L3_out_dist_RREADY;
  (* RS_HS = "m_axi_L3_out_dist_R.data" *)input [1:0] m_axi_L3_out_dist_RRESP;
  (* RS_HS = "m_axi_L3_out_dist_R.valid" *)input m_axi_L3_out_dist_RVALID;
  (* RS_HS = "m_axi_L3_out_dist_W.data" *)output [31:0] m_axi_L3_out_dist_WDATA;
  (* RS_HS = "m_axi_L3_out_dist_W.data" *)output m_axi_L3_out_dist_WLAST;
  (* RS_HS = "m_axi_L3_out_dist_W.ready" *)input m_axi_L3_out_dist_WREADY;
  (* RS_HS = "m_axi_L3_out_dist_W.data" *)output [3:0] m_axi_L3_out_dist_WSTRB;
  (* RS_HS = "m_axi_L3_out_dist_W.valid" *)output m_axi_L3_out_dist_WVALID;
  (* RS_HS = "m_axi_L3_out_id_AR.data" *)output [63:0] m_axi_L3_out_id_ARADDR;
  (* RS_HS = "m_axi_L3_out_id_AR.data" *)output [1:0] m_axi_L3_out_id_ARBURST;
  (* RS_HS = "m_axi_L3_out_id_AR.data" *)output [3:0] m_axi_L3_out_id_ARCACHE;
  (* RS_HS = "m_axi_L3_out_id_AR.data" *)output [0:0] m_axi_L3_out_id_ARID;
  (* RS_HS = "m_axi_L3_out_id_AR.data" *)output [7:0] m_axi_L3_out_id_ARLEN;
  (* RS_HS = "m_axi_L3_out_id_AR.data" *)output m_axi_L3_out_id_ARLOCK;
  (* RS_HS = "m_axi_L3_out_id_AR.data" *)output [2:0] m_axi_L3_out_id_ARPROT;
  (* RS_HS = "m_axi_L3_out_id_AR.data" *)output [3:0] m_axi_L3_out_id_ARQOS;
  (* RS_HS = "m_axi_L3_out_id_AR.ready" *)input m_axi_L3_out_id_ARREADY;
  (* RS_HS = "m_axi_L3_out_id_AR.data" *)output [2:0] m_axi_L3_out_id_ARSIZE;
  (* RS_HS = "m_axi_L3_out_id_AR.valid" *)output m_axi_L3_out_id_ARVALID;
  (* RS_HS = "m_axi_L3_out_id_AW.data" *)output [63:0] m_axi_L3_out_id_AWADDR;
  (* RS_HS = "m_axi_L3_out_id_AW.data" *)output [1:0] m_axi_L3_out_id_AWBURST;
  (* RS_HS = "m_axi_L3_out_id_AW.data" *)output [3:0] m_axi_L3_out_id_AWCACHE;
  (* RS_HS = "m_axi_L3_out_id_AW.data" *)output [0:0] m_axi_L3_out_id_AWID;
  (* RS_HS = "m_axi_L3_out_id_AW.data" *)output [7:0] m_axi_L3_out_id_AWLEN;
  (* RS_HS = "m_axi_L3_out_id_AW.data" *)output m_axi_L3_out_id_AWLOCK;
  (* RS_HS = "m_axi_L3_out_id_AW.data" *)output [2:0] m_axi_L3_out_id_AWPROT;
  (* RS_HS = "m_axi_L3_out_id_AW.data" *)output [3:0] m_axi_L3_out_id_AWQOS;
  (* RS_HS = "m_axi_L3_out_id_AW.ready" *)input m_axi_L3_out_id_AWREADY;
  (* RS_HS = "m_axi_L3_out_id_AW.data" *)output [2:0] m_axi_L3_out_id_AWSIZE;
  (* RS_HS = "m_axi_L3_out_id_AW.valid" *)output m_axi_L3_out_id_AWVALID;
  (* RS_HS = "m_axi_L3_out_id_B.data" *)input [0:0] m_axi_L3_out_id_BID;
  (* RS_HS = "m_axi_L3_out_id_B.ready" *)output m_axi_L3_out_id_BREADY;
  (* RS_HS = "m_axi_L3_out_id_B.data" *)input [1:0] m_axi_L3_out_id_BRESP;
  (* RS_HS = "m_axi_L3_out_id_B.valid" *)input m_axi_L3_out_id_BVALID;
  (* RS_HS = "m_axi_L3_out_id_R.data" *)input [31:0] m_axi_L3_out_id_RDATA;
  (* RS_HS = "m_axi_L3_out_id_R.data" *)input [0:0] m_axi_L3_out_id_RID;
  (* RS_HS = "m_axi_L3_out_id_R.data" *)input m_axi_L3_out_id_RLAST;
  (* RS_HS = "m_axi_L3_out_id_R.ready" *)output m_axi_L3_out_id_RREADY;
  (* RS_HS = "m_axi_L3_out_id_R.data" *)input [1:0] m_axi_L3_out_id_RRESP;
  (* RS_HS = "m_axi_L3_out_id_R.valid" *)input m_axi_L3_out_id_RVALID;
  (* RS_HS = "m_axi_L3_out_id_W.data" *)output [31:0] m_axi_L3_out_id_WDATA;
  (* RS_HS = "m_axi_L3_out_id_W.data" *)output m_axi_L3_out_id_WLAST;
  (* RS_HS = "m_axi_L3_out_id_W.ready" *)input m_axi_L3_out_id_WREADY;
  (* RS_HS = "m_axi_L3_out_id_W.data" *)output [3:0] m_axi_L3_out_id_WSTRB;
  (* RS_HS = "m_axi_L3_out_id_W.valid" *)output m_axi_L3_out_id_WVALID;
  (* RS_HS = "m_axi_in_0_AR.data" *)output [63:0] m_axi_in_0_ARADDR;
  (* RS_HS = "m_axi_in_0_AR.data" *)output [1:0] m_axi_in_0_ARBURST;
  (* RS_HS = "m_axi_in_0_AR.data" *)output [3:0] m_axi_in_0_ARCACHE;
  (* RS_HS = "m_axi_in_0_AR.data" *)output [0:0] m_axi_in_0_ARID;
  (* RS_HS = "m_axi_in_0_AR.data" *)output [7:0] m_axi_in_0_ARLEN;
  (* RS_HS = "m_axi_in_0_AR.data" *)output m_axi_in_0_ARLOCK;
  (* RS_HS = "m_axi_in_0_AR.data" *)output [2:0] m_axi_in_0_ARPROT;
  (* RS_HS = "m_axi_in_0_AR.data" *)output [3:0] m_axi_in_0_ARQOS;
  (* RS_HS = "m_axi_in_0_AR.ready" *)input m_axi_in_0_ARREADY;
  (* RS_HS = "m_axi_in_0_AR.data" *)output [2:0] m_axi_in_0_ARSIZE;
  (* RS_HS = "m_axi_in_0_AR.valid" *)output m_axi_in_0_ARVALID;
  (* RS_HS = "m_axi_in_0_AW.data" *)output [63:0] m_axi_in_0_AWADDR;
  (* RS_HS = "m_axi_in_0_AW.data" *)output [1:0] m_axi_in_0_AWBURST;
  (* RS_HS = "m_axi_in_0_AW.data" *)output [3:0] m_axi_in_0_AWCACHE;
  (* RS_HS = "m_axi_in_0_AW.data" *)output [0:0] m_axi_in_0_AWID;
  (* RS_HS = "m_axi_in_0_AW.data" *)output [7:0] m_axi_in_0_AWLEN;
  (* RS_HS = "m_axi_in_0_AW.data" *)output m_axi_in_0_AWLOCK;
  (* RS_HS = "m_axi_in_0_AW.data" *)output [2:0] m_axi_in_0_AWPROT;
  (* RS_HS = "m_axi_in_0_AW.data" *)output [3:0] m_axi_in_0_AWQOS;
  (* RS_HS = "m_axi_in_0_AW.ready" *)input m_axi_in_0_AWREADY;
  (* RS_HS = "m_axi_in_0_AW.data" *)output [2:0] m_axi_in_0_AWSIZE;
  (* RS_HS = "m_axi_in_0_AW.valid" *)output m_axi_in_0_AWVALID;
  (* RS_HS = "m_axi_in_0_B.data" *)input [0:0] m_axi_in_0_BID;
  (* RS_HS = "m_axi_in_0_B.ready" *)output m_axi_in_0_BREADY;
  (* RS_HS = "m_axi_in_0_B.data" *)input [1:0] m_axi_in_0_BRESP;
  (* RS_HS = "m_axi_in_0_B.valid" *)input m_axi_in_0_BVALID;
  (* RS_HS = "m_axi_in_0_R.data" *)input [255:0] m_axi_in_0_RDATA;
  (* RS_HS = "m_axi_in_0_R.data" *)input [0:0] m_axi_in_0_RID;
  (* RS_HS = "m_axi_in_0_R.data" *)input m_axi_in_0_RLAST;
  (* RS_HS = "m_axi_in_0_R.ready" *)output m_axi_in_0_RREADY;
  (* RS_HS = "m_axi_in_0_R.data" *)input [1:0] m_axi_in_0_RRESP;
  (* RS_HS = "m_axi_in_0_R.valid" *)input m_axi_in_0_RVALID;
  (* RS_HS = "m_axi_in_0_W.data" *)output [255:0] m_axi_in_0_WDATA;
  (* RS_HS = "m_axi_in_0_W.data" *)output m_axi_in_0_WLAST;
  (* RS_HS = "m_axi_in_0_W.ready" *)input m_axi_in_0_WREADY;
  (* RS_HS = "m_axi_in_0_W.data" *)output [31:0] m_axi_in_0_WSTRB;
  (* RS_HS = "m_axi_in_0_W.valid" *)output m_axi_in_0_WVALID;
  (* RS_HS = "m_axi_in_1_AR.data" *)output [63:0] m_axi_in_1_ARADDR;
  (* RS_HS = "m_axi_in_1_AR.data" *)output [1:0] m_axi_in_1_ARBURST;
  (* RS_HS = "m_axi_in_1_AR.data" *)output [3:0] m_axi_in_1_ARCACHE;
  (* RS_HS = "m_axi_in_1_AR.data" *)output [0:0] m_axi_in_1_ARID;
  (* RS_HS = "m_axi_in_1_AR.data" *)output [7:0] m_axi_in_1_ARLEN;
  (* RS_HS = "m_axi_in_1_AR.data" *)output m_axi_in_1_ARLOCK;
  (* RS_HS = "m_axi_in_1_AR.data" *)output [2:0] m_axi_in_1_ARPROT;
  (* RS_HS = "m_axi_in_1_AR.data" *)output [3:0] m_axi_in_1_ARQOS;
  (* RS_HS = "m_axi_in_1_AR.ready" *)input m_axi_in_1_ARREADY;
  (* RS_HS = "m_axi_in_1_AR.data" *)output [2:0] m_axi_in_1_ARSIZE;
  (* RS_HS = "m_axi_in_1_AR.valid" *)output m_axi_in_1_ARVALID;
  (* RS_HS = "m_axi_in_1_AW.data" *)output [63:0] m_axi_in_1_AWADDR;
  (* RS_HS = "m_axi_in_1_AW.data" *)output [1:0] m_axi_in_1_AWBURST;
  (* RS_HS = "m_axi_in_1_AW.data" *)output [3:0] m_axi_in_1_AWCACHE;
  (* RS_HS = "m_axi_in_1_AW.data" *)output [0:0] m_axi_in_1_AWID;
  (* RS_HS = "m_axi_in_1_AW.data" *)output [7:0] m_axi_in_1_AWLEN;
  (* RS_HS = "m_axi_in_1_AW.data" *)output m_axi_in_1_AWLOCK;
  (* RS_HS = "m_axi_in_1_AW.data" *)output [2:0] m_axi_in_1_AWPROT;
  (* RS_HS = "m_axi_in_1_AW.data" *)output [3:0] m_axi_in_1_AWQOS;
  (* RS_HS = "m_axi_in_1_AW.ready" *)input m_axi_in_1_AWREADY;
  (* RS_HS = "m_axi_in_1_AW.data" *)output [2:0] m_axi_in_1_AWSIZE;
  (* RS_HS = "m_axi_in_1_AW.valid" *)output m_axi_in_1_AWVALID;
  (* RS_HS = "m_axi_in_1_B.data" *)input [0:0] m_axi_in_1_BID;
  (* RS_HS = "m_axi_in_1_B.ready" *)output m_axi_in_1_BREADY;
  (* RS_HS = "m_axi_in_1_B.data" *)input [1:0] m_axi_in_1_BRESP;
  (* RS_HS = "m_axi_in_1_B.valid" *)input m_axi_in_1_BVALID;
  (* RS_HS = "m_axi_in_1_R.data" *)input [255:0] m_axi_in_1_RDATA;
  (* RS_HS = "m_axi_in_1_R.data" *)input [0:0] m_axi_in_1_RID;
  (* RS_HS = "m_axi_in_1_R.data" *)input m_axi_in_1_RLAST;
  (* RS_HS = "m_axi_in_1_R.ready" *)output m_axi_in_1_RREADY;
  (* RS_HS = "m_axi_in_1_R.data" *)input [1:0] m_axi_in_1_RRESP;
  (* RS_HS = "m_axi_in_1_R.valid" *)input m_axi_in_1_RVALID;
  (* RS_HS = "m_axi_in_1_W.data" *)output [255:0] m_axi_in_1_WDATA;
  (* RS_HS = "m_axi_in_1_W.data" *)output m_axi_in_1_WLAST;
  (* RS_HS = "m_axi_in_1_W.ready" *)input m_axi_in_1_WREADY;
  (* RS_HS = "m_axi_in_1_W.data" *)output [31:0] m_axi_in_1_WSTRB;
  (* RS_HS = "m_axi_in_1_W.valid" *)output m_axi_in_1_WVALID;
  (* RS_HS = "m_axi_in_10_AR.data" *)output [63:0] m_axi_in_10_ARADDR;
  (* RS_HS = "m_axi_in_10_AR.data" *)output [1:0] m_axi_in_10_ARBURST;
  (* RS_HS = "m_axi_in_10_AR.data" *)output [3:0] m_axi_in_10_ARCACHE;
  (* RS_HS = "m_axi_in_10_AR.data" *)output [0:0] m_axi_in_10_ARID;
  (* RS_HS = "m_axi_in_10_AR.data" *)output [7:0] m_axi_in_10_ARLEN;
  (* RS_HS = "m_axi_in_10_AR.data" *)output m_axi_in_10_ARLOCK;
  (* RS_HS = "m_axi_in_10_AR.data" *)output [2:0] m_axi_in_10_ARPROT;
  (* RS_HS = "m_axi_in_10_AR.data" *)output [3:0] m_axi_in_10_ARQOS;
  (* RS_HS = "m_axi_in_10_AR.ready" *)input m_axi_in_10_ARREADY;
  (* RS_HS = "m_axi_in_10_AR.data" *)output [2:0] m_axi_in_10_ARSIZE;
  (* RS_HS = "m_axi_in_10_AR.valid" *)output m_axi_in_10_ARVALID;
  (* RS_HS = "m_axi_in_10_AW.data" *)output [63:0] m_axi_in_10_AWADDR;
  (* RS_HS = "m_axi_in_10_AW.data" *)output [1:0] m_axi_in_10_AWBURST;
  (* RS_HS = "m_axi_in_10_AW.data" *)output [3:0] m_axi_in_10_AWCACHE;
  (* RS_HS = "m_axi_in_10_AW.data" *)output [0:0] m_axi_in_10_AWID;
  (* RS_HS = "m_axi_in_10_AW.data" *)output [7:0] m_axi_in_10_AWLEN;
  (* RS_HS = "m_axi_in_10_AW.data" *)output m_axi_in_10_AWLOCK;
  (* RS_HS = "m_axi_in_10_AW.data" *)output [2:0] m_axi_in_10_AWPROT;
  (* RS_HS = "m_axi_in_10_AW.data" *)output [3:0] m_axi_in_10_AWQOS;
  (* RS_HS = "m_axi_in_10_AW.ready" *)input m_axi_in_10_AWREADY;
  (* RS_HS = "m_axi_in_10_AW.data" *)output [2:0] m_axi_in_10_AWSIZE;
  (* RS_HS = "m_axi_in_10_AW.valid" *)output m_axi_in_10_AWVALID;
  (* RS_HS = "m_axi_in_10_B.data" *)input [0:0] m_axi_in_10_BID;
  (* RS_HS = "m_axi_in_10_B.ready" *)output m_axi_in_10_BREADY;
  (* RS_HS = "m_axi_in_10_B.data" *)input [1:0] m_axi_in_10_BRESP;
  (* RS_HS = "m_axi_in_10_B.valid" *)input m_axi_in_10_BVALID;
  (* RS_HS = "m_axi_in_10_R.data" *)input [255:0] m_axi_in_10_RDATA;
  (* RS_HS = "m_axi_in_10_R.data" *)input [0:0] m_axi_in_10_RID;
  (* RS_HS = "m_axi_in_10_R.data" *)input m_axi_in_10_RLAST;
  (* RS_HS = "m_axi_in_10_R.ready" *)output m_axi_in_10_RREADY;
  (* RS_HS = "m_axi_in_10_R.data" *)input [1:0] m_axi_in_10_RRESP;
  (* RS_HS = "m_axi_in_10_R.valid" *)input m_axi_in_10_RVALID;
  (* RS_HS = "m_axi_in_10_W.data" *)output [255:0] m_axi_in_10_WDATA;
  (* RS_HS = "m_axi_in_10_W.data" *)output m_axi_in_10_WLAST;
  (* RS_HS = "m_axi_in_10_W.ready" *)input m_axi_in_10_WREADY;
  (* RS_HS = "m_axi_in_10_W.data" *)output [31:0] m_axi_in_10_WSTRB;
  (* RS_HS = "m_axi_in_10_W.valid" *)output m_axi_in_10_WVALID;
  (* RS_HS = "m_axi_in_11_AR.data" *)output [63:0] m_axi_in_11_ARADDR;
  (* RS_HS = "m_axi_in_11_AR.data" *)output [1:0] m_axi_in_11_ARBURST;
  (* RS_HS = "m_axi_in_11_AR.data" *)output [3:0] m_axi_in_11_ARCACHE;
  (* RS_HS = "m_axi_in_11_AR.data" *)output [0:0] m_axi_in_11_ARID;
  (* RS_HS = "m_axi_in_11_AR.data" *)output [7:0] m_axi_in_11_ARLEN;
  (* RS_HS = "m_axi_in_11_AR.data" *)output m_axi_in_11_ARLOCK;
  (* RS_HS = "m_axi_in_11_AR.data" *)output [2:0] m_axi_in_11_ARPROT;
  (* RS_HS = "m_axi_in_11_AR.data" *)output [3:0] m_axi_in_11_ARQOS;
  (* RS_HS = "m_axi_in_11_AR.ready" *)input m_axi_in_11_ARREADY;
  (* RS_HS = "m_axi_in_11_AR.data" *)output [2:0] m_axi_in_11_ARSIZE;
  (* RS_HS = "m_axi_in_11_AR.valid" *)output m_axi_in_11_ARVALID;
  (* RS_HS = "m_axi_in_11_AW.data" *)output [63:0] m_axi_in_11_AWADDR;
  (* RS_HS = "m_axi_in_11_AW.data" *)output [1:0] m_axi_in_11_AWBURST;
  (* RS_HS = "m_axi_in_11_AW.data" *)output [3:0] m_axi_in_11_AWCACHE;
  (* RS_HS = "m_axi_in_11_AW.data" *)output [0:0] m_axi_in_11_AWID;
  (* RS_HS = "m_axi_in_11_AW.data" *)output [7:0] m_axi_in_11_AWLEN;
  (* RS_HS = "m_axi_in_11_AW.data" *)output m_axi_in_11_AWLOCK;
  (* RS_HS = "m_axi_in_11_AW.data" *)output [2:0] m_axi_in_11_AWPROT;
  (* RS_HS = "m_axi_in_11_AW.data" *)output [3:0] m_axi_in_11_AWQOS;
  (* RS_HS = "m_axi_in_11_AW.ready" *)input m_axi_in_11_AWREADY;
  (* RS_HS = "m_axi_in_11_AW.data" *)output [2:0] m_axi_in_11_AWSIZE;
  (* RS_HS = "m_axi_in_11_AW.valid" *)output m_axi_in_11_AWVALID;
  (* RS_HS = "m_axi_in_11_B.data" *)input [0:0] m_axi_in_11_BID;
  (* RS_HS = "m_axi_in_11_B.ready" *)output m_axi_in_11_BREADY;
  (* RS_HS = "m_axi_in_11_B.data" *)input [1:0] m_axi_in_11_BRESP;
  (* RS_HS = "m_axi_in_11_B.valid" *)input m_axi_in_11_BVALID;
  (* RS_HS = "m_axi_in_11_R.data" *)input [255:0] m_axi_in_11_RDATA;
  (* RS_HS = "m_axi_in_11_R.data" *)input [0:0] m_axi_in_11_RID;
  (* RS_HS = "m_axi_in_11_R.data" *)input m_axi_in_11_RLAST;
  (* RS_HS = "m_axi_in_11_R.ready" *)output m_axi_in_11_RREADY;
  (* RS_HS = "m_axi_in_11_R.data" *)input [1:0] m_axi_in_11_RRESP;
  (* RS_HS = "m_axi_in_11_R.valid" *)input m_axi_in_11_RVALID;
  (* RS_HS = "m_axi_in_11_W.data" *)output [255:0] m_axi_in_11_WDATA;
  (* RS_HS = "m_axi_in_11_W.data" *)output m_axi_in_11_WLAST;
  (* RS_HS = "m_axi_in_11_W.ready" *)input m_axi_in_11_WREADY;
  (* RS_HS = "m_axi_in_11_W.data" *)output [31:0] m_axi_in_11_WSTRB;
  (* RS_HS = "m_axi_in_11_W.valid" *)output m_axi_in_11_WVALID;
  (* RS_HS = "m_axi_in_12_AR.data" *)output [63:0] m_axi_in_12_ARADDR;
  (* RS_HS = "m_axi_in_12_AR.data" *)output [1:0] m_axi_in_12_ARBURST;
  (* RS_HS = "m_axi_in_12_AR.data" *)output [3:0] m_axi_in_12_ARCACHE;
  (* RS_HS = "m_axi_in_12_AR.data" *)output [0:0] m_axi_in_12_ARID;
  (* RS_HS = "m_axi_in_12_AR.data" *)output [7:0] m_axi_in_12_ARLEN;
  (* RS_HS = "m_axi_in_12_AR.data" *)output m_axi_in_12_ARLOCK;
  (* RS_HS = "m_axi_in_12_AR.data" *)output [2:0] m_axi_in_12_ARPROT;
  (* RS_HS = "m_axi_in_12_AR.data" *)output [3:0] m_axi_in_12_ARQOS;
  (* RS_HS = "m_axi_in_12_AR.ready" *)input m_axi_in_12_ARREADY;
  (* RS_HS = "m_axi_in_12_AR.data" *)output [2:0] m_axi_in_12_ARSIZE;
  (* RS_HS = "m_axi_in_12_AR.valid" *)output m_axi_in_12_ARVALID;
  (* RS_HS = "m_axi_in_12_AW.data" *)output [63:0] m_axi_in_12_AWADDR;
  (* RS_HS = "m_axi_in_12_AW.data" *)output [1:0] m_axi_in_12_AWBURST;
  (* RS_HS = "m_axi_in_12_AW.data" *)output [3:0] m_axi_in_12_AWCACHE;
  (* RS_HS = "m_axi_in_12_AW.data" *)output [0:0] m_axi_in_12_AWID;
  (* RS_HS = "m_axi_in_12_AW.data" *)output [7:0] m_axi_in_12_AWLEN;
  (* RS_HS = "m_axi_in_12_AW.data" *)output m_axi_in_12_AWLOCK;
  (* RS_HS = "m_axi_in_12_AW.data" *)output [2:0] m_axi_in_12_AWPROT;
  (* RS_HS = "m_axi_in_12_AW.data" *)output [3:0] m_axi_in_12_AWQOS;
  (* RS_HS = "m_axi_in_12_AW.ready" *)input m_axi_in_12_AWREADY;
  (* RS_HS = "m_axi_in_12_AW.data" *)output [2:0] m_axi_in_12_AWSIZE;
  (* RS_HS = "m_axi_in_12_AW.valid" *)output m_axi_in_12_AWVALID;
  (* RS_HS = "m_axi_in_12_B.data" *)input [0:0] m_axi_in_12_BID;
  (* RS_HS = "m_axi_in_12_B.ready" *)output m_axi_in_12_BREADY;
  (* RS_HS = "m_axi_in_12_B.data" *)input [1:0] m_axi_in_12_BRESP;
  (* RS_HS = "m_axi_in_12_B.valid" *)input m_axi_in_12_BVALID;
  (* RS_HS = "m_axi_in_12_R.data" *)input [255:0] m_axi_in_12_RDATA;
  (* RS_HS = "m_axi_in_12_R.data" *)input [0:0] m_axi_in_12_RID;
  (* RS_HS = "m_axi_in_12_R.data" *)input m_axi_in_12_RLAST;
  (* RS_HS = "m_axi_in_12_R.ready" *)output m_axi_in_12_RREADY;
  (* RS_HS = "m_axi_in_12_R.data" *)input [1:0] m_axi_in_12_RRESP;
  (* RS_HS = "m_axi_in_12_R.valid" *)input m_axi_in_12_RVALID;
  (* RS_HS = "m_axi_in_12_W.data" *)output [255:0] m_axi_in_12_WDATA;
  (* RS_HS = "m_axi_in_12_W.data" *)output m_axi_in_12_WLAST;
  (* RS_HS = "m_axi_in_12_W.ready" *)input m_axi_in_12_WREADY;
  (* RS_HS = "m_axi_in_12_W.data" *)output [31:0] m_axi_in_12_WSTRB;
  (* RS_HS = "m_axi_in_12_W.valid" *)output m_axi_in_12_WVALID;
  (* RS_HS = "m_axi_in_13_AR.data" *)output [63:0] m_axi_in_13_ARADDR;
  (* RS_HS = "m_axi_in_13_AR.data" *)output [1:0] m_axi_in_13_ARBURST;
  (* RS_HS = "m_axi_in_13_AR.data" *)output [3:0] m_axi_in_13_ARCACHE;
  (* RS_HS = "m_axi_in_13_AR.data" *)output [0:0] m_axi_in_13_ARID;
  (* RS_HS = "m_axi_in_13_AR.data" *)output [7:0] m_axi_in_13_ARLEN;
  (* RS_HS = "m_axi_in_13_AR.data" *)output m_axi_in_13_ARLOCK;
  (* RS_HS = "m_axi_in_13_AR.data" *)output [2:0] m_axi_in_13_ARPROT;
  (* RS_HS = "m_axi_in_13_AR.data" *)output [3:0] m_axi_in_13_ARQOS;
  (* RS_HS = "m_axi_in_13_AR.ready" *)input m_axi_in_13_ARREADY;
  (* RS_HS = "m_axi_in_13_AR.data" *)output [2:0] m_axi_in_13_ARSIZE;
  (* RS_HS = "m_axi_in_13_AR.valid" *)output m_axi_in_13_ARVALID;
  (* RS_HS = "m_axi_in_13_AW.data" *)output [63:0] m_axi_in_13_AWADDR;
  (* RS_HS = "m_axi_in_13_AW.data" *)output [1:0] m_axi_in_13_AWBURST;
  (* RS_HS = "m_axi_in_13_AW.data" *)output [3:0] m_axi_in_13_AWCACHE;
  (* RS_HS = "m_axi_in_13_AW.data" *)output [0:0] m_axi_in_13_AWID;
  (* RS_HS = "m_axi_in_13_AW.data" *)output [7:0] m_axi_in_13_AWLEN;
  (* RS_HS = "m_axi_in_13_AW.data" *)output m_axi_in_13_AWLOCK;
  (* RS_HS = "m_axi_in_13_AW.data" *)output [2:0] m_axi_in_13_AWPROT;
  (* RS_HS = "m_axi_in_13_AW.data" *)output [3:0] m_axi_in_13_AWQOS;
  (* RS_HS = "m_axi_in_13_AW.ready" *)input m_axi_in_13_AWREADY;
  (* RS_HS = "m_axi_in_13_AW.data" *)output [2:0] m_axi_in_13_AWSIZE;
  (* RS_HS = "m_axi_in_13_AW.valid" *)output m_axi_in_13_AWVALID;
  (* RS_HS = "m_axi_in_13_B.data" *)input [0:0] m_axi_in_13_BID;
  (* RS_HS = "m_axi_in_13_B.ready" *)output m_axi_in_13_BREADY;
  (* RS_HS = "m_axi_in_13_B.data" *)input [1:0] m_axi_in_13_BRESP;
  (* RS_HS = "m_axi_in_13_B.valid" *)input m_axi_in_13_BVALID;
  (* RS_HS = "m_axi_in_13_R.data" *)input [255:0] m_axi_in_13_RDATA;
  (* RS_HS = "m_axi_in_13_R.data" *)input [0:0] m_axi_in_13_RID;
  (* RS_HS = "m_axi_in_13_R.data" *)input m_axi_in_13_RLAST;
  (* RS_HS = "m_axi_in_13_R.ready" *)output m_axi_in_13_RREADY;
  (* RS_HS = "m_axi_in_13_R.data" *)input [1:0] m_axi_in_13_RRESP;
  (* RS_HS = "m_axi_in_13_R.valid" *)input m_axi_in_13_RVALID;
  (* RS_HS = "m_axi_in_13_W.data" *)output [255:0] m_axi_in_13_WDATA;
  (* RS_HS = "m_axi_in_13_W.data" *)output m_axi_in_13_WLAST;
  (* RS_HS = "m_axi_in_13_W.ready" *)input m_axi_in_13_WREADY;
  (* RS_HS = "m_axi_in_13_W.data" *)output [31:0] m_axi_in_13_WSTRB;
  (* RS_HS = "m_axi_in_13_W.valid" *)output m_axi_in_13_WVALID;
  (* RS_HS = "m_axi_in_14_AR.data" *)output [63:0] m_axi_in_14_ARADDR;
  (* RS_HS = "m_axi_in_14_AR.data" *)output [1:0] m_axi_in_14_ARBURST;
  (* RS_HS = "m_axi_in_14_AR.data" *)output [3:0] m_axi_in_14_ARCACHE;
  (* RS_HS = "m_axi_in_14_AR.data" *)output [0:0] m_axi_in_14_ARID;
  (* RS_HS = "m_axi_in_14_AR.data" *)output [7:0] m_axi_in_14_ARLEN;
  (* RS_HS = "m_axi_in_14_AR.data" *)output m_axi_in_14_ARLOCK;
  (* RS_HS = "m_axi_in_14_AR.data" *)output [2:0] m_axi_in_14_ARPROT;
  (* RS_HS = "m_axi_in_14_AR.data" *)output [3:0] m_axi_in_14_ARQOS;
  (* RS_HS = "m_axi_in_14_AR.ready" *)input m_axi_in_14_ARREADY;
  (* RS_HS = "m_axi_in_14_AR.data" *)output [2:0] m_axi_in_14_ARSIZE;
  (* RS_HS = "m_axi_in_14_AR.valid" *)output m_axi_in_14_ARVALID;
  (* RS_HS = "m_axi_in_14_AW.data" *)output [63:0] m_axi_in_14_AWADDR;
  (* RS_HS = "m_axi_in_14_AW.data" *)output [1:0] m_axi_in_14_AWBURST;
  (* RS_HS = "m_axi_in_14_AW.data" *)output [3:0] m_axi_in_14_AWCACHE;
  (* RS_HS = "m_axi_in_14_AW.data" *)output [0:0] m_axi_in_14_AWID;
  (* RS_HS = "m_axi_in_14_AW.data" *)output [7:0] m_axi_in_14_AWLEN;
  (* RS_HS = "m_axi_in_14_AW.data" *)output m_axi_in_14_AWLOCK;
  (* RS_HS = "m_axi_in_14_AW.data" *)output [2:0] m_axi_in_14_AWPROT;
  (* RS_HS = "m_axi_in_14_AW.data" *)output [3:0] m_axi_in_14_AWQOS;
  (* RS_HS = "m_axi_in_14_AW.ready" *)input m_axi_in_14_AWREADY;
  (* RS_HS = "m_axi_in_14_AW.data" *)output [2:0] m_axi_in_14_AWSIZE;
  (* RS_HS = "m_axi_in_14_AW.valid" *)output m_axi_in_14_AWVALID;
  (* RS_HS = "m_axi_in_14_B.data" *)input [0:0] m_axi_in_14_BID;
  (* RS_HS = "m_axi_in_14_B.ready" *)output m_axi_in_14_BREADY;
  (* RS_HS = "m_axi_in_14_B.data" *)input [1:0] m_axi_in_14_BRESP;
  (* RS_HS = "m_axi_in_14_B.valid" *)input m_axi_in_14_BVALID;
  (* RS_HS = "m_axi_in_14_R.data" *)input [255:0] m_axi_in_14_RDATA;
  (* RS_HS = "m_axi_in_14_R.data" *)input [0:0] m_axi_in_14_RID;
  (* RS_HS = "m_axi_in_14_R.data" *)input m_axi_in_14_RLAST;
  (* RS_HS = "m_axi_in_14_R.ready" *)output m_axi_in_14_RREADY;
  (* RS_HS = "m_axi_in_14_R.data" *)input [1:0] m_axi_in_14_RRESP;
  (* RS_HS = "m_axi_in_14_R.valid" *)input m_axi_in_14_RVALID;
  (* RS_HS = "m_axi_in_14_W.data" *)output [255:0] m_axi_in_14_WDATA;
  (* RS_HS = "m_axi_in_14_W.data" *)output m_axi_in_14_WLAST;
  (* RS_HS = "m_axi_in_14_W.ready" *)input m_axi_in_14_WREADY;
  (* RS_HS = "m_axi_in_14_W.data" *)output [31:0] m_axi_in_14_WSTRB;
  (* RS_HS = "m_axi_in_14_W.valid" *)output m_axi_in_14_WVALID;
  (* RS_HS = "m_axi_in_15_AR.data" *)output [63:0] m_axi_in_15_ARADDR;
  (* RS_HS = "m_axi_in_15_AR.data" *)output [1:0] m_axi_in_15_ARBURST;
  (* RS_HS = "m_axi_in_15_AR.data" *)output [3:0] m_axi_in_15_ARCACHE;
  (* RS_HS = "m_axi_in_15_AR.data" *)output [0:0] m_axi_in_15_ARID;
  (* RS_HS = "m_axi_in_15_AR.data" *)output [7:0] m_axi_in_15_ARLEN;
  (* RS_HS = "m_axi_in_15_AR.data" *)output m_axi_in_15_ARLOCK;
  (* RS_HS = "m_axi_in_15_AR.data" *)output [2:0] m_axi_in_15_ARPROT;
  (* RS_HS = "m_axi_in_15_AR.data" *)output [3:0] m_axi_in_15_ARQOS;
  (* RS_HS = "m_axi_in_15_AR.ready" *)input m_axi_in_15_ARREADY;
  (* RS_HS = "m_axi_in_15_AR.data" *)output [2:0] m_axi_in_15_ARSIZE;
  (* RS_HS = "m_axi_in_15_AR.valid" *)output m_axi_in_15_ARVALID;
  (* RS_HS = "m_axi_in_15_AW.data" *)output [63:0] m_axi_in_15_AWADDR;
  (* RS_HS = "m_axi_in_15_AW.data" *)output [1:0] m_axi_in_15_AWBURST;
  (* RS_HS = "m_axi_in_15_AW.data" *)output [3:0] m_axi_in_15_AWCACHE;
  (* RS_HS = "m_axi_in_15_AW.data" *)output [0:0] m_axi_in_15_AWID;
  (* RS_HS = "m_axi_in_15_AW.data" *)output [7:0] m_axi_in_15_AWLEN;
  (* RS_HS = "m_axi_in_15_AW.data" *)output m_axi_in_15_AWLOCK;
  (* RS_HS = "m_axi_in_15_AW.data" *)output [2:0] m_axi_in_15_AWPROT;
  (* RS_HS = "m_axi_in_15_AW.data" *)output [3:0] m_axi_in_15_AWQOS;
  (* RS_HS = "m_axi_in_15_AW.ready" *)input m_axi_in_15_AWREADY;
  (* RS_HS = "m_axi_in_15_AW.data" *)output [2:0] m_axi_in_15_AWSIZE;
  (* RS_HS = "m_axi_in_15_AW.valid" *)output m_axi_in_15_AWVALID;
  (* RS_HS = "m_axi_in_15_B.data" *)input [0:0] m_axi_in_15_BID;
  (* RS_HS = "m_axi_in_15_B.ready" *)output m_axi_in_15_BREADY;
  (* RS_HS = "m_axi_in_15_B.data" *)input [1:0] m_axi_in_15_BRESP;
  (* RS_HS = "m_axi_in_15_B.valid" *)input m_axi_in_15_BVALID;
  (* RS_HS = "m_axi_in_15_R.data" *)input [255:0] m_axi_in_15_RDATA;
  (* RS_HS = "m_axi_in_15_R.data" *)input [0:0] m_axi_in_15_RID;
  (* RS_HS = "m_axi_in_15_R.data" *)input m_axi_in_15_RLAST;
  (* RS_HS = "m_axi_in_15_R.ready" *)output m_axi_in_15_RREADY;
  (* RS_HS = "m_axi_in_15_R.data" *)input [1:0] m_axi_in_15_RRESP;
  (* RS_HS = "m_axi_in_15_R.valid" *)input m_axi_in_15_RVALID;
  (* RS_HS = "m_axi_in_15_W.data" *)output [255:0] m_axi_in_15_WDATA;
  (* RS_HS = "m_axi_in_15_W.data" *)output m_axi_in_15_WLAST;
  (* RS_HS = "m_axi_in_15_W.ready" *)input m_axi_in_15_WREADY;
  (* RS_HS = "m_axi_in_15_W.data" *)output [31:0] m_axi_in_15_WSTRB;
  (* RS_HS = "m_axi_in_15_W.valid" *)output m_axi_in_15_WVALID;
  (* RS_HS = "m_axi_in_16_AR.data" *)output [63:0] m_axi_in_16_ARADDR;
  (* RS_HS = "m_axi_in_16_AR.data" *)output [1:0] m_axi_in_16_ARBURST;
  (* RS_HS = "m_axi_in_16_AR.data" *)output [3:0] m_axi_in_16_ARCACHE;
  (* RS_HS = "m_axi_in_16_AR.data" *)output [0:0] m_axi_in_16_ARID;
  (* RS_HS = "m_axi_in_16_AR.data" *)output [7:0] m_axi_in_16_ARLEN;
  (* RS_HS = "m_axi_in_16_AR.data" *)output m_axi_in_16_ARLOCK;
  (* RS_HS = "m_axi_in_16_AR.data" *)output [2:0] m_axi_in_16_ARPROT;
  (* RS_HS = "m_axi_in_16_AR.data" *)output [3:0] m_axi_in_16_ARQOS;
  (* RS_HS = "m_axi_in_16_AR.ready" *)input m_axi_in_16_ARREADY;
  (* RS_HS = "m_axi_in_16_AR.data" *)output [2:0] m_axi_in_16_ARSIZE;
  (* RS_HS = "m_axi_in_16_AR.valid" *)output m_axi_in_16_ARVALID;
  (* RS_HS = "m_axi_in_16_AW.data" *)output [63:0] m_axi_in_16_AWADDR;
  (* RS_HS = "m_axi_in_16_AW.data" *)output [1:0] m_axi_in_16_AWBURST;
  (* RS_HS = "m_axi_in_16_AW.data" *)output [3:0] m_axi_in_16_AWCACHE;
  (* RS_HS = "m_axi_in_16_AW.data" *)output [0:0] m_axi_in_16_AWID;
  (* RS_HS = "m_axi_in_16_AW.data" *)output [7:0] m_axi_in_16_AWLEN;
  (* RS_HS = "m_axi_in_16_AW.data" *)output m_axi_in_16_AWLOCK;
  (* RS_HS = "m_axi_in_16_AW.data" *)output [2:0] m_axi_in_16_AWPROT;
  (* RS_HS = "m_axi_in_16_AW.data" *)output [3:0] m_axi_in_16_AWQOS;
  (* RS_HS = "m_axi_in_16_AW.ready" *)input m_axi_in_16_AWREADY;
  (* RS_HS = "m_axi_in_16_AW.data" *)output [2:0] m_axi_in_16_AWSIZE;
  (* RS_HS = "m_axi_in_16_AW.valid" *)output m_axi_in_16_AWVALID;
  (* RS_HS = "m_axi_in_16_B.data" *)input [0:0] m_axi_in_16_BID;
  (* RS_HS = "m_axi_in_16_B.ready" *)output m_axi_in_16_BREADY;
  (* RS_HS = "m_axi_in_16_B.data" *)input [1:0] m_axi_in_16_BRESP;
  (* RS_HS = "m_axi_in_16_B.valid" *)input m_axi_in_16_BVALID;
  (* RS_HS = "m_axi_in_16_R.data" *)input [255:0] m_axi_in_16_RDATA;
  (* RS_HS = "m_axi_in_16_R.data" *)input [0:0] m_axi_in_16_RID;
  (* RS_HS = "m_axi_in_16_R.data" *)input m_axi_in_16_RLAST;
  (* RS_HS = "m_axi_in_16_R.ready" *)output m_axi_in_16_RREADY;
  (* RS_HS = "m_axi_in_16_R.data" *)input [1:0] m_axi_in_16_RRESP;
  (* RS_HS = "m_axi_in_16_R.valid" *)input m_axi_in_16_RVALID;
  (* RS_HS = "m_axi_in_16_W.data" *)output [255:0] m_axi_in_16_WDATA;
  (* RS_HS = "m_axi_in_16_W.data" *)output m_axi_in_16_WLAST;
  (* RS_HS = "m_axi_in_16_W.ready" *)input m_axi_in_16_WREADY;
  (* RS_HS = "m_axi_in_16_W.data" *)output [31:0] m_axi_in_16_WSTRB;
  (* RS_HS = "m_axi_in_16_W.valid" *)output m_axi_in_16_WVALID;
  (* RS_HS = "m_axi_in_17_AR.data" *)output [63:0] m_axi_in_17_ARADDR;
  (* RS_HS = "m_axi_in_17_AR.data" *)output [1:0] m_axi_in_17_ARBURST;
  (* RS_HS = "m_axi_in_17_AR.data" *)output [3:0] m_axi_in_17_ARCACHE;
  (* RS_HS = "m_axi_in_17_AR.data" *)output [0:0] m_axi_in_17_ARID;
  (* RS_HS = "m_axi_in_17_AR.data" *)output [7:0] m_axi_in_17_ARLEN;
  (* RS_HS = "m_axi_in_17_AR.data" *)output m_axi_in_17_ARLOCK;
  (* RS_HS = "m_axi_in_17_AR.data" *)output [2:0] m_axi_in_17_ARPROT;
  (* RS_HS = "m_axi_in_17_AR.data" *)output [3:0] m_axi_in_17_ARQOS;
  (* RS_HS = "m_axi_in_17_AR.ready" *)input m_axi_in_17_ARREADY;
  (* RS_HS = "m_axi_in_17_AR.data" *)output [2:0] m_axi_in_17_ARSIZE;
  (* RS_HS = "m_axi_in_17_AR.valid" *)output m_axi_in_17_ARVALID;
  (* RS_HS = "m_axi_in_17_AW.data" *)output [63:0] m_axi_in_17_AWADDR;
  (* RS_HS = "m_axi_in_17_AW.data" *)output [1:0] m_axi_in_17_AWBURST;
  (* RS_HS = "m_axi_in_17_AW.data" *)output [3:0] m_axi_in_17_AWCACHE;
  (* RS_HS = "m_axi_in_17_AW.data" *)output [0:0] m_axi_in_17_AWID;
  (* RS_HS = "m_axi_in_17_AW.data" *)output [7:0] m_axi_in_17_AWLEN;
  (* RS_HS = "m_axi_in_17_AW.data" *)output m_axi_in_17_AWLOCK;
  (* RS_HS = "m_axi_in_17_AW.data" *)output [2:0] m_axi_in_17_AWPROT;
  (* RS_HS = "m_axi_in_17_AW.data" *)output [3:0] m_axi_in_17_AWQOS;
  (* RS_HS = "m_axi_in_17_AW.ready" *)input m_axi_in_17_AWREADY;
  (* RS_HS = "m_axi_in_17_AW.data" *)output [2:0] m_axi_in_17_AWSIZE;
  (* RS_HS = "m_axi_in_17_AW.valid" *)output m_axi_in_17_AWVALID;
  (* RS_HS = "m_axi_in_17_B.data" *)input [0:0] m_axi_in_17_BID;
  (* RS_HS = "m_axi_in_17_B.ready" *)output m_axi_in_17_BREADY;
  (* RS_HS = "m_axi_in_17_B.data" *)input [1:0] m_axi_in_17_BRESP;
  (* RS_HS = "m_axi_in_17_B.valid" *)input m_axi_in_17_BVALID;
  (* RS_HS = "m_axi_in_17_R.data" *)input [255:0] m_axi_in_17_RDATA;
  (* RS_HS = "m_axi_in_17_R.data" *)input [0:0] m_axi_in_17_RID;
  (* RS_HS = "m_axi_in_17_R.data" *)input m_axi_in_17_RLAST;
  (* RS_HS = "m_axi_in_17_R.ready" *)output m_axi_in_17_RREADY;
  (* RS_HS = "m_axi_in_17_R.data" *)input [1:0] m_axi_in_17_RRESP;
  (* RS_HS = "m_axi_in_17_R.valid" *)input m_axi_in_17_RVALID;
  (* RS_HS = "m_axi_in_17_W.data" *)output [255:0] m_axi_in_17_WDATA;
  (* RS_HS = "m_axi_in_17_W.data" *)output m_axi_in_17_WLAST;
  (* RS_HS = "m_axi_in_17_W.ready" *)input m_axi_in_17_WREADY;
  (* RS_HS = "m_axi_in_17_W.data" *)output [31:0] m_axi_in_17_WSTRB;
  (* RS_HS = "m_axi_in_17_W.valid" *)output m_axi_in_17_WVALID;
  (* RS_HS = "m_axi_in_18_AR.data" *)output [63:0] m_axi_in_18_ARADDR;
  (* RS_HS = "m_axi_in_18_AR.data" *)output [1:0] m_axi_in_18_ARBURST;
  (* RS_HS = "m_axi_in_18_AR.data" *)output [3:0] m_axi_in_18_ARCACHE;
  (* RS_HS = "m_axi_in_18_AR.data" *)output [0:0] m_axi_in_18_ARID;
  (* RS_HS = "m_axi_in_18_AR.data" *)output [7:0] m_axi_in_18_ARLEN;
  (* RS_HS = "m_axi_in_18_AR.data" *)output m_axi_in_18_ARLOCK;
  (* RS_HS = "m_axi_in_18_AR.data" *)output [2:0] m_axi_in_18_ARPROT;
  (* RS_HS = "m_axi_in_18_AR.data" *)output [3:0] m_axi_in_18_ARQOS;
  (* RS_HS = "m_axi_in_18_AR.ready" *)input m_axi_in_18_ARREADY;
  (* RS_HS = "m_axi_in_18_AR.data" *)output [2:0] m_axi_in_18_ARSIZE;
  (* RS_HS = "m_axi_in_18_AR.valid" *)output m_axi_in_18_ARVALID;
  (* RS_HS = "m_axi_in_18_AW.data" *)output [63:0] m_axi_in_18_AWADDR;
  (* RS_HS = "m_axi_in_18_AW.data" *)output [1:0] m_axi_in_18_AWBURST;
  (* RS_HS = "m_axi_in_18_AW.data" *)output [3:0] m_axi_in_18_AWCACHE;
  (* RS_HS = "m_axi_in_18_AW.data" *)output [0:0] m_axi_in_18_AWID;
  (* RS_HS = "m_axi_in_18_AW.data" *)output [7:0] m_axi_in_18_AWLEN;
  (* RS_HS = "m_axi_in_18_AW.data" *)output m_axi_in_18_AWLOCK;
  (* RS_HS = "m_axi_in_18_AW.data" *)output [2:0] m_axi_in_18_AWPROT;
  (* RS_HS = "m_axi_in_18_AW.data" *)output [3:0] m_axi_in_18_AWQOS;
  (* RS_HS = "m_axi_in_18_AW.ready" *)input m_axi_in_18_AWREADY;
  (* RS_HS = "m_axi_in_18_AW.data" *)output [2:0] m_axi_in_18_AWSIZE;
  (* RS_HS = "m_axi_in_18_AW.valid" *)output m_axi_in_18_AWVALID;
  (* RS_HS = "m_axi_in_18_B.data" *)input [0:0] m_axi_in_18_BID;
  (* RS_HS = "m_axi_in_18_B.ready" *)output m_axi_in_18_BREADY;
  (* RS_HS = "m_axi_in_18_B.data" *)input [1:0] m_axi_in_18_BRESP;
  (* RS_HS = "m_axi_in_18_B.valid" *)input m_axi_in_18_BVALID;
  (* RS_HS = "m_axi_in_18_R.data" *)input [255:0] m_axi_in_18_RDATA;
  (* RS_HS = "m_axi_in_18_R.data" *)input [0:0] m_axi_in_18_RID;
  (* RS_HS = "m_axi_in_18_R.data" *)input m_axi_in_18_RLAST;
  (* RS_HS = "m_axi_in_18_R.ready" *)output m_axi_in_18_RREADY;
  (* RS_HS = "m_axi_in_18_R.data" *)input [1:0] m_axi_in_18_RRESP;
  (* RS_HS = "m_axi_in_18_R.valid" *)input m_axi_in_18_RVALID;
  (* RS_HS = "m_axi_in_18_W.data" *)output [255:0] m_axi_in_18_WDATA;
  (* RS_HS = "m_axi_in_18_W.data" *)output m_axi_in_18_WLAST;
  (* RS_HS = "m_axi_in_18_W.ready" *)input m_axi_in_18_WREADY;
  (* RS_HS = "m_axi_in_18_W.data" *)output [31:0] m_axi_in_18_WSTRB;
  (* RS_HS = "m_axi_in_18_W.valid" *)output m_axi_in_18_WVALID;
  (* RS_HS = "m_axi_in_19_AR.data" *)output [63:0] m_axi_in_19_ARADDR;
  (* RS_HS = "m_axi_in_19_AR.data" *)output [1:0] m_axi_in_19_ARBURST;
  (* RS_HS = "m_axi_in_19_AR.data" *)output [3:0] m_axi_in_19_ARCACHE;
  (* RS_HS = "m_axi_in_19_AR.data" *)output [0:0] m_axi_in_19_ARID;
  (* RS_HS = "m_axi_in_19_AR.data" *)output [7:0] m_axi_in_19_ARLEN;
  (* RS_HS = "m_axi_in_19_AR.data" *)output m_axi_in_19_ARLOCK;
  (* RS_HS = "m_axi_in_19_AR.data" *)output [2:0] m_axi_in_19_ARPROT;
  (* RS_HS = "m_axi_in_19_AR.data" *)output [3:0] m_axi_in_19_ARQOS;
  (* RS_HS = "m_axi_in_19_AR.ready" *)input m_axi_in_19_ARREADY;
  (* RS_HS = "m_axi_in_19_AR.data" *)output [2:0] m_axi_in_19_ARSIZE;
  (* RS_HS = "m_axi_in_19_AR.valid" *)output m_axi_in_19_ARVALID;
  (* RS_HS = "m_axi_in_19_AW.data" *)output [63:0] m_axi_in_19_AWADDR;
  (* RS_HS = "m_axi_in_19_AW.data" *)output [1:0] m_axi_in_19_AWBURST;
  (* RS_HS = "m_axi_in_19_AW.data" *)output [3:0] m_axi_in_19_AWCACHE;
  (* RS_HS = "m_axi_in_19_AW.data" *)output [0:0] m_axi_in_19_AWID;
  (* RS_HS = "m_axi_in_19_AW.data" *)output [7:0] m_axi_in_19_AWLEN;
  (* RS_HS = "m_axi_in_19_AW.data" *)output m_axi_in_19_AWLOCK;
  (* RS_HS = "m_axi_in_19_AW.data" *)output [2:0] m_axi_in_19_AWPROT;
  (* RS_HS = "m_axi_in_19_AW.data" *)output [3:0] m_axi_in_19_AWQOS;
  (* RS_HS = "m_axi_in_19_AW.ready" *)input m_axi_in_19_AWREADY;
  (* RS_HS = "m_axi_in_19_AW.data" *)output [2:0] m_axi_in_19_AWSIZE;
  (* RS_HS = "m_axi_in_19_AW.valid" *)output m_axi_in_19_AWVALID;
  (* RS_HS = "m_axi_in_19_B.data" *)input [0:0] m_axi_in_19_BID;
  (* RS_HS = "m_axi_in_19_B.ready" *)output m_axi_in_19_BREADY;
  (* RS_HS = "m_axi_in_19_B.data" *)input [1:0] m_axi_in_19_BRESP;
  (* RS_HS = "m_axi_in_19_B.valid" *)input m_axi_in_19_BVALID;
  (* RS_HS = "m_axi_in_19_R.data" *)input [255:0] m_axi_in_19_RDATA;
  (* RS_HS = "m_axi_in_19_R.data" *)input [0:0] m_axi_in_19_RID;
  (* RS_HS = "m_axi_in_19_R.data" *)input m_axi_in_19_RLAST;
  (* RS_HS = "m_axi_in_19_R.ready" *)output m_axi_in_19_RREADY;
  (* RS_HS = "m_axi_in_19_R.data" *)input [1:0] m_axi_in_19_RRESP;
  (* RS_HS = "m_axi_in_19_R.valid" *)input m_axi_in_19_RVALID;
  (* RS_HS = "m_axi_in_19_W.data" *)output [255:0] m_axi_in_19_WDATA;
  (* RS_HS = "m_axi_in_19_W.data" *)output m_axi_in_19_WLAST;
  (* RS_HS = "m_axi_in_19_W.ready" *)input m_axi_in_19_WREADY;
  (* RS_HS = "m_axi_in_19_W.data" *)output [31:0] m_axi_in_19_WSTRB;
  (* RS_HS = "m_axi_in_19_W.valid" *)output m_axi_in_19_WVALID;
  (* RS_HS = "m_axi_in_2_AR.data" *)output [63:0] m_axi_in_2_ARADDR;
  (* RS_HS = "m_axi_in_2_AR.data" *)output [1:0] m_axi_in_2_ARBURST;
  (* RS_HS = "m_axi_in_2_AR.data" *)output [3:0] m_axi_in_2_ARCACHE;
  (* RS_HS = "m_axi_in_2_AR.data" *)output [0:0] m_axi_in_2_ARID;
  (* RS_HS = "m_axi_in_2_AR.data" *)output [7:0] m_axi_in_2_ARLEN;
  (* RS_HS = "m_axi_in_2_AR.data" *)output m_axi_in_2_ARLOCK;
  (* RS_HS = "m_axi_in_2_AR.data" *)output [2:0] m_axi_in_2_ARPROT;
  (* RS_HS = "m_axi_in_2_AR.data" *)output [3:0] m_axi_in_2_ARQOS;
  (* RS_HS = "m_axi_in_2_AR.ready" *)input m_axi_in_2_ARREADY;
  (* RS_HS = "m_axi_in_2_AR.data" *)output [2:0] m_axi_in_2_ARSIZE;
  (* RS_HS = "m_axi_in_2_AR.valid" *)output m_axi_in_2_ARVALID;
  (* RS_HS = "m_axi_in_2_AW.data" *)output [63:0] m_axi_in_2_AWADDR;
  (* RS_HS = "m_axi_in_2_AW.data" *)output [1:0] m_axi_in_2_AWBURST;
  (* RS_HS = "m_axi_in_2_AW.data" *)output [3:0] m_axi_in_2_AWCACHE;
  (* RS_HS = "m_axi_in_2_AW.data" *)output [0:0] m_axi_in_2_AWID;
  (* RS_HS = "m_axi_in_2_AW.data" *)output [7:0] m_axi_in_2_AWLEN;
  (* RS_HS = "m_axi_in_2_AW.data" *)output m_axi_in_2_AWLOCK;
  (* RS_HS = "m_axi_in_2_AW.data" *)output [2:0] m_axi_in_2_AWPROT;
  (* RS_HS = "m_axi_in_2_AW.data" *)output [3:0] m_axi_in_2_AWQOS;
  (* RS_HS = "m_axi_in_2_AW.ready" *)input m_axi_in_2_AWREADY;
  (* RS_HS = "m_axi_in_2_AW.data" *)output [2:0] m_axi_in_2_AWSIZE;
  (* RS_HS = "m_axi_in_2_AW.valid" *)output m_axi_in_2_AWVALID;
  (* RS_HS = "m_axi_in_2_B.data" *)input [0:0] m_axi_in_2_BID;
  (* RS_HS = "m_axi_in_2_B.ready" *)output m_axi_in_2_BREADY;
  (* RS_HS = "m_axi_in_2_B.data" *)input [1:0] m_axi_in_2_BRESP;
  (* RS_HS = "m_axi_in_2_B.valid" *)input m_axi_in_2_BVALID;
  (* RS_HS = "m_axi_in_2_R.data" *)input [255:0] m_axi_in_2_RDATA;
  (* RS_HS = "m_axi_in_2_R.data" *)input [0:0] m_axi_in_2_RID;
  (* RS_HS = "m_axi_in_2_R.data" *)input m_axi_in_2_RLAST;
  (* RS_HS = "m_axi_in_2_R.ready" *)output m_axi_in_2_RREADY;
  (* RS_HS = "m_axi_in_2_R.data" *)input [1:0] m_axi_in_2_RRESP;
  (* RS_HS = "m_axi_in_2_R.valid" *)input m_axi_in_2_RVALID;
  (* RS_HS = "m_axi_in_2_W.data" *)output [255:0] m_axi_in_2_WDATA;
  (* RS_HS = "m_axi_in_2_W.data" *)output m_axi_in_2_WLAST;
  (* RS_HS = "m_axi_in_2_W.ready" *)input m_axi_in_2_WREADY;
  (* RS_HS = "m_axi_in_2_W.data" *)output [31:0] m_axi_in_2_WSTRB;
  (* RS_HS = "m_axi_in_2_W.valid" *)output m_axi_in_2_WVALID;
  (* RS_HS = "m_axi_in_20_AR.data" *)output [63:0] m_axi_in_20_ARADDR;
  (* RS_HS = "m_axi_in_20_AR.data" *)output [1:0] m_axi_in_20_ARBURST;
  (* RS_HS = "m_axi_in_20_AR.data" *)output [3:0] m_axi_in_20_ARCACHE;
  (* RS_HS = "m_axi_in_20_AR.data" *)output [0:0] m_axi_in_20_ARID;
  (* RS_HS = "m_axi_in_20_AR.data" *)output [7:0] m_axi_in_20_ARLEN;
  (* RS_HS = "m_axi_in_20_AR.data" *)output m_axi_in_20_ARLOCK;
  (* RS_HS = "m_axi_in_20_AR.data" *)output [2:0] m_axi_in_20_ARPROT;
  (* RS_HS = "m_axi_in_20_AR.data" *)output [3:0] m_axi_in_20_ARQOS;
  (* RS_HS = "m_axi_in_20_AR.ready" *)input m_axi_in_20_ARREADY;
  (* RS_HS = "m_axi_in_20_AR.data" *)output [2:0] m_axi_in_20_ARSIZE;
  (* RS_HS = "m_axi_in_20_AR.valid" *)output m_axi_in_20_ARVALID;
  (* RS_HS = "m_axi_in_20_AW.data" *)output [63:0] m_axi_in_20_AWADDR;
  (* RS_HS = "m_axi_in_20_AW.data" *)output [1:0] m_axi_in_20_AWBURST;
  (* RS_HS = "m_axi_in_20_AW.data" *)output [3:0] m_axi_in_20_AWCACHE;
  (* RS_HS = "m_axi_in_20_AW.data" *)output [0:0] m_axi_in_20_AWID;
  (* RS_HS = "m_axi_in_20_AW.data" *)output [7:0] m_axi_in_20_AWLEN;
  (* RS_HS = "m_axi_in_20_AW.data" *)output m_axi_in_20_AWLOCK;
  (* RS_HS = "m_axi_in_20_AW.data" *)output [2:0] m_axi_in_20_AWPROT;
  (* RS_HS = "m_axi_in_20_AW.data" *)output [3:0] m_axi_in_20_AWQOS;
  (* RS_HS = "m_axi_in_20_AW.ready" *)input m_axi_in_20_AWREADY;
  (* RS_HS = "m_axi_in_20_AW.data" *)output [2:0] m_axi_in_20_AWSIZE;
  (* RS_HS = "m_axi_in_20_AW.valid" *)output m_axi_in_20_AWVALID;
  (* RS_HS = "m_axi_in_20_B.data" *)input [0:0] m_axi_in_20_BID;
  (* RS_HS = "m_axi_in_20_B.ready" *)output m_axi_in_20_BREADY;
  (* RS_HS = "m_axi_in_20_B.data" *)input [1:0] m_axi_in_20_BRESP;
  (* RS_HS = "m_axi_in_20_B.valid" *)input m_axi_in_20_BVALID;
  (* RS_HS = "m_axi_in_20_R.data" *)input [255:0] m_axi_in_20_RDATA;
  (* RS_HS = "m_axi_in_20_R.data" *)input [0:0] m_axi_in_20_RID;
  (* RS_HS = "m_axi_in_20_R.data" *)input m_axi_in_20_RLAST;
  (* RS_HS = "m_axi_in_20_R.ready" *)output m_axi_in_20_RREADY;
  (* RS_HS = "m_axi_in_20_R.data" *)input [1:0] m_axi_in_20_RRESP;
  (* RS_HS = "m_axi_in_20_R.valid" *)input m_axi_in_20_RVALID;
  (* RS_HS = "m_axi_in_20_W.data" *)output [255:0] m_axi_in_20_WDATA;
  (* RS_HS = "m_axi_in_20_W.data" *)output m_axi_in_20_WLAST;
  (* RS_HS = "m_axi_in_20_W.ready" *)input m_axi_in_20_WREADY;
  (* RS_HS = "m_axi_in_20_W.data" *)output [31:0] m_axi_in_20_WSTRB;
  (* RS_HS = "m_axi_in_20_W.valid" *)output m_axi_in_20_WVALID;
  (* RS_HS = "m_axi_in_21_AR.data" *)output [63:0] m_axi_in_21_ARADDR;
  (* RS_HS = "m_axi_in_21_AR.data" *)output [1:0] m_axi_in_21_ARBURST;
  (* RS_HS = "m_axi_in_21_AR.data" *)output [3:0] m_axi_in_21_ARCACHE;
  (* RS_HS = "m_axi_in_21_AR.data" *)output [0:0] m_axi_in_21_ARID;
  (* RS_HS = "m_axi_in_21_AR.data" *)output [7:0] m_axi_in_21_ARLEN;
  (* RS_HS = "m_axi_in_21_AR.data" *)output m_axi_in_21_ARLOCK;
  (* RS_HS = "m_axi_in_21_AR.data" *)output [2:0] m_axi_in_21_ARPROT;
  (* RS_HS = "m_axi_in_21_AR.data" *)output [3:0] m_axi_in_21_ARQOS;
  (* RS_HS = "m_axi_in_21_AR.ready" *)input m_axi_in_21_ARREADY;
  (* RS_HS = "m_axi_in_21_AR.data" *)output [2:0] m_axi_in_21_ARSIZE;
  (* RS_HS = "m_axi_in_21_AR.valid" *)output m_axi_in_21_ARVALID;
  (* RS_HS = "m_axi_in_21_AW.data" *)output [63:0] m_axi_in_21_AWADDR;
  (* RS_HS = "m_axi_in_21_AW.data" *)output [1:0] m_axi_in_21_AWBURST;
  (* RS_HS = "m_axi_in_21_AW.data" *)output [3:0] m_axi_in_21_AWCACHE;
  (* RS_HS = "m_axi_in_21_AW.data" *)output [0:0] m_axi_in_21_AWID;
  (* RS_HS = "m_axi_in_21_AW.data" *)output [7:0] m_axi_in_21_AWLEN;
  (* RS_HS = "m_axi_in_21_AW.data" *)output m_axi_in_21_AWLOCK;
  (* RS_HS = "m_axi_in_21_AW.data" *)output [2:0] m_axi_in_21_AWPROT;
  (* RS_HS = "m_axi_in_21_AW.data" *)output [3:0] m_axi_in_21_AWQOS;
  (* RS_HS = "m_axi_in_21_AW.ready" *)input m_axi_in_21_AWREADY;
  (* RS_HS = "m_axi_in_21_AW.data" *)output [2:0] m_axi_in_21_AWSIZE;
  (* RS_HS = "m_axi_in_21_AW.valid" *)output m_axi_in_21_AWVALID;
  (* RS_HS = "m_axi_in_21_B.data" *)input [0:0] m_axi_in_21_BID;
  (* RS_HS = "m_axi_in_21_B.ready" *)output m_axi_in_21_BREADY;
  (* RS_HS = "m_axi_in_21_B.data" *)input [1:0] m_axi_in_21_BRESP;
  (* RS_HS = "m_axi_in_21_B.valid" *)input m_axi_in_21_BVALID;
  (* RS_HS = "m_axi_in_21_R.data" *)input [255:0] m_axi_in_21_RDATA;
  (* RS_HS = "m_axi_in_21_R.data" *)input [0:0] m_axi_in_21_RID;
  (* RS_HS = "m_axi_in_21_R.data" *)input m_axi_in_21_RLAST;
  (* RS_HS = "m_axi_in_21_R.ready" *)output m_axi_in_21_RREADY;
  (* RS_HS = "m_axi_in_21_R.data" *)input [1:0] m_axi_in_21_RRESP;
  (* RS_HS = "m_axi_in_21_R.valid" *)input m_axi_in_21_RVALID;
  (* RS_HS = "m_axi_in_21_W.data" *)output [255:0] m_axi_in_21_WDATA;
  (* RS_HS = "m_axi_in_21_W.data" *)output m_axi_in_21_WLAST;
  (* RS_HS = "m_axi_in_21_W.ready" *)input m_axi_in_21_WREADY;
  (* RS_HS = "m_axi_in_21_W.data" *)output [31:0] m_axi_in_21_WSTRB;
  (* RS_HS = "m_axi_in_21_W.valid" *)output m_axi_in_21_WVALID;
  (* RS_HS = "m_axi_in_22_AR.data" *)output [63:0] m_axi_in_22_ARADDR;
  (* RS_HS = "m_axi_in_22_AR.data" *)output [1:0] m_axi_in_22_ARBURST;
  (* RS_HS = "m_axi_in_22_AR.data" *)output [3:0] m_axi_in_22_ARCACHE;
  (* RS_HS = "m_axi_in_22_AR.data" *)output [0:0] m_axi_in_22_ARID;
  (* RS_HS = "m_axi_in_22_AR.data" *)output [7:0] m_axi_in_22_ARLEN;
  (* RS_HS = "m_axi_in_22_AR.data" *)output m_axi_in_22_ARLOCK;
  (* RS_HS = "m_axi_in_22_AR.data" *)output [2:0] m_axi_in_22_ARPROT;
  (* RS_HS = "m_axi_in_22_AR.data" *)output [3:0] m_axi_in_22_ARQOS;
  (* RS_HS = "m_axi_in_22_AR.ready" *)input m_axi_in_22_ARREADY;
  (* RS_HS = "m_axi_in_22_AR.data" *)output [2:0] m_axi_in_22_ARSIZE;
  (* RS_HS = "m_axi_in_22_AR.valid" *)output m_axi_in_22_ARVALID;
  (* RS_HS = "m_axi_in_22_AW.data" *)output [63:0] m_axi_in_22_AWADDR;
  (* RS_HS = "m_axi_in_22_AW.data" *)output [1:0] m_axi_in_22_AWBURST;
  (* RS_HS = "m_axi_in_22_AW.data" *)output [3:0] m_axi_in_22_AWCACHE;
  (* RS_HS = "m_axi_in_22_AW.data" *)output [0:0] m_axi_in_22_AWID;
  (* RS_HS = "m_axi_in_22_AW.data" *)output [7:0] m_axi_in_22_AWLEN;
  (* RS_HS = "m_axi_in_22_AW.data" *)output m_axi_in_22_AWLOCK;
  (* RS_HS = "m_axi_in_22_AW.data" *)output [2:0] m_axi_in_22_AWPROT;
  (* RS_HS = "m_axi_in_22_AW.data" *)output [3:0] m_axi_in_22_AWQOS;
  (* RS_HS = "m_axi_in_22_AW.ready" *)input m_axi_in_22_AWREADY;
  (* RS_HS = "m_axi_in_22_AW.data" *)output [2:0] m_axi_in_22_AWSIZE;
  (* RS_HS = "m_axi_in_22_AW.valid" *)output m_axi_in_22_AWVALID;
  (* RS_HS = "m_axi_in_22_B.data" *)input [0:0] m_axi_in_22_BID;
  (* RS_HS = "m_axi_in_22_B.ready" *)output m_axi_in_22_BREADY;
  (* RS_HS = "m_axi_in_22_B.data" *)input [1:0] m_axi_in_22_BRESP;
  (* RS_HS = "m_axi_in_22_B.valid" *)input m_axi_in_22_BVALID;
  (* RS_HS = "m_axi_in_22_R.data" *)input [255:0] m_axi_in_22_RDATA;
  (* RS_HS = "m_axi_in_22_R.data" *)input [0:0] m_axi_in_22_RID;
  (* RS_HS = "m_axi_in_22_R.data" *)input m_axi_in_22_RLAST;
  (* RS_HS = "m_axi_in_22_R.ready" *)output m_axi_in_22_RREADY;
  (* RS_HS = "m_axi_in_22_R.data" *)input [1:0] m_axi_in_22_RRESP;
  (* RS_HS = "m_axi_in_22_R.valid" *)input m_axi_in_22_RVALID;
  (* RS_HS = "m_axi_in_22_W.data" *)output [255:0] m_axi_in_22_WDATA;
  (* RS_HS = "m_axi_in_22_W.data" *)output m_axi_in_22_WLAST;
  (* RS_HS = "m_axi_in_22_W.ready" *)input m_axi_in_22_WREADY;
  (* RS_HS = "m_axi_in_22_W.data" *)output [31:0] m_axi_in_22_WSTRB;
  (* RS_HS = "m_axi_in_22_W.valid" *)output m_axi_in_22_WVALID;
  (* RS_HS = "m_axi_in_23_AR.data" *)output [63:0] m_axi_in_23_ARADDR;
  (* RS_HS = "m_axi_in_23_AR.data" *)output [1:0] m_axi_in_23_ARBURST;
  (* RS_HS = "m_axi_in_23_AR.data" *)output [3:0] m_axi_in_23_ARCACHE;
  (* RS_HS = "m_axi_in_23_AR.data" *)output [0:0] m_axi_in_23_ARID;
  (* RS_HS = "m_axi_in_23_AR.data" *)output [7:0] m_axi_in_23_ARLEN;
  (* RS_HS = "m_axi_in_23_AR.data" *)output m_axi_in_23_ARLOCK;
  (* RS_HS = "m_axi_in_23_AR.data" *)output [2:0] m_axi_in_23_ARPROT;
  (* RS_HS = "m_axi_in_23_AR.data" *)output [3:0] m_axi_in_23_ARQOS;
  (* RS_HS = "m_axi_in_23_AR.ready" *)input m_axi_in_23_ARREADY;
  (* RS_HS = "m_axi_in_23_AR.data" *)output [2:0] m_axi_in_23_ARSIZE;
  (* RS_HS = "m_axi_in_23_AR.valid" *)output m_axi_in_23_ARVALID;
  (* RS_HS = "m_axi_in_23_AW.data" *)output [63:0] m_axi_in_23_AWADDR;
  (* RS_HS = "m_axi_in_23_AW.data" *)output [1:0] m_axi_in_23_AWBURST;
  (* RS_HS = "m_axi_in_23_AW.data" *)output [3:0] m_axi_in_23_AWCACHE;
  (* RS_HS = "m_axi_in_23_AW.data" *)output [0:0] m_axi_in_23_AWID;
  (* RS_HS = "m_axi_in_23_AW.data" *)output [7:0] m_axi_in_23_AWLEN;
  (* RS_HS = "m_axi_in_23_AW.data" *)output m_axi_in_23_AWLOCK;
  (* RS_HS = "m_axi_in_23_AW.data" *)output [2:0] m_axi_in_23_AWPROT;
  (* RS_HS = "m_axi_in_23_AW.data" *)output [3:0] m_axi_in_23_AWQOS;
  (* RS_HS = "m_axi_in_23_AW.ready" *)input m_axi_in_23_AWREADY;
  (* RS_HS = "m_axi_in_23_AW.data" *)output [2:0] m_axi_in_23_AWSIZE;
  (* RS_HS = "m_axi_in_23_AW.valid" *)output m_axi_in_23_AWVALID;
  (* RS_HS = "m_axi_in_23_B.data" *)input [0:0] m_axi_in_23_BID;
  (* RS_HS = "m_axi_in_23_B.ready" *)output m_axi_in_23_BREADY;
  (* RS_HS = "m_axi_in_23_B.data" *)input [1:0] m_axi_in_23_BRESP;
  (* RS_HS = "m_axi_in_23_B.valid" *)input m_axi_in_23_BVALID;
  (* RS_HS = "m_axi_in_23_R.data" *)input [255:0] m_axi_in_23_RDATA;
  (* RS_HS = "m_axi_in_23_R.data" *)input [0:0] m_axi_in_23_RID;
  (* RS_HS = "m_axi_in_23_R.data" *)input m_axi_in_23_RLAST;
  (* RS_HS = "m_axi_in_23_R.ready" *)output m_axi_in_23_RREADY;
  (* RS_HS = "m_axi_in_23_R.data" *)input [1:0] m_axi_in_23_RRESP;
  (* RS_HS = "m_axi_in_23_R.valid" *)input m_axi_in_23_RVALID;
  (* RS_HS = "m_axi_in_23_W.data" *)output [255:0] m_axi_in_23_WDATA;
  (* RS_HS = "m_axi_in_23_W.data" *)output m_axi_in_23_WLAST;
  (* RS_HS = "m_axi_in_23_W.ready" *)input m_axi_in_23_WREADY;
  (* RS_HS = "m_axi_in_23_W.data" *)output [31:0] m_axi_in_23_WSTRB;
  (* RS_HS = "m_axi_in_23_W.valid" *)output m_axi_in_23_WVALID;
  (* RS_HS = "m_axi_in_24_AR.data" *)output [63:0] m_axi_in_24_ARADDR;
  (* RS_HS = "m_axi_in_24_AR.data" *)output [1:0] m_axi_in_24_ARBURST;
  (* RS_HS = "m_axi_in_24_AR.data" *)output [3:0] m_axi_in_24_ARCACHE;
  (* RS_HS = "m_axi_in_24_AR.data" *)output [0:0] m_axi_in_24_ARID;
  (* RS_HS = "m_axi_in_24_AR.data" *)output [7:0] m_axi_in_24_ARLEN;
  (* RS_HS = "m_axi_in_24_AR.data" *)output m_axi_in_24_ARLOCK;
  (* RS_HS = "m_axi_in_24_AR.data" *)output [2:0] m_axi_in_24_ARPROT;
  (* RS_HS = "m_axi_in_24_AR.data" *)output [3:0] m_axi_in_24_ARQOS;
  (* RS_HS = "m_axi_in_24_AR.ready" *)input m_axi_in_24_ARREADY;
  (* RS_HS = "m_axi_in_24_AR.data" *)output [2:0] m_axi_in_24_ARSIZE;
  (* RS_HS = "m_axi_in_24_AR.valid" *)output m_axi_in_24_ARVALID;
  (* RS_HS = "m_axi_in_24_AW.data" *)output [63:0] m_axi_in_24_AWADDR;
  (* RS_HS = "m_axi_in_24_AW.data" *)output [1:0] m_axi_in_24_AWBURST;
  (* RS_HS = "m_axi_in_24_AW.data" *)output [3:0] m_axi_in_24_AWCACHE;
  (* RS_HS = "m_axi_in_24_AW.data" *)output [0:0] m_axi_in_24_AWID;
  (* RS_HS = "m_axi_in_24_AW.data" *)output [7:0] m_axi_in_24_AWLEN;
  (* RS_HS = "m_axi_in_24_AW.data" *)output m_axi_in_24_AWLOCK;
  (* RS_HS = "m_axi_in_24_AW.data" *)output [2:0] m_axi_in_24_AWPROT;
  (* RS_HS = "m_axi_in_24_AW.data" *)output [3:0] m_axi_in_24_AWQOS;
  (* RS_HS = "m_axi_in_24_AW.ready" *)input m_axi_in_24_AWREADY;
  (* RS_HS = "m_axi_in_24_AW.data" *)output [2:0] m_axi_in_24_AWSIZE;
  (* RS_HS = "m_axi_in_24_AW.valid" *)output m_axi_in_24_AWVALID;
  (* RS_HS = "m_axi_in_24_B.data" *)input [0:0] m_axi_in_24_BID;
  (* RS_HS = "m_axi_in_24_B.ready" *)output m_axi_in_24_BREADY;
  (* RS_HS = "m_axi_in_24_B.data" *)input [1:0] m_axi_in_24_BRESP;
  (* RS_HS = "m_axi_in_24_B.valid" *)input m_axi_in_24_BVALID;
  (* RS_HS = "m_axi_in_24_R.data" *)input [255:0] m_axi_in_24_RDATA;
  (* RS_HS = "m_axi_in_24_R.data" *)input [0:0] m_axi_in_24_RID;
  (* RS_HS = "m_axi_in_24_R.data" *)input m_axi_in_24_RLAST;
  (* RS_HS = "m_axi_in_24_R.ready" *)output m_axi_in_24_RREADY;
  (* RS_HS = "m_axi_in_24_R.data" *)input [1:0] m_axi_in_24_RRESP;
  (* RS_HS = "m_axi_in_24_R.valid" *)input m_axi_in_24_RVALID;
  (* RS_HS = "m_axi_in_24_W.data" *)output [255:0] m_axi_in_24_WDATA;
  (* RS_HS = "m_axi_in_24_W.data" *)output m_axi_in_24_WLAST;
  (* RS_HS = "m_axi_in_24_W.ready" *)input m_axi_in_24_WREADY;
  (* RS_HS = "m_axi_in_24_W.data" *)output [31:0] m_axi_in_24_WSTRB;
  (* RS_HS = "m_axi_in_24_W.valid" *)output m_axi_in_24_WVALID;
  (* RS_HS = "m_axi_in_25_AR.data" *)output [63:0] m_axi_in_25_ARADDR;
  (* RS_HS = "m_axi_in_25_AR.data" *)output [1:0] m_axi_in_25_ARBURST;
  (* RS_HS = "m_axi_in_25_AR.data" *)output [3:0] m_axi_in_25_ARCACHE;
  (* RS_HS = "m_axi_in_25_AR.data" *)output [0:0] m_axi_in_25_ARID;
  (* RS_HS = "m_axi_in_25_AR.data" *)output [7:0] m_axi_in_25_ARLEN;
  (* RS_HS = "m_axi_in_25_AR.data" *)output m_axi_in_25_ARLOCK;
  (* RS_HS = "m_axi_in_25_AR.data" *)output [2:0] m_axi_in_25_ARPROT;
  (* RS_HS = "m_axi_in_25_AR.data" *)output [3:0] m_axi_in_25_ARQOS;
  (* RS_HS = "m_axi_in_25_AR.ready" *)input m_axi_in_25_ARREADY;
  (* RS_HS = "m_axi_in_25_AR.data" *)output [2:0] m_axi_in_25_ARSIZE;
  (* RS_HS = "m_axi_in_25_AR.valid" *)output m_axi_in_25_ARVALID;
  (* RS_HS = "m_axi_in_25_AW.data" *)output [63:0] m_axi_in_25_AWADDR;
  (* RS_HS = "m_axi_in_25_AW.data" *)output [1:0] m_axi_in_25_AWBURST;
  (* RS_HS = "m_axi_in_25_AW.data" *)output [3:0] m_axi_in_25_AWCACHE;
  (* RS_HS = "m_axi_in_25_AW.data" *)output [0:0] m_axi_in_25_AWID;
  (* RS_HS = "m_axi_in_25_AW.data" *)output [7:0] m_axi_in_25_AWLEN;
  (* RS_HS = "m_axi_in_25_AW.data" *)output m_axi_in_25_AWLOCK;
  (* RS_HS = "m_axi_in_25_AW.data" *)output [2:0] m_axi_in_25_AWPROT;
  (* RS_HS = "m_axi_in_25_AW.data" *)output [3:0] m_axi_in_25_AWQOS;
  (* RS_HS = "m_axi_in_25_AW.ready" *)input m_axi_in_25_AWREADY;
  (* RS_HS = "m_axi_in_25_AW.data" *)output [2:0] m_axi_in_25_AWSIZE;
  (* RS_HS = "m_axi_in_25_AW.valid" *)output m_axi_in_25_AWVALID;
  (* RS_HS = "m_axi_in_25_B.data" *)input [0:0] m_axi_in_25_BID;
  (* RS_HS = "m_axi_in_25_B.ready" *)output m_axi_in_25_BREADY;
  (* RS_HS = "m_axi_in_25_B.data" *)input [1:0] m_axi_in_25_BRESP;
  (* RS_HS = "m_axi_in_25_B.valid" *)input m_axi_in_25_BVALID;
  (* RS_HS = "m_axi_in_25_R.data" *)input [255:0] m_axi_in_25_RDATA;
  (* RS_HS = "m_axi_in_25_R.data" *)input [0:0] m_axi_in_25_RID;
  (* RS_HS = "m_axi_in_25_R.data" *)input m_axi_in_25_RLAST;
  (* RS_HS = "m_axi_in_25_R.ready" *)output m_axi_in_25_RREADY;
  (* RS_HS = "m_axi_in_25_R.data" *)input [1:0] m_axi_in_25_RRESP;
  (* RS_HS = "m_axi_in_25_R.valid" *)input m_axi_in_25_RVALID;
  (* RS_HS = "m_axi_in_25_W.data" *)output [255:0] m_axi_in_25_WDATA;
  (* RS_HS = "m_axi_in_25_W.data" *)output m_axi_in_25_WLAST;
  (* RS_HS = "m_axi_in_25_W.ready" *)input m_axi_in_25_WREADY;
  (* RS_HS = "m_axi_in_25_W.data" *)output [31:0] m_axi_in_25_WSTRB;
  (* RS_HS = "m_axi_in_25_W.valid" *)output m_axi_in_25_WVALID;
  (* RS_HS = "m_axi_in_26_AR.data" *)output [63:0] m_axi_in_26_ARADDR;
  (* RS_HS = "m_axi_in_26_AR.data" *)output [1:0] m_axi_in_26_ARBURST;
  (* RS_HS = "m_axi_in_26_AR.data" *)output [3:0] m_axi_in_26_ARCACHE;
  (* RS_HS = "m_axi_in_26_AR.data" *)output [0:0] m_axi_in_26_ARID;
  (* RS_HS = "m_axi_in_26_AR.data" *)output [7:0] m_axi_in_26_ARLEN;
  (* RS_HS = "m_axi_in_26_AR.data" *)output m_axi_in_26_ARLOCK;
  (* RS_HS = "m_axi_in_26_AR.data" *)output [2:0] m_axi_in_26_ARPROT;
  (* RS_HS = "m_axi_in_26_AR.data" *)output [3:0] m_axi_in_26_ARQOS;
  (* RS_HS = "m_axi_in_26_AR.ready" *)input m_axi_in_26_ARREADY;
  (* RS_HS = "m_axi_in_26_AR.data" *)output [2:0] m_axi_in_26_ARSIZE;
  (* RS_HS = "m_axi_in_26_AR.valid" *)output m_axi_in_26_ARVALID;
  (* RS_HS = "m_axi_in_26_AW.data" *)output [63:0] m_axi_in_26_AWADDR;
  (* RS_HS = "m_axi_in_26_AW.data" *)output [1:0] m_axi_in_26_AWBURST;
  (* RS_HS = "m_axi_in_26_AW.data" *)output [3:0] m_axi_in_26_AWCACHE;
  (* RS_HS = "m_axi_in_26_AW.data" *)output [0:0] m_axi_in_26_AWID;
  (* RS_HS = "m_axi_in_26_AW.data" *)output [7:0] m_axi_in_26_AWLEN;
  (* RS_HS = "m_axi_in_26_AW.data" *)output m_axi_in_26_AWLOCK;
  (* RS_HS = "m_axi_in_26_AW.data" *)output [2:0] m_axi_in_26_AWPROT;
  (* RS_HS = "m_axi_in_26_AW.data" *)output [3:0] m_axi_in_26_AWQOS;
  (* RS_HS = "m_axi_in_26_AW.ready" *)input m_axi_in_26_AWREADY;
  (* RS_HS = "m_axi_in_26_AW.data" *)output [2:0] m_axi_in_26_AWSIZE;
  (* RS_HS = "m_axi_in_26_AW.valid" *)output m_axi_in_26_AWVALID;
  (* RS_HS = "m_axi_in_26_B.data" *)input [0:0] m_axi_in_26_BID;
  (* RS_HS = "m_axi_in_26_B.ready" *)output m_axi_in_26_BREADY;
  (* RS_HS = "m_axi_in_26_B.data" *)input [1:0] m_axi_in_26_BRESP;
  (* RS_HS = "m_axi_in_26_B.valid" *)input m_axi_in_26_BVALID;
  (* RS_HS = "m_axi_in_26_R.data" *)input [255:0] m_axi_in_26_RDATA;
  (* RS_HS = "m_axi_in_26_R.data" *)input [0:0] m_axi_in_26_RID;
  (* RS_HS = "m_axi_in_26_R.data" *)input m_axi_in_26_RLAST;
  (* RS_HS = "m_axi_in_26_R.ready" *)output m_axi_in_26_RREADY;
  (* RS_HS = "m_axi_in_26_R.data" *)input [1:0] m_axi_in_26_RRESP;
  (* RS_HS = "m_axi_in_26_R.valid" *)input m_axi_in_26_RVALID;
  (* RS_HS = "m_axi_in_26_W.data" *)output [255:0] m_axi_in_26_WDATA;
  (* RS_HS = "m_axi_in_26_W.data" *)output m_axi_in_26_WLAST;
  (* RS_HS = "m_axi_in_26_W.ready" *)input m_axi_in_26_WREADY;
  (* RS_HS = "m_axi_in_26_W.data" *)output [31:0] m_axi_in_26_WSTRB;
  (* RS_HS = "m_axi_in_26_W.valid" *)output m_axi_in_26_WVALID;
  (* RS_HS = "m_axi_in_3_AR.data" *)output [63:0] m_axi_in_3_ARADDR;
  (* RS_HS = "m_axi_in_3_AR.data" *)output [1:0] m_axi_in_3_ARBURST;
  (* RS_HS = "m_axi_in_3_AR.data" *)output [3:0] m_axi_in_3_ARCACHE;
  (* RS_HS = "m_axi_in_3_AR.data" *)output [0:0] m_axi_in_3_ARID;
  (* RS_HS = "m_axi_in_3_AR.data" *)output [7:0] m_axi_in_3_ARLEN;
  (* RS_HS = "m_axi_in_3_AR.data" *)output m_axi_in_3_ARLOCK;
  (* RS_HS = "m_axi_in_3_AR.data" *)output [2:0] m_axi_in_3_ARPROT;
  (* RS_HS = "m_axi_in_3_AR.data" *)output [3:0] m_axi_in_3_ARQOS;
  (* RS_HS = "m_axi_in_3_AR.ready" *)input m_axi_in_3_ARREADY;
  (* RS_HS = "m_axi_in_3_AR.data" *)output [2:0] m_axi_in_3_ARSIZE;
  (* RS_HS = "m_axi_in_3_AR.valid" *)output m_axi_in_3_ARVALID;
  (* RS_HS = "m_axi_in_3_AW.data" *)output [63:0] m_axi_in_3_AWADDR;
  (* RS_HS = "m_axi_in_3_AW.data" *)output [1:0] m_axi_in_3_AWBURST;
  (* RS_HS = "m_axi_in_3_AW.data" *)output [3:0] m_axi_in_3_AWCACHE;
  (* RS_HS = "m_axi_in_3_AW.data" *)output [0:0] m_axi_in_3_AWID;
  (* RS_HS = "m_axi_in_3_AW.data" *)output [7:0] m_axi_in_3_AWLEN;
  (* RS_HS = "m_axi_in_3_AW.data" *)output m_axi_in_3_AWLOCK;
  (* RS_HS = "m_axi_in_3_AW.data" *)output [2:0] m_axi_in_3_AWPROT;
  (* RS_HS = "m_axi_in_3_AW.data" *)output [3:0] m_axi_in_3_AWQOS;
  (* RS_HS = "m_axi_in_3_AW.ready" *)input m_axi_in_3_AWREADY;
  (* RS_HS = "m_axi_in_3_AW.data" *)output [2:0] m_axi_in_3_AWSIZE;
  (* RS_HS = "m_axi_in_3_AW.valid" *)output m_axi_in_3_AWVALID;
  (* RS_HS = "m_axi_in_3_B.data" *)input [0:0] m_axi_in_3_BID;
  (* RS_HS = "m_axi_in_3_B.ready" *)output m_axi_in_3_BREADY;
  (* RS_HS = "m_axi_in_3_B.data" *)input [1:0] m_axi_in_3_BRESP;
  (* RS_HS = "m_axi_in_3_B.valid" *)input m_axi_in_3_BVALID;
  (* RS_HS = "m_axi_in_3_R.data" *)input [255:0] m_axi_in_3_RDATA;
  (* RS_HS = "m_axi_in_3_R.data" *)input [0:0] m_axi_in_3_RID;
  (* RS_HS = "m_axi_in_3_R.data" *)input m_axi_in_3_RLAST;
  (* RS_HS = "m_axi_in_3_R.ready" *)output m_axi_in_3_RREADY;
  (* RS_HS = "m_axi_in_3_R.data" *)input [1:0] m_axi_in_3_RRESP;
  (* RS_HS = "m_axi_in_3_R.valid" *)input m_axi_in_3_RVALID;
  (* RS_HS = "m_axi_in_3_W.data" *)output [255:0] m_axi_in_3_WDATA;
  (* RS_HS = "m_axi_in_3_W.data" *)output m_axi_in_3_WLAST;
  (* RS_HS = "m_axi_in_3_W.ready" *)input m_axi_in_3_WREADY;
  (* RS_HS = "m_axi_in_3_W.data" *)output [31:0] m_axi_in_3_WSTRB;
  (* RS_HS = "m_axi_in_3_W.valid" *)output m_axi_in_3_WVALID;
  (* RS_HS = "m_axi_in_4_AR.data" *)output [63:0] m_axi_in_4_ARADDR;
  (* RS_HS = "m_axi_in_4_AR.data" *)output [1:0] m_axi_in_4_ARBURST;
  (* RS_HS = "m_axi_in_4_AR.data" *)output [3:0] m_axi_in_4_ARCACHE;
  (* RS_HS = "m_axi_in_4_AR.data" *)output [0:0] m_axi_in_4_ARID;
  (* RS_HS = "m_axi_in_4_AR.data" *)output [7:0] m_axi_in_4_ARLEN;
  (* RS_HS = "m_axi_in_4_AR.data" *)output m_axi_in_4_ARLOCK;
  (* RS_HS = "m_axi_in_4_AR.data" *)output [2:0] m_axi_in_4_ARPROT;
  (* RS_HS = "m_axi_in_4_AR.data" *)output [3:0] m_axi_in_4_ARQOS;
  (* RS_HS = "m_axi_in_4_AR.ready" *)input m_axi_in_4_ARREADY;
  (* RS_HS = "m_axi_in_4_AR.data" *)output [2:0] m_axi_in_4_ARSIZE;
  (* RS_HS = "m_axi_in_4_AR.valid" *)output m_axi_in_4_ARVALID;
  (* RS_HS = "m_axi_in_4_AW.data" *)output [63:0] m_axi_in_4_AWADDR;
  (* RS_HS = "m_axi_in_4_AW.data" *)output [1:0] m_axi_in_4_AWBURST;
  (* RS_HS = "m_axi_in_4_AW.data" *)output [3:0] m_axi_in_4_AWCACHE;
  (* RS_HS = "m_axi_in_4_AW.data" *)output [0:0] m_axi_in_4_AWID;
  (* RS_HS = "m_axi_in_4_AW.data" *)output [7:0] m_axi_in_4_AWLEN;
  (* RS_HS = "m_axi_in_4_AW.data" *)output m_axi_in_4_AWLOCK;
  (* RS_HS = "m_axi_in_4_AW.data" *)output [2:0] m_axi_in_4_AWPROT;
  (* RS_HS = "m_axi_in_4_AW.data" *)output [3:0] m_axi_in_4_AWQOS;
  (* RS_HS = "m_axi_in_4_AW.ready" *)input m_axi_in_4_AWREADY;
  (* RS_HS = "m_axi_in_4_AW.data" *)output [2:0] m_axi_in_4_AWSIZE;
  (* RS_HS = "m_axi_in_4_AW.valid" *)output m_axi_in_4_AWVALID;
  (* RS_HS = "m_axi_in_4_B.data" *)input [0:0] m_axi_in_4_BID;
  (* RS_HS = "m_axi_in_4_B.ready" *)output m_axi_in_4_BREADY;
  (* RS_HS = "m_axi_in_4_B.data" *)input [1:0] m_axi_in_4_BRESP;
  (* RS_HS = "m_axi_in_4_B.valid" *)input m_axi_in_4_BVALID;
  (* RS_HS = "m_axi_in_4_R.data" *)input [255:0] m_axi_in_4_RDATA;
  (* RS_HS = "m_axi_in_4_R.data" *)input [0:0] m_axi_in_4_RID;
  (* RS_HS = "m_axi_in_4_R.data" *)input m_axi_in_4_RLAST;
  (* RS_HS = "m_axi_in_4_R.ready" *)output m_axi_in_4_RREADY;
  (* RS_HS = "m_axi_in_4_R.data" *)input [1:0] m_axi_in_4_RRESP;
  (* RS_HS = "m_axi_in_4_R.valid" *)input m_axi_in_4_RVALID;
  (* RS_HS = "m_axi_in_4_W.data" *)output [255:0] m_axi_in_4_WDATA;
  (* RS_HS = "m_axi_in_4_W.data" *)output m_axi_in_4_WLAST;
  (* RS_HS = "m_axi_in_4_W.ready" *)input m_axi_in_4_WREADY;
  (* RS_HS = "m_axi_in_4_W.data" *)output [31:0] m_axi_in_4_WSTRB;
  (* RS_HS = "m_axi_in_4_W.valid" *)output m_axi_in_4_WVALID;
  (* RS_HS = "m_axi_in_5_AR.data" *)output [63:0] m_axi_in_5_ARADDR;
  (* RS_HS = "m_axi_in_5_AR.data" *)output [1:0] m_axi_in_5_ARBURST;
  (* RS_HS = "m_axi_in_5_AR.data" *)output [3:0] m_axi_in_5_ARCACHE;
  (* RS_HS = "m_axi_in_5_AR.data" *)output [0:0] m_axi_in_5_ARID;
  (* RS_HS = "m_axi_in_5_AR.data" *)output [7:0] m_axi_in_5_ARLEN;
  (* RS_HS = "m_axi_in_5_AR.data" *)output m_axi_in_5_ARLOCK;
  (* RS_HS = "m_axi_in_5_AR.data" *)output [2:0] m_axi_in_5_ARPROT;
  (* RS_HS = "m_axi_in_5_AR.data" *)output [3:0] m_axi_in_5_ARQOS;
  (* RS_HS = "m_axi_in_5_AR.ready" *)input m_axi_in_5_ARREADY;
  (* RS_HS = "m_axi_in_5_AR.data" *)output [2:0] m_axi_in_5_ARSIZE;
  (* RS_HS = "m_axi_in_5_AR.valid" *)output m_axi_in_5_ARVALID;
  (* RS_HS = "m_axi_in_5_AW.data" *)output [63:0] m_axi_in_5_AWADDR;
  (* RS_HS = "m_axi_in_5_AW.data" *)output [1:0] m_axi_in_5_AWBURST;
  (* RS_HS = "m_axi_in_5_AW.data" *)output [3:0] m_axi_in_5_AWCACHE;
  (* RS_HS = "m_axi_in_5_AW.data" *)output [0:0] m_axi_in_5_AWID;
  (* RS_HS = "m_axi_in_5_AW.data" *)output [7:0] m_axi_in_5_AWLEN;
  (* RS_HS = "m_axi_in_5_AW.data" *)output m_axi_in_5_AWLOCK;
  (* RS_HS = "m_axi_in_5_AW.data" *)output [2:0] m_axi_in_5_AWPROT;
  (* RS_HS = "m_axi_in_5_AW.data" *)output [3:0] m_axi_in_5_AWQOS;
  (* RS_HS = "m_axi_in_5_AW.ready" *)input m_axi_in_5_AWREADY;
  (* RS_HS = "m_axi_in_5_AW.data" *)output [2:0] m_axi_in_5_AWSIZE;
  (* RS_HS = "m_axi_in_5_AW.valid" *)output m_axi_in_5_AWVALID;
  (* RS_HS = "m_axi_in_5_B.data" *)input [0:0] m_axi_in_5_BID;
  (* RS_HS = "m_axi_in_5_B.ready" *)output m_axi_in_5_BREADY;
  (* RS_HS = "m_axi_in_5_B.data" *)input [1:0] m_axi_in_5_BRESP;
  (* RS_HS = "m_axi_in_5_B.valid" *)input m_axi_in_5_BVALID;
  (* RS_HS = "m_axi_in_5_R.data" *)input [255:0] m_axi_in_5_RDATA;
  (* RS_HS = "m_axi_in_5_R.data" *)input [0:0] m_axi_in_5_RID;
  (* RS_HS = "m_axi_in_5_R.data" *)input m_axi_in_5_RLAST;
  (* RS_HS = "m_axi_in_5_R.ready" *)output m_axi_in_5_RREADY;
  (* RS_HS = "m_axi_in_5_R.data" *)input [1:0] m_axi_in_5_RRESP;
  (* RS_HS = "m_axi_in_5_R.valid" *)input m_axi_in_5_RVALID;
  (* RS_HS = "m_axi_in_5_W.data" *)output [255:0] m_axi_in_5_WDATA;
  (* RS_HS = "m_axi_in_5_W.data" *)output m_axi_in_5_WLAST;
  (* RS_HS = "m_axi_in_5_W.ready" *)input m_axi_in_5_WREADY;
  (* RS_HS = "m_axi_in_5_W.data" *)output [31:0] m_axi_in_5_WSTRB;
  (* RS_HS = "m_axi_in_5_W.valid" *)output m_axi_in_5_WVALID;
  (* RS_HS = "m_axi_in_6_AR.data" *)output [63:0] m_axi_in_6_ARADDR;
  (* RS_HS = "m_axi_in_6_AR.data" *)output [1:0] m_axi_in_6_ARBURST;
  (* RS_HS = "m_axi_in_6_AR.data" *)output [3:0] m_axi_in_6_ARCACHE;
  (* RS_HS = "m_axi_in_6_AR.data" *)output [0:0] m_axi_in_6_ARID;
  (* RS_HS = "m_axi_in_6_AR.data" *)output [7:0] m_axi_in_6_ARLEN;
  (* RS_HS = "m_axi_in_6_AR.data" *)output m_axi_in_6_ARLOCK;
  (* RS_HS = "m_axi_in_6_AR.data" *)output [2:0] m_axi_in_6_ARPROT;
  (* RS_HS = "m_axi_in_6_AR.data" *)output [3:0] m_axi_in_6_ARQOS;
  (* RS_HS = "m_axi_in_6_AR.ready" *)input m_axi_in_6_ARREADY;
  (* RS_HS = "m_axi_in_6_AR.data" *)output [2:0] m_axi_in_6_ARSIZE;
  (* RS_HS = "m_axi_in_6_AR.valid" *)output m_axi_in_6_ARVALID;
  (* RS_HS = "m_axi_in_6_AW.data" *)output [63:0] m_axi_in_6_AWADDR;
  (* RS_HS = "m_axi_in_6_AW.data" *)output [1:0] m_axi_in_6_AWBURST;
  (* RS_HS = "m_axi_in_6_AW.data" *)output [3:0] m_axi_in_6_AWCACHE;
  (* RS_HS = "m_axi_in_6_AW.data" *)output [0:0] m_axi_in_6_AWID;
  (* RS_HS = "m_axi_in_6_AW.data" *)output [7:0] m_axi_in_6_AWLEN;
  (* RS_HS = "m_axi_in_6_AW.data" *)output m_axi_in_6_AWLOCK;
  (* RS_HS = "m_axi_in_6_AW.data" *)output [2:0] m_axi_in_6_AWPROT;
  (* RS_HS = "m_axi_in_6_AW.data" *)output [3:0] m_axi_in_6_AWQOS;
  (* RS_HS = "m_axi_in_6_AW.ready" *)input m_axi_in_6_AWREADY;
  (* RS_HS = "m_axi_in_6_AW.data" *)output [2:0] m_axi_in_6_AWSIZE;
  (* RS_HS = "m_axi_in_6_AW.valid" *)output m_axi_in_6_AWVALID;
  (* RS_HS = "m_axi_in_6_B.data" *)input [0:0] m_axi_in_6_BID;
  (* RS_HS = "m_axi_in_6_B.ready" *)output m_axi_in_6_BREADY;
  (* RS_HS = "m_axi_in_6_B.data" *)input [1:0] m_axi_in_6_BRESP;
  (* RS_HS = "m_axi_in_6_B.valid" *)input m_axi_in_6_BVALID;
  (* RS_HS = "m_axi_in_6_R.data" *)input [255:0] m_axi_in_6_RDATA;
  (* RS_HS = "m_axi_in_6_R.data" *)input [0:0] m_axi_in_6_RID;
  (* RS_HS = "m_axi_in_6_R.data" *)input m_axi_in_6_RLAST;
  (* RS_HS = "m_axi_in_6_R.ready" *)output m_axi_in_6_RREADY;
  (* RS_HS = "m_axi_in_6_R.data" *)input [1:0] m_axi_in_6_RRESP;
  (* RS_HS = "m_axi_in_6_R.valid" *)input m_axi_in_6_RVALID;
  (* RS_HS = "m_axi_in_6_W.data" *)output [255:0] m_axi_in_6_WDATA;
  (* RS_HS = "m_axi_in_6_W.data" *)output m_axi_in_6_WLAST;
  (* RS_HS = "m_axi_in_6_W.ready" *)input m_axi_in_6_WREADY;
  (* RS_HS = "m_axi_in_6_W.data" *)output [31:0] m_axi_in_6_WSTRB;
  (* RS_HS = "m_axi_in_6_W.valid" *)output m_axi_in_6_WVALID;
  (* RS_HS = "m_axi_in_7_AR.data" *)output [63:0] m_axi_in_7_ARADDR;
  (* RS_HS = "m_axi_in_7_AR.data" *)output [1:0] m_axi_in_7_ARBURST;
  (* RS_HS = "m_axi_in_7_AR.data" *)output [3:0] m_axi_in_7_ARCACHE;
  (* RS_HS = "m_axi_in_7_AR.data" *)output [0:0] m_axi_in_7_ARID;
  (* RS_HS = "m_axi_in_7_AR.data" *)output [7:0] m_axi_in_7_ARLEN;
  (* RS_HS = "m_axi_in_7_AR.data" *)output m_axi_in_7_ARLOCK;
  (* RS_HS = "m_axi_in_7_AR.data" *)output [2:0] m_axi_in_7_ARPROT;
  (* RS_HS = "m_axi_in_7_AR.data" *)output [3:0] m_axi_in_7_ARQOS;
  (* RS_HS = "m_axi_in_7_AR.ready" *)input m_axi_in_7_ARREADY;
  (* RS_HS = "m_axi_in_7_AR.data" *)output [2:0] m_axi_in_7_ARSIZE;
  (* RS_HS = "m_axi_in_7_AR.valid" *)output m_axi_in_7_ARVALID;
  (* RS_HS = "m_axi_in_7_AW.data" *)output [63:0] m_axi_in_7_AWADDR;
  (* RS_HS = "m_axi_in_7_AW.data" *)output [1:0] m_axi_in_7_AWBURST;
  (* RS_HS = "m_axi_in_7_AW.data" *)output [3:0] m_axi_in_7_AWCACHE;
  (* RS_HS = "m_axi_in_7_AW.data" *)output [0:0] m_axi_in_7_AWID;
  (* RS_HS = "m_axi_in_7_AW.data" *)output [7:0] m_axi_in_7_AWLEN;
  (* RS_HS = "m_axi_in_7_AW.data" *)output m_axi_in_7_AWLOCK;
  (* RS_HS = "m_axi_in_7_AW.data" *)output [2:0] m_axi_in_7_AWPROT;
  (* RS_HS = "m_axi_in_7_AW.data" *)output [3:0] m_axi_in_7_AWQOS;
  (* RS_HS = "m_axi_in_7_AW.ready" *)input m_axi_in_7_AWREADY;
  (* RS_HS = "m_axi_in_7_AW.data" *)output [2:0] m_axi_in_7_AWSIZE;
  (* RS_HS = "m_axi_in_7_AW.valid" *)output m_axi_in_7_AWVALID;
  (* RS_HS = "m_axi_in_7_B.data" *)input [0:0] m_axi_in_7_BID;
  (* RS_HS = "m_axi_in_7_B.ready" *)output m_axi_in_7_BREADY;
  (* RS_HS = "m_axi_in_7_B.data" *)input [1:0] m_axi_in_7_BRESP;
  (* RS_HS = "m_axi_in_7_B.valid" *)input m_axi_in_7_BVALID;
  (* RS_HS = "m_axi_in_7_R.data" *)input [255:0] m_axi_in_7_RDATA;
  (* RS_HS = "m_axi_in_7_R.data" *)input [0:0] m_axi_in_7_RID;
  (* RS_HS = "m_axi_in_7_R.data" *)input m_axi_in_7_RLAST;
  (* RS_HS = "m_axi_in_7_R.ready" *)output m_axi_in_7_RREADY;
  (* RS_HS = "m_axi_in_7_R.data" *)input [1:0] m_axi_in_7_RRESP;
  (* RS_HS = "m_axi_in_7_R.valid" *)input m_axi_in_7_RVALID;
  (* RS_HS = "m_axi_in_7_W.data" *)output [255:0] m_axi_in_7_WDATA;
  (* RS_HS = "m_axi_in_7_W.data" *)output m_axi_in_7_WLAST;
  (* RS_HS = "m_axi_in_7_W.ready" *)input m_axi_in_7_WREADY;
  (* RS_HS = "m_axi_in_7_W.data" *)output [31:0] m_axi_in_7_WSTRB;
  (* RS_HS = "m_axi_in_7_W.valid" *)output m_axi_in_7_WVALID;
  (* RS_HS = "m_axi_in_8_AR.data" *)output [63:0] m_axi_in_8_ARADDR;
  (* RS_HS = "m_axi_in_8_AR.data" *)output [1:0] m_axi_in_8_ARBURST;
  (* RS_HS = "m_axi_in_8_AR.data" *)output [3:0] m_axi_in_8_ARCACHE;
  (* RS_HS = "m_axi_in_8_AR.data" *)output [0:0] m_axi_in_8_ARID;
  (* RS_HS = "m_axi_in_8_AR.data" *)output [7:0] m_axi_in_8_ARLEN;
  (* RS_HS = "m_axi_in_8_AR.data" *)output m_axi_in_8_ARLOCK;
  (* RS_HS = "m_axi_in_8_AR.data" *)output [2:0] m_axi_in_8_ARPROT;
  (* RS_HS = "m_axi_in_8_AR.data" *)output [3:0] m_axi_in_8_ARQOS;
  (* RS_HS = "m_axi_in_8_AR.ready" *)input m_axi_in_8_ARREADY;
  (* RS_HS = "m_axi_in_8_AR.data" *)output [2:0] m_axi_in_8_ARSIZE;
  (* RS_HS = "m_axi_in_8_AR.valid" *)output m_axi_in_8_ARVALID;
  (* RS_HS = "m_axi_in_8_AW.data" *)output [63:0] m_axi_in_8_AWADDR;
  (* RS_HS = "m_axi_in_8_AW.data" *)output [1:0] m_axi_in_8_AWBURST;
  (* RS_HS = "m_axi_in_8_AW.data" *)output [3:0] m_axi_in_8_AWCACHE;
  (* RS_HS = "m_axi_in_8_AW.data" *)output [0:0] m_axi_in_8_AWID;
  (* RS_HS = "m_axi_in_8_AW.data" *)output [7:0] m_axi_in_8_AWLEN;
  (* RS_HS = "m_axi_in_8_AW.data" *)output m_axi_in_8_AWLOCK;
  (* RS_HS = "m_axi_in_8_AW.data" *)output [2:0] m_axi_in_8_AWPROT;
  (* RS_HS = "m_axi_in_8_AW.data" *)output [3:0] m_axi_in_8_AWQOS;
  (* RS_HS = "m_axi_in_8_AW.ready" *)input m_axi_in_8_AWREADY;
  (* RS_HS = "m_axi_in_8_AW.data" *)output [2:0] m_axi_in_8_AWSIZE;
  (* RS_HS = "m_axi_in_8_AW.valid" *)output m_axi_in_8_AWVALID;
  (* RS_HS = "m_axi_in_8_B.data" *)input [0:0] m_axi_in_8_BID;
  (* RS_HS = "m_axi_in_8_B.ready" *)output m_axi_in_8_BREADY;
  (* RS_HS = "m_axi_in_8_B.data" *)input [1:0] m_axi_in_8_BRESP;
  (* RS_HS = "m_axi_in_8_B.valid" *)input m_axi_in_8_BVALID;
  (* RS_HS = "m_axi_in_8_R.data" *)input [255:0] m_axi_in_8_RDATA;
  (* RS_HS = "m_axi_in_8_R.data" *)input [0:0] m_axi_in_8_RID;
  (* RS_HS = "m_axi_in_8_R.data" *)input m_axi_in_8_RLAST;
  (* RS_HS = "m_axi_in_8_R.ready" *)output m_axi_in_8_RREADY;
  (* RS_HS = "m_axi_in_8_R.data" *)input [1:0] m_axi_in_8_RRESP;
  (* RS_HS = "m_axi_in_8_R.valid" *)input m_axi_in_8_RVALID;
  (* RS_HS = "m_axi_in_8_W.data" *)output [255:0] m_axi_in_8_WDATA;
  (* RS_HS = "m_axi_in_8_W.data" *)output m_axi_in_8_WLAST;
  (* RS_HS = "m_axi_in_8_W.ready" *)input m_axi_in_8_WREADY;
  (* RS_HS = "m_axi_in_8_W.data" *)output [31:0] m_axi_in_8_WSTRB;
  (* RS_HS = "m_axi_in_8_W.valid" *)output m_axi_in_8_WVALID;
  (* RS_HS = "m_axi_in_9_AR.data" *)output [63:0] m_axi_in_9_ARADDR;
  (* RS_HS = "m_axi_in_9_AR.data" *)output [1:0] m_axi_in_9_ARBURST;
  (* RS_HS = "m_axi_in_9_AR.data" *)output [3:0] m_axi_in_9_ARCACHE;
  (* RS_HS = "m_axi_in_9_AR.data" *)output [0:0] m_axi_in_9_ARID;
  (* RS_HS = "m_axi_in_9_AR.data" *)output [7:0] m_axi_in_9_ARLEN;
  (* RS_HS = "m_axi_in_9_AR.data" *)output m_axi_in_9_ARLOCK;
  (* RS_HS = "m_axi_in_9_AR.data" *)output [2:0] m_axi_in_9_ARPROT;
  (* RS_HS = "m_axi_in_9_AR.data" *)output [3:0] m_axi_in_9_ARQOS;
  (* RS_HS = "m_axi_in_9_AR.ready" *)input m_axi_in_9_ARREADY;
  (* RS_HS = "m_axi_in_9_AR.data" *)output [2:0] m_axi_in_9_ARSIZE;
  (* RS_HS = "m_axi_in_9_AR.valid" *)output m_axi_in_9_ARVALID;
  (* RS_HS = "m_axi_in_9_AW.data" *)output [63:0] m_axi_in_9_AWADDR;
  (* RS_HS = "m_axi_in_9_AW.data" *)output [1:0] m_axi_in_9_AWBURST;
  (* RS_HS = "m_axi_in_9_AW.data" *)output [3:0] m_axi_in_9_AWCACHE;
  (* RS_HS = "m_axi_in_9_AW.data" *)output [0:0] m_axi_in_9_AWID;
  (* RS_HS = "m_axi_in_9_AW.data" *)output [7:0] m_axi_in_9_AWLEN;
  (* RS_HS = "m_axi_in_9_AW.data" *)output m_axi_in_9_AWLOCK;
  (* RS_HS = "m_axi_in_9_AW.data" *)output [2:0] m_axi_in_9_AWPROT;
  (* RS_HS = "m_axi_in_9_AW.data" *)output [3:0] m_axi_in_9_AWQOS;
  (* RS_HS = "m_axi_in_9_AW.ready" *)input m_axi_in_9_AWREADY;
  (* RS_HS = "m_axi_in_9_AW.data" *)output [2:0] m_axi_in_9_AWSIZE;
  (* RS_HS = "m_axi_in_9_AW.valid" *)output m_axi_in_9_AWVALID;
  (* RS_HS = "m_axi_in_9_B.data" *)input [0:0] m_axi_in_9_BID;
  (* RS_HS = "m_axi_in_9_B.ready" *)output m_axi_in_9_BREADY;
  (* RS_HS = "m_axi_in_9_B.data" *)input [1:0] m_axi_in_9_BRESP;
  (* RS_HS = "m_axi_in_9_B.valid" *)input m_axi_in_9_BVALID;
  (* RS_HS = "m_axi_in_9_R.data" *)input [255:0] m_axi_in_9_RDATA;
  (* RS_HS = "m_axi_in_9_R.data" *)input [0:0] m_axi_in_9_RID;
  (* RS_HS = "m_axi_in_9_R.data" *)input m_axi_in_9_RLAST;
  (* RS_HS = "m_axi_in_9_R.ready" *)output m_axi_in_9_RREADY;
  (* RS_HS = "m_axi_in_9_R.data" *)input [1:0] m_axi_in_9_RRESP;
  (* RS_HS = "m_axi_in_9_R.valid" *)input m_axi_in_9_RVALID;
  (* RS_HS = "m_axi_in_9_W.data" *)output [255:0] m_axi_in_9_WDATA;
  (* RS_HS = "m_axi_in_9_W.data" *)output m_axi_in_9_WLAST;
  (* RS_HS = "m_axi_in_9_W.ready" *)input m_axi_in_9_WREADY;
  (* RS_HS = "m_axi_in_9_W.data" *)output [31:0] m_axi_in_9_WSTRB;
  (* RS_HS = "m_axi_in_9_W.valid" *)output m_axi_in_9_WVALID;
  wire ap_start;
  wire [63:0] in_0;
  wire [63:0] in_1;
  wire [63:0] in_2;
  wire [63:0] in_3;
  wire [63:0] in_4;
  wire [63:0] in_5;
  wire [63:0] in_6;
  wire [63:0] in_7;
  wire [63:0] in_8;
  wire [63:0] in_9;
  wire [63:0] in_10;
  wire [63:0] in_11;
  wire [63:0] in_12;
  wire [63:0] in_13;
  wire [63:0] in_14;
  wire [63:0] in_15;
  wire [63:0] in_16;
  wire [63:0] in_17;
  wire [63:0] in_18;
  wire [63:0] in_19;
  wire [63:0] in_20;
  wire [63:0] in_21;
  wire [63:0] in_22;
  wire [63:0] in_23;
  wire [63:0] in_24;
  wire [63:0] in_25;
  wire [63:0] in_26;
  wire [63:0] L3_out_dist;
  wire [63:0] L3_out_id;
  wire [65:0] L1_out_dist_0__dout;
  wire L1_out_dist_0__empty_n;
  wire L1_out_dist_0__read;
  wire [65:0] L1_out_dist_0__din;
  wire L1_out_dist_0__full_n;
  wire L1_out_dist_0__write;
  wire [65:0] L1_out_dist_1__dout;
  wire L1_out_dist_1__empty_n;
  wire L1_out_dist_1__read;
  wire [65:0] L1_out_dist_1__din;
  wire L1_out_dist_1__full_n;
  wire L1_out_dist_1__write;
  wire [65:0] L1_out_dist_2__dout;
  wire L1_out_dist_2__empty_n;
  wire L1_out_dist_2__read;
  wire [65:0] L1_out_dist_2__din;
  wire L1_out_dist_2__full_n;
  wire L1_out_dist_2__write;
  wire [65:0] L1_out_dist_3__dout;
  wire L1_out_dist_3__empty_n;
  wire L1_out_dist_3__read;
  wire [65:0] L1_out_dist_3__din;
  wire L1_out_dist_3__full_n;
  wire L1_out_dist_3__write;
  wire [65:0] L1_out_dist_4__dout;
  wire L1_out_dist_4__empty_n;
  wire L1_out_dist_4__read;
  wire [65:0] L1_out_dist_4__din;
  wire L1_out_dist_4__full_n;
  wire L1_out_dist_4__write;
  wire [65:0] L1_out_dist_5__dout;
  wire L1_out_dist_5__empty_n;
  wire L1_out_dist_5__read;
  wire [65:0] L1_out_dist_5__din;
  wire L1_out_dist_5__full_n;
  wire L1_out_dist_5__write;
  wire [65:0] L1_out_dist_6__dout;
  wire L1_out_dist_6__empty_n;
  wire L1_out_dist_6__read;
  wire [65:0] L1_out_dist_6__din;
  wire L1_out_dist_6__full_n;
  wire L1_out_dist_6__write;
  wire [65:0] L1_out_dist_7__dout;
  wire L1_out_dist_7__empty_n;
  wire L1_out_dist_7__read;
  wire [65:0] L1_out_dist_7__din;
  wire L1_out_dist_7__full_n;
  wire L1_out_dist_7__write;
  wire [65:0] L1_out_dist_8__dout;
  wire L1_out_dist_8__empty_n;
  wire L1_out_dist_8__read;
  wire [65:0] L1_out_dist_8__din;
  wire L1_out_dist_8__full_n;
  wire L1_out_dist_8__write;
  wire [65:0] L1_out_id_0__dout;
  wire L1_out_id_0__empty_n;
  wire L1_out_id_0__read;
  wire [65:0] L1_out_id_0__din;
  wire L1_out_id_0__full_n;
  wire L1_out_id_0__write;
  wire [65:0] L1_out_id_1__dout;
  wire L1_out_id_1__empty_n;
  wire L1_out_id_1__read;
  wire [65:0] L1_out_id_1__din;
  wire L1_out_id_1__full_n;
  wire L1_out_id_1__write;
  wire [65:0] L1_out_id_2__dout;
  wire L1_out_id_2__empty_n;
  wire L1_out_id_2__read;
  wire [65:0] L1_out_id_2__din;
  wire L1_out_id_2__full_n;
  wire L1_out_id_2__write;
  wire [65:0] L1_out_id_3__dout;
  wire L1_out_id_3__empty_n;
  wire L1_out_id_3__read;
  wire [65:0] L1_out_id_3__din;
  wire L1_out_id_3__full_n;
  wire L1_out_id_3__write;
  wire [65:0] L1_out_id_4__dout;
  wire L1_out_id_4__empty_n;
  wire L1_out_id_4__read;
  wire [65:0] L1_out_id_4__din;
  wire L1_out_id_4__full_n;
  wire L1_out_id_4__write;
  wire [65:0] L1_out_id_5__dout;
  wire L1_out_id_5__empty_n;
  wire L1_out_id_5__read;
  wire [65:0] L1_out_id_5__din;
  wire L1_out_id_5__full_n;
  wire L1_out_id_5__write;
  wire [65:0] L1_out_id_6__dout;
  wire L1_out_id_6__empty_n;
  wire L1_out_id_6__read;
  wire [65:0] L1_out_id_6__din;
  wire L1_out_id_6__full_n;
  wire L1_out_id_6__write;
  wire [65:0] L1_out_id_7__dout;
  wire L1_out_id_7__empty_n;
  wire L1_out_id_7__read;
  wire [65:0] L1_out_id_7__din;
  wire L1_out_id_7__full_n;
  wire L1_out_id_7__write;
  wire [65:0] L1_out_id_8__dout;
  wire L1_out_id_8__empty_n;
  wire L1_out_id_8__read;
  wire [65:0] L1_out_id_8__din;
  wire L1_out_id_8__full_n;
  wire L1_out_id_8__write;
  wire [65:0] L2_out_dist0__dout;
  wire L2_out_dist0__empty_n;
  wire L2_out_dist0__read;
  wire [65:0] L2_out_dist0__din;
  wire L2_out_dist0__full_n;
  wire L2_out_dist0__write;
  wire [65:0] L2_out_dist1__dout;
  wire L2_out_dist1__empty_n;
  wire L2_out_dist1__read;
  wire [65:0] L2_out_dist1__din;
  wire L2_out_dist1__full_n;
  wire L2_out_dist1__write;
  wire [65:0] L2_out_dist2__dout;
  wire L2_out_dist2__empty_n;
  wire L2_out_dist2__read;
  wire [65:0] L2_out_dist2__din;
  wire L2_out_dist2__full_n;
  wire L2_out_dist2__write;
  wire [65:0] L2_out_id0__dout;
  wire L2_out_id0__empty_n;
  wire L2_out_id0__read;
  wire [65:0] L2_out_id0__din;
  wire L2_out_id0__full_n;
  wire L2_out_id0__write;
  wire [65:0] L2_out_id1__dout;
  wire L2_out_id1__empty_n;
  wire L2_out_id1__read;
  wire [65:0] L2_out_id1__din;
  wire L2_out_id1__full_n;
  wire L2_out_id1__write;
  wire [65:0] L2_out_id2__dout;
  wire L2_out_id2__empty_n;
  wire L2_out_id2__read;
  wire [65:0] L2_out_id2__din;
  wire L2_out_id2__full_n;
  wire L2_out_id2__write;
  wire [65:0] L3_out_dist_stream__dout;
  wire L3_out_dist_stream__empty_n;
  wire L3_out_dist_stream__read;
  wire [65:0] L3_out_dist_stream__din;
  wire L3_out_dist_stream__full_n;
  wire L3_out_dist_stream__write;
  wire [65:0] L3_out_id_stream__dout;
  wire L3_out_id_stream__empty_n;
  wire L3_out_id_stream__read;
  wire [65:0] L3_out_id_stream__din;
  wire L3_out_id_stream__full_n;
  wire L3_out_id_stream__write;
  wire [65:0] out_dist_0__dout;
  wire out_dist_0__empty_n;
  wire out_dist_0__read;
  wire [65:0] out_dist_0__din;
  wire out_dist_0__full_n;
  wire out_dist_0__write;
  wire [65:0] out_dist_10__dout;
  wire out_dist_10__empty_n;
  wire out_dist_10__read;
  wire [65:0] out_dist_10__din;
  wire out_dist_10__full_n;
  wire out_dist_10__write;
  wire [65:0] out_dist_11__dout;
  wire out_dist_11__empty_n;
  wire out_dist_11__read;
  wire [65:0] out_dist_11__din;
  wire out_dist_11__full_n;
  wire out_dist_11__write;
  wire [65:0] out_dist_12__dout;
  wire out_dist_12__empty_n;
  wire out_dist_12__read;
  wire [65:0] out_dist_12__din;
  wire out_dist_12__full_n;
  wire out_dist_12__write;
  wire [65:0] out_dist_13__dout;
  wire out_dist_13__empty_n;
  wire out_dist_13__read;
  wire [65:0] out_dist_13__din;
  wire out_dist_13__full_n;
  wire out_dist_13__write;
  wire [65:0] out_dist_14__dout;
  wire out_dist_14__empty_n;
  wire out_dist_14__read;
  wire [65:0] out_dist_14__din;
  wire out_dist_14__full_n;
  wire out_dist_14__write;
  wire [65:0] out_dist_15__dout;
  wire out_dist_15__empty_n;
  wire out_dist_15__read;
  wire [65:0] out_dist_15__din;
  wire out_dist_15__full_n;
  wire out_dist_15__write;
  wire [65:0] out_dist_16__dout;
  wire out_dist_16__empty_n;
  wire out_dist_16__read;
  wire [65:0] out_dist_16__din;
  wire out_dist_16__full_n;
  wire out_dist_16__write;
  wire [65:0] out_dist_17__dout;
  wire out_dist_17__empty_n;
  wire out_dist_17__read;
  wire [65:0] out_dist_17__din;
  wire out_dist_17__full_n;
  wire out_dist_17__write;
  wire [65:0] out_dist_18__dout;
  wire out_dist_18__empty_n;
  wire out_dist_18__read;
  wire [65:0] out_dist_18__din;
  wire out_dist_18__full_n;
  wire out_dist_18__write;
  wire [65:0] out_dist_19__dout;
  wire out_dist_19__empty_n;
  wire out_dist_19__read;
  wire [65:0] out_dist_19__din;
  wire out_dist_19__full_n;
  wire out_dist_19__write;
  wire [65:0] out_dist_1__dout;
  wire out_dist_1__empty_n;
  wire out_dist_1__read;
  wire [65:0] out_dist_1__din;
  wire out_dist_1__full_n;
  wire out_dist_1__write;
  wire [65:0] out_dist_20__dout;
  wire out_dist_20__empty_n;
  wire out_dist_20__read;
  wire [65:0] out_dist_20__din;
  wire out_dist_20__full_n;
  wire out_dist_20__write;
  wire [65:0] out_dist_21__dout;
  wire out_dist_21__empty_n;
  wire out_dist_21__read;
  wire [65:0] out_dist_21__din;
  wire out_dist_21__full_n;
  wire out_dist_21__write;
  wire [65:0] out_dist_22__dout;
  wire out_dist_22__empty_n;
  wire out_dist_22__read;
  wire [65:0] out_dist_22__din;
  wire out_dist_22__full_n;
  wire out_dist_22__write;
  wire [65:0] out_dist_23__dout;
  wire out_dist_23__empty_n;
  wire out_dist_23__read;
  wire [65:0] out_dist_23__din;
  wire out_dist_23__full_n;
  wire out_dist_23__write;
  wire [65:0] out_dist_24__dout;
  wire out_dist_24__empty_n;
  wire out_dist_24__read;
  wire [65:0] out_dist_24__din;
  wire out_dist_24__full_n;
  wire out_dist_24__write;
  wire [65:0] out_dist_25__dout;
  wire out_dist_25__empty_n;
  wire out_dist_25__read;
  wire [65:0] out_dist_25__din;
  wire out_dist_25__full_n;
  wire out_dist_25__write;
  wire [65:0] out_dist_26__dout;
  wire out_dist_26__empty_n;
  wire out_dist_26__read;
  wire [65:0] out_dist_26__din;
  wire out_dist_26__full_n;
  wire out_dist_26__write;
  wire [65:0] out_dist_2__dout;
  wire out_dist_2__empty_n;
  wire out_dist_2__read;
  wire [65:0] out_dist_2__din;
  wire out_dist_2__full_n;
  wire out_dist_2__write;
  wire [65:0] out_dist_3__dout;
  wire out_dist_3__empty_n;
  wire out_dist_3__read;
  wire [65:0] out_dist_3__din;
  wire out_dist_3__full_n;
  wire out_dist_3__write;
  wire [65:0] out_dist_4__dout;
  wire out_dist_4__empty_n;
  wire out_dist_4__read;
  wire [65:0] out_dist_4__din;
  wire out_dist_4__full_n;
  wire out_dist_4__write;
  wire [65:0] out_dist_5__dout;
  wire out_dist_5__empty_n;
  wire out_dist_5__read;
  wire [65:0] out_dist_5__din;
  wire out_dist_5__full_n;
  wire out_dist_5__write;
  wire [65:0] out_dist_6__dout;
  wire out_dist_6__empty_n;
  wire out_dist_6__read;
  wire [65:0] out_dist_6__din;
  wire out_dist_6__full_n;
  wire out_dist_6__write;
  wire [65:0] out_dist_7__dout;
  wire out_dist_7__empty_n;
  wire out_dist_7__read;
  wire [65:0] out_dist_7__din;
  wire out_dist_7__full_n;
  wire out_dist_7__write;
  wire [65:0] out_dist_8__dout;
  wire out_dist_8__empty_n;
  wire out_dist_8__read;
  wire [65:0] out_dist_8__din;
  wire out_dist_8__full_n;
  wire out_dist_8__write;
  wire [65:0] out_dist_9__dout;
  wire out_dist_9__empty_n;
  wire out_dist_9__read;
  wire [65:0] out_dist_9__din;
  wire out_dist_9__full_n;
  wire out_dist_9__write;
  wire [65:0] out_id_0__dout;
  wire out_id_0__empty_n;
  wire out_id_0__read;
  wire [65:0] out_id_0__din;
  wire out_id_0__full_n;
  wire out_id_0__write;
  wire [65:0] out_id_10__dout;
  wire out_id_10__empty_n;
  wire out_id_10__read;
  wire [65:0] out_id_10__din;
  wire out_id_10__full_n;
  wire out_id_10__write;
  wire [65:0] out_id_11__dout;
  wire out_id_11__empty_n;
  wire out_id_11__read;
  wire [65:0] out_id_11__din;
  wire out_id_11__full_n;
  wire out_id_11__write;
  wire [65:0] out_id_12__dout;
  wire out_id_12__empty_n;
  wire out_id_12__read;
  wire [65:0] out_id_12__din;
  wire out_id_12__full_n;
  wire out_id_12__write;
  wire [65:0] out_id_13__dout;
  wire out_id_13__empty_n;
  wire out_id_13__read;
  wire [65:0] out_id_13__din;
  wire out_id_13__full_n;
  wire out_id_13__write;
  wire [65:0] out_id_14__dout;
  wire out_id_14__empty_n;
  wire out_id_14__read;
  wire [65:0] out_id_14__din;
  wire out_id_14__full_n;
  wire out_id_14__write;
  wire [65:0] out_id_15__dout;
  wire out_id_15__empty_n;
  wire out_id_15__read;
  wire [65:0] out_id_15__din;
  wire out_id_15__full_n;
  wire out_id_15__write;
  wire [65:0] out_id_16__dout;
  wire out_id_16__empty_n;
  wire out_id_16__read;
  wire [65:0] out_id_16__din;
  wire out_id_16__full_n;
  wire out_id_16__write;
  wire [65:0] out_id_17__dout;
  wire out_id_17__empty_n;
  wire out_id_17__read;
  wire [65:0] out_id_17__din;
  wire out_id_17__full_n;
  wire out_id_17__write;
  wire [65:0] out_id_18__dout;
  wire out_id_18__empty_n;
  wire out_id_18__read;
  wire [65:0] out_id_18__din;
  wire out_id_18__full_n;
  wire out_id_18__write;
  wire [65:0] out_id_19__dout;
  wire out_id_19__empty_n;
  wire out_id_19__read;
  wire [65:0] out_id_19__din;
  wire out_id_19__full_n;
  wire out_id_19__write;
  wire [65:0] out_id_1__dout;
  wire out_id_1__empty_n;
  wire out_id_1__read;
  wire [65:0] out_id_1__din;
  wire out_id_1__full_n;
  wire out_id_1__write;
  wire [65:0] out_id_20__dout;
  wire out_id_20__empty_n;
  wire out_id_20__read;
  wire [65:0] out_id_20__din;
  wire out_id_20__full_n;
  wire out_id_20__write;
  wire [65:0] out_id_21__dout;
  wire out_id_21__empty_n;
  wire out_id_21__read;
  wire [65:0] out_id_21__din;
  wire out_id_21__full_n;
  wire out_id_21__write;
  wire [65:0] out_id_22__dout;
  wire out_id_22__empty_n;
  wire out_id_22__read;
  wire [65:0] out_id_22__din;
  wire out_id_22__full_n;
  wire out_id_22__write;
  wire [65:0] out_id_23__dout;
  wire out_id_23__empty_n;
  wire out_id_23__read;
  wire [65:0] out_id_23__din;
  wire out_id_23__full_n;
  wire out_id_23__write;
  wire [65:0] out_id_24__dout;
  wire out_id_24__empty_n;
  wire out_id_24__read;
  wire [65:0] out_id_24__din;
  wire out_id_24__full_n;
  wire out_id_24__write;
  wire [65:0] out_id_25__dout;
  wire out_id_25__empty_n;
  wire out_id_25__read;
  wire [65:0] out_id_25__din;
  wire out_id_25__full_n;
  wire out_id_25__write;
  wire [65:0] out_id_26__dout;
  wire out_id_26__empty_n;
  wire out_id_26__read;
  wire [65:0] out_id_26__din;
  wire out_id_26__full_n;
  wire out_id_26__write;
  wire [65:0] out_id_2__dout;
  wire out_id_2__empty_n;
  wire out_id_2__read;
  wire [65:0] out_id_2__din;
  wire out_id_2__full_n;
  wire out_id_2__write;
  wire [65:0] out_id_3__dout;
  wire out_id_3__empty_n;
  wire out_id_3__read;
  wire [65:0] out_id_3__din;
  wire out_id_3__full_n;
  wire out_id_3__write;
  wire [65:0] out_id_4__dout;
  wire out_id_4__empty_n;
  wire out_id_4__read;
  wire [65:0] out_id_4__din;
  wire out_id_4__full_n;
  wire out_id_4__write;
  wire [65:0] out_id_5__dout;
  wire out_id_5__empty_n;
  wire out_id_5__read;
  wire [65:0] out_id_5__din;
  wire out_id_5__full_n;
  wire out_id_5__write;
  wire [65:0] out_id_6__dout;
  wire out_id_6__empty_n;
  wire out_id_6__read;
  wire [65:0] out_id_6__din;
  wire out_id_6__full_n;
  wire out_id_6__write;
  wire [65:0] out_id_7__dout;
  wire out_id_7__empty_n;
  wire out_id_7__read;
  wire [65:0] out_id_7__din;
  wire out_id_7__full_n;
  wire out_id_7__write;
  wire [65:0] out_id_8__dout;
  wire out_id_8__empty_n;
  wire out_id_8__read;
  wire [65:0] out_id_8__din;
  wire out_id_8__full_n;
  wire out_id_8__write;
  wire [65:0] out_id_9__dout;
  wire out_id_9__empty_n;
  wire out_id_9__read;
  wire [65:0] out_id_9__din;
  wire out_id_9__full_n;
  wire out_id_9__write;
  wire krnl_globalSort_L1_L2_0__ap_start;
  wire krnl_globalSort_L1_L2_0__ap_ready;
  wire krnl_globalSort_L1_L2_0__ap_done;
  wire krnl_globalSort_L1_L2_0__ap_idle;
  wire krnl_globalSort_L1_L2_1__ap_start;
  wire krnl_globalSort_L1_L2_1__ap_ready;
  wire krnl_globalSort_L1_L2_1__ap_done;
  wire krnl_globalSort_L1_L2_1__ap_idle;
  wire krnl_globalSort_L1_L2_2__ap_start;
  wire krnl_globalSort_L1_L2_2__ap_ready;
  wire krnl_globalSort_L1_L2_2__ap_done;
  wire krnl_globalSort_L1_L2_2__ap_idle;
  wire krnl_globalSort_L1_L2_3__ap_start;
  wire krnl_globalSort_L1_L2_3__ap_ready;
  wire krnl_globalSort_L1_L2_3__ap_done;
  wire krnl_globalSort_L1_L2_3__ap_idle;
  wire krnl_globalSort_L1_L2_4__ap_start;
  wire krnl_globalSort_L1_L2_4__ap_ready;
  wire krnl_globalSort_L1_L2_4__ap_done;
  wire krnl_globalSort_L1_L2_4__ap_idle;
  wire krnl_globalSort_L1_L2_5__ap_start;
  wire krnl_globalSort_L1_L2_5__ap_ready;
  wire krnl_globalSort_L1_L2_5__ap_done;
  wire krnl_globalSort_L1_L2_5__ap_idle;
  wire krnl_globalSort_L1_L2_6__ap_start;
  wire krnl_globalSort_L1_L2_6__ap_ready;
  wire krnl_globalSort_L1_L2_6__ap_done;
  wire krnl_globalSort_L1_L2_6__ap_idle;
  wire krnl_globalSort_L1_L2_7__ap_start;
  wire krnl_globalSort_L1_L2_7__ap_ready;
  wire krnl_globalSort_L1_L2_7__ap_done;
  wire krnl_globalSort_L1_L2_7__ap_idle;
  wire krnl_globalSort_L1_L2_8__ap_start;
  wire krnl_globalSort_L1_L2_8__ap_ready;
  wire krnl_globalSort_L1_L2_8__ap_done;
  wire krnl_globalSort_L1_L2_8__ap_idle;
  wire krnl_globalSort_L1_L2_9__ap_start;
  wire krnl_globalSort_L1_L2_9__ap_ready;
  wire krnl_globalSort_L1_L2_9__ap_done;
  wire krnl_globalSort_L1_L2_9__ap_idle;
  wire krnl_globalSort_L1_L2_10__ap_start;
  wire krnl_globalSort_L1_L2_10__ap_ready;
  wire krnl_globalSort_L1_L2_10__ap_done;
  wire krnl_globalSort_L1_L2_10__ap_idle;
  wire krnl_globalSort_L1_L2_11__ap_start;
  wire krnl_globalSort_L1_L2_11__ap_ready;
  wire krnl_globalSort_L1_L2_11__ap_done;
  wire krnl_globalSort_L1_L2_11__ap_idle;
  wire krnl_globalSort_L1_L2_12__ap_start;
  wire krnl_globalSort_L1_L2_12__ap_ready;
  wire krnl_globalSort_L1_L2_12__ap_done;
  wire krnl_globalSort_L1_L2_12__ap_idle;
  wire [63:0] krnl_output_dist_id_0___L3_out_dist__q0;
  wire [63:0] L3_out_dist_read_addr__din;
  wire L3_out_dist_read_addr__full_n;
  wire L3_out_dist_read_addr__write;
  wire [31:0] L3_out_dist_read_data__dout;
  wire L3_out_dist_read_data__empty_n;
  wire L3_out_dist_read_data__read;
  wire [63:0] L3_out_dist_write_addr__din;
  wire L3_out_dist_write_addr__full_n;
  wire L3_out_dist_write_addr__write;
  wire [31:0] L3_out_dist_write_data__din;
  wire L3_out_dist_write_data__full_n;
  wire L3_out_dist_write_data__write;
  wire [7:0] L3_out_dist_write_resp__dout;
  wire L3_out_dist_write_resp__empty_n;
  wire L3_out_dist_write_resp__read;
  wire [63:0] krnl_output_dist_id_0___L3_out_id__q0;
  wire [63:0] L3_out_id_read_addr__din;
  wire L3_out_id_read_addr__full_n;
  wire L3_out_id_read_addr__write;
  wire [31:0] L3_out_id_read_data__dout;
  wire L3_out_id_read_data__empty_n;
  wire L3_out_id_read_data__read;
  wire [63:0] L3_out_id_write_addr__din;
  wire L3_out_id_write_addr__full_n;
  wire L3_out_id_write_addr__write;
  wire [31:0] L3_out_id_write_data__din;
  wire L3_out_id_write_data__full_n;
  wire L3_out_id_write_data__write;
  wire [7:0] L3_out_id_write_resp__dout;
  wire L3_out_id_write_resp__empty_n;
  wire L3_out_id_write_resp__read;
  wire krnl_output_dist_id_0__ap_start;
  wire krnl_output_dist_id_0__ap_ready;
  wire krnl_output_dist_id_0__ap_done;
  wire krnl_output_dist_id_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_0_0___in_0__q0;
  wire [63:0] in_0_read_addr__din;
  wire in_0_read_addr__full_n;
  wire in_0_read_addr__write;
  wire [255:0] in_0_read_data__dout;
  wire in_0_read_data__empty_n;
  wire in_0_read_data__read;
  wire [63:0] in_0_write_addr__din;
  wire in_0_write_addr__full_n;
  wire in_0_write_addr__write;
  wire [255:0] in_0_write_data__din;
  wire in_0_write_data__full_n;
  wire in_0_write_data__write;
  wire [7:0] in_0_write_resp__dout;
  wire in_0_write_resp__empty_n;
  wire in_0_write_resp__read;
  wire krnl_partialKnn_wrapper_0_0__ap_start;
  wire krnl_partialKnn_wrapper_0_0__ap_ready;
  wire krnl_partialKnn_wrapper_0_0__ap_done;
  wire krnl_partialKnn_wrapper_0_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_1_0___in_1__q0;
  wire [63:0] in_1_read_addr__din;
  wire in_1_read_addr__full_n;
  wire in_1_read_addr__write;
  wire [255:0] in_1_read_data__dout;
  wire in_1_read_data__empty_n;
  wire in_1_read_data__read;
  wire [63:0] in_1_write_addr__din;
  wire in_1_write_addr__full_n;
  wire in_1_write_addr__write;
  wire [255:0] in_1_write_data__din;
  wire in_1_write_data__full_n;
  wire in_1_write_data__write;
  wire [7:0] in_1_write_resp__dout;
  wire in_1_write_resp__empty_n;
  wire in_1_write_resp__read;
  wire krnl_partialKnn_wrapper_1_0__ap_start;
  wire krnl_partialKnn_wrapper_1_0__ap_ready;
  wire krnl_partialKnn_wrapper_1_0__ap_done;
  wire krnl_partialKnn_wrapper_1_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_10_0___in_10__q0;
  wire [63:0] in_10_read_addr__din;
  wire in_10_read_addr__full_n;
  wire in_10_read_addr__write;
  wire [255:0] in_10_read_data__dout;
  wire in_10_read_data__empty_n;
  wire in_10_read_data__read;
  wire [63:0] in_10_write_addr__din;
  wire in_10_write_addr__full_n;
  wire in_10_write_addr__write;
  wire [255:0] in_10_write_data__din;
  wire in_10_write_data__full_n;
  wire in_10_write_data__write;
  wire [7:0] in_10_write_resp__dout;
  wire in_10_write_resp__empty_n;
  wire in_10_write_resp__read;
  wire krnl_partialKnn_wrapper_10_0__ap_start;
  wire krnl_partialKnn_wrapper_10_0__ap_ready;
  wire krnl_partialKnn_wrapper_10_0__ap_done;
  wire krnl_partialKnn_wrapper_10_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_11_0___in_11__q0;
  wire [63:0] in_11_read_addr__din;
  wire in_11_read_addr__full_n;
  wire in_11_read_addr__write;
  wire [255:0] in_11_read_data__dout;
  wire in_11_read_data__empty_n;
  wire in_11_read_data__read;
  wire [63:0] in_11_write_addr__din;
  wire in_11_write_addr__full_n;
  wire in_11_write_addr__write;
  wire [255:0] in_11_write_data__din;
  wire in_11_write_data__full_n;
  wire in_11_write_data__write;
  wire [7:0] in_11_write_resp__dout;
  wire in_11_write_resp__empty_n;
  wire in_11_write_resp__read;
  wire krnl_partialKnn_wrapper_11_0__ap_start;
  wire krnl_partialKnn_wrapper_11_0__ap_ready;
  wire krnl_partialKnn_wrapper_11_0__ap_done;
  wire krnl_partialKnn_wrapper_11_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_12_0___in_12__q0;
  wire [63:0] in_12_read_addr__din;
  wire in_12_read_addr__full_n;
  wire in_12_read_addr__write;
  wire [255:0] in_12_read_data__dout;
  wire in_12_read_data__empty_n;
  wire in_12_read_data__read;
  wire [63:0] in_12_write_addr__din;
  wire in_12_write_addr__full_n;
  wire in_12_write_addr__write;
  wire [255:0] in_12_write_data__din;
  wire in_12_write_data__full_n;
  wire in_12_write_data__write;
  wire [7:0] in_12_write_resp__dout;
  wire in_12_write_resp__empty_n;
  wire in_12_write_resp__read;
  wire krnl_partialKnn_wrapper_12_0__ap_start;
  wire krnl_partialKnn_wrapper_12_0__ap_ready;
  wire krnl_partialKnn_wrapper_12_0__ap_done;
  wire krnl_partialKnn_wrapper_12_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_13_0___in_13__q0;
  wire [63:0] in_13_read_addr__din;
  wire in_13_read_addr__full_n;
  wire in_13_read_addr__write;
  wire [255:0] in_13_read_data__dout;
  wire in_13_read_data__empty_n;
  wire in_13_read_data__read;
  wire [63:0] in_13_write_addr__din;
  wire in_13_write_addr__full_n;
  wire in_13_write_addr__write;
  wire [255:0] in_13_write_data__din;
  wire in_13_write_data__full_n;
  wire in_13_write_data__write;
  wire [7:0] in_13_write_resp__dout;
  wire in_13_write_resp__empty_n;
  wire in_13_write_resp__read;
  wire krnl_partialKnn_wrapper_13_0__ap_start;
  wire krnl_partialKnn_wrapper_13_0__ap_ready;
  wire krnl_partialKnn_wrapper_13_0__ap_done;
  wire krnl_partialKnn_wrapper_13_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_14_0___in_14__q0;
  wire [63:0] in_14_read_addr__din;
  wire in_14_read_addr__full_n;
  wire in_14_read_addr__write;
  wire [255:0] in_14_read_data__dout;
  wire in_14_read_data__empty_n;
  wire in_14_read_data__read;
  wire [63:0] in_14_write_addr__din;
  wire in_14_write_addr__full_n;
  wire in_14_write_addr__write;
  wire [255:0] in_14_write_data__din;
  wire in_14_write_data__full_n;
  wire in_14_write_data__write;
  wire [7:0] in_14_write_resp__dout;
  wire in_14_write_resp__empty_n;
  wire in_14_write_resp__read;
  wire krnl_partialKnn_wrapper_14_0__ap_start;
  wire krnl_partialKnn_wrapper_14_0__ap_ready;
  wire krnl_partialKnn_wrapper_14_0__ap_done;
  wire krnl_partialKnn_wrapper_14_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_15_0___in_15__q0;
  wire [63:0] in_15_read_addr__din;
  wire in_15_read_addr__full_n;
  wire in_15_read_addr__write;
  wire [255:0] in_15_read_data__dout;
  wire in_15_read_data__empty_n;
  wire in_15_read_data__read;
  wire [63:0] in_15_write_addr__din;
  wire in_15_write_addr__full_n;
  wire in_15_write_addr__write;
  wire [255:0] in_15_write_data__din;
  wire in_15_write_data__full_n;
  wire in_15_write_data__write;
  wire [7:0] in_15_write_resp__dout;
  wire in_15_write_resp__empty_n;
  wire in_15_write_resp__read;
  wire krnl_partialKnn_wrapper_15_0__ap_start;
  wire krnl_partialKnn_wrapper_15_0__ap_ready;
  wire krnl_partialKnn_wrapper_15_0__ap_done;
  wire krnl_partialKnn_wrapper_15_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_16_0___in_16__q0;
  wire [63:0] in_16_read_addr__din;
  wire in_16_read_addr__full_n;
  wire in_16_read_addr__write;
  wire [255:0] in_16_read_data__dout;
  wire in_16_read_data__empty_n;
  wire in_16_read_data__read;
  wire [63:0] in_16_write_addr__din;
  wire in_16_write_addr__full_n;
  wire in_16_write_addr__write;
  wire [255:0] in_16_write_data__din;
  wire in_16_write_data__full_n;
  wire in_16_write_data__write;
  wire [7:0] in_16_write_resp__dout;
  wire in_16_write_resp__empty_n;
  wire in_16_write_resp__read;
  wire krnl_partialKnn_wrapper_16_0__ap_start;
  wire krnl_partialKnn_wrapper_16_0__ap_ready;
  wire krnl_partialKnn_wrapper_16_0__ap_done;
  wire krnl_partialKnn_wrapper_16_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_17_0___in_17__q0;
  wire [63:0] in_17_read_addr__din;
  wire in_17_read_addr__full_n;
  wire in_17_read_addr__write;
  wire [255:0] in_17_read_data__dout;
  wire in_17_read_data__empty_n;
  wire in_17_read_data__read;
  wire [63:0] in_17_write_addr__din;
  wire in_17_write_addr__full_n;
  wire in_17_write_addr__write;
  wire [255:0] in_17_write_data__din;
  wire in_17_write_data__full_n;
  wire in_17_write_data__write;
  wire [7:0] in_17_write_resp__dout;
  wire in_17_write_resp__empty_n;
  wire in_17_write_resp__read;
  wire krnl_partialKnn_wrapper_17_0__ap_start;
  wire krnl_partialKnn_wrapper_17_0__ap_ready;
  wire krnl_partialKnn_wrapper_17_0__ap_done;
  wire krnl_partialKnn_wrapper_17_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_18_0___in_18__q0;
  wire [63:0] in_18_read_addr__din;
  wire in_18_read_addr__full_n;
  wire in_18_read_addr__write;
  wire [255:0] in_18_read_data__dout;
  wire in_18_read_data__empty_n;
  wire in_18_read_data__read;
  wire [63:0] in_18_write_addr__din;
  wire in_18_write_addr__full_n;
  wire in_18_write_addr__write;
  wire [255:0] in_18_write_data__din;
  wire in_18_write_data__full_n;
  wire in_18_write_data__write;
  wire [7:0] in_18_write_resp__dout;
  wire in_18_write_resp__empty_n;
  wire in_18_write_resp__read;
  wire krnl_partialKnn_wrapper_18_0__ap_start;
  wire krnl_partialKnn_wrapper_18_0__ap_ready;
  wire krnl_partialKnn_wrapper_18_0__ap_done;
  wire krnl_partialKnn_wrapper_18_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_19_0___in_19__q0;
  wire [63:0] in_19_read_addr__din;
  wire in_19_read_addr__full_n;
  wire in_19_read_addr__write;
  wire [255:0] in_19_read_data__dout;
  wire in_19_read_data__empty_n;
  wire in_19_read_data__read;
  wire [63:0] in_19_write_addr__din;
  wire in_19_write_addr__full_n;
  wire in_19_write_addr__write;
  wire [255:0] in_19_write_data__din;
  wire in_19_write_data__full_n;
  wire in_19_write_data__write;
  wire [7:0] in_19_write_resp__dout;
  wire in_19_write_resp__empty_n;
  wire in_19_write_resp__read;
  wire krnl_partialKnn_wrapper_19_0__ap_start;
  wire krnl_partialKnn_wrapper_19_0__ap_ready;
  wire krnl_partialKnn_wrapper_19_0__ap_done;
  wire krnl_partialKnn_wrapper_19_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_2_0___in_2__q0;
  wire [63:0] in_2_read_addr__din;
  wire in_2_read_addr__full_n;
  wire in_2_read_addr__write;
  wire [255:0] in_2_read_data__dout;
  wire in_2_read_data__empty_n;
  wire in_2_read_data__read;
  wire [63:0] in_2_write_addr__din;
  wire in_2_write_addr__full_n;
  wire in_2_write_addr__write;
  wire [255:0] in_2_write_data__din;
  wire in_2_write_data__full_n;
  wire in_2_write_data__write;
  wire [7:0] in_2_write_resp__dout;
  wire in_2_write_resp__empty_n;
  wire in_2_write_resp__read;
  wire krnl_partialKnn_wrapper_2_0__ap_start;
  wire krnl_partialKnn_wrapper_2_0__ap_ready;
  wire krnl_partialKnn_wrapper_2_0__ap_done;
  wire krnl_partialKnn_wrapper_2_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_20_0___in_20__q0;
  wire [63:0] in_20_read_addr__din;
  wire in_20_read_addr__full_n;
  wire in_20_read_addr__write;
  wire [255:0] in_20_read_data__dout;
  wire in_20_read_data__empty_n;
  wire in_20_read_data__read;
  wire [63:0] in_20_write_addr__din;
  wire in_20_write_addr__full_n;
  wire in_20_write_addr__write;
  wire [255:0] in_20_write_data__din;
  wire in_20_write_data__full_n;
  wire in_20_write_data__write;
  wire [7:0] in_20_write_resp__dout;
  wire in_20_write_resp__empty_n;
  wire in_20_write_resp__read;
  wire krnl_partialKnn_wrapper_20_0__ap_start;
  wire krnl_partialKnn_wrapper_20_0__ap_ready;
  wire krnl_partialKnn_wrapper_20_0__ap_done;
  wire krnl_partialKnn_wrapper_20_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_21_0___in_21__q0;
  wire [63:0] in_21_read_addr__din;
  wire in_21_read_addr__full_n;
  wire in_21_read_addr__write;
  wire [255:0] in_21_read_data__dout;
  wire in_21_read_data__empty_n;
  wire in_21_read_data__read;
  wire [63:0] in_21_write_addr__din;
  wire in_21_write_addr__full_n;
  wire in_21_write_addr__write;
  wire [255:0] in_21_write_data__din;
  wire in_21_write_data__full_n;
  wire in_21_write_data__write;
  wire [7:0] in_21_write_resp__dout;
  wire in_21_write_resp__empty_n;
  wire in_21_write_resp__read;
  wire krnl_partialKnn_wrapper_21_0__ap_start;
  wire krnl_partialKnn_wrapper_21_0__ap_ready;
  wire krnl_partialKnn_wrapper_21_0__ap_done;
  wire krnl_partialKnn_wrapper_21_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_22_0___in_22__q0;
  wire [63:0] in_22_read_addr__din;
  wire in_22_read_addr__full_n;
  wire in_22_read_addr__write;
  wire [255:0] in_22_read_data__dout;
  wire in_22_read_data__empty_n;
  wire in_22_read_data__read;
  wire [63:0] in_22_write_addr__din;
  wire in_22_write_addr__full_n;
  wire in_22_write_addr__write;
  wire [255:0] in_22_write_data__din;
  wire in_22_write_data__full_n;
  wire in_22_write_data__write;
  wire [7:0] in_22_write_resp__dout;
  wire in_22_write_resp__empty_n;
  wire in_22_write_resp__read;
  wire krnl_partialKnn_wrapper_22_0__ap_start;
  wire krnl_partialKnn_wrapper_22_0__ap_ready;
  wire krnl_partialKnn_wrapper_22_0__ap_done;
  wire krnl_partialKnn_wrapper_22_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_23_0___in_23__q0;
  wire [63:0] in_23_read_addr__din;
  wire in_23_read_addr__full_n;
  wire in_23_read_addr__write;
  wire [255:0] in_23_read_data__dout;
  wire in_23_read_data__empty_n;
  wire in_23_read_data__read;
  wire [63:0] in_23_write_addr__din;
  wire in_23_write_addr__full_n;
  wire in_23_write_addr__write;
  wire [255:0] in_23_write_data__din;
  wire in_23_write_data__full_n;
  wire in_23_write_data__write;
  wire [7:0] in_23_write_resp__dout;
  wire in_23_write_resp__empty_n;
  wire in_23_write_resp__read;
  wire krnl_partialKnn_wrapper_23_0__ap_start;
  wire krnl_partialKnn_wrapper_23_0__ap_ready;
  wire krnl_partialKnn_wrapper_23_0__ap_done;
  wire krnl_partialKnn_wrapper_23_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_24_0___in_24__q0;
  wire [63:0] in_24_read_addr__din;
  wire in_24_read_addr__full_n;
  wire in_24_read_addr__write;
  wire [255:0] in_24_read_data__dout;
  wire in_24_read_data__empty_n;
  wire in_24_read_data__read;
  wire [63:0] in_24_write_addr__din;
  wire in_24_write_addr__full_n;
  wire in_24_write_addr__write;
  wire [255:0] in_24_write_data__din;
  wire in_24_write_data__full_n;
  wire in_24_write_data__write;
  wire [7:0] in_24_write_resp__dout;
  wire in_24_write_resp__empty_n;
  wire in_24_write_resp__read;
  wire krnl_partialKnn_wrapper_24_0__ap_start;
  wire krnl_partialKnn_wrapper_24_0__ap_ready;
  wire krnl_partialKnn_wrapper_24_0__ap_done;
  wire krnl_partialKnn_wrapper_24_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_25_0___in_25__q0;
  wire [63:0] in_25_read_addr__din;
  wire in_25_read_addr__full_n;
  wire in_25_read_addr__write;
  wire [255:0] in_25_read_data__dout;
  wire in_25_read_data__empty_n;
  wire in_25_read_data__read;
  wire [63:0] in_25_write_addr__din;
  wire in_25_write_addr__full_n;
  wire in_25_write_addr__write;
  wire [255:0] in_25_write_data__din;
  wire in_25_write_data__full_n;
  wire in_25_write_data__write;
  wire [7:0] in_25_write_resp__dout;
  wire in_25_write_resp__empty_n;
  wire in_25_write_resp__read;
  wire krnl_partialKnn_wrapper_25_0__ap_start;
  wire krnl_partialKnn_wrapper_25_0__ap_ready;
  wire krnl_partialKnn_wrapper_25_0__ap_done;
  wire krnl_partialKnn_wrapper_25_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_26_0___in_26__q0;
  wire [63:0] in_26_read_addr__din;
  wire in_26_read_addr__full_n;
  wire in_26_read_addr__write;
  wire [255:0] in_26_read_data__dout;
  wire in_26_read_data__empty_n;
  wire in_26_read_data__read;
  wire [63:0] in_26_write_addr__din;
  wire in_26_write_addr__full_n;
  wire in_26_write_addr__write;
  wire [255:0] in_26_write_data__din;
  wire in_26_write_data__full_n;
  wire in_26_write_data__write;
  wire [7:0] in_26_write_resp__dout;
  wire in_26_write_resp__empty_n;
  wire in_26_write_resp__read;
  wire krnl_partialKnn_wrapper_26_0__ap_start;
  wire krnl_partialKnn_wrapper_26_0__ap_ready;
  wire krnl_partialKnn_wrapper_26_0__ap_done;
  wire krnl_partialKnn_wrapper_26_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_3_0___in_3__q0;
  wire [63:0] in_3_read_addr__din;
  wire in_3_read_addr__full_n;
  wire in_3_read_addr__write;
  wire [255:0] in_3_read_data__dout;
  wire in_3_read_data__empty_n;
  wire in_3_read_data__read;
  wire [63:0] in_3_write_addr__din;
  wire in_3_write_addr__full_n;
  wire in_3_write_addr__write;
  wire [255:0] in_3_write_data__din;
  wire in_3_write_data__full_n;
  wire in_3_write_data__write;
  wire [7:0] in_3_write_resp__dout;
  wire in_3_write_resp__empty_n;
  wire in_3_write_resp__read;
  wire krnl_partialKnn_wrapper_3_0__ap_start;
  wire krnl_partialKnn_wrapper_3_0__ap_ready;
  wire krnl_partialKnn_wrapper_3_0__ap_done;
  wire krnl_partialKnn_wrapper_3_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_4_0___in_4__q0;
  wire [63:0] in_4_read_addr__din;
  wire in_4_read_addr__full_n;
  wire in_4_read_addr__write;
  wire [255:0] in_4_read_data__dout;
  wire in_4_read_data__empty_n;
  wire in_4_read_data__read;
  wire [63:0] in_4_write_addr__din;
  wire in_4_write_addr__full_n;
  wire in_4_write_addr__write;
  wire [255:0] in_4_write_data__din;
  wire in_4_write_data__full_n;
  wire in_4_write_data__write;
  wire [7:0] in_4_write_resp__dout;
  wire in_4_write_resp__empty_n;
  wire in_4_write_resp__read;
  wire krnl_partialKnn_wrapper_4_0__ap_start;
  wire krnl_partialKnn_wrapper_4_0__ap_ready;
  wire krnl_partialKnn_wrapper_4_0__ap_done;
  wire krnl_partialKnn_wrapper_4_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_5_0___in_5__q0;
  wire [63:0] in_5_read_addr__din;
  wire in_5_read_addr__full_n;
  wire in_5_read_addr__write;
  wire [255:0] in_5_read_data__dout;
  wire in_5_read_data__empty_n;
  wire in_5_read_data__read;
  wire [63:0] in_5_write_addr__din;
  wire in_5_write_addr__full_n;
  wire in_5_write_addr__write;
  wire [255:0] in_5_write_data__din;
  wire in_5_write_data__full_n;
  wire in_5_write_data__write;
  wire [7:0] in_5_write_resp__dout;
  wire in_5_write_resp__empty_n;
  wire in_5_write_resp__read;
  wire krnl_partialKnn_wrapper_5_0__ap_start;
  wire krnl_partialKnn_wrapper_5_0__ap_ready;
  wire krnl_partialKnn_wrapper_5_0__ap_done;
  wire krnl_partialKnn_wrapper_5_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_6_0___in_6__q0;
  wire [63:0] in_6_read_addr__din;
  wire in_6_read_addr__full_n;
  wire in_6_read_addr__write;
  wire [255:0] in_6_read_data__dout;
  wire in_6_read_data__empty_n;
  wire in_6_read_data__read;
  wire [63:0] in_6_write_addr__din;
  wire in_6_write_addr__full_n;
  wire in_6_write_addr__write;
  wire [255:0] in_6_write_data__din;
  wire in_6_write_data__full_n;
  wire in_6_write_data__write;
  wire [7:0] in_6_write_resp__dout;
  wire in_6_write_resp__empty_n;
  wire in_6_write_resp__read;
  wire krnl_partialKnn_wrapper_6_0__ap_start;
  wire krnl_partialKnn_wrapper_6_0__ap_ready;
  wire krnl_partialKnn_wrapper_6_0__ap_done;
  wire krnl_partialKnn_wrapper_6_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_7_0___in_7__q0;
  wire [63:0] in_7_read_addr__din;
  wire in_7_read_addr__full_n;
  wire in_7_read_addr__write;
  wire [255:0] in_7_read_data__dout;
  wire in_7_read_data__empty_n;
  wire in_7_read_data__read;
  wire [63:0] in_7_write_addr__din;
  wire in_7_write_addr__full_n;
  wire in_7_write_addr__write;
  wire [255:0] in_7_write_data__din;
  wire in_7_write_data__full_n;
  wire in_7_write_data__write;
  wire [7:0] in_7_write_resp__dout;
  wire in_7_write_resp__empty_n;
  wire in_7_write_resp__read;
  wire krnl_partialKnn_wrapper_7_0__ap_start;
  wire krnl_partialKnn_wrapper_7_0__ap_ready;
  wire krnl_partialKnn_wrapper_7_0__ap_done;
  wire krnl_partialKnn_wrapper_7_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_8_0___in_8__q0;
  wire [63:0] in_8_read_addr__din;
  wire in_8_read_addr__full_n;
  wire in_8_read_addr__write;
  wire [255:0] in_8_read_data__dout;
  wire in_8_read_data__empty_n;
  wire in_8_read_data__read;
  wire [63:0] in_8_write_addr__din;
  wire in_8_write_addr__full_n;
  wire in_8_write_addr__write;
  wire [255:0] in_8_write_data__din;
  wire in_8_write_data__full_n;
  wire in_8_write_data__write;
  wire [7:0] in_8_write_resp__dout;
  wire in_8_write_resp__empty_n;
  wire in_8_write_resp__read;
  wire krnl_partialKnn_wrapper_8_0__ap_start;
  wire krnl_partialKnn_wrapper_8_0__ap_ready;
  wire krnl_partialKnn_wrapper_8_0__ap_done;
  wire krnl_partialKnn_wrapper_8_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_9_0___in_9__q0;
  wire [63:0] in_9_read_addr__din;
  wire in_9_read_addr__full_n;
  wire in_9_read_addr__write;
  wire [255:0] in_9_read_data__dout;
  wire in_9_read_data__empty_n;
  wire in_9_read_data__read;
  wire [63:0] in_9_write_addr__din;
  wire in_9_write_addr__full_n;
  wire in_9_write_addr__write;
  wire [255:0] in_9_write_data__din;
  wire in_9_write_data__full_n;
  wire in_9_write_data__write;
  wire [7:0] in_9_write_resp__dout;
  wire in_9_write_resp__empty_n;
  wire in_9_write_resp__read;
  wire krnl_partialKnn_wrapper_9_0__ap_start;
  wire krnl_partialKnn_wrapper_9_0__ap_ready;
  wire krnl_partialKnn_wrapper_9_0__ap_done;
  wire krnl_partialKnn_wrapper_9_0__ap_idle;
  wire ap_rst_n_inv;
  wire ap_done;
  wire ap_idle;
  wire ap_ready;

  Knn_control_s_axi
  #(
    .C_S_AXI_ADDR_WIDTH(C_S_AXI_CONTROL_ADDR_WIDTH),
    .C_S_AXI_DATA_WIDTH(C_S_AXI_CONTROL_DATA_WIDTH)
  )
  control_s_axi_U
  (
    .AWVALID(s_axi_control_AWVALID),
    .AWREADY(s_axi_control_AWREADY),
    .AWADDR(s_axi_control_AWADDR),
    .WVALID(s_axi_control_WVALID),
    .WREADY(s_axi_control_WREADY),
    .WDATA(s_axi_control_WDATA),
    .WSTRB(s_axi_control_WSTRB),
    .ARVALID(s_axi_control_ARVALID),
    .ARREADY(s_axi_control_ARREADY),
    .ARADDR(s_axi_control_ARADDR),
    .RVALID(s_axi_control_RVALID),
    .RREADY(s_axi_control_RREADY),
    .RDATA(s_axi_control_RDATA),
    .RRESP(s_axi_control_RRESP),
    .BVALID(s_axi_control_BVALID),
    .BREADY(s_axi_control_BREADY),
    .BRESP(s_axi_control_BRESP),
    .ACLK(ap_clk),
    .ARESET(ap_rst_n_inv),
    .ACLK_EN(1'b1),
    .in_0(in_0),
    .in_1(in_1),
    .in_2(in_2),
    .in_3(in_3),
    .in_4(in_4),
    .in_5(in_5),
    .in_6(in_6),
    .in_7(in_7),
    .in_8(in_8),
    .in_9(in_9),
    .in_10(in_10),
    .in_11(in_11),
    .in_12(in_12),
    .in_13(in_13),
    .in_14(in_14),
    .in_15(in_15),
    .in_16(in_16),
    .in_17(in_17),
    .in_18(in_18),
    .in_19(in_19),
    .in_20(in_20),
    .in_21(in_21),
    .in_22(in_22),
    .in_23(in_23),
    .in_24(in_24),
    .in_25(in_25),
    .in_26(in_26),
    .L3_out_dist(L3_out_dist),
    .L3_out_id(L3_out_id),
    .ap_start(ap_start),
    .interrupt(interrupt),
    .ap_ready(ap_ready),
    .ap_done(ap_done),
    .ap_idle(ap_idle)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_dist_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_dist_0__dout),
    .if_empty_n(L1_out_dist_0__empty_n),
    .if_read(L1_out_dist_0__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_dist_0__din),
    .if_full_n(L1_out_dist_0__full_n),
    .if_write(L1_out_dist_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_dist_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_dist_1__dout),
    .if_empty_n(L1_out_dist_1__empty_n),
    .if_read(L1_out_dist_1__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_dist_1__din),
    .if_full_n(L1_out_dist_1__full_n),
    .if_write(L1_out_dist_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_dist_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_dist_2__dout),
    .if_empty_n(L1_out_dist_2__empty_n),
    .if_read(L1_out_dist_2__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_dist_2__din),
    .if_full_n(L1_out_dist_2__full_n),
    .if_write(L1_out_dist_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_dist_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_dist_3__dout),
    .if_empty_n(L1_out_dist_3__empty_n),
    .if_read(L1_out_dist_3__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_dist_3__din),
    .if_full_n(L1_out_dist_3__full_n),
    .if_write(L1_out_dist_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_dist_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_dist_4__dout),
    .if_empty_n(L1_out_dist_4__empty_n),
    .if_read(L1_out_dist_4__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_dist_4__din),
    .if_full_n(L1_out_dist_4__full_n),
    .if_write(L1_out_dist_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_dist_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_dist_5__dout),
    .if_empty_n(L1_out_dist_5__empty_n),
    .if_read(L1_out_dist_5__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_dist_5__din),
    .if_full_n(L1_out_dist_5__full_n),
    .if_write(L1_out_dist_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_dist_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_dist_6__dout),
    .if_empty_n(L1_out_dist_6__empty_n),
    .if_read(L1_out_dist_6__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_dist_6__din),
    .if_full_n(L1_out_dist_6__full_n),
    .if_write(L1_out_dist_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_dist_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_dist_7__dout),
    .if_empty_n(L1_out_dist_7__empty_n),
    .if_read(L1_out_dist_7__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_dist_7__din),
    .if_full_n(L1_out_dist_7__full_n),
    .if_write(L1_out_dist_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_dist_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_dist_8__dout),
    .if_empty_n(L1_out_dist_8__empty_n),
    .if_read(L1_out_dist_8__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_dist_8__din),
    .if_full_n(L1_out_dist_8__full_n),
    .if_write(L1_out_dist_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_id_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_id_0__dout),
    .if_empty_n(L1_out_id_0__empty_n),
    .if_read(L1_out_id_0__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_id_0__din),
    .if_full_n(L1_out_id_0__full_n),
    .if_write(L1_out_id_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_id_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_id_1__dout),
    .if_empty_n(L1_out_id_1__empty_n),
    .if_read(L1_out_id_1__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_id_1__din),
    .if_full_n(L1_out_id_1__full_n),
    .if_write(L1_out_id_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_id_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_id_2__dout),
    .if_empty_n(L1_out_id_2__empty_n),
    .if_read(L1_out_id_2__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_id_2__din),
    .if_full_n(L1_out_id_2__full_n),
    .if_write(L1_out_id_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_id_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_id_3__dout),
    .if_empty_n(L1_out_id_3__empty_n),
    .if_read(L1_out_id_3__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_id_3__din),
    .if_full_n(L1_out_id_3__full_n),
    .if_write(L1_out_id_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_id_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_id_4__dout),
    .if_empty_n(L1_out_id_4__empty_n),
    .if_read(L1_out_id_4__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_id_4__din),
    .if_full_n(L1_out_id_4__full_n),
    .if_write(L1_out_id_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_id_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_id_5__dout),
    .if_empty_n(L1_out_id_5__empty_n),
    .if_read(L1_out_id_5__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_id_5__din),
    .if_full_n(L1_out_id_5__full_n),
    .if_write(L1_out_id_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_id_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_id_6__dout),
    .if_empty_n(L1_out_id_6__empty_n),
    .if_read(L1_out_id_6__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_id_6__din),
    .if_full_n(L1_out_id_6__full_n),
    .if_write(L1_out_id_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_id_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_id_7__dout),
    .if_empty_n(L1_out_id_7__empty_n),
    .if_read(L1_out_id_7__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_id_7__din),
    .if_full_n(L1_out_id_7__full_n),
    .if_write(L1_out_id_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L1_out_id_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L1_out_id_8__dout),
    .if_empty_n(L1_out_id_8__empty_n),
    .if_read(L1_out_id_8__read),
    .if_read_ce(1'b1),
    .if_din(L1_out_id_8__din),
    .if_full_n(L1_out_id_8__full_n),
    .if_write(L1_out_id_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L2_out_dist0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L2_out_dist0__dout),
    .if_empty_n(L2_out_dist0__empty_n),
    .if_read(L2_out_dist0__read),
    .if_read_ce(1'b1),
    .if_din(L2_out_dist0__din),
    .if_full_n(L2_out_dist0__full_n),
    .if_write(L2_out_dist0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L2_out_dist1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L2_out_dist1__dout),
    .if_empty_n(L2_out_dist1__empty_n),
    .if_read(L2_out_dist1__read),
    .if_read_ce(1'b1),
    .if_din(L2_out_dist1__din),
    .if_full_n(L2_out_dist1__full_n),
    .if_write(L2_out_dist1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L2_out_dist2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L2_out_dist2__dout),
    .if_empty_n(L2_out_dist2__empty_n),
    .if_read(L2_out_dist2__read),
    .if_read_ce(1'b1),
    .if_din(L2_out_dist2__din),
    .if_full_n(L2_out_dist2__full_n),
    .if_write(L2_out_dist2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L2_out_id0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L2_out_id0__dout),
    .if_empty_n(L2_out_id0__empty_n),
    .if_read(L2_out_id0__read),
    .if_read_ce(1'b1),
    .if_din(L2_out_id0__din),
    .if_full_n(L2_out_id0__full_n),
    .if_write(L2_out_id0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L2_out_id1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L2_out_id1__dout),
    .if_empty_n(L2_out_id1__empty_n),
    .if_read(L2_out_id1__read),
    .if_read_ce(1'b1),
    .if_din(L2_out_id1__din),
    .if_full_n(L2_out_id1__full_n),
    .if_write(L2_out_id1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L2_out_id2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L2_out_id2__dout),
    .if_empty_n(L2_out_id2__empty_n),
    .if_read(L2_out_id2__read),
    .if_read_ce(1'b1),
    .if_din(L2_out_id2__din),
    .if_full_n(L2_out_id2__full_n),
    .if_write(L2_out_id2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L3_out_dist_stream
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L3_out_dist_stream__dout),
    .if_empty_n(L3_out_dist_stream__empty_n),
    .if_read(L3_out_dist_stream__read),
    .if_read_ce(1'b1),
    .if_din(L3_out_dist_stream__din),
    .if_full_n(L3_out_dist_stream__full_n),
    .if_write(L3_out_dist_stream__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  L3_out_id_stream
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(L3_out_id_stream__dout),
    .if_empty_n(L3_out_id_stream__empty_n),
    .if_read(L3_out_id_stream__read),
    .if_read_ce(1'b1),
    .if_din(L3_out_id_stream__din),
    .if_full_n(L3_out_id_stream__full_n),
    .if_write(L3_out_id_stream__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_0__dout),
    .if_empty_n(out_dist_0__empty_n),
    .if_read(out_dist_0__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_0__din),
    .if_full_n(out_dist_0__full_n),
    .if_write(out_dist_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_10__dout),
    .if_empty_n(out_dist_10__empty_n),
    .if_read(out_dist_10__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_10__din),
    .if_full_n(out_dist_10__full_n),
    .if_write(out_dist_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_11__dout),
    .if_empty_n(out_dist_11__empty_n),
    .if_read(out_dist_11__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_11__din),
    .if_full_n(out_dist_11__full_n),
    .if_write(out_dist_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_12__dout),
    .if_empty_n(out_dist_12__empty_n),
    .if_read(out_dist_12__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_12__din),
    .if_full_n(out_dist_12__full_n),
    .if_write(out_dist_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_13__dout),
    .if_empty_n(out_dist_13__empty_n),
    .if_read(out_dist_13__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_13__din),
    .if_full_n(out_dist_13__full_n),
    .if_write(out_dist_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_14__dout),
    .if_empty_n(out_dist_14__empty_n),
    .if_read(out_dist_14__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_14__din),
    .if_full_n(out_dist_14__full_n),
    .if_write(out_dist_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_15__dout),
    .if_empty_n(out_dist_15__empty_n),
    .if_read(out_dist_15__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_15__din),
    .if_full_n(out_dist_15__full_n),
    .if_write(out_dist_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_16__dout),
    .if_empty_n(out_dist_16__empty_n),
    .if_read(out_dist_16__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_16__din),
    .if_full_n(out_dist_16__full_n),
    .if_write(out_dist_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_17__dout),
    .if_empty_n(out_dist_17__empty_n),
    .if_read(out_dist_17__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_17__din),
    .if_full_n(out_dist_17__full_n),
    .if_write(out_dist_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_18
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_18__dout),
    .if_empty_n(out_dist_18__empty_n),
    .if_read(out_dist_18__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_18__din),
    .if_full_n(out_dist_18__full_n),
    .if_write(out_dist_18__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_19
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_19__dout),
    .if_empty_n(out_dist_19__empty_n),
    .if_read(out_dist_19__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_19__din),
    .if_full_n(out_dist_19__full_n),
    .if_write(out_dist_19__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_1__dout),
    .if_empty_n(out_dist_1__empty_n),
    .if_read(out_dist_1__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_1__din),
    .if_full_n(out_dist_1__full_n),
    .if_write(out_dist_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_20
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_20__dout),
    .if_empty_n(out_dist_20__empty_n),
    .if_read(out_dist_20__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_20__din),
    .if_full_n(out_dist_20__full_n),
    .if_write(out_dist_20__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_21
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_21__dout),
    .if_empty_n(out_dist_21__empty_n),
    .if_read(out_dist_21__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_21__din),
    .if_full_n(out_dist_21__full_n),
    .if_write(out_dist_21__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_22
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_22__dout),
    .if_empty_n(out_dist_22__empty_n),
    .if_read(out_dist_22__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_22__din),
    .if_full_n(out_dist_22__full_n),
    .if_write(out_dist_22__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_23
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_23__dout),
    .if_empty_n(out_dist_23__empty_n),
    .if_read(out_dist_23__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_23__din),
    .if_full_n(out_dist_23__full_n),
    .if_write(out_dist_23__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_24
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_24__dout),
    .if_empty_n(out_dist_24__empty_n),
    .if_read(out_dist_24__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_24__din),
    .if_full_n(out_dist_24__full_n),
    .if_write(out_dist_24__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_25
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_25__dout),
    .if_empty_n(out_dist_25__empty_n),
    .if_read(out_dist_25__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_25__din),
    .if_full_n(out_dist_25__full_n),
    .if_write(out_dist_25__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_26
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_26__dout),
    .if_empty_n(out_dist_26__empty_n),
    .if_read(out_dist_26__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_26__din),
    .if_full_n(out_dist_26__full_n),
    .if_write(out_dist_26__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_2__dout),
    .if_empty_n(out_dist_2__empty_n),
    .if_read(out_dist_2__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_2__din),
    .if_full_n(out_dist_2__full_n),
    .if_write(out_dist_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_3__dout),
    .if_empty_n(out_dist_3__empty_n),
    .if_read(out_dist_3__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_3__din),
    .if_full_n(out_dist_3__full_n),
    .if_write(out_dist_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_4__dout),
    .if_empty_n(out_dist_4__empty_n),
    .if_read(out_dist_4__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_4__din),
    .if_full_n(out_dist_4__full_n),
    .if_write(out_dist_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_5__dout),
    .if_empty_n(out_dist_5__empty_n),
    .if_read(out_dist_5__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_5__din),
    .if_full_n(out_dist_5__full_n),
    .if_write(out_dist_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_6__dout),
    .if_empty_n(out_dist_6__empty_n),
    .if_read(out_dist_6__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_6__din),
    .if_full_n(out_dist_6__full_n),
    .if_write(out_dist_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_7__dout),
    .if_empty_n(out_dist_7__empty_n),
    .if_read(out_dist_7__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_7__din),
    .if_full_n(out_dist_7__full_n),
    .if_write(out_dist_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_8__dout),
    .if_empty_n(out_dist_8__empty_n),
    .if_read(out_dist_8__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_8__din),
    .if_full_n(out_dist_8__full_n),
    .if_write(out_dist_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_dist_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_dist_9__dout),
    .if_empty_n(out_dist_9__empty_n),
    .if_read(out_dist_9__read),
    .if_read_ce(1'b1),
    .if_din(out_dist_9__din),
    .if_full_n(out_dist_9__full_n),
    .if_write(out_dist_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_0
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_0__dout),
    .if_empty_n(out_id_0__empty_n),
    .if_read(out_id_0__read),
    .if_read_ce(1'b1),
    .if_din(out_id_0__din),
    .if_full_n(out_id_0__full_n),
    .if_write(out_id_0__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_10
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_10__dout),
    .if_empty_n(out_id_10__empty_n),
    .if_read(out_id_10__read),
    .if_read_ce(1'b1),
    .if_din(out_id_10__din),
    .if_full_n(out_id_10__full_n),
    .if_write(out_id_10__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_11
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_11__dout),
    .if_empty_n(out_id_11__empty_n),
    .if_read(out_id_11__read),
    .if_read_ce(1'b1),
    .if_din(out_id_11__din),
    .if_full_n(out_id_11__full_n),
    .if_write(out_id_11__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_12
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_12__dout),
    .if_empty_n(out_id_12__empty_n),
    .if_read(out_id_12__read),
    .if_read_ce(1'b1),
    .if_din(out_id_12__din),
    .if_full_n(out_id_12__full_n),
    .if_write(out_id_12__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_13
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_13__dout),
    .if_empty_n(out_id_13__empty_n),
    .if_read(out_id_13__read),
    .if_read_ce(1'b1),
    .if_din(out_id_13__din),
    .if_full_n(out_id_13__full_n),
    .if_write(out_id_13__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_14
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_14__dout),
    .if_empty_n(out_id_14__empty_n),
    .if_read(out_id_14__read),
    .if_read_ce(1'b1),
    .if_din(out_id_14__din),
    .if_full_n(out_id_14__full_n),
    .if_write(out_id_14__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_15
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_15__dout),
    .if_empty_n(out_id_15__empty_n),
    .if_read(out_id_15__read),
    .if_read_ce(1'b1),
    .if_din(out_id_15__din),
    .if_full_n(out_id_15__full_n),
    .if_write(out_id_15__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_16
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_16__dout),
    .if_empty_n(out_id_16__empty_n),
    .if_read(out_id_16__read),
    .if_read_ce(1'b1),
    .if_din(out_id_16__din),
    .if_full_n(out_id_16__full_n),
    .if_write(out_id_16__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_17
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_17__dout),
    .if_empty_n(out_id_17__empty_n),
    .if_read(out_id_17__read),
    .if_read_ce(1'b1),
    .if_din(out_id_17__din),
    .if_full_n(out_id_17__full_n),
    .if_write(out_id_17__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_18
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_18__dout),
    .if_empty_n(out_id_18__empty_n),
    .if_read(out_id_18__read),
    .if_read_ce(1'b1),
    .if_din(out_id_18__din),
    .if_full_n(out_id_18__full_n),
    .if_write(out_id_18__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_19
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_19__dout),
    .if_empty_n(out_id_19__empty_n),
    .if_read(out_id_19__read),
    .if_read_ce(1'b1),
    .if_din(out_id_19__din),
    .if_full_n(out_id_19__full_n),
    .if_write(out_id_19__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_1
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_1__dout),
    .if_empty_n(out_id_1__empty_n),
    .if_read(out_id_1__read),
    .if_read_ce(1'b1),
    .if_din(out_id_1__din),
    .if_full_n(out_id_1__full_n),
    .if_write(out_id_1__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_20
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_20__dout),
    .if_empty_n(out_id_20__empty_n),
    .if_read(out_id_20__read),
    .if_read_ce(1'b1),
    .if_din(out_id_20__din),
    .if_full_n(out_id_20__full_n),
    .if_write(out_id_20__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_21
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_21__dout),
    .if_empty_n(out_id_21__empty_n),
    .if_read(out_id_21__read),
    .if_read_ce(1'b1),
    .if_din(out_id_21__din),
    .if_full_n(out_id_21__full_n),
    .if_write(out_id_21__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_22
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_22__dout),
    .if_empty_n(out_id_22__empty_n),
    .if_read(out_id_22__read),
    .if_read_ce(1'b1),
    .if_din(out_id_22__din),
    .if_full_n(out_id_22__full_n),
    .if_write(out_id_22__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_23
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_23__dout),
    .if_empty_n(out_id_23__empty_n),
    .if_read(out_id_23__read),
    .if_read_ce(1'b1),
    .if_din(out_id_23__din),
    .if_full_n(out_id_23__full_n),
    .if_write(out_id_23__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_24
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_24__dout),
    .if_empty_n(out_id_24__empty_n),
    .if_read(out_id_24__read),
    .if_read_ce(1'b1),
    .if_din(out_id_24__din),
    .if_full_n(out_id_24__full_n),
    .if_write(out_id_24__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_25
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_25__dout),
    .if_empty_n(out_id_25__empty_n),
    .if_read(out_id_25__read),
    .if_read_ce(1'b1),
    .if_din(out_id_25__din),
    .if_full_n(out_id_25__full_n),
    .if_write(out_id_25__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_26
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_26__dout),
    .if_empty_n(out_id_26__empty_n),
    .if_read(out_id_26__read),
    .if_read_ce(1'b1),
    .if_din(out_id_26__din),
    .if_full_n(out_id_26__full_n),
    .if_write(out_id_26__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_2
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_2__dout),
    .if_empty_n(out_id_2__empty_n),
    .if_read(out_id_2__read),
    .if_read_ce(1'b1),
    .if_din(out_id_2__din),
    .if_full_n(out_id_2__full_n),
    .if_write(out_id_2__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_3
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_3__dout),
    .if_empty_n(out_id_3__empty_n),
    .if_read(out_id_3__read),
    .if_read_ce(1'b1),
    .if_din(out_id_3__din),
    .if_full_n(out_id_3__full_n),
    .if_write(out_id_3__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_4
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_4__dout),
    .if_empty_n(out_id_4__empty_n),
    .if_read(out_id_4__read),
    .if_read_ce(1'b1),
    .if_din(out_id_4__din),
    .if_full_n(out_id_4__full_n),
    .if_write(out_id_4__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_5
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_5__dout),
    .if_empty_n(out_id_5__empty_n),
    .if_read(out_id_5__read),
    .if_read_ce(1'b1),
    .if_din(out_id_5__din),
    .if_full_n(out_id_5__full_n),
    .if_write(out_id_5__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_6
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_6__dout),
    .if_empty_n(out_id_6__empty_n),
    .if_read(out_id_6__read),
    .if_read_ce(1'b1),
    .if_din(out_id_6__din),
    .if_full_n(out_id_6__full_n),
    .if_write(out_id_6__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_7
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_7__dout),
    .if_empty_n(out_id_7__empty_n),
    .if_read(out_id_7__read),
    .if_read_ce(1'b1),
    .if_din(out_id_7__din),
    .if_full_n(out_id_7__full_n),
    .if_write(out_id_7__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_8
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_8__dout),
    .if_empty_n(out_id_8__empty_n),
    .if_read(out_id_8__read),
    .if_read_ce(1'b1),
    .if_din(out_id_8__din),
    .if_full_n(out_id_8__full_n),
    .if_write(out_id_8__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) fifo
  #(
    .DATA_WIDTH(66),
    .ADDR_WIDTH(1),
    .DEPTH(2)
  )
  out_id_9
  (
    .clk(ap_clk),
    .reset(~ap_rst_n),
    .if_dout(out_id_9__dout),
    .if_empty_n(out_id_9__empty_n),
    .if_read(out_id_9__read),
    .if_read_ce(1'b1),
    .if_din(out_id_9__din),
    .if_full_n(out_id_9__full_n),
    .if_write(out_id_9__write),
    .if_write_ce(1'b1)
  );


  (* keep_hierarchy = "yes" *) krnl_globalSort_L1_L2
  krnl_globalSort_L1_L2_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_globalSort_L1_L2_0__ap_start),
    .ap_done(krnl_globalSort_L1_L2_0__ap_done),
    .ap_idle(krnl_globalSort_L1_L2_0__ap_idle),
    .ap_ready(krnl_globalSort_L1_L2_0__ap_ready),
    .out_dist_din(L1_out_dist_0__din),
    .out_dist_full_n(L1_out_dist_0__full_n),
    .out_dist_write(L1_out_dist_0__write),
    .out_id_din(L1_out_id_0__din),
    .out_id_full_n(L1_out_id_0__full_n),
    .out_id_write(L1_out_id_0__write),
    .in_dist0_s_dout(out_dist_0__dout),
    .in_dist0_peek_dout(out_dist_0__dout),
    .in_dist0_s_empty_n(out_dist_0__empty_n),
    .in_dist0_peek_empty_n(out_dist_0__empty_n),
    .in_dist0_s_read(out_dist_0__read),
    .in_dist0_peek_read(),
    .in_dist1_s_dout(out_dist_1__dout),
    .in_dist1_peek_dout(out_dist_1__dout),
    .in_dist1_s_empty_n(out_dist_1__empty_n),
    .in_dist1_peek_empty_n(out_dist_1__empty_n),
    .in_dist1_s_read(out_dist_1__read),
    .in_dist1_peek_read(),
    .in_dist2_s_dout(out_dist_2__dout),
    .in_dist2_peek_dout(out_dist_2__dout),
    .in_dist2_s_empty_n(out_dist_2__empty_n),
    .in_dist2_peek_empty_n(out_dist_2__empty_n),
    .in_dist2_s_read(out_dist_2__read),
    .in_dist2_peek_read(),
    .in_id0_s_dout(out_id_0__dout),
    .in_id0_peek_dout(out_id_0__dout),
    .in_id0_s_empty_n(out_id_0__empty_n),
    .in_id0_peek_empty_n(out_id_0__empty_n),
    .in_id0_s_read(out_id_0__read),
    .in_id0_peek_read(),
    .in_id1_s_dout(out_id_1__dout),
    .in_id1_peek_dout(out_id_1__dout),
    .in_id1_s_empty_n(out_id_1__empty_n),
    .in_id1_peek_empty_n(out_id_1__empty_n),
    .in_id1_s_read(out_id_1__read),
    .in_id1_peek_read(),
    .in_id2_s_dout(out_id_2__dout),
    .in_id2_peek_dout(out_id_2__dout),
    .in_id2_s_empty_n(out_id_2__empty_n),
    .in_id2_peek_empty_n(out_id_2__empty_n),
    .in_id2_s_read(out_id_2__read),
    .in_id2_peek_read()
  );


  (* keep_hierarchy = "yes" *) krnl_globalSort_L1_L2
  krnl_globalSort_L1_L2_1
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_globalSort_L1_L2_1__ap_start),
    .ap_done(krnl_globalSort_L1_L2_1__ap_done),
    .ap_idle(krnl_globalSort_L1_L2_1__ap_idle),
    .ap_ready(krnl_globalSort_L1_L2_1__ap_ready),
    .out_dist_din(L1_out_dist_1__din),
    .out_dist_full_n(L1_out_dist_1__full_n),
    .out_dist_write(L1_out_dist_1__write),
    .out_id_din(L1_out_id_1__din),
    .out_id_full_n(L1_out_id_1__full_n),
    .out_id_write(L1_out_id_1__write),
    .in_dist0_s_dout(out_dist_3__dout),
    .in_dist0_peek_dout(out_dist_3__dout),
    .in_dist0_s_empty_n(out_dist_3__empty_n),
    .in_dist0_peek_empty_n(out_dist_3__empty_n),
    .in_dist0_s_read(out_dist_3__read),
    .in_dist0_peek_read(),
    .in_dist1_s_dout(out_dist_4__dout),
    .in_dist1_peek_dout(out_dist_4__dout),
    .in_dist1_s_empty_n(out_dist_4__empty_n),
    .in_dist1_peek_empty_n(out_dist_4__empty_n),
    .in_dist1_s_read(out_dist_4__read),
    .in_dist1_peek_read(),
    .in_dist2_s_dout(out_dist_5__dout),
    .in_dist2_peek_dout(out_dist_5__dout),
    .in_dist2_s_empty_n(out_dist_5__empty_n),
    .in_dist2_peek_empty_n(out_dist_5__empty_n),
    .in_dist2_s_read(out_dist_5__read),
    .in_dist2_peek_read(),
    .in_id0_s_dout(out_id_3__dout),
    .in_id0_peek_dout(out_id_3__dout),
    .in_id0_s_empty_n(out_id_3__empty_n),
    .in_id0_peek_empty_n(out_id_3__empty_n),
    .in_id0_s_read(out_id_3__read),
    .in_id0_peek_read(),
    .in_id1_s_dout(out_id_4__dout),
    .in_id1_peek_dout(out_id_4__dout),
    .in_id1_s_empty_n(out_id_4__empty_n),
    .in_id1_peek_empty_n(out_id_4__empty_n),
    .in_id1_s_read(out_id_4__read),
    .in_id1_peek_read(),
    .in_id2_s_dout(out_id_5__dout),
    .in_id2_peek_dout(out_id_5__dout),
    .in_id2_s_empty_n(out_id_5__empty_n),
    .in_id2_peek_empty_n(out_id_5__empty_n),
    .in_id2_s_read(out_id_5__read),
    .in_id2_peek_read()
  );


  (* keep_hierarchy = "yes" *) krnl_globalSort_L1_L2
  krnl_globalSort_L1_L2_2
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_globalSort_L1_L2_2__ap_start),
    .ap_done(krnl_globalSort_L1_L2_2__ap_done),
    .ap_idle(krnl_globalSort_L1_L2_2__ap_idle),
    .ap_ready(krnl_globalSort_L1_L2_2__ap_ready),
    .out_dist_din(L1_out_dist_2__din),
    .out_dist_full_n(L1_out_dist_2__full_n),
    .out_dist_write(L1_out_dist_2__write),
    .out_id_din(L1_out_id_2__din),
    .out_id_full_n(L1_out_id_2__full_n),
    .out_id_write(L1_out_id_2__write),
    .in_dist0_s_dout(out_dist_6__dout),
    .in_dist0_peek_dout(out_dist_6__dout),
    .in_dist0_s_empty_n(out_dist_6__empty_n),
    .in_dist0_peek_empty_n(out_dist_6__empty_n),
    .in_dist0_s_read(out_dist_6__read),
    .in_dist0_peek_read(),
    .in_dist1_s_dout(out_dist_7__dout),
    .in_dist1_peek_dout(out_dist_7__dout),
    .in_dist1_s_empty_n(out_dist_7__empty_n),
    .in_dist1_peek_empty_n(out_dist_7__empty_n),
    .in_dist1_s_read(out_dist_7__read),
    .in_dist1_peek_read(),
    .in_dist2_s_dout(out_dist_8__dout),
    .in_dist2_peek_dout(out_dist_8__dout),
    .in_dist2_s_empty_n(out_dist_8__empty_n),
    .in_dist2_peek_empty_n(out_dist_8__empty_n),
    .in_dist2_s_read(out_dist_8__read),
    .in_dist2_peek_read(),
    .in_id0_s_dout(out_id_6__dout),
    .in_id0_peek_dout(out_id_6__dout),
    .in_id0_s_empty_n(out_id_6__empty_n),
    .in_id0_peek_empty_n(out_id_6__empty_n),
    .in_id0_s_read(out_id_6__read),
    .in_id0_peek_read(),
    .in_id1_s_dout(out_id_7__dout),
    .in_id1_peek_dout(out_id_7__dout),
    .in_id1_s_empty_n(out_id_7__empty_n),
    .in_id1_peek_empty_n(out_id_7__empty_n),
    .in_id1_s_read(out_id_7__read),
    .in_id1_peek_read(),
    .in_id2_s_dout(out_id_8__dout),
    .in_id2_peek_dout(out_id_8__dout),
    .in_id2_s_empty_n(out_id_8__empty_n),
    .in_id2_peek_empty_n(out_id_8__empty_n),
    .in_id2_s_read(out_id_8__read),
    .in_id2_peek_read()
  );


  (* keep_hierarchy = "yes" *) krnl_globalSort_L1_L2
  krnl_globalSort_L1_L2_3
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_globalSort_L1_L2_3__ap_start),
    .ap_done(krnl_globalSort_L1_L2_3__ap_done),
    .ap_idle(krnl_globalSort_L1_L2_3__ap_idle),
    .ap_ready(krnl_globalSort_L1_L2_3__ap_ready),
    .out_dist_din(L1_out_dist_3__din),
    .out_dist_full_n(L1_out_dist_3__full_n),
    .out_dist_write(L1_out_dist_3__write),
    .out_id_din(L1_out_id_3__din),
    .out_id_full_n(L1_out_id_3__full_n),
    .out_id_write(L1_out_id_3__write),
    .in_dist1_s_dout(out_dist_10__dout),
    .in_dist1_peek_dout(out_dist_10__dout),
    .in_dist1_s_empty_n(out_dist_10__empty_n),
    .in_dist1_peek_empty_n(out_dist_10__empty_n),
    .in_dist1_s_read(out_dist_10__read),
    .in_dist1_peek_read(),
    .in_dist2_s_dout(out_dist_11__dout),
    .in_dist2_peek_dout(out_dist_11__dout),
    .in_dist2_s_empty_n(out_dist_11__empty_n),
    .in_dist2_peek_empty_n(out_dist_11__empty_n),
    .in_dist2_s_read(out_dist_11__read),
    .in_dist2_peek_read(),
    .in_dist0_s_dout(out_dist_9__dout),
    .in_dist0_peek_dout(out_dist_9__dout),
    .in_dist0_s_empty_n(out_dist_9__empty_n),
    .in_dist0_peek_empty_n(out_dist_9__empty_n),
    .in_dist0_s_read(out_dist_9__read),
    .in_dist0_peek_read(),
    .in_id1_s_dout(out_id_10__dout),
    .in_id1_peek_dout(out_id_10__dout),
    .in_id1_s_empty_n(out_id_10__empty_n),
    .in_id1_peek_empty_n(out_id_10__empty_n),
    .in_id1_s_read(out_id_10__read),
    .in_id1_peek_read(),
    .in_id2_s_dout(out_id_11__dout),
    .in_id2_peek_dout(out_id_11__dout),
    .in_id2_s_empty_n(out_id_11__empty_n),
    .in_id2_peek_empty_n(out_id_11__empty_n),
    .in_id2_s_read(out_id_11__read),
    .in_id2_peek_read(),
    .in_id0_s_dout(out_id_9__dout),
    .in_id0_peek_dout(out_id_9__dout),
    .in_id0_s_empty_n(out_id_9__empty_n),
    .in_id0_peek_empty_n(out_id_9__empty_n),
    .in_id0_s_read(out_id_9__read),
    .in_id0_peek_read()
  );


  (* keep_hierarchy = "yes" *) krnl_globalSort_L1_L2
  krnl_globalSort_L1_L2_4
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_globalSort_L1_L2_4__ap_start),
    .ap_done(krnl_globalSort_L1_L2_4__ap_done),
    .ap_idle(krnl_globalSort_L1_L2_4__ap_idle),
    .ap_ready(krnl_globalSort_L1_L2_4__ap_ready),
    .out_dist_din(L1_out_dist_4__din),
    .out_dist_full_n(L1_out_dist_4__full_n),
    .out_dist_write(L1_out_dist_4__write),
    .out_id_din(L1_out_id_4__din),
    .out_id_full_n(L1_out_id_4__full_n),
    .out_id_write(L1_out_id_4__write),
    .in_dist0_s_dout(out_dist_12__dout),
    .in_dist0_peek_dout(out_dist_12__dout),
    .in_dist0_s_empty_n(out_dist_12__empty_n),
    .in_dist0_peek_empty_n(out_dist_12__empty_n),
    .in_dist0_s_read(out_dist_12__read),
    .in_dist0_peek_read(),
    .in_dist1_s_dout(out_dist_13__dout),
    .in_dist1_peek_dout(out_dist_13__dout),
    .in_dist1_s_empty_n(out_dist_13__empty_n),
    .in_dist1_peek_empty_n(out_dist_13__empty_n),
    .in_dist1_s_read(out_dist_13__read),
    .in_dist1_peek_read(),
    .in_dist2_s_dout(out_dist_14__dout),
    .in_dist2_peek_dout(out_dist_14__dout),
    .in_dist2_s_empty_n(out_dist_14__empty_n),
    .in_dist2_peek_empty_n(out_dist_14__empty_n),
    .in_dist2_s_read(out_dist_14__read),
    .in_dist2_peek_read(),
    .in_id0_s_dout(out_id_12__dout),
    .in_id0_peek_dout(out_id_12__dout),
    .in_id0_s_empty_n(out_id_12__empty_n),
    .in_id0_peek_empty_n(out_id_12__empty_n),
    .in_id0_s_read(out_id_12__read),
    .in_id0_peek_read(),
    .in_id1_s_dout(out_id_13__dout),
    .in_id1_peek_dout(out_id_13__dout),
    .in_id1_s_empty_n(out_id_13__empty_n),
    .in_id1_peek_empty_n(out_id_13__empty_n),
    .in_id1_s_read(out_id_13__read),
    .in_id1_peek_read(),
    .in_id2_s_dout(out_id_14__dout),
    .in_id2_peek_dout(out_id_14__dout),
    .in_id2_s_empty_n(out_id_14__empty_n),
    .in_id2_peek_empty_n(out_id_14__empty_n),
    .in_id2_s_read(out_id_14__read),
    .in_id2_peek_read()
  );


  (* keep_hierarchy = "yes" *) krnl_globalSort_L1_L2
  krnl_globalSort_L1_L2_5
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_globalSort_L1_L2_5__ap_start),
    .ap_done(krnl_globalSort_L1_L2_5__ap_done),
    .ap_idle(krnl_globalSort_L1_L2_5__ap_idle),
    .ap_ready(krnl_globalSort_L1_L2_5__ap_ready),
    .out_dist_din(L1_out_dist_5__din),
    .out_dist_full_n(L1_out_dist_5__full_n),
    .out_dist_write(L1_out_dist_5__write),
    .out_id_din(L1_out_id_5__din),
    .out_id_full_n(L1_out_id_5__full_n),
    .out_id_write(L1_out_id_5__write),
    .in_dist0_s_dout(out_dist_15__dout),
    .in_dist0_peek_dout(out_dist_15__dout),
    .in_dist0_s_empty_n(out_dist_15__empty_n),
    .in_dist0_peek_empty_n(out_dist_15__empty_n),
    .in_dist0_s_read(out_dist_15__read),
    .in_dist0_peek_read(),
    .in_dist1_s_dout(out_dist_16__dout),
    .in_dist1_peek_dout(out_dist_16__dout),
    .in_dist1_s_empty_n(out_dist_16__empty_n),
    .in_dist1_peek_empty_n(out_dist_16__empty_n),
    .in_dist1_s_read(out_dist_16__read),
    .in_dist1_peek_read(),
    .in_dist2_s_dout(out_dist_17__dout),
    .in_dist2_peek_dout(out_dist_17__dout),
    .in_dist2_s_empty_n(out_dist_17__empty_n),
    .in_dist2_peek_empty_n(out_dist_17__empty_n),
    .in_dist2_s_read(out_dist_17__read),
    .in_dist2_peek_read(),
    .in_id0_s_dout(out_id_15__dout),
    .in_id0_peek_dout(out_id_15__dout),
    .in_id0_s_empty_n(out_id_15__empty_n),
    .in_id0_peek_empty_n(out_id_15__empty_n),
    .in_id0_s_read(out_id_15__read),
    .in_id0_peek_read(),
    .in_id1_s_dout(out_id_16__dout),
    .in_id1_peek_dout(out_id_16__dout),
    .in_id1_s_empty_n(out_id_16__empty_n),
    .in_id1_peek_empty_n(out_id_16__empty_n),
    .in_id1_s_read(out_id_16__read),
    .in_id1_peek_read(),
    .in_id2_s_dout(out_id_17__dout),
    .in_id2_peek_dout(out_id_17__dout),
    .in_id2_s_empty_n(out_id_17__empty_n),
    .in_id2_peek_empty_n(out_id_17__empty_n),
    .in_id2_s_read(out_id_17__read),
    .in_id2_peek_read()
  );


  (* keep_hierarchy = "yes" *) krnl_globalSort_L1_L2
  krnl_globalSort_L1_L2_6
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_globalSort_L1_L2_6__ap_start),
    .ap_done(krnl_globalSort_L1_L2_6__ap_done),
    .ap_idle(krnl_globalSort_L1_L2_6__ap_idle),
    .ap_ready(krnl_globalSort_L1_L2_6__ap_ready),
    .out_dist_din(L1_out_dist_6__din),
    .out_dist_full_n(L1_out_dist_6__full_n),
    .out_dist_write(L1_out_dist_6__write),
    .out_id_din(L1_out_id_6__din),
    .out_id_full_n(L1_out_id_6__full_n),
    .out_id_write(L1_out_id_6__write),
    .in_dist0_s_dout(out_dist_18__dout),
    .in_dist0_peek_dout(out_dist_18__dout),
    .in_dist0_s_empty_n(out_dist_18__empty_n),
    .in_dist0_peek_empty_n(out_dist_18__empty_n),
    .in_dist0_s_read(out_dist_18__read),
    .in_dist0_peek_read(),
    .in_dist1_s_dout(out_dist_19__dout),
    .in_dist1_peek_dout(out_dist_19__dout),
    .in_dist1_s_empty_n(out_dist_19__empty_n),
    .in_dist1_peek_empty_n(out_dist_19__empty_n),
    .in_dist1_s_read(out_dist_19__read),
    .in_dist1_peek_read(),
    .in_dist2_s_dout(out_dist_20__dout),
    .in_dist2_peek_dout(out_dist_20__dout),
    .in_dist2_s_empty_n(out_dist_20__empty_n),
    .in_dist2_peek_empty_n(out_dist_20__empty_n),
    .in_dist2_s_read(out_dist_20__read),
    .in_dist2_peek_read(),
    .in_id0_s_dout(out_id_18__dout),
    .in_id0_peek_dout(out_id_18__dout),
    .in_id0_s_empty_n(out_id_18__empty_n),
    .in_id0_peek_empty_n(out_id_18__empty_n),
    .in_id0_s_read(out_id_18__read),
    .in_id0_peek_read(),
    .in_id1_s_dout(out_id_19__dout),
    .in_id1_peek_dout(out_id_19__dout),
    .in_id1_s_empty_n(out_id_19__empty_n),
    .in_id1_peek_empty_n(out_id_19__empty_n),
    .in_id1_s_read(out_id_19__read),
    .in_id1_peek_read(),
    .in_id2_s_dout(out_id_20__dout),
    .in_id2_peek_dout(out_id_20__dout),
    .in_id2_s_empty_n(out_id_20__empty_n),
    .in_id2_peek_empty_n(out_id_20__empty_n),
    .in_id2_s_read(out_id_20__read),
    .in_id2_peek_read()
  );


  (* keep_hierarchy = "yes" *) krnl_globalSort_L1_L2
  krnl_globalSort_L1_L2_7
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_globalSort_L1_L2_7__ap_start),
    .ap_done(krnl_globalSort_L1_L2_7__ap_done),
    .ap_idle(krnl_globalSort_L1_L2_7__ap_idle),
    .ap_ready(krnl_globalSort_L1_L2_7__ap_ready),
    .out_dist_din(L1_out_dist_7__din),
    .out_dist_full_n(L1_out_dist_7__full_n),
    .out_dist_write(L1_out_dist_7__write),
    .out_id_din(L1_out_id_7__din),
    .out_id_full_n(L1_out_id_7__full_n),
    .out_id_write(L1_out_id_7__write),
    .in_dist0_s_dout(out_dist_21__dout),
    .in_dist0_peek_dout(out_dist_21__dout),
    .in_dist0_s_empty_n(out_dist_21__empty_n),
    .in_dist0_peek_empty_n(out_dist_21__empty_n),
    .in_dist0_s_read(out_dist_21__read),
    .in_dist0_peek_read(),
    .in_dist1_s_dout(out_dist_22__dout),
    .in_dist1_peek_dout(out_dist_22__dout),
    .in_dist1_s_empty_n(out_dist_22__empty_n),
    .in_dist1_peek_empty_n(out_dist_22__empty_n),
    .in_dist1_s_read(out_dist_22__read),
    .in_dist1_peek_read(),
    .in_dist2_s_dout(out_dist_23__dout),
    .in_dist2_peek_dout(out_dist_23__dout),
    .in_dist2_s_empty_n(out_dist_23__empty_n),
    .in_dist2_peek_empty_n(out_dist_23__empty_n),
    .in_dist2_s_read(out_dist_23__read),
    .in_dist2_peek_read(),
    .in_id0_s_dout(out_id_21__dout),
    .in_id0_peek_dout(out_id_21__dout),
    .in_id0_s_empty_n(out_id_21__empty_n),
    .in_id0_peek_empty_n(out_id_21__empty_n),
    .in_id0_s_read(out_id_21__read),
    .in_id0_peek_read(),
    .in_id1_s_dout(out_id_22__dout),
    .in_id1_peek_dout(out_id_22__dout),
    .in_id1_s_empty_n(out_id_22__empty_n),
    .in_id1_peek_empty_n(out_id_22__empty_n),
    .in_id1_s_read(out_id_22__read),
    .in_id1_peek_read(),
    .in_id2_s_dout(out_id_23__dout),
    .in_id2_peek_dout(out_id_23__dout),
    .in_id2_s_empty_n(out_id_23__empty_n),
    .in_id2_peek_empty_n(out_id_23__empty_n),
    .in_id2_s_read(out_id_23__read),
    .in_id2_peek_read()
  );


  (* keep_hierarchy = "yes" *) krnl_globalSort_L1_L2
  krnl_globalSort_L1_L2_8
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_globalSort_L1_L2_8__ap_start),
    .ap_done(krnl_globalSort_L1_L2_8__ap_done),
    .ap_idle(krnl_globalSort_L1_L2_8__ap_idle),
    .ap_ready(krnl_globalSort_L1_L2_8__ap_ready),
    .out_dist_din(L1_out_dist_8__din),
    .out_dist_full_n(L1_out_dist_8__full_n),
    .out_dist_write(L1_out_dist_8__write),
    .out_id_din(L1_out_id_8__din),
    .out_id_full_n(L1_out_id_8__full_n),
    .out_id_write(L1_out_id_8__write),
    .in_dist0_s_dout(out_dist_24__dout),
    .in_dist0_peek_dout(out_dist_24__dout),
    .in_dist0_s_empty_n(out_dist_24__empty_n),
    .in_dist0_peek_empty_n(out_dist_24__empty_n),
    .in_dist0_s_read(out_dist_24__read),
    .in_dist0_peek_read(),
    .in_dist1_s_dout(out_dist_25__dout),
    .in_dist1_peek_dout(out_dist_25__dout),
    .in_dist1_s_empty_n(out_dist_25__empty_n),
    .in_dist1_peek_empty_n(out_dist_25__empty_n),
    .in_dist1_s_read(out_dist_25__read),
    .in_dist1_peek_read(),
    .in_dist2_s_dout(out_dist_26__dout),
    .in_dist2_peek_dout(out_dist_26__dout),
    .in_dist2_s_empty_n(out_dist_26__empty_n),
    .in_dist2_peek_empty_n(out_dist_26__empty_n),
    .in_dist2_s_read(out_dist_26__read),
    .in_dist2_peek_read(),
    .in_id0_s_dout(out_id_24__dout),
    .in_id0_peek_dout(out_id_24__dout),
    .in_id0_s_empty_n(out_id_24__empty_n),
    .in_id0_peek_empty_n(out_id_24__empty_n),
    .in_id0_s_read(out_id_24__read),
    .in_id0_peek_read(),
    .in_id1_s_dout(out_id_25__dout),
    .in_id1_peek_dout(out_id_25__dout),
    .in_id1_s_empty_n(out_id_25__empty_n),
    .in_id1_peek_empty_n(out_id_25__empty_n),
    .in_id1_s_read(out_id_25__read),
    .in_id1_peek_read(),
    .in_id2_s_dout(out_id_26__dout),
    .in_id2_peek_dout(out_id_26__dout),
    .in_id2_s_empty_n(out_id_26__empty_n),
    .in_id2_peek_empty_n(out_id_26__empty_n),
    .in_id2_s_read(out_id_26__read),
    .in_id2_peek_read()
  );


  (* keep_hierarchy = "yes" *) krnl_globalSort_L1_L2
  krnl_globalSort_L1_L2_9
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_globalSort_L1_L2_9__ap_start),
    .ap_done(krnl_globalSort_L1_L2_9__ap_done),
    .ap_idle(krnl_globalSort_L1_L2_9__ap_idle),
    .ap_ready(krnl_globalSort_L1_L2_9__ap_ready),
    .in_dist0_s_dout(L1_out_dist_0__dout),
    .in_dist0_peek_dout(L1_out_dist_0__dout),
    .in_dist0_s_empty_n(L1_out_dist_0__empty_n),
    .in_dist0_peek_empty_n(L1_out_dist_0__empty_n),
    .in_dist0_s_read(L1_out_dist_0__read),
    .in_dist0_peek_read(),
    .in_dist1_s_dout(L1_out_dist_1__dout),
    .in_dist1_peek_dout(L1_out_dist_1__dout),
    .in_dist1_s_empty_n(L1_out_dist_1__empty_n),
    .in_dist1_peek_empty_n(L1_out_dist_1__empty_n),
    .in_dist1_s_read(L1_out_dist_1__read),
    .in_dist1_peek_read(),
    .in_dist2_s_dout(L1_out_dist_2__dout),
    .in_dist2_peek_dout(L1_out_dist_2__dout),
    .in_dist2_s_empty_n(L1_out_dist_2__empty_n),
    .in_dist2_peek_empty_n(L1_out_dist_2__empty_n),
    .in_dist2_s_read(L1_out_dist_2__read),
    .in_dist2_peek_read(),
    .in_id0_s_dout(L1_out_id_0__dout),
    .in_id0_peek_dout(L1_out_id_0__dout),
    .in_id0_s_empty_n(L1_out_id_0__empty_n),
    .in_id0_peek_empty_n(L1_out_id_0__empty_n),
    .in_id0_s_read(L1_out_id_0__read),
    .in_id0_peek_read(),
    .in_id1_s_dout(L1_out_id_1__dout),
    .in_id1_peek_dout(L1_out_id_1__dout),
    .in_id1_s_empty_n(L1_out_id_1__empty_n),
    .in_id1_peek_empty_n(L1_out_id_1__empty_n),
    .in_id1_s_read(L1_out_id_1__read),
    .in_id1_peek_read(),
    .in_id2_s_dout(L1_out_id_2__dout),
    .in_id2_peek_dout(L1_out_id_2__dout),
    .in_id2_s_empty_n(L1_out_id_2__empty_n),
    .in_id2_peek_empty_n(L1_out_id_2__empty_n),
    .in_id2_s_read(L1_out_id_2__read),
    .in_id2_peek_read(),
    .out_dist_din(L2_out_dist0__din),
    .out_dist_full_n(L2_out_dist0__full_n),
    .out_dist_write(L2_out_dist0__write),
    .out_id_din(L2_out_id0__din),
    .out_id_full_n(L2_out_id0__full_n),
    .out_id_write(L2_out_id0__write)
  );


  (* keep_hierarchy = "yes" *) krnl_globalSort_L1_L2
  krnl_globalSort_L1_L2_10
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_globalSort_L1_L2_10__ap_start),
    .ap_done(krnl_globalSort_L1_L2_10__ap_done),
    .ap_idle(krnl_globalSort_L1_L2_10__ap_idle),
    .ap_ready(krnl_globalSort_L1_L2_10__ap_ready),
    .in_dist0_s_dout(L1_out_dist_3__dout),
    .in_dist0_peek_dout(L1_out_dist_3__dout),
    .in_dist0_s_empty_n(L1_out_dist_3__empty_n),
    .in_dist0_peek_empty_n(L1_out_dist_3__empty_n),
    .in_dist0_s_read(L1_out_dist_3__read),
    .in_dist0_peek_read(),
    .in_dist1_s_dout(L1_out_dist_4__dout),
    .in_dist1_peek_dout(L1_out_dist_4__dout),
    .in_dist1_s_empty_n(L1_out_dist_4__empty_n),
    .in_dist1_peek_empty_n(L1_out_dist_4__empty_n),
    .in_dist1_s_read(L1_out_dist_4__read),
    .in_dist1_peek_read(),
    .in_dist2_s_dout(L1_out_dist_5__dout),
    .in_dist2_peek_dout(L1_out_dist_5__dout),
    .in_dist2_s_empty_n(L1_out_dist_5__empty_n),
    .in_dist2_peek_empty_n(L1_out_dist_5__empty_n),
    .in_dist2_s_read(L1_out_dist_5__read),
    .in_dist2_peek_read(),
    .in_id0_s_dout(L1_out_id_3__dout),
    .in_id0_peek_dout(L1_out_id_3__dout),
    .in_id0_s_empty_n(L1_out_id_3__empty_n),
    .in_id0_peek_empty_n(L1_out_id_3__empty_n),
    .in_id0_s_read(L1_out_id_3__read),
    .in_id0_peek_read(),
    .in_id1_s_dout(L1_out_id_4__dout),
    .in_id1_peek_dout(L1_out_id_4__dout),
    .in_id1_s_empty_n(L1_out_id_4__empty_n),
    .in_id1_peek_empty_n(L1_out_id_4__empty_n),
    .in_id1_s_read(L1_out_id_4__read),
    .in_id1_peek_read(),
    .in_id2_s_dout(L1_out_id_5__dout),
    .in_id2_peek_dout(L1_out_id_5__dout),
    .in_id2_s_empty_n(L1_out_id_5__empty_n),
    .in_id2_peek_empty_n(L1_out_id_5__empty_n),
    .in_id2_s_read(L1_out_id_5__read),
    .in_id2_peek_read(),
    .out_dist_din(L2_out_dist1__din),
    .out_dist_full_n(L2_out_dist1__full_n),
    .out_dist_write(L2_out_dist1__write),
    .out_id_din(L2_out_id1__din),
    .out_id_full_n(L2_out_id1__full_n),
    .out_id_write(L2_out_id1__write)
  );


  (* keep_hierarchy = "yes" *) krnl_globalSort_L1_L2
  krnl_globalSort_L1_L2_11
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_globalSort_L1_L2_11__ap_start),
    .ap_done(krnl_globalSort_L1_L2_11__ap_done),
    .ap_idle(krnl_globalSort_L1_L2_11__ap_idle),
    .ap_ready(krnl_globalSort_L1_L2_11__ap_ready),
    .in_dist0_s_dout(L1_out_dist_6__dout),
    .in_dist0_peek_dout(L1_out_dist_6__dout),
    .in_dist0_s_empty_n(L1_out_dist_6__empty_n),
    .in_dist0_peek_empty_n(L1_out_dist_6__empty_n),
    .in_dist0_s_read(L1_out_dist_6__read),
    .in_dist0_peek_read(),
    .in_dist1_s_dout(L1_out_dist_7__dout),
    .in_dist1_peek_dout(L1_out_dist_7__dout),
    .in_dist1_s_empty_n(L1_out_dist_7__empty_n),
    .in_dist1_peek_empty_n(L1_out_dist_7__empty_n),
    .in_dist1_s_read(L1_out_dist_7__read),
    .in_dist1_peek_read(),
    .in_dist2_s_dout(L1_out_dist_8__dout),
    .in_dist2_peek_dout(L1_out_dist_8__dout),
    .in_dist2_s_empty_n(L1_out_dist_8__empty_n),
    .in_dist2_peek_empty_n(L1_out_dist_8__empty_n),
    .in_dist2_s_read(L1_out_dist_8__read),
    .in_dist2_peek_read(),
    .in_id0_s_dout(L1_out_id_6__dout),
    .in_id0_peek_dout(L1_out_id_6__dout),
    .in_id0_s_empty_n(L1_out_id_6__empty_n),
    .in_id0_peek_empty_n(L1_out_id_6__empty_n),
    .in_id0_s_read(L1_out_id_6__read),
    .in_id0_peek_read(),
    .in_id1_s_dout(L1_out_id_7__dout),
    .in_id1_peek_dout(L1_out_id_7__dout),
    .in_id1_s_empty_n(L1_out_id_7__empty_n),
    .in_id1_peek_empty_n(L1_out_id_7__empty_n),
    .in_id1_s_read(L1_out_id_7__read),
    .in_id1_peek_read(),
    .in_id2_s_dout(L1_out_id_8__dout),
    .in_id2_peek_dout(L1_out_id_8__dout),
    .in_id2_s_empty_n(L1_out_id_8__empty_n),
    .in_id2_peek_empty_n(L1_out_id_8__empty_n),
    .in_id2_s_read(L1_out_id_8__read),
    .in_id2_peek_read(),
    .out_dist_din(L2_out_dist2__din),
    .out_dist_full_n(L2_out_dist2__full_n),
    .out_dist_write(L2_out_dist2__write),
    .out_id_din(L2_out_id2__din),
    .out_id_full_n(L2_out_id2__full_n),
    .out_id_write(L2_out_id2__write)
  );


  (* keep_hierarchy = "yes" *) krnl_globalSort_L1_L2
  krnl_globalSort_L1_L2_12
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_globalSort_L1_L2_12__ap_start),
    .ap_done(krnl_globalSort_L1_L2_12__ap_done),
    .ap_idle(krnl_globalSort_L1_L2_12__ap_idle),
    .ap_ready(krnl_globalSort_L1_L2_12__ap_ready),
    .in_dist0_s_dout(L2_out_dist0__dout),
    .in_dist0_peek_dout(L2_out_dist0__dout),
    .in_dist0_s_empty_n(L2_out_dist0__empty_n),
    .in_dist0_peek_empty_n(L2_out_dist0__empty_n),
    .in_dist0_s_read(L2_out_dist0__read),
    .in_dist0_peek_read(),
    .in_dist1_s_dout(L2_out_dist1__dout),
    .in_dist1_peek_dout(L2_out_dist1__dout),
    .in_dist1_s_empty_n(L2_out_dist1__empty_n),
    .in_dist1_peek_empty_n(L2_out_dist1__empty_n),
    .in_dist1_s_read(L2_out_dist1__read),
    .in_dist1_peek_read(),
    .in_dist2_s_dout(L2_out_dist2__dout),
    .in_dist2_peek_dout(L2_out_dist2__dout),
    .in_dist2_s_empty_n(L2_out_dist2__empty_n),
    .in_dist2_peek_empty_n(L2_out_dist2__empty_n),
    .in_dist2_s_read(L2_out_dist2__read),
    .in_dist2_peek_read(),
    .in_id0_s_dout(L2_out_id0__dout),
    .in_id0_peek_dout(L2_out_id0__dout),
    .in_id0_s_empty_n(L2_out_id0__empty_n),
    .in_id0_peek_empty_n(L2_out_id0__empty_n),
    .in_id0_s_read(L2_out_id0__read),
    .in_id0_peek_read(),
    .in_id1_s_dout(L2_out_id1__dout),
    .in_id1_peek_dout(L2_out_id1__dout),
    .in_id1_s_empty_n(L2_out_id1__empty_n),
    .in_id1_peek_empty_n(L2_out_id1__empty_n),
    .in_id1_s_read(L2_out_id1__read),
    .in_id1_peek_read(),
    .in_id2_s_dout(L2_out_id2__dout),
    .in_id2_peek_dout(L2_out_id2__dout),
    .in_id2_s_empty_n(L2_out_id2__empty_n),
    .in_id2_peek_empty_n(L2_out_id2__empty_n),
    .in_id2_s_read(L2_out_id2__read),
    .in_id2_peek_read(),
    .out_dist_din(L3_out_dist_stream__din),
    .out_dist_full_n(L3_out_dist_stream__full_n),
    .out_dist_write(L3_out_dist_stream__write),
    .out_id_din(L3_out_id_stream__din),
    .out_id_full_n(L3_out_id_stream__full_n),
    .out_id_write(L3_out_id_stream__write)
  );


  (* keep_hierarchy = "yes" *) krnl_output_dist_id
  krnl_output_dist_id_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_output_dist_id_0__ap_start),
    .ap_done(krnl_output_dist_id_0__ap_done),
    .ap_idle(krnl_output_dist_id_0__ap_idle),
    .ap_ready(krnl_output_dist_id_0__ap_ready),
    .output_knnDist_read_addr_s_din(L3_out_dist_read_addr__din),
    .output_knnDist_read_addr_s_full_n(L3_out_dist_read_addr__full_n),
    .output_knnDist_read_addr_s_write(L3_out_dist_read_addr__write),
    .output_knnDist_read_addr_offset(krnl_output_dist_id_0___L3_out_dist__q0),
    .output_knnDist_read_data_s_dout({1'b0, L3_out_dist_read_data__dout}),
    .output_knnDist_read_data_peek_dout({1'b0, L3_out_dist_read_data__dout}),
    .output_knnDist_read_data_s_empty_n(L3_out_dist_read_data__empty_n),
    .output_knnDist_read_data_peek_empty_n(L3_out_dist_read_data__empty_n),
    .output_knnDist_read_data_s_read(L3_out_dist_read_data__read),
    .output_knnDist_read_data_peek_read(),
    .output_knnDist_write_addr_s_din(L3_out_dist_write_addr__din),
    .output_knnDist_write_addr_s_full_n(L3_out_dist_write_addr__full_n),
    .output_knnDist_write_addr_s_write(L3_out_dist_write_addr__write),
    .output_knnDist_write_addr_offset(krnl_output_dist_id_0___L3_out_dist__q0),
    .output_knnDist_write_data_din(L3_out_dist_write_data__din),
    .output_knnDist_write_data_full_n(L3_out_dist_write_data__full_n),
    .output_knnDist_write_data_write(L3_out_dist_write_data__write),
    .output_knnDist_write_resp_s_dout({1'b0, L3_out_dist_write_resp__dout}),
    .output_knnDist_write_resp_peek_dout({1'b0, L3_out_dist_write_resp__dout}),
    .output_knnDist_write_resp_s_empty_n(L3_out_dist_write_resp__empty_n),
    .output_knnDist_write_resp_peek_empty_n(L3_out_dist_write_resp__empty_n),
    .output_knnDist_write_resp_s_read(L3_out_dist_write_resp__read),
    .output_knnDist_write_resp_peek_read(),
    .in_dist_s_dout(L3_out_dist_stream__dout),
    .in_dist_peek_dout(L3_out_dist_stream__dout),
    .in_dist_s_empty_n(L3_out_dist_stream__empty_n),
    .in_dist_peek_empty_n(L3_out_dist_stream__empty_n),
    .in_dist_s_read(L3_out_dist_stream__read),
    .in_dist_peek_read(),
    .output_knnId_read_addr_s_din(L3_out_id_read_addr__din),
    .output_knnId_read_addr_s_full_n(L3_out_id_read_addr__full_n),
    .output_knnId_read_addr_s_write(L3_out_id_read_addr__write),
    .output_knnId_read_addr_offset(krnl_output_dist_id_0___L3_out_id__q0),
    .output_knnId_read_data_s_dout({1'b0, L3_out_id_read_data__dout}),
    .output_knnId_read_data_peek_dout({1'b0, L3_out_id_read_data__dout}),
    .output_knnId_read_data_s_empty_n(L3_out_id_read_data__empty_n),
    .output_knnId_read_data_peek_empty_n(L3_out_id_read_data__empty_n),
    .output_knnId_read_data_s_read(L3_out_id_read_data__read),
    .output_knnId_read_data_peek_read(),
    .output_knnId_write_addr_s_din(L3_out_id_write_addr__din),
    .output_knnId_write_addr_s_full_n(L3_out_id_write_addr__full_n),
    .output_knnId_write_addr_s_write(L3_out_id_write_addr__write),
    .output_knnId_write_addr_offset(krnl_output_dist_id_0___L3_out_id__q0),
    .output_knnId_write_data_din(L3_out_id_write_data__din),
    .output_knnId_write_data_full_n(L3_out_id_write_data__full_n),
    .output_knnId_write_data_write(L3_out_id_write_data__write),
    .output_knnId_write_resp_s_dout({1'b0, L3_out_id_write_resp__dout}),
    .output_knnId_write_resp_peek_dout({1'b0, L3_out_id_write_resp__dout}),
    .output_knnId_write_resp_s_empty_n(L3_out_id_write_resp__empty_n),
    .output_knnId_write_resp_peek_empty_n(L3_out_id_write_resp__empty_n),
    .output_knnId_write_resp_s_read(L3_out_id_write_resp__read),
    .output_knnId_write_resp_peek_read(),
    .in_id_s_dout(L3_out_id_stream__dout),
    .in_id_peek_dout(L3_out_id_stream__dout),
    .in_id_s_empty_n(L3_out_id_stream__empty_n),
    .in_id_peek_empty_n(L3_out_id_stream__empty_n),
    .in_id_s_read(L3_out_id_stream__read),
    .in_id_peek_read()
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_0
  krnl_partialKnn_wrapper_0_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_0_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_0_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_0_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_0_0__ap_ready),
    .start_id_0(64'd0),
    .searchSpace_0_read_addr_s_din(in_0_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_0_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_0_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_0_0___in_0__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_0_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_0_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_0_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_0_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_0_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_0_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_0_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_0_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_0_0___in_0__q0),
    .searchSpace_0_write_data_din(in_0_write_data__din),
    .searchSpace_0_write_data_full_n(in_0_write_data__full_n),
    .searchSpace_0_write_data_write(in_0_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_0_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_0_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_0_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_0_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_0_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_0__din),
    .out_dist_full_n(out_dist_0__full_n),
    .out_dist_write(out_dist_0__write),
    .out_id_din(out_id_0__din),
    .out_id_full_n(out_id_0__full_n),
    .out_id_write(out_id_0__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_1
  krnl_partialKnn_wrapper_1_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_1_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_1_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_1_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_1_0__ap_ready),
    .start_id_0(64'd8192),
    .searchSpace_0_read_addr_s_din(in_1_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_1_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_1_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_1_0___in_1__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_1_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_1_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_1_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_1_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_1_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_1_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_1_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_1_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_1_0___in_1__q0),
    .searchSpace_0_write_data_din(in_1_write_data__din),
    .searchSpace_0_write_data_full_n(in_1_write_data__full_n),
    .searchSpace_0_write_data_write(in_1_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_1_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_1_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_1_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_1_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_1_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_1__din),
    .out_dist_full_n(out_dist_1__full_n),
    .out_dist_write(out_dist_1__write),
    .out_id_din(out_id_1__din),
    .out_id_full_n(out_id_1__full_n),
    .out_id_write(out_id_1__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_10
  krnl_partialKnn_wrapper_10_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_10_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_10_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_10_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_10_0__ap_ready),
    .start_id_0(64'd81920),
    .searchSpace_0_read_addr_s_din(in_10_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_10_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_10_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_10_0___in_10__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_10_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_10_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_10_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_10_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_10_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_10_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_10_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_10_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_10_0___in_10__q0),
    .searchSpace_0_write_data_din(in_10_write_data__din),
    .searchSpace_0_write_data_full_n(in_10_write_data__full_n),
    .searchSpace_0_write_data_write(in_10_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_10_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_10_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_10_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_10_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_10_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_10__din),
    .out_dist_full_n(out_dist_10__full_n),
    .out_dist_write(out_dist_10__write),
    .out_id_din(out_id_10__din),
    .out_id_full_n(out_id_10__full_n),
    .out_id_write(out_id_10__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_11
  krnl_partialKnn_wrapper_11_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_11_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_11_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_11_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_11_0__ap_ready),
    .start_id_0(64'd90112),
    .searchSpace_0_read_addr_s_din(in_11_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_11_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_11_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_11_0___in_11__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_11_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_11_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_11_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_11_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_11_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_11_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_11_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_11_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_11_0___in_11__q0),
    .searchSpace_0_write_data_din(in_11_write_data__din),
    .searchSpace_0_write_data_full_n(in_11_write_data__full_n),
    .searchSpace_0_write_data_write(in_11_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_11_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_11_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_11_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_11_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_11_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_11__din),
    .out_dist_full_n(out_dist_11__full_n),
    .out_dist_write(out_dist_11__write),
    .out_id_din(out_id_11__din),
    .out_id_full_n(out_id_11__full_n),
    .out_id_write(out_id_11__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_12
  krnl_partialKnn_wrapper_12_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_12_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_12_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_12_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_12_0__ap_ready),
    .start_id_0(64'd98304),
    .searchSpace_0_read_addr_s_din(in_12_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_12_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_12_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_12_0___in_12__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_12_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_12_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_12_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_12_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_12_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_12_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_12_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_12_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_12_0___in_12__q0),
    .searchSpace_0_write_data_din(in_12_write_data__din),
    .searchSpace_0_write_data_full_n(in_12_write_data__full_n),
    .searchSpace_0_write_data_write(in_12_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_12_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_12_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_12_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_12_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_12_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_12__din),
    .out_dist_full_n(out_dist_12__full_n),
    .out_dist_write(out_dist_12__write),
    .out_id_din(out_id_12__din),
    .out_id_full_n(out_id_12__full_n),
    .out_id_write(out_id_12__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_13
  krnl_partialKnn_wrapper_13_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_13_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_13_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_13_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_13_0__ap_ready),
    .start_id_0(64'd106496),
    .searchSpace_0_read_addr_s_din(in_13_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_13_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_13_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_13_0___in_13__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_13_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_13_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_13_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_13_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_13_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_13_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_13_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_13_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_13_0___in_13__q0),
    .searchSpace_0_write_data_din(in_13_write_data__din),
    .searchSpace_0_write_data_full_n(in_13_write_data__full_n),
    .searchSpace_0_write_data_write(in_13_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_13_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_13_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_13_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_13_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_13_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_13__din),
    .out_dist_full_n(out_dist_13__full_n),
    .out_dist_write(out_dist_13__write),
    .out_id_din(out_id_13__din),
    .out_id_full_n(out_id_13__full_n),
    .out_id_write(out_id_13__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_14
  krnl_partialKnn_wrapper_14_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_14_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_14_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_14_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_14_0__ap_ready),
    .start_id_0(64'd114688),
    .searchSpace_0_read_addr_s_din(in_14_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_14_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_14_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_14_0___in_14__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_14_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_14_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_14_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_14_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_14_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_14_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_14_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_14_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_14_0___in_14__q0),
    .searchSpace_0_write_data_din(in_14_write_data__din),
    .searchSpace_0_write_data_full_n(in_14_write_data__full_n),
    .searchSpace_0_write_data_write(in_14_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_14_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_14_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_14_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_14_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_14_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_14__din),
    .out_dist_full_n(out_dist_14__full_n),
    .out_dist_write(out_dist_14__write),
    .out_id_din(out_id_14__din),
    .out_id_full_n(out_id_14__full_n),
    .out_id_write(out_id_14__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_15
  krnl_partialKnn_wrapper_15_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_15_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_15_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_15_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_15_0__ap_ready),
    .start_id_0(64'd122880),
    .searchSpace_0_read_addr_s_din(in_15_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_15_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_15_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_15_0___in_15__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_15_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_15_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_15_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_15_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_15_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_15_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_15_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_15_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_15_0___in_15__q0),
    .searchSpace_0_write_data_din(in_15_write_data__din),
    .searchSpace_0_write_data_full_n(in_15_write_data__full_n),
    .searchSpace_0_write_data_write(in_15_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_15_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_15_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_15_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_15_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_15_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_15__din),
    .out_dist_full_n(out_dist_15__full_n),
    .out_dist_write(out_dist_15__write),
    .out_id_din(out_id_15__din),
    .out_id_full_n(out_id_15__full_n),
    .out_id_write(out_id_15__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_16
  krnl_partialKnn_wrapper_16_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_16_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_16_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_16_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_16_0__ap_ready),
    .start_id_0(64'd131072),
    .searchSpace_0_read_addr_s_din(in_16_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_16_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_16_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_16_0___in_16__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_16_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_16_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_16_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_16_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_16_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_16_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_16_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_16_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_16_0___in_16__q0),
    .searchSpace_0_write_data_din(in_16_write_data__din),
    .searchSpace_0_write_data_full_n(in_16_write_data__full_n),
    .searchSpace_0_write_data_write(in_16_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_16_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_16_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_16_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_16_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_16_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_16__din),
    .out_dist_full_n(out_dist_16__full_n),
    .out_dist_write(out_dist_16__write),
    .out_id_din(out_id_16__din),
    .out_id_full_n(out_id_16__full_n),
    .out_id_write(out_id_16__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_17
  krnl_partialKnn_wrapper_17_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_17_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_17_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_17_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_17_0__ap_ready),
    .start_id_0(64'd139264),
    .searchSpace_0_read_addr_s_din(in_17_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_17_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_17_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_17_0___in_17__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_17_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_17_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_17_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_17_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_17_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_17_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_17_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_17_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_17_0___in_17__q0),
    .searchSpace_0_write_data_din(in_17_write_data__din),
    .searchSpace_0_write_data_full_n(in_17_write_data__full_n),
    .searchSpace_0_write_data_write(in_17_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_17_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_17_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_17_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_17_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_17_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_17__din),
    .out_dist_full_n(out_dist_17__full_n),
    .out_dist_write(out_dist_17__write),
    .out_id_din(out_id_17__din),
    .out_id_full_n(out_id_17__full_n),
    .out_id_write(out_id_17__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_18
  krnl_partialKnn_wrapper_18_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_18_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_18_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_18_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_18_0__ap_ready),
    .start_id_0(64'd147456),
    .searchSpace_0_read_addr_s_din(in_18_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_18_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_18_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_18_0___in_18__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_18_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_18_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_18_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_18_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_18_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_18_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_18_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_18_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_18_0___in_18__q0),
    .searchSpace_0_write_data_din(in_18_write_data__din),
    .searchSpace_0_write_data_full_n(in_18_write_data__full_n),
    .searchSpace_0_write_data_write(in_18_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_18_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_18_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_18_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_18_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_18_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_18__din),
    .out_dist_full_n(out_dist_18__full_n),
    .out_dist_write(out_dist_18__write),
    .out_id_din(out_id_18__din),
    .out_id_full_n(out_id_18__full_n),
    .out_id_write(out_id_18__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_19
  krnl_partialKnn_wrapper_19_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_19_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_19_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_19_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_19_0__ap_ready),
    .start_id_0(64'd155648),
    .searchSpace_0_read_addr_s_din(in_19_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_19_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_19_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_19_0___in_19__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_19_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_19_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_19_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_19_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_19_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_19_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_19_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_19_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_19_0___in_19__q0),
    .searchSpace_0_write_data_din(in_19_write_data__din),
    .searchSpace_0_write_data_full_n(in_19_write_data__full_n),
    .searchSpace_0_write_data_write(in_19_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_19_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_19_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_19_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_19_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_19_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_19__din),
    .out_dist_full_n(out_dist_19__full_n),
    .out_dist_write(out_dist_19__write),
    .out_id_din(out_id_19__din),
    .out_id_full_n(out_id_19__full_n),
    .out_id_write(out_id_19__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_2
  krnl_partialKnn_wrapper_2_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_2_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_2_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_2_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_2_0__ap_ready),
    .start_id_0(64'd16384),
    .searchSpace_0_read_addr_s_din(in_2_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_2_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_2_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_2_0___in_2__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_2_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_2_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_2_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_2_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_2_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_2_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_2_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_2_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_2_0___in_2__q0),
    .searchSpace_0_write_data_din(in_2_write_data__din),
    .searchSpace_0_write_data_full_n(in_2_write_data__full_n),
    .searchSpace_0_write_data_write(in_2_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_2_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_2_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_2_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_2_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_2_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_2__din),
    .out_dist_full_n(out_dist_2__full_n),
    .out_dist_write(out_dist_2__write),
    .out_id_din(out_id_2__din),
    .out_id_full_n(out_id_2__full_n),
    .out_id_write(out_id_2__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_20
  krnl_partialKnn_wrapper_20_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_20_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_20_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_20_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_20_0__ap_ready),
    .start_id_0(64'd163840),
    .searchSpace_0_read_addr_s_din(in_20_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_20_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_20_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_20_0___in_20__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_20_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_20_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_20_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_20_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_20_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_20_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_20_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_20_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_20_0___in_20__q0),
    .searchSpace_0_write_data_din(in_20_write_data__din),
    .searchSpace_0_write_data_full_n(in_20_write_data__full_n),
    .searchSpace_0_write_data_write(in_20_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_20_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_20_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_20_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_20_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_20_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_20__din),
    .out_dist_full_n(out_dist_20__full_n),
    .out_dist_write(out_dist_20__write),
    .out_id_din(out_id_20__din),
    .out_id_full_n(out_id_20__full_n),
    .out_id_write(out_id_20__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_21
  krnl_partialKnn_wrapper_21_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_21_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_21_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_21_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_21_0__ap_ready),
    .start_id_0(64'd172032),
    .searchSpace_0_read_addr_s_din(in_21_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_21_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_21_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_21_0___in_21__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_21_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_21_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_21_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_21_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_21_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_21_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_21_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_21_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_21_0___in_21__q0),
    .searchSpace_0_write_data_din(in_21_write_data__din),
    .searchSpace_0_write_data_full_n(in_21_write_data__full_n),
    .searchSpace_0_write_data_write(in_21_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_21_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_21_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_21_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_21_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_21_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_21__din),
    .out_dist_full_n(out_dist_21__full_n),
    .out_dist_write(out_dist_21__write),
    .out_id_din(out_id_21__din),
    .out_id_full_n(out_id_21__full_n),
    .out_id_write(out_id_21__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_22
  krnl_partialKnn_wrapper_22_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_22_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_22_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_22_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_22_0__ap_ready),
    .start_id_0(64'd180224),
    .searchSpace_0_read_addr_s_din(in_22_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_22_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_22_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_22_0___in_22__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_22_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_22_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_22_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_22_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_22_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_22_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_22_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_22_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_22_0___in_22__q0),
    .searchSpace_0_write_data_din(in_22_write_data__din),
    .searchSpace_0_write_data_full_n(in_22_write_data__full_n),
    .searchSpace_0_write_data_write(in_22_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_22_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_22_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_22_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_22_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_22_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_22__din),
    .out_dist_full_n(out_dist_22__full_n),
    .out_dist_write(out_dist_22__write),
    .out_id_din(out_id_22__din),
    .out_id_full_n(out_id_22__full_n),
    .out_id_write(out_id_22__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_23
  krnl_partialKnn_wrapper_23_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_23_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_23_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_23_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_23_0__ap_ready),
    .start_id_0(64'd188416),
    .searchSpace_0_read_addr_s_din(in_23_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_23_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_23_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_23_0___in_23__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_23_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_23_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_23_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_23_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_23_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_23_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_23_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_23_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_23_0___in_23__q0),
    .searchSpace_0_write_data_din(in_23_write_data__din),
    .searchSpace_0_write_data_full_n(in_23_write_data__full_n),
    .searchSpace_0_write_data_write(in_23_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_23_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_23_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_23_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_23_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_23_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_23__din),
    .out_dist_full_n(out_dist_23__full_n),
    .out_dist_write(out_dist_23__write),
    .out_id_din(out_id_23__din),
    .out_id_full_n(out_id_23__full_n),
    .out_id_write(out_id_23__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_24
  krnl_partialKnn_wrapper_24_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_24_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_24_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_24_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_24_0__ap_ready),
    .start_id_0(64'd196608),
    .searchSpace_0_read_addr_s_din(in_24_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_24_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_24_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_24_0___in_24__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_24_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_24_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_24_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_24_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_24_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_24_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_24_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_24_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_24_0___in_24__q0),
    .searchSpace_0_write_data_din(in_24_write_data__din),
    .searchSpace_0_write_data_full_n(in_24_write_data__full_n),
    .searchSpace_0_write_data_write(in_24_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_24_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_24_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_24_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_24_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_24_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_24__din),
    .out_dist_full_n(out_dist_24__full_n),
    .out_dist_write(out_dist_24__write),
    .out_id_din(out_id_24__din),
    .out_id_full_n(out_id_24__full_n),
    .out_id_write(out_id_24__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_25
  krnl_partialKnn_wrapper_25_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_25_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_25_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_25_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_25_0__ap_ready),
    .start_id_0(64'd204800),
    .searchSpace_0_read_addr_s_din(in_25_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_25_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_25_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_25_0___in_25__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_25_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_25_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_25_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_25_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_25_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_25_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_25_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_25_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_25_0___in_25__q0),
    .searchSpace_0_write_data_din(in_25_write_data__din),
    .searchSpace_0_write_data_full_n(in_25_write_data__full_n),
    .searchSpace_0_write_data_write(in_25_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_25_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_25_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_25_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_25_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_25_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_25__din),
    .out_dist_full_n(out_dist_25__full_n),
    .out_dist_write(out_dist_25__write),
    .out_id_din(out_id_25__din),
    .out_id_full_n(out_id_25__full_n),
    .out_id_write(out_id_25__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_26
  krnl_partialKnn_wrapper_26_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_26_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_26_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_26_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_26_0__ap_ready),
    .start_id_0(64'd212992),
    .searchSpace_0_read_addr_s_din(in_26_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_26_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_26_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_26_0___in_26__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_26_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_26_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_26_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_26_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_26_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_26_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_26_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_26_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_26_0___in_26__q0),
    .searchSpace_0_write_data_din(in_26_write_data__din),
    .searchSpace_0_write_data_full_n(in_26_write_data__full_n),
    .searchSpace_0_write_data_write(in_26_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_26_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_26_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_26_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_26_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_26_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_26__din),
    .out_dist_full_n(out_dist_26__full_n),
    .out_dist_write(out_dist_26__write),
    .out_id_din(out_id_26__din),
    .out_id_full_n(out_id_26__full_n),
    .out_id_write(out_id_26__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_3
  krnl_partialKnn_wrapper_3_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_3_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_3_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_3_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_3_0__ap_ready),
    .start_id_0(64'd24576),
    .searchSpace_0_read_addr_s_din(in_3_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_3_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_3_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_3_0___in_3__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_3_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_3_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_3_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_3_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_3_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_3_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_3_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_3_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_3_0___in_3__q0),
    .searchSpace_0_write_data_din(in_3_write_data__din),
    .searchSpace_0_write_data_full_n(in_3_write_data__full_n),
    .searchSpace_0_write_data_write(in_3_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_3_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_3_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_3_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_3_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_3_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_3__din),
    .out_dist_full_n(out_dist_3__full_n),
    .out_dist_write(out_dist_3__write),
    .out_id_din(out_id_3__din),
    .out_id_full_n(out_id_3__full_n),
    .out_id_write(out_id_3__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_4
  krnl_partialKnn_wrapper_4_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_4_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_4_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_4_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_4_0__ap_ready),
    .start_id_0(64'd32768),
    .searchSpace_0_read_addr_s_din(in_4_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_4_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_4_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_4_0___in_4__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_4_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_4_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_4_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_4_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_4_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_4_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_4_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_4_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_4_0___in_4__q0),
    .searchSpace_0_write_data_din(in_4_write_data__din),
    .searchSpace_0_write_data_full_n(in_4_write_data__full_n),
    .searchSpace_0_write_data_write(in_4_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_4_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_4_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_4_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_4_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_4_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_4__din),
    .out_dist_full_n(out_dist_4__full_n),
    .out_dist_write(out_dist_4__write),
    .out_id_din(out_id_4__din),
    .out_id_full_n(out_id_4__full_n),
    .out_id_write(out_id_4__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_5
  krnl_partialKnn_wrapper_5_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_5_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_5_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_5_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_5_0__ap_ready),
    .start_id_0(64'd40960),
    .searchSpace_0_read_addr_s_din(in_5_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_5_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_5_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_5_0___in_5__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_5_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_5_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_5_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_5_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_5_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_5_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_5_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_5_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_5_0___in_5__q0),
    .searchSpace_0_write_data_din(in_5_write_data__din),
    .searchSpace_0_write_data_full_n(in_5_write_data__full_n),
    .searchSpace_0_write_data_write(in_5_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_5_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_5_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_5_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_5_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_5_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_5__din),
    .out_dist_full_n(out_dist_5__full_n),
    .out_dist_write(out_dist_5__write),
    .out_id_din(out_id_5__din),
    .out_id_full_n(out_id_5__full_n),
    .out_id_write(out_id_5__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_6
  krnl_partialKnn_wrapper_6_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_6_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_6_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_6_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_6_0__ap_ready),
    .start_id_0(64'd49152),
    .searchSpace_0_read_addr_s_din(in_6_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_6_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_6_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_6_0___in_6__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_6_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_6_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_6_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_6_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_6_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_6_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_6_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_6_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_6_0___in_6__q0),
    .searchSpace_0_write_data_din(in_6_write_data__din),
    .searchSpace_0_write_data_full_n(in_6_write_data__full_n),
    .searchSpace_0_write_data_write(in_6_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_6_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_6_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_6_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_6_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_6_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_6__din),
    .out_dist_full_n(out_dist_6__full_n),
    .out_dist_write(out_dist_6__write),
    .out_id_din(out_id_6__din),
    .out_id_full_n(out_id_6__full_n),
    .out_id_write(out_id_6__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_7
  krnl_partialKnn_wrapper_7_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_7_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_7_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_7_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_7_0__ap_ready),
    .start_id_0(64'd57344),
    .searchSpace_0_read_addr_s_din(in_7_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_7_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_7_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_7_0___in_7__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_7_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_7_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_7_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_7_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_7_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_7_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_7_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_7_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_7_0___in_7__q0),
    .searchSpace_0_write_data_din(in_7_write_data__din),
    .searchSpace_0_write_data_full_n(in_7_write_data__full_n),
    .searchSpace_0_write_data_write(in_7_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_7_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_7_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_7_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_7_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_7_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_7__din),
    .out_dist_full_n(out_dist_7__full_n),
    .out_dist_write(out_dist_7__write),
    .out_id_din(out_id_7__din),
    .out_id_full_n(out_id_7__full_n),
    .out_id_write(out_id_7__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_8
  krnl_partialKnn_wrapper_8_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_8_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_8_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_8_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_8_0__ap_ready),
    .start_id_0(64'd65536),
    .searchSpace_0_read_addr_s_din(in_8_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_8_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_8_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_8_0___in_8__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_8_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_8_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_8_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_8_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_8_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_8_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_8_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_8_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_8_0___in_8__q0),
    .searchSpace_0_write_data_din(in_8_write_data__din),
    .searchSpace_0_write_data_full_n(in_8_write_data__full_n),
    .searchSpace_0_write_data_write(in_8_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_8_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_8_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_8_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_8_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_8_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_8__din),
    .out_dist_full_n(out_dist_8__full_n),
    .out_dist_write(out_dist_8__write),
    .out_id_din(out_id_8__din),
    .out_id_full_n(out_id_8__full_n),
    .out_id_write(out_id_8__write)
  );


  (* keep_hierarchy = "yes" *) krnl_partialKnn_wrapper_9
  krnl_partialKnn_wrapper_9_0
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(krnl_partialKnn_wrapper_9_0__ap_start),
    .ap_done(krnl_partialKnn_wrapper_9_0__ap_done),
    .ap_idle(krnl_partialKnn_wrapper_9_0__ap_idle),
    .ap_ready(krnl_partialKnn_wrapper_9_0__ap_ready),
    .start_id_0(64'd73728),
    .searchSpace_0_read_addr_s_din(in_9_read_addr__din),
    .searchSpace_0_read_addr_s_full_n(in_9_read_addr__full_n),
    .searchSpace_0_read_addr_s_write(in_9_read_addr__write),
    .searchSpace_0_read_addr_offset(krnl_partialKnn_wrapper_9_0___in_9__q0),
    .searchSpace_0_read_data_s_dout({1'b0, in_9_read_data__dout}),
    .searchSpace_0_read_data_peek_dout({1'b0, in_9_read_data__dout}),
    .searchSpace_0_read_data_s_empty_n(in_9_read_data__empty_n),
    .searchSpace_0_read_data_peek_empty_n(in_9_read_data__empty_n),
    .searchSpace_0_read_data_s_read(in_9_read_data__read),
    .searchSpace_0_read_data_peek_read(),
    .searchSpace_0_write_addr_s_din(in_9_write_addr__din),
    .searchSpace_0_write_addr_s_full_n(in_9_write_addr__full_n),
    .searchSpace_0_write_addr_s_write(in_9_write_addr__write),
    .searchSpace_0_write_addr_offset(krnl_partialKnn_wrapper_9_0___in_9__q0),
    .searchSpace_0_write_data_din(in_9_write_data__din),
    .searchSpace_0_write_data_full_n(in_9_write_data__full_n),
    .searchSpace_0_write_data_write(in_9_write_data__write),
    .searchSpace_0_write_resp_s_dout({1'b0, in_9_write_resp__dout}),
    .searchSpace_0_write_resp_peek_dout({1'b0, in_9_write_resp__dout}),
    .searchSpace_0_write_resp_s_empty_n(in_9_write_resp__empty_n),
    .searchSpace_0_write_resp_peek_empty_n(in_9_write_resp__empty_n),
    .searchSpace_0_write_resp_s_read(in_9_write_resp__read),
    .searchSpace_0_write_resp_peek_read(),
    .out_dist_din(out_dist_9__din),
    .out_dist_full_n(out_dist_9__full_n),
    .out_dist_write(out_dist_9__write),
    .out_id_din(out_id_9__din),
    .out_id_full_n(out_id_9__full_n),
    .out_id_write(out_id_9__write)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(32),
    .DataWidthBytesLog(2),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(255)
  )
  L3_out_dist__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_L3_out_dist_ARADDR),
    .m_axi_ARBURST(m_axi_L3_out_dist_ARBURST),
    .m_axi_ARCACHE(m_axi_L3_out_dist_ARCACHE),
    .m_axi_ARID(m_axi_L3_out_dist_ARID),
    .m_axi_ARLEN(m_axi_L3_out_dist_ARLEN),
    .m_axi_ARLOCK(m_axi_L3_out_dist_ARLOCK),
    .m_axi_ARPROT(m_axi_L3_out_dist_ARPROT),
    .m_axi_ARQOS(m_axi_L3_out_dist_ARQOS),
    .m_axi_ARREADY(m_axi_L3_out_dist_ARREADY),
    .m_axi_ARSIZE(m_axi_L3_out_dist_ARSIZE),
    .m_axi_ARVALID(m_axi_L3_out_dist_ARVALID),
    .m_axi_AWADDR(m_axi_L3_out_dist_AWADDR),
    .m_axi_AWBURST(m_axi_L3_out_dist_AWBURST),
    .m_axi_AWCACHE(m_axi_L3_out_dist_AWCACHE),
    .m_axi_AWID(m_axi_L3_out_dist_AWID),
    .m_axi_AWLEN(m_axi_L3_out_dist_AWLEN),
    .m_axi_AWLOCK(m_axi_L3_out_dist_AWLOCK),
    .m_axi_AWPROT(m_axi_L3_out_dist_AWPROT),
    .m_axi_AWQOS(m_axi_L3_out_dist_AWQOS),
    .m_axi_AWREADY(m_axi_L3_out_dist_AWREADY),
    .m_axi_AWSIZE(m_axi_L3_out_dist_AWSIZE),
    .m_axi_AWVALID(m_axi_L3_out_dist_AWVALID),
    .m_axi_BID(m_axi_L3_out_dist_BID),
    .m_axi_BREADY(m_axi_L3_out_dist_BREADY),
    .m_axi_BRESP(m_axi_L3_out_dist_BRESP),
    .m_axi_BVALID(m_axi_L3_out_dist_BVALID),
    .m_axi_RDATA(m_axi_L3_out_dist_RDATA),
    .m_axi_RID(m_axi_L3_out_dist_RID),
    .m_axi_RLAST(m_axi_L3_out_dist_RLAST),
    .m_axi_RREADY(m_axi_L3_out_dist_RREADY),
    .m_axi_RRESP(m_axi_L3_out_dist_RRESP),
    .m_axi_RVALID(m_axi_L3_out_dist_RVALID),
    .m_axi_WDATA(m_axi_L3_out_dist_WDATA),
    .m_axi_WLAST(m_axi_L3_out_dist_WLAST),
    .m_axi_WREADY(m_axi_L3_out_dist_WREADY),
    .m_axi_WSTRB(m_axi_L3_out_dist_WSTRB),
    .m_axi_WVALID(m_axi_L3_out_dist_WVALID),
    .read_addr_din(L3_out_dist_read_addr__din),
    .read_addr_full_n(L3_out_dist_read_addr__full_n),
    .read_addr_write(L3_out_dist_read_addr__write),
    .read_data_dout(L3_out_dist_read_data__dout),
    .read_data_empty_n(L3_out_dist_read_data__empty_n),
    .read_data_read(L3_out_dist_read_data__read),
    .write_addr_din(L3_out_dist_write_addr__din),
    .write_addr_full_n(L3_out_dist_write_addr__full_n),
    .write_addr_write(L3_out_dist_write_addr__write),
    .write_data_din(L3_out_dist_write_data__din),
    .write_data_full_n(L3_out_dist_write_data__full_n),
    .write_data_write(L3_out_dist_write_data__write),
    .write_resp_dout(L3_out_dist_write_resp__dout),
    .write_resp_empty_n(L3_out_dist_write_resp__empty_n),
    .write_resp_read(L3_out_dist_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(32),
    .DataWidthBytesLog(2),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(255)
  )
  L3_out_id__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_L3_out_id_ARADDR),
    .m_axi_ARBURST(m_axi_L3_out_id_ARBURST),
    .m_axi_ARCACHE(m_axi_L3_out_id_ARCACHE),
    .m_axi_ARID(m_axi_L3_out_id_ARID),
    .m_axi_ARLEN(m_axi_L3_out_id_ARLEN),
    .m_axi_ARLOCK(m_axi_L3_out_id_ARLOCK),
    .m_axi_ARPROT(m_axi_L3_out_id_ARPROT),
    .m_axi_ARQOS(m_axi_L3_out_id_ARQOS),
    .m_axi_ARREADY(m_axi_L3_out_id_ARREADY),
    .m_axi_ARSIZE(m_axi_L3_out_id_ARSIZE),
    .m_axi_ARVALID(m_axi_L3_out_id_ARVALID),
    .m_axi_AWADDR(m_axi_L3_out_id_AWADDR),
    .m_axi_AWBURST(m_axi_L3_out_id_AWBURST),
    .m_axi_AWCACHE(m_axi_L3_out_id_AWCACHE),
    .m_axi_AWID(m_axi_L3_out_id_AWID),
    .m_axi_AWLEN(m_axi_L3_out_id_AWLEN),
    .m_axi_AWLOCK(m_axi_L3_out_id_AWLOCK),
    .m_axi_AWPROT(m_axi_L3_out_id_AWPROT),
    .m_axi_AWQOS(m_axi_L3_out_id_AWQOS),
    .m_axi_AWREADY(m_axi_L3_out_id_AWREADY),
    .m_axi_AWSIZE(m_axi_L3_out_id_AWSIZE),
    .m_axi_AWVALID(m_axi_L3_out_id_AWVALID),
    .m_axi_BID(m_axi_L3_out_id_BID),
    .m_axi_BREADY(m_axi_L3_out_id_BREADY),
    .m_axi_BRESP(m_axi_L3_out_id_BRESP),
    .m_axi_BVALID(m_axi_L3_out_id_BVALID),
    .m_axi_RDATA(m_axi_L3_out_id_RDATA),
    .m_axi_RID(m_axi_L3_out_id_RID),
    .m_axi_RLAST(m_axi_L3_out_id_RLAST),
    .m_axi_RREADY(m_axi_L3_out_id_RREADY),
    .m_axi_RRESP(m_axi_L3_out_id_RRESP),
    .m_axi_RVALID(m_axi_L3_out_id_RVALID),
    .m_axi_WDATA(m_axi_L3_out_id_WDATA),
    .m_axi_WLAST(m_axi_L3_out_id_WLAST),
    .m_axi_WREADY(m_axi_L3_out_id_WREADY),
    .m_axi_WSTRB(m_axi_L3_out_id_WSTRB),
    .m_axi_WVALID(m_axi_L3_out_id_WVALID),
    .read_addr_din(L3_out_id_read_addr__din),
    .read_addr_full_n(L3_out_id_read_addr__full_n),
    .read_addr_write(L3_out_id_read_addr__write),
    .read_data_dout(L3_out_id_read_data__dout),
    .read_data_empty_n(L3_out_id_read_data__empty_n),
    .read_data_read(L3_out_id_read_data__read),
    .write_addr_din(L3_out_id_write_addr__din),
    .write_addr_full_n(L3_out_id_write_addr__full_n),
    .write_addr_write(L3_out_id_write_addr__write),
    .write_data_din(L3_out_id_write_data__din),
    .write_data_full_n(L3_out_id_write_data__full_n),
    .write_data_write(L3_out_id_write_data__write),
    .write_resp_dout(L3_out_id_write_resp__dout),
    .write_resp_empty_n(L3_out_id_write_resp__empty_n),
    .write_resp_read(L3_out_id_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_0__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_0_ARADDR),
    .m_axi_ARBURST(m_axi_in_0_ARBURST),
    .m_axi_ARCACHE(m_axi_in_0_ARCACHE),
    .m_axi_ARID(m_axi_in_0_ARID),
    .m_axi_ARLEN(m_axi_in_0_ARLEN),
    .m_axi_ARLOCK(m_axi_in_0_ARLOCK),
    .m_axi_ARPROT(m_axi_in_0_ARPROT),
    .m_axi_ARQOS(m_axi_in_0_ARQOS),
    .m_axi_ARREADY(m_axi_in_0_ARREADY),
    .m_axi_ARSIZE(m_axi_in_0_ARSIZE),
    .m_axi_ARVALID(m_axi_in_0_ARVALID),
    .m_axi_AWADDR(m_axi_in_0_AWADDR),
    .m_axi_AWBURST(m_axi_in_0_AWBURST),
    .m_axi_AWCACHE(m_axi_in_0_AWCACHE),
    .m_axi_AWID(m_axi_in_0_AWID),
    .m_axi_AWLEN(m_axi_in_0_AWLEN),
    .m_axi_AWLOCK(m_axi_in_0_AWLOCK),
    .m_axi_AWPROT(m_axi_in_0_AWPROT),
    .m_axi_AWQOS(m_axi_in_0_AWQOS),
    .m_axi_AWREADY(m_axi_in_0_AWREADY),
    .m_axi_AWSIZE(m_axi_in_0_AWSIZE),
    .m_axi_AWVALID(m_axi_in_0_AWVALID),
    .m_axi_BID(m_axi_in_0_BID),
    .m_axi_BREADY(m_axi_in_0_BREADY),
    .m_axi_BRESP(m_axi_in_0_BRESP),
    .m_axi_BVALID(m_axi_in_0_BVALID),
    .m_axi_RDATA(m_axi_in_0_RDATA),
    .m_axi_RID(m_axi_in_0_RID),
    .m_axi_RLAST(m_axi_in_0_RLAST),
    .m_axi_RREADY(m_axi_in_0_RREADY),
    .m_axi_RRESP(m_axi_in_0_RRESP),
    .m_axi_RVALID(m_axi_in_0_RVALID),
    .m_axi_WDATA(m_axi_in_0_WDATA),
    .m_axi_WLAST(m_axi_in_0_WLAST),
    .m_axi_WREADY(m_axi_in_0_WREADY),
    .m_axi_WSTRB(m_axi_in_0_WSTRB),
    .m_axi_WVALID(m_axi_in_0_WVALID),
    .read_addr_din(in_0_read_addr__din),
    .read_addr_full_n(in_0_read_addr__full_n),
    .read_addr_write(in_0_read_addr__write),
    .read_data_dout(in_0_read_data__dout),
    .read_data_empty_n(in_0_read_data__empty_n),
    .read_data_read(in_0_read_data__read),
    .write_addr_din(in_0_write_addr__din),
    .write_addr_full_n(in_0_write_addr__full_n),
    .write_addr_write(in_0_write_addr__write),
    .write_data_din(in_0_write_data__din),
    .write_data_full_n(in_0_write_data__full_n),
    .write_data_write(in_0_write_data__write),
    .write_resp_dout(in_0_write_resp__dout),
    .write_resp_empty_n(in_0_write_resp__empty_n),
    .write_resp_read(in_0_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_1__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_1_ARADDR),
    .m_axi_ARBURST(m_axi_in_1_ARBURST),
    .m_axi_ARCACHE(m_axi_in_1_ARCACHE),
    .m_axi_ARID(m_axi_in_1_ARID),
    .m_axi_ARLEN(m_axi_in_1_ARLEN),
    .m_axi_ARLOCK(m_axi_in_1_ARLOCK),
    .m_axi_ARPROT(m_axi_in_1_ARPROT),
    .m_axi_ARQOS(m_axi_in_1_ARQOS),
    .m_axi_ARREADY(m_axi_in_1_ARREADY),
    .m_axi_ARSIZE(m_axi_in_1_ARSIZE),
    .m_axi_ARVALID(m_axi_in_1_ARVALID),
    .m_axi_AWADDR(m_axi_in_1_AWADDR),
    .m_axi_AWBURST(m_axi_in_1_AWBURST),
    .m_axi_AWCACHE(m_axi_in_1_AWCACHE),
    .m_axi_AWID(m_axi_in_1_AWID),
    .m_axi_AWLEN(m_axi_in_1_AWLEN),
    .m_axi_AWLOCK(m_axi_in_1_AWLOCK),
    .m_axi_AWPROT(m_axi_in_1_AWPROT),
    .m_axi_AWQOS(m_axi_in_1_AWQOS),
    .m_axi_AWREADY(m_axi_in_1_AWREADY),
    .m_axi_AWSIZE(m_axi_in_1_AWSIZE),
    .m_axi_AWVALID(m_axi_in_1_AWVALID),
    .m_axi_BID(m_axi_in_1_BID),
    .m_axi_BREADY(m_axi_in_1_BREADY),
    .m_axi_BRESP(m_axi_in_1_BRESP),
    .m_axi_BVALID(m_axi_in_1_BVALID),
    .m_axi_RDATA(m_axi_in_1_RDATA),
    .m_axi_RID(m_axi_in_1_RID),
    .m_axi_RLAST(m_axi_in_1_RLAST),
    .m_axi_RREADY(m_axi_in_1_RREADY),
    .m_axi_RRESP(m_axi_in_1_RRESP),
    .m_axi_RVALID(m_axi_in_1_RVALID),
    .m_axi_WDATA(m_axi_in_1_WDATA),
    .m_axi_WLAST(m_axi_in_1_WLAST),
    .m_axi_WREADY(m_axi_in_1_WREADY),
    .m_axi_WSTRB(m_axi_in_1_WSTRB),
    .m_axi_WVALID(m_axi_in_1_WVALID),
    .read_addr_din(in_1_read_addr__din),
    .read_addr_full_n(in_1_read_addr__full_n),
    .read_addr_write(in_1_read_addr__write),
    .read_data_dout(in_1_read_data__dout),
    .read_data_empty_n(in_1_read_data__empty_n),
    .read_data_read(in_1_read_data__read),
    .write_addr_din(in_1_write_addr__din),
    .write_addr_full_n(in_1_write_addr__full_n),
    .write_addr_write(in_1_write_addr__write),
    .write_data_din(in_1_write_data__din),
    .write_data_full_n(in_1_write_data__full_n),
    .write_data_write(in_1_write_data__write),
    .write_resp_dout(in_1_write_resp__dout),
    .write_resp_empty_n(in_1_write_resp__empty_n),
    .write_resp_read(in_1_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_10__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_10_ARADDR),
    .m_axi_ARBURST(m_axi_in_10_ARBURST),
    .m_axi_ARCACHE(m_axi_in_10_ARCACHE),
    .m_axi_ARID(m_axi_in_10_ARID),
    .m_axi_ARLEN(m_axi_in_10_ARLEN),
    .m_axi_ARLOCK(m_axi_in_10_ARLOCK),
    .m_axi_ARPROT(m_axi_in_10_ARPROT),
    .m_axi_ARQOS(m_axi_in_10_ARQOS),
    .m_axi_ARREADY(m_axi_in_10_ARREADY),
    .m_axi_ARSIZE(m_axi_in_10_ARSIZE),
    .m_axi_ARVALID(m_axi_in_10_ARVALID),
    .m_axi_AWADDR(m_axi_in_10_AWADDR),
    .m_axi_AWBURST(m_axi_in_10_AWBURST),
    .m_axi_AWCACHE(m_axi_in_10_AWCACHE),
    .m_axi_AWID(m_axi_in_10_AWID),
    .m_axi_AWLEN(m_axi_in_10_AWLEN),
    .m_axi_AWLOCK(m_axi_in_10_AWLOCK),
    .m_axi_AWPROT(m_axi_in_10_AWPROT),
    .m_axi_AWQOS(m_axi_in_10_AWQOS),
    .m_axi_AWREADY(m_axi_in_10_AWREADY),
    .m_axi_AWSIZE(m_axi_in_10_AWSIZE),
    .m_axi_AWVALID(m_axi_in_10_AWVALID),
    .m_axi_BID(m_axi_in_10_BID),
    .m_axi_BREADY(m_axi_in_10_BREADY),
    .m_axi_BRESP(m_axi_in_10_BRESP),
    .m_axi_BVALID(m_axi_in_10_BVALID),
    .m_axi_RDATA(m_axi_in_10_RDATA),
    .m_axi_RID(m_axi_in_10_RID),
    .m_axi_RLAST(m_axi_in_10_RLAST),
    .m_axi_RREADY(m_axi_in_10_RREADY),
    .m_axi_RRESP(m_axi_in_10_RRESP),
    .m_axi_RVALID(m_axi_in_10_RVALID),
    .m_axi_WDATA(m_axi_in_10_WDATA),
    .m_axi_WLAST(m_axi_in_10_WLAST),
    .m_axi_WREADY(m_axi_in_10_WREADY),
    .m_axi_WSTRB(m_axi_in_10_WSTRB),
    .m_axi_WVALID(m_axi_in_10_WVALID),
    .read_addr_din(in_10_read_addr__din),
    .read_addr_full_n(in_10_read_addr__full_n),
    .read_addr_write(in_10_read_addr__write),
    .read_data_dout(in_10_read_data__dout),
    .read_data_empty_n(in_10_read_data__empty_n),
    .read_data_read(in_10_read_data__read),
    .write_addr_din(in_10_write_addr__din),
    .write_addr_full_n(in_10_write_addr__full_n),
    .write_addr_write(in_10_write_addr__write),
    .write_data_din(in_10_write_data__din),
    .write_data_full_n(in_10_write_data__full_n),
    .write_data_write(in_10_write_data__write),
    .write_resp_dout(in_10_write_resp__dout),
    .write_resp_empty_n(in_10_write_resp__empty_n),
    .write_resp_read(in_10_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_11__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_11_ARADDR),
    .m_axi_ARBURST(m_axi_in_11_ARBURST),
    .m_axi_ARCACHE(m_axi_in_11_ARCACHE),
    .m_axi_ARID(m_axi_in_11_ARID),
    .m_axi_ARLEN(m_axi_in_11_ARLEN),
    .m_axi_ARLOCK(m_axi_in_11_ARLOCK),
    .m_axi_ARPROT(m_axi_in_11_ARPROT),
    .m_axi_ARQOS(m_axi_in_11_ARQOS),
    .m_axi_ARREADY(m_axi_in_11_ARREADY),
    .m_axi_ARSIZE(m_axi_in_11_ARSIZE),
    .m_axi_ARVALID(m_axi_in_11_ARVALID),
    .m_axi_AWADDR(m_axi_in_11_AWADDR),
    .m_axi_AWBURST(m_axi_in_11_AWBURST),
    .m_axi_AWCACHE(m_axi_in_11_AWCACHE),
    .m_axi_AWID(m_axi_in_11_AWID),
    .m_axi_AWLEN(m_axi_in_11_AWLEN),
    .m_axi_AWLOCK(m_axi_in_11_AWLOCK),
    .m_axi_AWPROT(m_axi_in_11_AWPROT),
    .m_axi_AWQOS(m_axi_in_11_AWQOS),
    .m_axi_AWREADY(m_axi_in_11_AWREADY),
    .m_axi_AWSIZE(m_axi_in_11_AWSIZE),
    .m_axi_AWVALID(m_axi_in_11_AWVALID),
    .m_axi_BID(m_axi_in_11_BID),
    .m_axi_BREADY(m_axi_in_11_BREADY),
    .m_axi_BRESP(m_axi_in_11_BRESP),
    .m_axi_BVALID(m_axi_in_11_BVALID),
    .m_axi_RDATA(m_axi_in_11_RDATA),
    .m_axi_RID(m_axi_in_11_RID),
    .m_axi_RLAST(m_axi_in_11_RLAST),
    .m_axi_RREADY(m_axi_in_11_RREADY),
    .m_axi_RRESP(m_axi_in_11_RRESP),
    .m_axi_RVALID(m_axi_in_11_RVALID),
    .m_axi_WDATA(m_axi_in_11_WDATA),
    .m_axi_WLAST(m_axi_in_11_WLAST),
    .m_axi_WREADY(m_axi_in_11_WREADY),
    .m_axi_WSTRB(m_axi_in_11_WSTRB),
    .m_axi_WVALID(m_axi_in_11_WVALID),
    .read_addr_din(in_11_read_addr__din),
    .read_addr_full_n(in_11_read_addr__full_n),
    .read_addr_write(in_11_read_addr__write),
    .read_data_dout(in_11_read_data__dout),
    .read_data_empty_n(in_11_read_data__empty_n),
    .read_data_read(in_11_read_data__read),
    .write_addr_din(in_11_write_addr__din),
    .write_addr_full_n(in_11_write_addr__full_n),
    .write_addr_write(in_11_write_addr__write),
    .write_data_din(in_11_write_data__din),
    .write_data_full_n(in_11_write_data__full_n),
    .write_data_write(in_11_write_data__write),
    .write_resp_dout(in_11_write_resp__dout),
    .write_resp_empty_n(in_11_write_resp__empty_n),
    .write_resp_read(in_11_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_12__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_12_ARADDR),
    .m_axi_ARBURST(m_axi_in_12_ARBURST),
    .m_axi_ARCACHE(m_axi_in_12_ARCACHE),
    .m_axi_ARID(m_axi_in_12_ARID),
    .m_axi_ARLEN(m_axi_in_12_ARLEN),
    .m_axi_ARLOCK(m_axi_in_12_ARLOCK),
    .m_axi_ARPROT(m_axi_in_12_ARPROT),
    .m_axi_ARQOS(m_axi_in_12_ARQOS),
    .m_axi_ARREADY(m_axi_in_12_ARREADY),
    .m_axi_ARSIZE(m_axi_in_12_ARSIZE),
    .m_axi_ARVALID(m_axi_in_12_ARVALID),
    .m_axi_AWADDR(m_axi_in_12_AWADDR),
    .m_axi_AWBURST(m_axi_in_12_AWBURST),
    .m_axi_AWCACHE(m_axi_in_12_AWCACHE),
    .m_axi_AWID(m_axi_in_12_AWID),
    .m_axi_AWLEN(m_axi_in_12_AWLEN),
    .m_axi_AWLOCK(m_axi_in_12_AWLOCK),
    .m_axi_AWPROT(m_axi_in_12_AWPROT),
    .m_axi_AWQOS(m_axi_in_12_AWQOS),
    .m_axi_AWREADY(m_axi_in_12_AWREADY),
    .m_axi_AWSIZE(m_axi_in_12_AWSIZE),
    .m_axi_AWVALID(m_axi_in_12_AWVALID),
    .m_axi_BID(m_axi_in_12_BID),
    .m_axi_BREADY(m_axi_in_12_BREADY),
    .m_axi_BRESP(m_axi_in_12_BRESP),
    .m_axi_BVALID(m_axi_in_12_BVALID),
    .m_axi_RDATA(m_axi_in_12_RDATA),
    .m_axi_RID(m_axi_in_12_RID),
    .m_axi_RLAST(m_axi_in_12_RLAST),
    .m_axi_RREADY(m_axi_in_12_RREADY),
    .m_axi_RRESP(m_axi_in_12_RRESP),
    .m_axi_RVALID(m_axi_in_12_RVALID),
    .m_axi_WDATA(m_axi_in_12_WDATA),
    .m_axi_WLAST(m_axi_in_12_WLAST),
    .m_axi_WREADY(m_axi_in_12_WREADY),
    .m_axi_WSTRB(m_axi_in_12_WSTRB),
    .m_axi_WVALID(m_axi_in_12_WVALID),
    .read_addr_din(in_12_read_addr__din),
    .read_addr_full_n(in_12_read_addr__full_n),
    .read_addr_write(in_12_read_addr__write),
    .read_data_dout(in_12_read_data__dout),
    .read_data_empty_n(in_12_read_data__empty_n),
    .read_data_read(in_12_read_data__read),
    .write_addr_din(in_12_write_addr__din),
    .write_addr_full_n(in_12_write_addr__full_n),
    .write_addr_write(in_12_write_addr__write),
    .write_data_din(in_12_write_data__din),
    .write_data_full_n(in_12_write_data__full_n),
    .write_data_write(in_12_write_data__write),
    .write_resp_dout(in_12_write_resp__dout),
    .write_resp_empty_n(in_12_write_resp__empty_n),
    .write_resp_read(in_12_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_13__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_13_ARADDR),
    .m_axi_ARBURST(m_axi_in_13_ARBURST),
    .m_axi_ARCACHE(m_axi_in_13_ARCACHE),
    .m_axi_ARID(m_axi_in_13_ARID),
    .m_axi_ARLEN(m_axi_in_13_ARLEN),
    .m_axi_ARLOCK(m_axi_in_13_ARLOCK),
    .m_axi_ARPROT(m_axi_in_13_ARPROT),
    .m_axi_ARQOS(m_axi_in_13_ARQOS),
    .m_axi_ARREADY(m_axi_in_13_ARREADY),
    .m_axi_ARSIZE(m_axi_in_13_ARSIZE),
    .m_axi_ARVALID(m_axi_in_13_ARVALID),
    .m_axi_AWADDR(m_axi_in_13_AWADDR),
    .m_axi_AWBURST(m_axi_in_13_AWBURST),
    .m_axi_AWCACHE(m_axi_in_13_AWCACHE),
    .m_axi_AWID(m_axi_in_13_AWID),
    .m_axi_AWLEN(m_axi_in_13_AWLEN),
    .m_axi_AWLOCK(m_axi_in_13_AWLOCK),
    .m_axi_AWPROT(m_axi_in_13_AWPROT),
    .m_axi_AWQOS(m_axi_in_13_AWQOS),
    .m_axi_AWREADY(m_axi_in_13_AWREADY),
    .m_axi_AWSIZE(m_axi_in_13_AWSIZE),
    .m_axi_AWVALID(m_axi_in_13_AWVALID),
    .m_axi_BID(m_axi_in_13_BID),
    .m_axi_BREADY(m_axi_in_13_BREADY),
    .m_axi_BRESP(m_axi_in_13_BRESP),
    .m_axi_BVALID(m_axi_in_13_BVALID),
    .m_axi_RDATA(m_axi_in_13_RDATA),
    .m_axi_RID(m_axi_in_13_RID),
    .m_axi_RLAST(m_axi_in_13_RLAST),
    .m_axi_RREADY(m_axi_in_13_RREADY),
    .m_axi_RRESP(m_axi_in_13_RRESP),
    .m_axi_RVALID(m_axi_in_13_RVALID),
    .m_axi_WDATA(m_axi_in_13_WDATA),
    .m_axi_WLAST(m_axi_in_13_WLAST),
    .m_axi_WREADY(m_axi_in_13_WREADY),
    .m_axi_WSTRB(m_axi_in_13_WSTRB),
    .m_axi_WVALID(m_axi_in_13_WVALID),
    .read_addr_din(in_13_read_addr__din),
    .read_addr_full_n(in_13_read_addr__full_n),
    .read_addr_write(in_13_read_addr__write),
    .read_data_dout(in_13_read_data__dout),
    .read_data_empty_n(in_13_read_data__empty_n),
    .read_data_read(in_13_read_data__read),
    .write_addr_din(in_13_write_addr__din),
    .write_addr_full_n(in_13_write_addr__full_n),
    .write_addr_write(in_13_write_addr__write),
    .write_data_din(in_13_write_data__din),
    .write_data_full_n(in_13_write_data__full_n),
    .write_data_write(in_13_write_data__write),
    .write_resp_dout(in_13_write_resp__dout),
    .write_resp_empty_n(in_13_write_resp__empty_n),
    .write_resp_read(in_13_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_14__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_14_ARADDR),
    .m_axi_ARBURST(m_axi_in_14_ARBURST),
    .m_axi_ARCACHE(m_axi_in_14_ARCACHE),
    .m_axi_ARID(m_axi_in_14_ARID),
    .m_axi_ARLEN(m_axi_in_14_ARLEN),
    .m_axi_ARLOCK(m_axi_in_14_ARLOCK),
    .m_axi_ARPROT(m_axi_in_14_ARPROT),
    .m_axi_ARQOS(m_axi_in_14_ARQOS),
    .m_axi_ARREADY(m_axi_in_14_ARREADY),
    .m_axi_ARSIZE(m_axi_in_14_ARSIZE),
    .m_axi_ARVALID(m_axi_in_14_ARVALID),
    .m_axi_AWADDR(m_axi_in_14_AWADDR),
    .m_axi_AWBURST(m_axi_in_14_AWBURST),
    .m_axi_AWCACHE(m_axi_in_14_AWCACHE),
    .m_axi_AWID(m_axi_in_14_AWID),
    .m_axi_AWLEN(m_axi_in_14_AWLEN),
    .m_axi_AWLOCK(m_axi_in_14_AWLOCK),
    .m_axi_AWPROT(m_axi_in_14_AWPROT),
    .m_axi_AWQOS(m_axi_in_14_AWQOS),
    .m_axi_AWREADY(m_axi_in_14_AWREADY),
    .m_axi_AWSIZE(m_axi_in_14_AWSIZE),
    .m_axi_AWVALID(m_axi_in_14_AWVALID),
    .m_axi_BID(m_axi_in_14_BID),
    .m_axi_BREADY(m_axi_in_14_BREADY),
    .m_axi_BRESP(m_axi_in_14_BRESP),
    .m_axi_BVALID(m_axi_in_14_BVALID),
    .m_axi_RDATA(m_axi_in_14_RDATA),
    .m_axi_RID(m_axi_in_14_RID),
    .m_axi_RLAST(m_axi_in_14_RLAST),
    .m_axi_RREADY(m_axi_in_14_RREADY),
    .m_axi_RRESP(m_axi_in_14_RRESP),
    .m_axi_RVALID(m_axi_in_14_RVALID),
    .m_axi_WDATA(m_axi_in_14_WDATA),
    .m_axi_WLAST(m_axi_in_14_WLAST),
    .m_axi_WREADY(m_axi_in_14_WREADY),
    .m_axi_WSTRB(m_axi_in_14_WSTRB),
    .m_axi_WVALID(m_axi_in_14_WVALID),
    .read_addr_din(in_14_read_addr__din),
    .read_addr_full_n(in_14_read_addr__full_n),
    .read_addr_write(in_14_read_addr__write),
    .read_data_dout(in_14_read_data__dout),
    .read_data_empty_n(in_14_read_data__empty_n),
    .read_data_read(in_14_read_data__read),
    .write_addr_din(in_14_write_addr__din),
    .write_addr_full_n(in_14_write_addr__full_n),
    .write_addr_write(in_14_write_addr__write),
    .write_data_din(in_14_write_data__din),
    .write_data_full_n(in_14_write_data__full_n),
    .write_data_write(in_14_write_data__write),
    .write_resp_dout(in_14_write_resp__dout),
    .write_resp_empty_n(in_14_write_resp__empty_n),
    .write_resp_read(in_14_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_15__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_15_ARADDR),
    .m_axi_ARBURST(m_axi_in_15_ARBURST),
    .m_axi_ARCACHE(m_axi_in_15_ARCACHE),
    .m_axi_ARID(m_axi_in_15_ARID),
    .m_axi_ARLEN(m_axi_in_15_ARLEN),
    .m_axi_ARLOCK(m_axi_in_15_ARLOCK),
    .m_axi_ARPROT(m_axi_in_15_ARPROT),
    .m_axi_ARQOS(m_axi_in_15_ARQOS),
    .m_axi_ARREADY(m_axi_in_15_ARREADY),
    .m_axi_ARSIZE(m_axi_in_15_ARSIZE),
    .m_axi_ARVALID(m_axi_in_15_ARVALID),
    .m_axi_AWADDR(m_axi_in_15_AWADDR),
    .m_axi_AWBURST(m_axi_in_15_AWBURST),
    .m_axi_AWCACHE(m_axi_in_15_AWCACHE),
    .m_axi_AWID(m_axi_in_15_AWID),
    .m_axi_AWLEN(m_axi_in_15_AWLEN),
    .m_axi_AWLOCK(m_axi_in_15_AWLOCK),
    .m_axi_AWPROT(m_axi_in_15_AWPROT),
    .m_axi_AWQOS(m_axi_in_15_AWQOS),
    .m_axi_AWREADY(m_axi_in_15_AWREADY),
    .m_axi_AWSIZE(m_axi_in_15_AWSIZE),
    .m_axi_AWVALID(m_axi_in_15_AWVALID),
    .m_axi_BID(m_axi_in_15_BID),
    .m_axi_BREADY(m_axi_in_15_BREADY),
    .m_axi_BRESP(m_axi_in_15_BRESP),
    .m_axi_BVALID(m_axi_in_15_BVALID),
    .m_axi_RDATA(m_axi_in_15_RDATA),
    .m_axi_RID(m_axi_in_15_RID),
    .m_axi_RLAST(m_axi_in_15_RLAST),
    .m_axi_RREADY(m_axi_in_15_RREADY),
    .m_axi_RRESP(m_axi_in_15_RRESP),
    .m_axi_RVALID(m_axi_in_15_RVALID),
    .m_axi_WDATA(m_axi_in_15_WDATA),
    .m_axi_WLAST(m_axi_in_15_WLAST),
    .m_axi_WREADY(m_axi_in_15_WREADY),
    .m_axi_WSTRB(m_axi_in_15_WSTRB),
    .m_axi_WVALID(m_axi_in_15_WVALID),
    .read_addr_din(in_15_read_addr__din),
    .read_addr_full_n(in_15_read_addr__full_n),
    .read_addr_write(in_15_read_addr__write),
    .read_data_dout(in_15_read_data__dout),
    .read_data_empty_n(in_15_read_data__empty_n),
    .read_data_read(in_15_read_data__read),
    .write_addr_din(in_15_write_addr__din),
    .write_addr_full_n(in_15_write_addr__full_n),
    .write_addr_write(in_15_write_addr__write),
    .write_data_din(in_15_write_data__din),
    .write_data_full_n(in_15_write_data__full_n),
    .write_data_write(in_15_write_data__write),
    .write_resp_dout(in_15_write_resp__dout),
    .write_resp_empty_n(in_15_write_resp__empty_n),
    .write_resp_read(in_15_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_16__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_16_ARADDR),
    .m_axi_ARBURST(m_axi_in_16_ARBURST),
    .m_axi_ARCACHE(m_axi_in_16_ARCACHE),
    .m_axi_ARID(m_axi_in_16_ARID),
    .m_axi_ARLEN(m_axi_in_16_ARLEN),
    .m_axi_ARLOCK(m_axi_in_16_ARLOCK),
    .m_axi_ARPROT(m_axi_in_16_ARPROT),
    .m_axi_ARQOS(m_axi_in_16_ARQOS),
    .m_axi_ARREADY(m_axi_in_16_ARREADY),
    .m_axi_ARSIZE(m_axi_in_16_ARSIZE),
    .m_axi_ARVALID(m_axi_in_16_ARVALID),
    .m_axi_AWADDR(m_axi_in_16_AWADDR),
    .m_axi_AWBURST(m_axi_in_16_AWBURST),
    .m_axi_AWCACHE(m_axi_in_16_AWCACHE),
    .m_axi_AWID(m_axi_in_16_AWID),
    .m_axi_AWLEN(m_axi_in_16_AWLEN),
    .m_axi_AWLOCK(m_axi_in_16_AWLOCK),
    .m_axi_AWPROT(m_axi_in_16_AWPROT),
    .m_axi_AWQOS(m_axi_in_16_AWQOS),
    .m_axi_AWREADY(m_axi_in_16_AWREADY),
    .m_axi_AWSIZE(m_axi_in_16_AWSIZE),
    .m_axi_AWVALID(m_axi_in_16_AWVALID),
    .m_axi_BID(m_axi_in_16_BID),
    .m_axi_BREADY(m_axi_in_16_BREADY),
    .m_axi_BRESP(m_axi_in_16_BRESP),
    .m_axi_BVALID(m_axi_in_16_BVALID),
    .m_axi_RDATA(m_axi_in_16_RDATA),
    .m_axi_RID(m_axi_in_16_RID),
    .m_axi_RLAST(m_axi_in_16_RLAST),
    .m_axi_RREADY(m_axi_in_16_RREADY),
    .m_axi_RRESP(m_axi_in_16_RRESP),
    .m_axi_RVALID(m_axi_in_16_RVALID),
    .m_axi_WDATA(m_axi_in_16_WDATA),
    .m_axi_WLAST(m_axi_in_16_WLAST),
    .m_axi_WREADY(m_axi_in_16_WREADY),
    .m_axi_WSTRB(m_axi_in_16_WSTRB),
    .m_axi_WVALID(m_axi_in_16_WVALID),
    .read_addr_din(in_16_read_addr__din),
    .read_addr_full_n(in_16_read_addr__full_n),
    .read_addr_write(in_16_read_addr__write),
    .read_data_dout(in_16_read_data__dout),
    .read_data_empty_n(in_16_read_data__empty_n),
    .read_data_read(in_16_read_data__read),
    .write_addr_din(in_16_write_addr__din),
    .write_addr_full_n(in_16_write_addr__full_n),
    .write_addr_write(in_16_write_addr__write),
    .write_data_din(in_16_write_data__din),
    .write_data_full_n(in_16_write_data__full_n),
    .write_data_write(in_16_write_data__write),
    .write_resp_dout(in_16_write_resp__dout),
    .write_resp_empty_n(in_16_write_resp__empty_n),
    .write_resp_read(in_16_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_17__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_17_ARADDR),
    .m_axi_ARBURST(m_axi_in_17_ARBURST),
    .m_axi_ARCACHE(m_axi_in_17_ARCACHE),
    .m_axi_ARID(m_axi_in_17_ARID),
    .m_axi_ARLEN(m_axi_in_17_ARLEN),
    .m_axi_ARLOCK(m_axi_in_17_ARLOCK),
    .m_axi_ARPROT(m_axi_in_17_ARPROT),
    .m_axi_ARQOS(m_axi_in_17_ARQOS),
    .m_axi_ARREADY(m_axi_in_17_ARREADY),
    .m_axi_ARSIZE(m_axi_in_17_ARSIZE),
    .m_axi_ARVALID(m_axi_in_17_ARVALID),
    .m_axi_AWADDR(m_axi_in_17_AWADDR),
    .m_axi_AWBURST(m_axi_in_17_AWBURST),
    .m_axi_AWCACHE(m_axi_in_17_AWCACHE),
    .m_axi_AWID(m_axi_in_17_AWID),
    .m_axi_AWLEN(m_axi_in_17_AWLEN),
    .m_axi_AWLOCK(m_axi_in_17_AWLOCK),
    .m_axi_AWPROT(m_axi_in_17_AWPROT),
    .m_axi_AWQOS(m_axi_in_17_AWQOS),
    .m_axi_AWREADY(m_axi_in_17_AWREADY),
    .m_axi_AWSIZE(m_axi_in_17_AWSIZE),
    .m_axi_AWVALID(m_axi_in_17_AWVALID),
    .m_axi_BID(m_axi_in_17_BID),
    .m_axi_BREADY(m_axi_in_17_BREADY),
    .m_axi_BRESP(m_axi_in_17_BRESP),
    .m_axi_BVALID(m_axi_in_17_BVALID),
    .m_axi_RDATA(m_axi_in_17_RDATA),
    .m_axi_RID(m_axi_in_17_RID),
    .m_axi_RLAST(m_axi_in_17_RLAST),
    .m_axi_RREADY(m_axi_in_17_RREADY),
    .m_axi_RRESP(m_axi_in_17_RRESP),
    .m_axi_RVALID(m_axi_in_17_RVALID),
    .m_axi_WDATA(m_axi_in_17_WDATA),
    .m_axi_WLAST(m_axi_in_17_WLAST),
    .m_axi_WREADY(m_axi_in_17_WREADY),
    .m_axi_WSTRB(m_axi_in_17_WSTRB),
    .m_axi_WVALID(m_axi_in_17_WVALID),
    .read_addr_din(in_17_read_addr__din),
    .read_addr_full_n(in_17_read_addr__full_n),
    .read_addr_write(in_17_read_addr__write),
    .read_data_dout(in_17_read_data__dout),
    .read_data_empty_n(in_17_read_data__empty_n),
    .read_data_read(in_17_read_data__read),
    .write_addr_din(in_17_write_addr__din),
    .write_addr_full_n(in_17_write_addr__full_n),
    .write_addr_write(in_17_write_addr__write),
    .write_data_din(in_17_write_data__din),
    .write_data_full_n(in_17_write_data__full_n),
    .write_data_write(in_17_write_data__write),
    .write_resp_dout(in_17_write_resp__dout),
    .write_resp_empty_n(in_17_write_resp__empty_n),
    .write_resp_read(in_17_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_18__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_18_ARADDR),
    .m_axi_ARBURST(m_axi_in_18_ARBURST),
    .m_axi_ARCACHE(m_axi_in_18_ARCACHE),
    .m_axi_ARID(m_axi_in_18_ARID),
    .m_axi_ARLEN(m_axi_in_18_ARLEN),
    .m_axi_ARLOCK(m_axi_in_18_ARLOCK),
    .m_axi_ARPROT(m_axi_in_18_ARPROT),
    .m_axi_ARQOS(m_axi_in_18_ARQOS),
    .m_axi_ARREADY(m_axi_in_18_ARREADY),
    .m_axi_ARSIZE(m_axi_in_18_ARSIZE),
    .m_axi_ARVALID(m_axi_in_18_ARVALID),
    .m_axi_AWADDR(m_axi_in_18_AWADDR),
    .m_axi_AWBURST(m_axi_in_18_AWBURST),
    .m_axi_AWCACHE(m_axi_in_18_AWCACHE),
    .m_axi_AWID(m_axi_in_18_AWID),
    .m_axi_AWLEN(m_axi_in_18_AWLEN),
    .m_axi_AWLOCK(m_axi_in_18_AWLOCK),
    .m_axi_AWPROT(m_axi_in_18_AWPROT),
    .m_axi_AWQOS(m_axi_in_18_AWQOS),
    .m_axi_AWREADY(m_axi_in_18_AWREADY),
    .m_axi_AWSIZE(m_axi_in_18_AWSIZE),
    .m_axi_AWVALID(m_axi_in_18_AWVALID),
    .m_axi_BID(m_axi_in_18_BID),
    .m_axi_BREADY(m_axi_in_18_BREADY),
    .m_axi_BRESP(m_axi_in_18_BRESP),
    .m_axi_BVALID(m_axi_in_18_BVALID),
    .m_axi_RDATA(m_axi_in_18_RDATA),
    .m_axi_RID(m_axi_in_18_RID),
    .m_axi_RLAST(m_axi_in_18_RLAST),
    .m_axi_RREADY(m_axi_in_18_RREADY),
    .m_axi_RRESP(m_axi_in_18_RRESP),
    .m_axi_RVALID(m_axi_in_18_RVALID),
    .m_axi_WDATA(m_axi_in_18_WDATA),
    .m_axi_WLAST(m_axi_in_18_WLAST),
    .m_axi_WREADY(m_axi_in_18_WREADY),
    .m_axi_WSTRB(m_axi_in_18_WSTRB),
    .m_axi_WVALID(m_axi_in_18_WVALID),
    .read_addr_din(in_18_read_addr__din),
    .read_addr_full_n(in_18_read_addr__full_n),
    .read_addr_write(in_18_read_addr__write),
    .read_data_dout(in_18_read_data__dout),
    .read_data_empty_n(in_18_read_data__empty_n),
    .read_data_read(in_18_read_data__read),
    .write_addr_din(in_18_write_addr__din),
    .write_addr_full_n(in_18_write_addr__full_n),
    .write_addr_write(in_18_write_addr__write),
    .write_data_din(in_18_write_data__din),
    .write_data_full_n(in_18_write_data__full_n),
    .write_data_write(in_18_write_data__write),
    .write_resp_dout(in_18_write_resp__dout),
    .write_resp_empty_n(in_18_write_resp__empty_n),
    .write_resp_read(in_18_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_19__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_19_ARADDR),
    .m_axi_ARBURST(m_axi_in_19_ARBURST),
    .m_axi_ARCACHE(m_axi_in_19_ARCACHE),
    .m_axi_ARID(m_axi_in_19_ARID),
    .m_axi_ARLEN(m_axi_in_19_ARLEN),
    .m_axi_ARLOCK(m_axi_in_19_ARLOCK),
    .m_axi_ARPROT(m_axi_in_19_ARPROT),
    .m_axi_ARQOS(m_axi_in_19_ARQOS),
    .m_axi_ARREADY(m_axi_in_19_ARREADY),
    .m_axi_ARSIZE(m_axi_in_19_ARSIZE),
    .m_axi_ARVALID(m_axi_in_19_ARVALID),
    .m_axi_AWADDR(m_axi_in_19_AWADDR),
    .m_axi_AWBURST(m_axi_in_19_AWBURST),
    .m_axi_AWCACHE(m_axi_in_19_AWCACHE),
    .m_axi_AWID(m_axi_in_19_AWID),
    .m_axi_AWLEN(m_axi_in_19_AWLEN),
    .m_axi_AWLOCK(m_axi_in_19_AWLOCK),
    .m_axi_AWPROT(m_axi_in_19_AWPROT),
    .m_axi_AWQOS(m_axi_in_19_AWQOS),
    .m_axi_AWREADY(m_axi_in_19_AWREADY),
    .m_axi_AWSIZE(m_axi_in_19_AWSIZE),
    .m_axi_AWVALID(m_axi_in_19_AWVALID),
    .m_axi_BID(m_axi_in_19_BID),
    .m_axi_BREADY(m_axi_in_19_BREADY),
    .m_axi_BRESP(m_axi_in_19_BRESP),
    .m_axi_BVALID(m_axi_in_19_BVALID),
    .m_axi_RDATA(m_axi_in_19_RDATA),
    .m_axi_RID(m_axi_in_19_RID),
    .m_axi_RLAST(m_axi_in_19_RLAST),
    .m_axi_RREADY(m_axi_in_19_RREADY),
    .m_axi_RRESP(m_axi_in_19_RRESP),
    .m_axi_RVALID(m_axi_in_19_RVALID),
    .m_axi_WDATA(m_axi_in_19_WDATA),
    .m_axi_WLAST(m_axi_in_19_WLAST),
    .m_axi_WREADY(m_axi_in_19_WREADY),
    .m_axi_WSTRB(m_axi_in_19_WSTRB),
    .m_axi_WVALID(m_axi_in_19_WVALID),
    .read_addr_din(in_19_read_addr__din),
    .read_addr_full_n(in_19_read_addr__full_n),
    .read_addr_write(in_19_read_addr__write),
    .read_data_dout(in_19_read_data__dout),
    .read_data_empty_n(in_19_read_data__empty_n),
    .read_data_read(in_19_read_data__read),
    .write_addr_din(in_19_write_addr__din),
    .write_addr_full_n(in_19_write_addr__full_n),
    .write_addr_write(in_19_write_addr__write),
    .write_data_din(in_19_write_data__din),
    .write_data_full_n(in_19_write_data__full_n),
    .write_data_write(in_19_write_data__write),
    .write_resp_dout(in_19_write_resp__dout),
    .write_resp_empty_n(in_19_write_resp__empty_n),
    .write_resp_read(in_19_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_2__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_2_ARADDR),
    .m_axi_ARBURST(m_axi_in_2_ARBURST),
    .m_axi_ARCACHE(m_axi_in_2_ARCACHE),
    .m_axi_ARID(m_axi_in_2_ARID),
    .m_axi_ARLEN(m_axi_in_2_ARLEN),
    .m_axi_ARLOCK(m_axi_in_2_ARLOCK),
    .m_axi_ARPROT(m_axi_in_2_ARPROT),
    .m_axi_ARQOS(m_axi_in_2_ARQOS),
    .m_axi_ARREADY(m_axi_in_2_ARREADY),
    .m_axi_ARSIZE(m_axi_in_2_ARSIZE),
    .m_axi_ARVALID(m_axi_in_2_ARVALID),
    .m_axi_AWADDR(m_axi_in_2_AWADDR),
    .m_axi_AWBURST(m_axi_in_2_AWBURST),
    .m_axi_AWCACHE(m_axi_in_2_AWCACHE),
    .m_axi_AWID(m_axi_in_2_AWID),
    .m_axi_AWLEN(m_axi_in_2_AWLEN),
    .m_axi_AWLOCK(m_axi_in_2_AWLOCK),
    .m_axi_AWPROT(m_axi_in_2_AWPROT),
    .m_axi_AWQOS(m_axi_in_2_AWQOS),
    .m_axi_AWREADY(m_axi_in_2_AWREADY),
    .m_axi_AWSIZE(m_axi_in_2_AWSIZE),
    .m_axi_AWVALID(m_axi_in_2_AWVALID),
    .m_axi_BID(m_axi_in_2_BID),
    .m_axi_BREADY(m_axi_in_2_BREADY),
    .m_axi_BRESP(m_axi_in_2_BRESP),
    .m_axi_BVALID(m_axi_in_2_BVALID),
    .m_axi_RDATA(m_axi_in_2_RDATA),
    .m_axi_RID(m_axi_in_2_RID),
    .m_axi_RLAST(m_axi_in_2_RLAST),
    .m_axi_RREADY(m_axi_in_2_RREADY),
    .m_axi_RRESP(m_axi_in_2_RRESP),
    .m_axi_RVALID(m_axi_in_2_RVALID),
    .m_axi_WDATA(m_axi_in_2_WDATA),
    .m_axi_WLAST(m_axi_in_2_WLAST),
    .m_axi_WREADY(m_axi_in_2_WREADY),
    .m_axi_WSTRB(m_axi_in_2_WSTRB),
    .m_axi_WVALID(m_axi_in_2_WVALID),
    .read_addr_din(in_2_read_addr__din),
    .read_addr_full_n(in_2_read_addr__full_n),
    .read_addr_write(in_2_read_addr__write),
    .read_data_dout(in_2_read_data__dout),
    .read_data_empty_n(in_2_read_data__empty_n),
    .read_data_read(in_2_read_data__read),
    .write_addr_din(in_2_write_addr__din),
    .write_addr_full_n(in_2_write_addr__full_n),
    .write_addr_write(in_2_write_addr__write),
    .write_data_din(in_2_write_data__din),
    .write_data_full_n(in_2_write_data__full_n),
    .write_data_write(in_2_write_data__write),
    .write_resp_dout(in_2_write_resp__dout),
    .write_resp_empty_n(in_2_write_resp__empty_n),
    .write_resp_read(in_2_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_20__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_20_ARADDR),
    .m_axi_ARBURST(m_axi_in_20_ARBURST),
    .m_axi_ARCACHE(m_axi_in_20_ARCACHE),
    .m_axi_ARID(m_axi_in_20_ARID),
    .m_axi_ARLEN(m_axi_in_20_ARLEN),
    .m_axi_ARLOCK(m_axi_in_20_ARLOCK),
    .m_axi_ARPROT(m_axi_in_20_ARPROT),
    .m_axi_ARQOS(m_axi_in_20_ARQOS),
    .m_axi_ARREADY(m_axi_in_20_ARREADY),
    .m_axi_ARSIZE(m_axi_in_20_ARSIZE),
    .m_axi_ARVALID(m_axi_in_20_ARVALID),
    .m_axi_AWADDR(m_axi_in_20_AWADDR),
    .m_axi_AWBURST(m_axi_in_20_AWBURST),
    .m_axi_AWCACHE(m_axi_in_20_AWCACHE),
    .m_axi_AWID(m_axi_in_20_AWID),
    .m_axi_AWLEN(m_axi_in_20_AWLEN),
    .m_axi_AWLOCK(m_axi_in_20_AWLOCK),
    .m_axi_AWPROT(m_axi_in_20_AWPROT),
    .m_axi_AWQOS(m_axi_in_20_AWQOS),
    .m_axi_AWREADY(m_axi_in_20_AWREADY),
    .m_axi_AWSIZE(m_axi_in_20_AWSIZE),
    .m_axi_AWVALID(m_axi_in_20_AWVALID),
    .m_axi_BID(m_axi_in_20_BID),
    .m_axi_BREADY(m_axi_in_20_BREADY),
    .m_axi_BRESP(m_axi_in_20_BRESP),
    .m_axi_BVALID(m_axi_in_20_BVALID),
    .m_axi_RDATA(m_axi_in_20_RDATA),
    .m_axi_RID(m_axi_in_20_RID),
    .m_axi_RLAST(m_axi_in_20_RLAST),
    .m_axi_RREADY(m_axi_in_20_RREADY),
    .m_axi_RRESP(m_axi_in_20_RRESP),
    .m_axi_RVALID(m_axi_in_20_RVALID),
    .m_axi_WDATA(m_axi_in_20_WDATA),
    .m_axi_WLAST(m_axi_in_20_WLAST),
    .m_axi_WREADY(m_axi_in_20_WREADY),
    .m_axi_WSTRB(m_axi_in_20_WSTRB),
    .m_axi_WVALID(m_axi_in_20_WVALID),
    .read_addr_din(in_20_read_addr__din),
    .read_addr_full_n(in_20_read_addr__full_n),
    .read_addr_write(in_20_read_addr__write),
    .read_data_dout(in_20_read_data__dout),
    .read_data_empty_n(in_20_read_data__empty_n),
    .read_data_read(in_20_read_data__read),
    .write_addr_din(in_20_write_addr__din),
    .write_addr_full_n(in_20_write_addr__full_n),
    .write_addr_write(in_20_write_addr__write),
    .write_data_din(in_20_write_data__din),
    .write_data_full_n(in_20_write_data__full_n),
    .write_data_write(in_20_write_data__write),
    .write_resp_dout(in_20_write_resp__dout),
    .write_resp_empty_n(in_20_write_resp__empty_n),
    .write_resp_read(in_20_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_21__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_21_ARADDR),
    .m_axi_ARBURST(m_axi_in_21_ARBURST),
    .m_axi_ARCACHE(m_axi_in_21_ARCACHE),
    .m_axi_ARID(m_axi_in_21_ARID),
    .m_axi_ARLEN(m_axi_in_21_ARLEN),
    .m_axi_ARLOCK(m_axi_in_21_ARLOCK),
    .m_axi_ARPROT(m_axi_in_21_ARPROT),
    .m_axi_ARQOS(m_axi_in_21_ARQOS),
    .m_axi_ARREADY(m_axi_in_21_ARREADY),
    .m_axi_ARSIZE(m_axi_in_21_ARSIZE),
    .m_axi_ARVALID(m_axi_in_21_ARVALID),
    .m_axi_AWADDR(m_axi_in_21_AWADDR),
    .m_axi_AWBURST(m_axi_in_21_AWBURST),
    .m_axi_AWCACHE(m_axi_in_21_AWCACHE),
    .m_axi_AWID(m_axi_in_21_AWID),
    .m_axi_AWLEN(m_axi_in_21_AWLEN),
    .m_axi_AWLOCK(m_axi_in_21_AWLOCK),
    .m_axi_AWPROT(m_axi_in_21_AWPROT),
    .m_axi_AWQOS(m_axi_in_21_AWQOS),
    .m_axi_AWREADY(m_axi_in_21_AWREADY),
    .m_axi_AWSIZE(m_axi_in_21_AWSIZE),
    .m_axi_AWVALID(m_axi_in_21_AWVALID),
    .m_axi_BID(m_axi_in_21_BID),
    .m_axi_BREADY(m_axi_in_21_BREADY),
    .m_axi_BRESP(m_axi_in_21_BRESP),
    .m_axi_BVALID(m_axi_in_21_BVALID),
    .m_axi_RDATA(m_axi_in_21_RDATA),
    .m_axi_RID(m_axi_in_21_RID),
    .m_axi_RLAST(m_axi_in_21_RLAST),
    .m_axi_RREADY(m_axi_in_21_RREADY),
    .m_axi_RRESP(m_axi_in_21_RRESP),
    .m_axi_RVALID(m_axi_in_21_RVALID),
    .m_axi_WDATA(m_axi_in_21_WDATA),
    .m_axi_WLAST(m_axi_in_21_WLAST),
    .m_axi_WREADY(m_axi_in_21_WREADY),
    .m_axi_WSTRB(m_axi_in_21_WSTRB),
    .m_axi_WVALID(m_axi_in_21_WVALID),
    .read_addr_din(in_21_read_addr__din),
    .read_addr_full_n(in_21_read_addr__full_n),
    .read_addr_write(in_21_read_addr__write),
    .read_data_dout(in_21_read_data__dout),
    .read_data_empty_n(in_21_read_data__empty_n),
    .read_data_read(in_21_read_data__read),
    .write_addr_din(in_21_write_addr__din),
    .write_addr_full_n(in_21_write_addr__full_n),
    .write_addr_write(in_21_write_addr__write),
    .write_data_din(in_21_write_data__din),
    .write_data_full_n(in_21_write_data__full_n),
    .write_data_write(in_21_write_data__write),
    .write_resp_dout(in_21_write_resp__dout),
    .write_resp_empty_n(in_21_write_resp__empty_n),
    .write_resp_read(in_21_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_22__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_22_ARADDR),
    .m_axi_ARBURST(m_axi_in_22_ARBURST),
    .m_axi_ARCACHE(m_axi_in_22_ARCACHE),
    .m_axi_ARID(m_axi_in_22_ARID),
    .m_axi_ARLEN(m_axi_in_22_ARLEN),
    .m_axi_ARLOCK(m_axi_in_22_ARLOCK),
    .m_axi_ARPROT(m_axi_in_22_ARPROT),
    .m_axi_ARQOS(m_axi_in_22_ARQOS),
    .m_axi_ARREADY(m_axi_in_22_ARREADY),
    .m_axi_ARSIZE(m_axi_in_22_ARSIZE),
    .m_axi_ARVALID(m_axi_in_22_ARVALID),
    .m_axi_AWADDR(m_axi_in_22_AWADDR),
    .m_axi_AWBURST(m_axi_in_22_AWBURST),
    .m_axi_AWCACHE(m_axi_in_22_AWCACHE),
    .m_axi_AWID(m_axi_in_22_AWID),
    .m_axi_AWLEN(m_axi_in_22_AWLEN),
    .m_axi_AWLOCK(m_axi_in_22_AWLOCK),
    .m_axi_AWPROT(m_axi_in_22_AWPROT),
    .m_axi_AWQOS(m_axi_in_22_AWQOS),
    .m_axi_AWREADY(m_axi_in_22_AWREADY),
    .m_axi_AWSIZE(m_axi_in_22_AWSIZE),
    .m_axi_AWVALID(m_axi_in_22_AWVALID),
    .m_axi_BID(m_axi_in_22_BID),
    .m_axi_BREADY(m_axi_in_22_BREADY),
    .m_axi_BRESP(m_axi_in_22_BRESP),
    .m_axi_BVALID(m_axi_in_22_BVALID),
    .m_axi_RDATA(m_axi_in_22_RDATA),
    .m_axi_RID(m_axi_in_22_RID),
    .m_axi_RLAST(m_axi_in_22_RLAST),
    .m_axi_RREADY(m_axi_in_22_RREADY),
    .m_axi_RRESP(m_axi_in_22_RRESP),
    .m_axi_RVALID(m_axi_in_22_RVALID),
    .m_axi_WDATA(m_axi_in_22_WDATA),
    .m_axi_WLAST(m_axi_in_22_WLAST),
    .m_axi_WREADY(m_axi_in_22_WREADY),
    .m_axi_WSTRB(m_axi_in_22_WSTRB),
    .m_axi_WVALID(m_axi_in_22_WVALID),
    .read_addr_din(in_22_read_addr__din),
    .read_addr_full_n(in_22_read_addr__full_n),
    .read_addr_write(in_22_read_addr__write),
    .read_data_dout(in_22_read_data__dout),
    .read_data_empty_n(in_22_read_data__empty_n),
    .read_data_read(in_22_read_data__read),
    .write_addr_din(in_22_write_addr__din),
    .write_addr_full_n(in_22_write_addr__full_n),
    .write_addr_write(in_22_write_addr__write),
    .write_data_din(in_22_write_data__din),
    .write_data_full_n(in_22_write_data__full_n),
    .write_data_write(in_22_write_data__write),
    .write_resp_dout(in_22_write_resp__dout),
    .write_resp_empty_n(in_22_write_resp__empty_n),
    .write_resp_read(in_22_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_23__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_23_ARADDR),
    .m_axi_ARBURST(m_axi_in_23_ARBURST),
    .m_axi_ARCACHE(m_axi_in_23_ARCACHE),
    .m_axi_ARID(m_axi_in_23_ARID),
    .m_axi_ARLEN(m_axi_in_23_ARLEN),
    .m_axi_ARLOCK(m_axi_in_23_ARLOCK),
    .m_axi_ARPROT(m_axi_in_23_ARPROT),
    .m_axi_ARQOS(m_axi_in_23_ARQOS),
    .m_axi_ARREADY(m_axi_in_23_ARREADY),
    .m_axi_ARSIZE(m_axi_in_23_ARSIZE),
    .m_axi_ARVALID(m_axi_in_23_ARVALID),
    .m_axi_AWADDR(m_axi_in_23_AWADDR),
    .m_axi_AWBURST(m_axi_in_23_AWBURST),
    .m_axi_AWCACHE(m_axi_in_23_AWCACHE),
    .m_axi_AWID(m_axi_in_23_AWID),
    .m_axi_AWLEN(m_axi_in_23_AWLEN),
    .m_axi_AWLOCK(m_axi_in_23_AWLOCK),
    .m_axi_AWPROT(m_axi_in_23_AWPROT),
    .m_axi_AWQOS(m_axi_in_23_AWQOS),
    .m_axi_AWREADY(m_axi_in_23_AWREADY),
    .m_axi_AWSIZE(m_axi_in_23_AWSIZE),
    .m_axi_AWVALID(m_axi_in_23_AWVALID),
    .m_axi_BID(m_axi_in_23_BID),
    .m_axi_BREADY(m_axi_in_23_BREADY),
    .m_axi_BRESP(m_axi_in_23_BRESP),
    .m_axi_BVALID(m_axi_in_23_BVALID),
    .m_axi_RDATA(m_axi_in_23_RDATA),
    .m_axi_RID(m_axi_in_23_RID),
    .m_axi_RLAST(m_axi_in_23_RLAST),
    .m_axi_RREADY(m_axi_in_23_RREADY),
    .m_axi_RRESP(m_axi_in_23_RRESP),
    .m_axi_RVALID(m_axi_in_23_RVALID),
    .m_axi_WDATA(m_axi_in_23_WDATA),
    .m_axi_WLAST(m_axi_in_23_WLAST),
    .m_axi_WREADY(m_axi_in_23_WREADY),
    .m_axi_WSTRB(m_axi_in_23_WSTRB),
    .m_axi_WVALID(m_axi_in_23_WVALID),
    .read_addr_din(in_23_read_addr__din),
    .read_addr_full_n(in_23_read_addr__full_n),
    .read_addr_write(in_23_read_addr__write),
    .read_data_dout(in_23_read_data__dout),
    .read_data_empty_n(in_23_read_data__empty_n),
    .read_data_read(in_23_read_data__read),
    .write_addr_din(in_23_write_addr__din),
    .write_addr_full_n(in_23_write_addr__full_n),
    .write_addr_write(in_23_write_addr__write),
    .write_data_din(in_23_write_data__din),
    .write_data_full_n(in_23_write_data__full_n),
    .write_data_write(in_23_write_data__write),
    .write_resp_dout(in_23_write_resp__dout),
    .write_resp_empty_n(in_23_write_resp__empty_n),
    .write_resp_read(in_23_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_24__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_24_ARADDR),
    .m_axi_ARBURST(m_axi_in_24_ARBURST),
    .m_axi_ARCACHE(m_axi_in_24_ARCACHE),
    .m_axi_ARID(m_axi_in_24_ARID),
    .m_axi_ARLEN(m_axi_in_24_ARLEN),
    .m_axi_ARLOCK(m_axi_in_24_ARLOCK),
    .m_axi_ARPROT(m_axi_in_24_ARPROT),
    .m_axi_ARQOS(m_axi_in_24_ARQOS),
    .m_axi_ARREADY(m_axi_in_24_ARREADY),
    .m_axi_ARSIZE(m_axi_in_24_ARSIZE),
    .m_axi_ARVALID(m_axi_in_24_ARVALID),
    .m_axi_AWADDR(m_axi_in_24_AWADDR),
    .m_axi_AWBURST(m_axi_in_24_AWBURST),
    .m_axi_AWCACHE(m_axi_in_24_AWCACHE),
    .m_axi_AWID(m_axi_in_24_AWID),
    .m_axi_AWLEN(m_axi_in_24_AWLEN),
    .m_axi_AWLOCK(m_axi_in_24_AWLOCK),
    .m_axi_AWPROT(m_axi_in_24_AWPROT),
    .m_axi_AWQOS(m_axi_in_24_AWQOS),
    .m_axi_AWREADY(m_axi_in_24_AWREADY),
    .m_axi_AWSIZE(m_axi_in_24_AWSIZE),
    .m_axi_AWVALID(m_axi_in_24_AWVALID),
    .m_axi_BID(m_axi_in_24_BID),
    .m_axi_BREADY(m_axi_in_24_BREADY),
    .m_axi_BRESP(m_axi_in_24_BRESP),
    .m_axi_BVALID(m_axi_in_24_BVALID),
    .m_axi_RDATA(m_axi_in_24_RDATA),
    .m_axi_RID(m_axi_in_24_RID),
    .m_axi_RLAST(m_axi_in_24_RLAST),
    .m_axi_RREADY(m_axi_in_24_RREADY),
    .m_axi_RRESP(m_axi_in_24_RRESP),
    .m_axi_RVALID(m_axi_in_24_RVALID),
    .m_axi_WDATA(m_axi_in_24_WDATA),
    .m_axi_WLAST(m_axi_in_24_WLAST),
    .m_axi_WREADY(m_axi_in_24_WREADY),
    .m_axi_WSTRB(m_axi_in_24_WSTRB),
    .m_axi_WVALID(m_axi_in_24_WVALID),
    .read_addr_din(in_24_read_addr__din),
    .read_addr_full_n(in_24_read_addr__full_n),
    .read_addr_write(in_24_read_addr__write),
    .read_data_dout(in_24_read_data__dout),
    .read_data_empty_n(in_24_read_data__empty_n),
    .read_data_read(in_24_read_data__read),
    .write_addr_din(in_24_write_addr__din),
    .write_addr_full_n(in_24_write_addr__full_n),
    .write_addr_write(in_24_write_addr__write),
    .write_data_din(in_24_write_data__din),
    .write_data_full_n(in_24_write_data__full_n),
    .write_data_write(in_24_write_data__write),
    .write_resp_dout(in_24_write_resp__dout),
    .write_resp_empty_n(in_24_write_resp__empty_n),
    .write_resp_read(in_24_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_25__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_25_ARADDR),
    .m_axi_ARBURST(m_axi_in_25_ARBURST),
    .m_axi_ARCACHE(m_axi_in_25_ARCACHE),
    .m_axi_ARID(m_axi_in_25_ARID),
    .m_axi_ARLEN(m_axi_in_25_ARLEN),
    .m_axi_ARLOCK(m_axi_in_25_ARLOCK),
    .m_axi_ARPROT(m_axi_in_25_ARPROT),
    .m_axi_ARQOS(m_axi_in_25_ARQOS),
    .m_axi_ARREADY(m_axi_in_25_ARREADY),
    .m_axi_ARSIZE(m_axi_in_25_ARSIZE),
    .m_axi_ARVALID(m_axi_in_25_ARVALID),
    .m_axi_AWADDR(m_axi_in_25_AWADDR),
    .m_axi_AWBURST(m_axi_in_25_AWBURST),
    .m_axi_AWCACHE(m_axi_in_25_AWCACHE),
    .m_axi_AWID(m_axi_in_25_AWID),
    .m_axi_AWLEN(m_axi_in_25_AWLEN),
    .m_axi_AWLOCK(m_axi_in_25_AWLOCK),
    .m_axi_AWPROT(m_axi_in_25_AWPROT),
    .m_axi_AWQOS(m_axi_in_25_AWQOS),
    .m_axi_AWREADY(m_axi_in_25_AWREADY),
    .m_axi_AWSIZE(m_axi_in_25_AWSIZE),
    .m_axi_AWVALID(m_axi_in_25_AWVALID),
    .m_axi_BID(m_axi_in_25_BID),
    .m_axi_BREADY(m_axi_in_25_BREADY),
    .m_axi_BRESP(m_axi_in_25_BRESP),
    .m_axi_BVALID(m_axi_in_25_BVALID),
    .m_axi_RDATA(m_axi_in_25_RDATA),
    .m_axi_RID(m_axi_in_25_RID),
    .m_axi_RLAST(m_axi_in_25_RLAST),
    .m_axi_RREADY(m_axi_in_25_RREADY),
    .m_axi_RRESP(m_axi_in_25_RRESP),
    .m_axi_RVALID(m_axi_in_25_RVALID),
    .m_axi_WDATA(m_axi_in_25_WDATA),
    .m_axi_WLAST(m_axi_in_25_WLAST),
    .m_axi_WREADY(m_axi_in_25_WREADY),
    .m_axi_WSTRB(m_axi_in_25_WSTRB),
    .m_axi_WVALID(m_axi_in_25_WVALID),
    .read_addr_din(in_25_read_addr__din),
    .read_addr_full_n(in_25_read_addr__full_n),
    .read_addr_write(in_25_read_addr__write),
    .read_data_dout(in_25_read_data__dout),
    .read_data_empty_n(in_25_read_data__empty_n),
    .read_data_read(in_25_read_data__read),
    .write_addr_din(in_25_write_addr__din),
    .write_addr_full_n(in_25_write_addr__full_n),
    .write_addr_write(in_25_write_addr__write),
    .write_data_din(in_25_write_data__din),
    .write_data_full_n(in_25_write_data__full_n),
    .write_data_write(in_25_write_data__write),
    .write_resp_dout(in_25_write_resp__dout),
    .write_resp_empty_n(in_25_write_resp__empty_n),
    .write_resp_read(in_25_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_26__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_26_ARADDR),
    .m_axi_ARBURST(m_axi_in_26_ARBURST),
    .m_axi_ARCACHE(m_axi_in_26_ARCACHE),
    .m_axi_ARID(m_axi_in_26_ARID),
    .m_axi_ARLEN(m_axi_in_26_ARLEN),
    .m_axi_ARLOCK(m_axi_in_26_ARLOCK),
    .m_axi_ARPROT(m_axi_in_26_ARPROT),
    .m_axi_ARQOS(m_axi_in_26_ARQOS),
    .m_axi_ARREADY(m_axi_in_26_ARREADY),
    .m_axi_ARSIZE(m_axi_in_26_ARSIZE),
    .m_axi_ARVALID(m_axi_in_26_ARVALID),
    .m_axi_AWADDR(m_axi_in_26_AWADDR),
    .m_axi_AWBURST(m_axi_in_26_AWBURST),
    .m_axi_AWCACHE(m_axi_in_26_AWCACHE),
    .m_axi_AWID(m_axi_in_26_AWID),
    .m_axi_AWLEN(m_axi_in_26_AWLEN),
    .m_axi_AWLOCK(m_axi_in_26_AWLOCK),
    .m_axi_AWPROT(m_axi_in_26_AWPROT),
    .m_axi_AWQOS(m_axi_in_26_AWQOS),
    .m_axi_AWREADY(m_axi_in_26_AWREADY),
    .m_axi_AWSIZE(m_axi_in_26_AWSIZE),
    .m_axi_AWVALID(m_axi_in_26_AWVALID),
    .m_axi_BID(m_axi_in_26_BID),
    .m_axi_BREADY(m_axi_in_26_BREADY),
    .m_axi_BRESP(m_axi_in_26_BRESP),
    .m_axi_BVALID(m_axi_in_26_BVALID),
    .m_axi_RDATA(m_axi_in_26_RDATA),
    .m_axi_RID(m_axi_in_26_RID),
    .m_axi_RLAST(m_axi_in_26_RLAST),
    .m_axi_RREADY(m_axi_in_26_RREADY),
    .m_axi_RRESP(m_axi_in_26_RRESP),
    .m_axi_RVALID(m_axi_in_26_RVALID),
    .m_axi_WDATA(m_axi_in_26_WDATA),
    .m_axi_WLAST(m_axi_in_26_WLAST),
    .m_axi_WREADY(m_axi_in_26_WREADY),
    .m_axi_WSTRB(m_axi_in_26_WSTRB),
    .m_axi_WVALID(m_axi_in_26_WVALID),
    .read_addr_din(in_26_read_addr__din),
    .read_addr_full_n(in_26_read_addr__full_n),
    .read_addr_write(in_26_read_addr__write),
    .read_data_dout(in_26_read_data__dout),
    .read_data_empty_n(in_26_read_data__empty_n),
    .read_data_read(in_26_read_data__read),
    .write_addr_din(in_26_write_addr__din),
    .write_addr_full_n(in_26_write_addr__full_n),
    .write_addr_write(in_26_write_addr__write),
    .write_data_din(in_26_write_data__din),
    .write_data_full_n(in_26_write_data__full_n),
    .write_data_write(in_26_write_data__write),
    .write_resp_dout(in_26_write_resp__dout),
    .write_resp_empty_n(in_26_write_resp__empty_n),
    .write_resp_read(in_26_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_3__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_3_ARADDR),
    .m_axi_ARBURST(m_axi_in_3_ARBURST),
    .m_axi_ARCACHE(m_axi_in_3_ARCACHE),
    .m_axi_ARID(m_axi_in_3_ARID),
    .m_axi_ARLEN(m_axi_in_3_ARLEN),
    .m_axi_ARLOCK(m_axi_in_3_ARLOCK),
    .m_axi_ARPROT(m_axi_in_3_ARPROT),
    .m_axi_ARQOS(m_axi_in_3_ARQOS),
    .m_axi_ARREADY(m_axi_in_3_ARREADY),
    .m_axi_ARSIZE(m_axi_in_3_ARSIZE),
    .m_axi_ARVALID(m_axi_in_3_ARVALID),
    .m_axi_AWADDR(m_axi_in_3_AWADDR),
    .m_axi_AWBURST(m_axi_in_3_AWBURST),
    .m_axi_AWCACHE(m_axi_in_3_AWCACHE),
    .m_axi_AWID(m_axi_in_3_AWID),
    .m_axi_AWLEN(m_axi_in_3_AWLEN),
    .m_axi_AWLOCK(m_axi_in_3_AWLOCK),
    .m_axi_AWPROT(m_axi_in_3_AWPROT),
    .m_axi_AWQOS(m_axi_in_3_AWQOS),
    .m_axi_AWREADY(m_axi_in_3_AWREADY),
    .m_axi_AWSIZE(m_axi_in_3_AWSIZE),
    .m_axi_AWVALID(m_axi_in_3_AWVALID),
    .m_axi_BID(m_axi_in_3_BID),
    .m_axi_BREADY(m_axi_in_3_BREADY),
    .m_axi_BRESP(m_axi_in_3_BRESP),
    .m_axi_BVALID(m_axi_in_3_BVALID),
    .m_axi_RDATA(m_axi_in_3_RDATA),
    .m_axi_RID(m_axi_in_3_RID),
    .m_axi_RLAST(m_axi_in_3_RLAST),
    .m_axi_RREADY(m_axi_in_3_RREADY),
    .m_axi_RRESP(m_axi_in_3_RRESP),
    .m_axi_RVALID(m_axi_in_3_RVALID),
    .m_axi_WDATA(m_axi_in_3_WDATA),
    .m_axi_WLAST(m_axi_in_3_WLAST),
    .m_axi_WREADY(m_axi_in_3_WREADY),
    .m_axi_WSTRB(m_axi_in_3_WSTRB),
    .m_axi_WVALID(m_axi_in_3_WVALID),
    .read_addr_din(in_3_read_addr__din),
    .read_addr_full_n(in_3_read_addr__full_n),
    .read_addr_write(in_3_read_addr__write),
    .read_data_dout(in_3_read_data__dout),
    .read_data_empty_n(in_3_read_data__empty_n),
    .read_data_read(in_3_read_data__read),
    .write_addr_din(in_3_write_addr__din),
    .write_addr_full_n(in_3_write_addr__full_n),
    .write_addr_write(in_3_write_addr__write),
    .write_data_din(in_3_write_data__din),
    .write_data_full_n(in_3_write_data__full_n),
    .write_data_write(in_3_write_data__write),
    .write_resp_dout(in_3_write_resp__dout),
    .write_resp_empty_n(in_3_write_resp__empty_n),
    .write_resp_read(in_3_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_4__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_4_ARADDR),
    .m_axi_ARBURST(m_axi_in_4_ARBURST),
    .m_axi_ARCACHE(m_axi_in_4_ARCACHE),
    .m_axi_ARID(m_axi_in_4_ARID),
    .m_axi_ARLEN(m_axi_in_4_ARLEN),
    .m_axi_ARLOCK(m_axi_in_4_ARLOCK),
    .m_axi_ARPROT(m_axi_in_4_ARPROT),
    .m_axi_ARQOS(m_axi_in_4_ARQOS),
    .m_axi_ARREADY(m_axi_in_4_ARREADY),
    .m_axi_ARSIZE(m_axi_in_4_ARSIZE),
    .m_axi_ARVALID(m_axi_in_4_ARVALID),
    .m_axi_AWADDR(m_axi_in_4_AWADDR),
    .m_axi_AWBURST(m_axi_in_4_AWBURST),
    .m_axi_AWCACHE(m_axi_in_4_AWCACHE),
    .m_axi_AWID(m_axi_in_4_AWID),
    .m_axi_AWLEN(m_axi_in_4_AWLEN),
    .m_axi_AWLOCK(m_axi_in_4_AWLOCK),
    .m_axi_AWPROT(m_axi_in_4_AWPROT),
    .m_axi_AWQOS(m_axi_in_4_AWQOS),
    .m_axi_AWREADY(m_axi_in_4_AWREADY),
    .m_axi_AWSIZE(m_axi_in_4_AWSIZE),
    .m_axi_AWVALID(m_axi_in_4_AWVALID),
    .m_axi_BID(m_axi_in_4_BID),
    .m_axi_BREADY(m_axi_in_4_BREADY),
    .m_axi_BRESP(m_axi_in_4_BRESP),
    .m_axi_BVALID(m_axi_in_4_BVALID),
    .m_axi_RDATA(m_axi_in_4_RDATA),
    .m_axi_RID(m_axi_in_4_RID),
    .m_axi_RLAST(m_axi_in_4_RLAST),
    .m_axi_RREADY(m_axi_in_4_RREADY),
    .m_axi_RRESP(m_axi_in_4_RRESP),
    .m_axi_RVALID(m_axi_in_4_RVALID),
    .m_axi_WDATA(m_axi_in_4_WDATA),
    .m_axi_WLAST(m_axi_in_4_WLAST),
    .m_axi_WREADY(m_axi_in_4_WREADY),
    .m_axi_WSTRB(m_axi_in_4_WSTRB),
    .m_axi_WVALID(m_axi_in_4_WVALID),
    .read_addr_din(in_4_read_addr__din),
    .read_addr_full_n(in_4_read_addr__full_n),
    .read_addr_write(in_4_read_addr__write),
    .read_data_dout(in_4_read_data__dout),
    .read_data_empty_n(in_4_read_data__empty_n),
    .read_data_read(in_4_read_data__read),
    .write_addr_din(in_4_write_addr__din),
    .write_addr_full_n(in_4_write_addr__full_n),
    .write_addr_write(in_4_write_addr__write),
    .write_data_din(in_4_write_data__din),
    .write_data_full_n(in_4_write_data__full_n),
    .write_data_write(in_4_write_data__write),
    .write_resp_dout(in_4_write_resp__dout),
    .write_resp_empty_n(in_4_write_resp__empty_n),
    .write_resp_read(in_4_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_5__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_5_ARADDR),
    .m_axi_ARBURST(m_axi_in_5_ARBURST),
    .m_axi_ARCACHE(m_axi_in_5_ARCACHE),
    .m_axi_ARID(m_axi_in_5_ARID),
    .m_axi_ARLEN(m_axi_in_5_ARLEN),
    .m_axi_ARLOCK(m_axi_in_5_ARLOCK),
    .m_axi_ARPROT(m_axi_in_5_ARPROT),
    .m_axi_ARQOS(m_axi_in_5_ARQOS),
    .m_axi_ARREADY(m_axi_in_5_ARREADY),
    .m_axi_ARSIZE(m_axi_in_5_ARSIZE),
    .m_axi_ARVALID(m_axi_in_5_ARVALID),
    .m_axi_AWADDR(m_axi_in_5_AWADDR),
    .m_axi_AWBURST(m_axi_in_5_AWBURST),
    .m_axi_AWCACHE(m_axi_in_5_AWCACHE),
    .m_axi_AWID(m_axi_in_5_AWID),
    .m_axi_AWLEN(m_axi_in_5_AWLEN),
    .m_axi_AWLOCK(m_axi_in_5_AWLOCK),
    .m_axi_AWPROT(m_axi_in_5_AWPROT),
    .m_axi_AWQOS(m_axi_in_5_AWQOS),
    .m_axi_AWREADY(m_axi_in_5_AWREADY),
    .m_axi_AWSIZE(m_axi_in_5_AWSIZE),
    .m_axi_AWVALID(m_axi_in_5_AWVALID),
    .m_axi_BID(m_axi_in_5_BID),
    .m_axi_BREADY(m_axi_in_5_BREADY),
    .m_axi_BRESP(m_axi_in_5_BRESP),
    .m_axi_BVALID(m_axi_in_5_BVALID),
    .m_axi_RDATA(m_axi_in_5_RDATA),
    .m_axi_RID(m_axi_in_5_RID),
    .m_axi_RLAST(m_axi_in_5_RLAST),
    .m_axi_RREADY(m_axi_in_5_RREADY),
    .m_axi_RRESP(m_axi_in_5_RRESP),
    .m_axi_RVALID(m_axi_in_5_RVALID),
    .m_axi_WDATA(m_axi_in_5_WDATA),
    .m_axi_WLAST(m_axi_in_5_WLAST),
    .m_axi_WREADY(m_axi_in_5_WREADY),
    .m_axi_WSTRB(m_axi_in_5_WSTRB),
    .m_axi_WVALID(m_axi_in_5_WVALID),
    .read_addr_din(in_5_read_addr__din),
    .read_addr_full_n(in_5_read_addr__full_n),
    .read_addr_write(in_5_read_addr__write),
    .read_data_dout(in_5_read_data__dout),
    .read_data_empty_n(in_5_read_data__empty_n),
    .read_data_read(in_5_read_data__read),
    .write_addr_din(in_5_write_addr__din),
    .write_addr_full_n(in_5_write_addr__full_n),
    .write_addr_write(in_5_write_addr__write),
    .write_data_din(in_5_write_data__din),
    .write_data_full_n(in_5_write_data__full_n),
    .write_data_write(in_5_write_data__write),
    .write_resp_dout(in_5_write_resp__dout),
    .write_resp_empty_n(in_5_write_resp__empty_n),
    .write_resp_read(in_5_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_6__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_6_ARADDR),
    .m_axi_ARBURST(m_axi_in_6_ARBURST),
    .m_axi_ARCACHE(m_axi_in_6_ARCACHE),
    .m_axi_ARID(m_axi_in_6_ARID),
    .m_axi_ARLEN(m_axi_in_6_ARLEN),
    .m_axi_ARLOCK(m_axi_in_6_ARLOCK),
    .m_axi_ARPROT(m_axi_in_6_ARPROT),
    .m_axi_ARQOS(m_axi_in_6_ARQOS),
    .m_axi_ARREADY(m_axi_in_6_ARREADY),
    .m_axi_ARSIZE(m_axi_in_6_ARSIZE),
    .m_axi_ARVALID(m_axi_in_6_ARVALID),
    .m_axi_AWADDR(m_axi_in_6_AWADDR),
    .m_axi_AWBURST(m_axi_in_6_AWBURST),
    .m_axi_AWCACHE(m_axi_in_6_AWCACHE),
    .m_axi_AWID(m_axi_in_6_AWID),
    .m_axi_AWLEN(m_axi_in_6_AWLEN),
    .m_axi_AWLOCK(m_axi_in_6_AWLOCK),
    .m_axi_AWPROT(m_axi_in_6_AWPROT),
    .m_axi_AWQOS(m_axi_in_6_AWQOS),
    .m_axi_AWREADY(m_axi_in_6_AWREADY),
    .m_axi_AWSIZE(m_axi_in_6_AWSIZE),
    .m_axi_AWVALID(m_axi_in_6_AWVALID),
    .m_axi_BID(m_axi_in_6_BID),
    .m_axi_BREADY(m_axi_in_6_BREADY),
    .m_axi_BRESP(m_axi_in_6_BRESP),
    .m_axi_BVALID(m_axi_in_6_BVALID),
    .m_axi_RDATA(m_axi_in_6_RDATA),
    .m_axi_RID(m_axi_in_6_RID),
    .m_axi_RLAST(m_axi_in_6_RLAST),
    .m_axi_RREADY(m_axi_in_6_RREADY),
    .m_axi_RRESP(m_axi_in_6_RRESP),
    .m_axi_RVALID(m_axi_in_6_RVALID),
    .m_axi_WDATA(m_axi_in_6_WDATA),
    .m_axi_WLAST(m_axi_in_6_WLAST),
    .m_axi_WREADY(m_axi_in_6_WREADY),
    .m_axi_WSTRB(m_axi_in_6_WSTRB),
    .m_axi_WVALID(m_axi_in_6_WVALID),
    .read_addr_din(in_6_read_addr__din),
    .read_addr_full_n(in_6_read_addr__full_n),
    .read_addr_write(in_6_read_addr__write),
    .read_data_dout(in_6_read_data__dout),
    .read_data_empty_n(in_6_read_data__empty_n),
    .read_data_read(in_6_read_data__read),
    .write_addr_din(in_6_write_addr__din),
    .write_addr_full_n(in_6_write_addr__full_n),
    .write_addr_write(in_6_write_addr__write),
    .write_data_din(in_6_write_data__din),
    .write_data_full_n(in_6_write_data__full_n),
    .write_data_write(in_6_write_data__write),
    .write_resp_dout(in_6_write_resp__dout),
    .write_resp_empty_n(in_6_write_resp__empty_n),
    .write_resp_read(in_6_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_7__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_7_ARADDR),
    .m_axi_ARBURST(m_axi_in_7_ARBURST),
    .m_axi_ARCACHE(m_axi_in_7_ARCACHE),
    .m_axi_ARID(m_axi_in_7_ARID),
    .m_axi_ARLEN(m_axi_in_7_ARLEN),
    .m_axi_ARLOCK(m_axi_in_7_ARLOCK),
    .m_axi_ARPROT(m_axi_in_7_ARPROT),
    .m_axi_ARQOS(m_axi_in_7_ARQOS),
    .m_axi_ARREADY(m_axi_in_7_ARREADY),
    .m_axi_ARSIZE(m_axi_in_7_ARSIZE),
    .m_axi_ARVALID(m_axi_in_7_ARVALID),
    .m_axi_AWADDR(m_axi_in_7_AWADDR),
    .m_axi_AWBURST(m_axi_in_7_AWBURST),
    .m_axi_AWCACHE(m_axi_in_7_AWCACHE),
    .m_axi_AWID(m_axi_in_7_AWID),
    .m_axi_AWLEN(m_axi_in_7_AWLEN),
    .m_axi_AWLOCK(m_axi_in_7_AWLOCK),
    .m_axi_AWPROT(m_axi_in_7_AWPROT),
    .m_axi_AWQOS(m_axi_in_7_AWQOS),
    .m_axi_AWREADY(m_axi_in_7_AWREADY),
    .m_axi_AWSIZE(m_axi_in_7_AWSIZE),
    .m_axi_AWVALID(m_axi_in_7_AWVALID),
    .m_axi_BID(m_axi_in_7_BID),
    .m_axi_BREADY(m_axi_in_7_BREADY),
    .m_axi_BRESP(m_axi_in_7_BRESP),
    .m_axi_BVALID(m_axi_in_7_BVALID),
    .m_axi_RDATA(m_axi_in_7_RDATA),
    .m_axi_RID(m_axi_in_7_RID),
    .m_axi_RLAST(m_axi_in_7_RLAST),
    .m_axi_RREADY(m_axi_in_7_RREADY),
    .m_axi_RRESP(m_axi_in_7_RRESP),
    .m_axi_RVALID(m_axi_in_7_RVALID),
    .m_axi_WDATA(m_axi_in_7_WDATA),
    .m_axi_WLAST(m_axi_in_7_WLAST),
    .m_axi_WREADY(m_axi_in_7_WREADY),
    .m_axi_WSTRB(m_axi_in_7_WSTRB),
    .m_axi_WVALID(m_axi_in_7_WVALID),
    .read_addr_din(in_7_read_addr__din),
    .read_addr_full_n(in_7_read_addr__full_n),
    .read_addr_write(in_7_read_addr__write),
    .read_data_dout(in_7_read_data__dout),
    .read_data_empty_n(in_7_read_data__empty_n),
    .read_data_read(in_7_read_data__read),
    .write_addr_din(in_7_write_addr__din),
    .write_addr_full_n(in_7_write_addr__full_n),
    .write_addr_write(in_7_write_addr__write),
    .write_data_din(in_7_write_data__din),
    .write_data_full_n(in_7_write_data__full_n),
    .write_data_write(in_7_write_data__write),
    .write_resp_dout(in_7_write_resp__dout),
    .write_resp_empty_n(in_7_write_resp__empty_n),
    .write_resp_read(in_7_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_8__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_8_ARADDR),
    .m_axi_ARBURST(m_axi_in_8_ARBURST),
    .m_axi_ARCACHE(m_axi_in_8_ARCACHE),
    .m_axi_ARID(m_axi_in_8_ARID),
    .m_axi_ARLEN(m_axi_in_8_ARLEN),
    .m_axi_ARLOCK(m_axi_in_8_ARLOCK),
    .m_axi_ARPROT(m_axi_in_8_ARPROT),
    .m_axi_ARQOS(m_axi_in_8_ARQOS),
    .m_axi_ARREADY(m_axi_in_8_ARREADY),
    .m_axi_ARSIZE(m_axi_in_8_ARSIZE),
    .m_axi_ARVALID(m_axi_in_8_ARVALID),
    .m_axi_AWADDR(m_axi_in_8_AWADDR),
    .m_axi_AWBURST(m_axi_in_8_AWBURST),
    .m_axi_AWCACHE(m_axi_in_8_AWCACHE),
    .m_axi_AWID(m_axi_in_8_AWID),
    .m_axi_AWLEN(m_axi_in_8_AWLEN),
    .m_axi_AWLOCK(m_axi_in_8_AWLOCK),
    .m_axi_AWPROT(m_axi_in_8_AWPROT),
    .m_axi_AWQOS(m_axi_in_8_AWQOS),
    .m_axi_AWREADY(m_axi_in_8_AWREADY),
    .m_axi_AWSIZE(m_axi_in_8_AWSIZE),
    .m_axi_AWVALID(m_axi_in_8_AWVALID),
    .m_axi_BID(m_axi_in_8_BID),
    .m_axi_BREADY(m_axi_in_8_BREADY),
    .m_axi_BRESP(m_axi_in_8_BRESP),
    .m_axi_BVALID(m_axi_in_8_BVALID),
    .m_axi_RDATA(m_axi_in_8_RDATA),
    .m_axi_RID(m_axi_in_8_RID),
    .m_axi_RLAST(m_axi_in_8_RLAST),
    .m_axi_RREADY(m_axi_in_8_RREADY),
    .m_axi_RRESP(m_axi_in_8_RRESP),
    .m_axi_RVALID(m_axi_in_8_RVALID),
    .m_axi_WDATA(m_axi_in_8_WDATA),
    .m_axi_WLAST(m_axi_in_8_WLAST),
    .m_axi_WREADY(m_axi_in_8_WREADY),
    .m_axi_WSTRB(m_axi_in_8_WSTRB),
    .m_axi_WVALID(m_axi_in_8_WVALID),
    .read_addr_din(in_8_read_addr__din),
    .read_addr_full_n(in_8_read_addr__full_n),
    .read_addr_write(in_8_read_addr__write),
    .read_data_dout(in_8_read_data__dout),
    .read_data_empty_n(in_8_read_data__empty_n),
    .read_data_read(in_8_read_data__read),
    .write_addr_din(in_8_write_addr__din),
    .write_addr_full_n(in_8_write_addr__full_n),
    .write_addr_write(in_8_write_addr__write),
    .write_data_din(in_8_write_data__din),
    .write_data_full_n(in_8_write_data__full_n),
    .write_data_write(in_8_write_data__write),
    .write_resp_dout(in_8_write_resp__dout),
    .write_resp_empty_n(in_8_write_resp__empty_n),
    .write_resp_read(in_8_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) async_mmap
  #(
    .DataWidth(256),
    .DataWidthBytesLog(5),
    .AddrWidth(64),
    .WaitTimeWidth(2),
    .MaxWaitTime(3),
    .BurstLenWidth(9),
    .MaxBurstLen(31)
  )
  in_9__m_axi
  (
    .clk(ap_clk),
    .rst(~ap_rst_n),
    .m_axi_ARADDR(m_axi_in_9_ARADDR),
    .m_axi_ARBURST(m_axi_in_9_ARBURST),
    .m_axi_ARCACHE(m_axi_in_9_ARCACHE),
    .m_axi_ARID(m_axi_in_9_ARID),
    .m_axi_ARLEN(m_axi_in_9_ARLEN),
    .m_axi_ARLOCK(m_axi_in_9_ARLOCK),
    .m_axi_ARPROT(m_axi_in_9_ARPROT),
    .m_axi_ARQOS(m_axi_in_9_ARQOS),
    .m_axi_ARREADY(m_axi_in_9_ARREADY),
    .m_axi_ARSIZE(m_axi_in_9_ARSIZE),
    .m_axi_ARVALID(m_axi_in_9_ARVALID),
    .m_axi_AWADDR(m_axi_in_9_AWADDR),
    .m_axi_AWBURST(m_axi_in_9_AWBURST),
    .m_axi_AWCACHE(m_axi_in_9_AWCACHE),
    .m_axi_AWID(m_axi_in_9_AWID),
    .m_axi_AWLEN(m_axi_in_9_AWLEN),
    .m_axi_AWLOCK(m_axi_in_9_AWLOCK),
    .m_axi_AWPROT(m_axi_in_9_AWPROT),
    .m_axi_AWQOS(m_axi_in_9_AWQOS),
    .m_axi_AWREADY(m_axi_in_9_AWREADY),
    .m_axi_AWSIZE(m_axi_in_9_AWSIZE),
    .m_axi_AWVALID(m_axi_in_9_AWVALID),
    .m_axi_BID(m_axi_in_9_BID),
    .m_axi_BREADY(m_axi_in_9_BREADY),
    .m_axi_BRESP(m_axi_in_9_BRESP),
    .m_axi_BVALID(m_axi_in_9_BVALID),
    .m_axi_RDATA(m_axi_in_9_RDATA),
    .m_axi_RID(m_axi_in_9_RID),
    .m_axi_RLAST(m_axi_in_9_RLAST),
    .m_axi_RREADY(m_axi_in_9_RREADY),
    .m_axi_RRESP(m_axi_in_9_RRESP),
    .m_axi_RVALID(m_axi_in_9_RVALID),
    .m_axi_WDATA(m_axi_in_9_WDATA),
    .m_axi_WLAST(m_axi_in_9_WLAST),
    .m_axi_WREADY(m_axi_in_9_WREADY),
    .m_axi_WSTRB(m_axi_in_9_WSTRB),
    .m_axi_WVALID(m_axi_in_9_WVALID),
    .read_addr_din(in_9_read_addr__din),
    .read_addr_full_n(in_9_read_addr__full_n),
    .read_addr_write(in_9_read_addr__write),
    .read_data_dout(in_9_read_data__dout),
    .read_data_empty_n(in_9_read_data__empty_n),
    .read_data_read(in_9_read_data__read),
    .write_addr_din(in_9_write_addr__din),
    .write_addr_full_n(in_9_write_addr__full_n),
    .write_addr_write(in_9_write_addr__write),
    .write_data_din(in_9_write_data__din),
    .write_data_full_n(in_9_write_data__full_n),
    .write_data_write(in_9_write_data__write),
    .write_resp_dout(in_9_write_resp__dout),
    .write_resp_empty_n(in_9_write_resp__empty_n),
    .write_resp_read(in_9_write_resp__read)
  );


  (* keep_hierarchy = "yes" *) Knn_fsm
  __tapa_fsm_unit
  (
    .ap_clk(ap_clk),
    .ap_rst_n(ap_rst_n),
    .ap_start(ap_start),
    .ap_done(ap_done),
    .ap_idle(ap_idle),
    .ap_ready(ap_ready),
    .L3_out_dist(L3_out_dist),
    .L3_out_id(L3_out_id),
    .in_0(in_0),
    .in_1(in_1),
    .in_10(in_10),
    .in_11(in_11),
    .in_12(in_12),
    .in_13(in_13),
    .in_14(in_14),
    .in_15(in_15),
    .in_16(in_16),
    .in_17(in_17),
    .in_18(in_18),
    .in_19(in_19),
    .in_2(in_2),
    .in_20(in_20),
    .in_21(in_21),
    .in_22(in_22),
    .in_23(in_23),
    .in_24(in_24),
    .in_25(in_25),
    .in_26(in_26),
    .in_3(in_3),
    .in_4(in_4),
    .in_5(in_5),
    .in_6(in_6),
    .in_7(in_7),
    .in_8(in_8),
    .in_9(in_9),
    .krnl_globalSort_L1_L2_0__ap_start(krnl_globalSort_L1_L2_0__ap_start),
    .krnl_globalSort_L1_L2_0__ap_ready(krnl_globalSort_L1_L2_0__ap_ready),
    .krnl_globalSort_L1_L2_0__ap_done(krnl_globalSort_L1_L2_0__ap_done),
    .krnl_globalSort_L1_L2_0__ap_idle(krnl_globalSort_L1_L2_0__ap_idle),
    .krnl_globalSort_L1_L2_1__ap_start(krnl_globalSort_L1_L2_1__ap_start),
    .krnl_globalSort_L1_L2_1__ap_ready(krnl_globalSort_L1_L2_1__ap_ready),
    .krnl_globalSort_L1_L2_1__ap_done(krnl_globalSort_L1_L2_1__ap_done),
    .krnl_globalSort_L1_L2_1__ap_idle(krnl_globalSort_L1_L2_1__ap_idle),
    .krnl_globalSort_L1_L2_2__ap_start(krnl_globalSort_L1_L2_2__ap_start),
    .krnl_globalSort_L1_L2_2__ap_ready(krnl_globalSort_L1_L2_2__ap_ready),
    .krnl_globalSort_L1_L2_2__ap_done(krnl_globalSort_L1_L2_2__ap_done),
    .krnl_globalSort_L1_L2_2__ap_idle(krnl_globalSort_L1_L2_2__ap_idle),
    .krnl_globalSort_L1_L2_3__ap_start(krnl_globalSort_L1_L2_3__ap_start),
    .krnl_globalSort_L1_L2_3__ap_ready(krnl_globalSort_L1_L2_3__ap_ready),
    .krnl_globalSort_L1_L2_3__ap_done(krnl_globalSort_L1_L2_3__ap_done),
    .krnl_globalSort_L1_L2_3__ap_idle(krnl_globalSort_L1_L2_3__ap_idle),
    .krnl_globalSort_L1_L2_4__ap_start(krnl_globalSort_L1_L2_4__ap_start),
    .krnl_globalSort_L1_L2_4__ap_ready(krnl_globalSort_L1_L2_4__ap_ready),
    .krnl_globalSort_L1_L2_4__ap_done(krnl_globalSort_L1_L2_4__ap_done),
    .krnl_globalSort_L1_L2_4__ap_idle(krnl_globalSort_L1_L2_4__ap_idle),
    .krnl_globalSort_L1_L2_5__ap_start(krnl_globalSort_L1_L2_5__ap_start),
    .krnl_globalSort_L1_L2_5__ap_ready(krnl_globalSort_L1_L2_5__ap_ready),
    .krnl_globalSort_L1_L2_5__ap_done(krnl_globalSort_L1_L2_5__ap_done),
    .krnl_globalSort_L1_L2_5__ap_idle(krnl_globalSort_L1_L2_5__ap_idle),
    .krnl_globalSort_L1_L2_6__ap_start(krnl_globalSort_L1_L2_6__ap_start),
    .krnl_globalSort_L1_L2_6__ap_ready(krnl_globalSort_L1_L2_6__ap_ready),
    .krnl_globalSort_L1_L2_6__ap_done(krnl_globalSort_L1_L2_6__ap_done),
    .krnl_globalSort_L1_L2_6__ap_idle(krnl_globalSort_L1_L2_6__ap_idle),
    .krnl_globalSort_L1_L2_7__ap_start(krnl_globalSort_L1_L2_7__ap_start),
    .krnl_globalSort_L1_L2_7__ap_ready(krnl_globalSort_L1_L2_7__ap_ready),
    .krnl_globalSort_L1_L2_7__ap_done(krnl_globalSort_L1_L2_7__ap_done),
    .krnl_globalSort_L1_L2_7__ap_idle(krnl_globalSort_L1_L2_7__ap_idle),
    .krnl_globalSort_L1_L2_8__ap_start(krnl_globalSort_L1_L2_8__ap_start),
    .krnl_globalSort_L1_L2_8__ap_ready(krnl_globalSort_L1_L2_8__ap_ready),
    .krnl_globalSort_L1_L2_8__ap_done(krnl_globalSort_L1_L2_8__ap_done),
    .krnl_globalSort_L1_L2_8__ap_idle(krnl_globalSort_L1_L2_8__ap_idle),
    .krnl_globalSort_L1_L2_9__ap_start(krnl_globalSort_L1_L2_9__ap_start),
    .krnl_globalSort_L1_L2_9__ap_ready(krnl_globalSort_L1_L2_9__ap_ready),
    .krnl_globalSort_L1_L2_9__ap_done(krnl_globalSort_L1_L2_9__ap_done),
    .krnl_globalSort_L1_L2_9__ap_idle(krnl_globalSort_L1_L2_9__ap_idle),
    .krnl_globalSort_L1_L2_10__ap_start(krnl_globalSort_L1_L2_10__ap_start),
    .krnl_globalSort_L1_L2_10__ap_ready(krnl_globalSort_L1_L2_10__ap_ready),
    .krnl_globalSort_L1_L2_10__ap_done(krnl_globalSort_L1_L2_10__ap_done),
    .krnl_globalSort_L1_L2_10__ap_idle(krnl_globalSort_L1_L2_10__ap_idle),
    .krnl_globalSort_L1_L2_11__ap_start(krnl_globalSort_L1_L2_11__ap_start),
    .krnl_globalSort_L1_L2_11__ap_ready(krnl_globalSort_L1_L2_11__ap_ready),
    .krnl_globalSort_L1_L2_11__ap_done(krnl_globalSort_L1_L2_11__ap_done),
    .krnl_globalSort_L1_L2_11__ap_idle(krnl_globalSort_L1_L2_11__ap_idle),
    .krnl_globalSort_L1_L2_12__ap_start(krnl_globalSort_L1_L2_12__ap_start),
    .krnl_globalSort_L1_L2_12__ap_ready(krnl_globalSort_L1_L2_12__ap_ready),
    .krnl_globalSort_L1_L2_12__ap_done(krnl_globalSort_L1_L2_12__ap_done),
    .krnl_globalSort_L1_L2_12__ap_idle(krnl_globalSort_L1_L2_12__ap_idle),
    .krnl_output_dist_id_0___L3_out_dist__q0(krnl_output_dist_id_0___L3_out_dist__q0),
    .krnl_output_dist_id_0___L3_out_id__q0(krnl_output_dist_id_0___L3_out_id__q0),
    .krnl_output_dist_id_0__ap_start(krnl_output_dist_id_0__ap_start),
    .krnl_output_dist_id_0__ap_ready(krnl_output_dist_id_0__ap_ready),
    .krnl_output_dist_id_0__ap_done(krnl_output_dist_id_0__ap_done),
    .krnl_output_dist_id_0__ap_idle(krnl_output_dist_id_0__ap_idle),
    .krnl_partialKnn_wrapper_0_0___in_0__q0(krnl_partialKnn_wrapper_0_0___in_0__q0),
    .krnl_partialKnn_wrapper_0_0__ap_start(krnl_partialKnn_wrapper_0_0__ap_start),
    .krnl_partialKnn_wrapper_0_0__ap_ready(krnl_partialKnn_wrapper_0_0__ap_ready),
    .krnl_partialKnn_wrapper_0_0__ap_done(krnl_partialKnn_wrapper_0_0__ap_done),
    .krnl_partialKnn_wrapper_0_0__ap_idle(krnl_partialKnn_wrapper_0_0__ap_idle),
    .krnl_partialKnn_wrapper_1_0___in_1__q0(krnl_partialKnn_wrapper_1_0___in_1__q0),
    .krnl_partialKnn_wrapper_1_0__ap_start(krnl_partialKnn_wrapper_1_0__ap_start),
    .krnl_partialKnn_wrapper_1_0__ap_ready(krnl_partialKnn_wrapper_1_0__ap_ready),
    .krnl_partialKnn_wrapper_1_0__ap_done(krnl_partialKnn_wrapper_1_0__ap_done),
    .krnl_partialKnn_wrapper_1_0__ap_idle(krnl_partialKnn_wrapper_1_0__ap_idle),
    .krnl_partialKnn_wrapper_10_0___in_10__q0(krnl_partialKnn_wrapper_10_0___in_10__q0),
    .krnl_partialKnn_wrapper_10_0__ap_start(krnl_partialKnn_wrapper_10_0__ap_start),
    .krnl_partialKnn_wrapper_10_0__ap_ready(krnl_partialKnn_wrapper_10_0__ap_ready),
    .krnl_partialKnn_wrapper_10_0__ap_done(krnl_partialKnn_wrapper_10_0__ap_done),
    .krnl_partialKnn_wrapper_10_0__ap_idle(krnl_partialKnn_wrapper_10_0__ap_idle),
    .krnl_partialKnn_wrapper_11_0___in_11__q0(krnl_partialKnn_wrapper_11_0___in_11__q0),
    .krnl_partialKnn_wrapper_11_0__ap_start(krnl_partialKnn_wrapper_11_0__ap_start),
    .krnl_partialKnn_wrapper_11_0__ap_ready(krnl_partialKnn_wrapper_11_0__ap_ready),
    .krnl_partialKnn_wrapper_11_0__ap_done(krnl_partialKnn_wrapper_11_0__ap_done),
    .krnl_partialKnn_wrapper_11_0__ap_idle(krnl_partialKnn_wrapper_11_0__ap_idle),
    .krnl_partialKnn_wrapper_12_0___in_12__q0(krnl_partialKnn_wrapper_12_0___in_12__q0),
    .krnl_partialKnn_wrapper_12_0__ap_start(krnl_partialKnn_wrapper_12_0__ap_start),
    .krnl_partialKnn_wrapper_12_0__ap_ready(krnl_partialKnn_wrapper_12_0__ap_ready),
    .krnl_partialKnn_wrapper_12_0__ap_done(krnl_partialKnn_wrapper_12_0__ap_done),
    .krnl_partialKnn_wrapper_12_0__ap_idle(krnl_partialKnn_wrapper_12_0__ap_idle),
    .krnl_partialKnn_wrapper_13_0___in_13__q0(krnl_partialKnn_wrapper_13_0___in_13__q0),
    .krnl_partialKnn_wrapper_13_0__ap_start(krnl_partialKnn_wrapper_13_0__ap_start),
    .krnl_partialKnn_wrapper_13_0__ap_ready(krnl_partialKnn_wrapper_13_0__ap_ready),
    .krnl_partialKnn_wrapper_13_0__ap_done(krnl_partialKnn_wrapper_13_0__ap_done),
    .krnl_partialKnn_wrapper_13_0__ap_idle(krnl_partialKnn_wrapper_13_0__ap_idle),
    .krnl_partialKnn_wrapper_14_0___in_14__q0(krnl_partialKnn_wrapper_14_0___in_14__q0),
    .krnl_partialKnn_wrapper_14_0__ap_start(krnl_partialKnn_wrapper_14_0__ap_start),
    .krnl_partialKnn_wrapper_14_0__ap_ready(krnl_partialKnn_wrapper_14_0__ap_ready),
    .krnl_partialKnn_wrapper_14_0__ap_done(krnl_partialKnn_wrapper_14_0__ap_done),
    .krnl_partialKnn_wrapper_14_0__ap_idle(krnl_partialKnn_wrapper_14_0__ap_idle),
    .krnl_partialKnn_wrapper_15_0___in_15__q0(krnl_partialKnn_wrapper_15_0___in_15__q0),
    .krnl_partialKnn_wrapper_15_0__ap_start(krnl_partialKnn_wrapper_15_0__ap_start),
    .krnl_partialKnn_wrapper_15_0__ap_ready(krnl_partialKnn_wrapper_15_0__ap_ready),
    .krnl_partialKnn_wrapper_15_0__ap_done(krnl_partialKnn_wrapper_15_0__ap_done),
    .krnl_partialKnn_wrapper_15_0__ap_idle(krnl_partialKnn_wrapper_15_0__ap_idle),
    .krnl_partialKnn_wrapper_16_0___in_16__q0(krnl_partialKnn_wrapper_16_0___in_16__q0),
    .krnl_partialKnn_wrapper_16_0__ap_start(krnl_partialKnn_wrapper_16_0__ap_start),
    .krnl_partialKnn_wrapper_16_0__ap_ready(krnl_partialKnn_wrapper_16_0__ap_ready),
    .krnl_partialKnn_wrapper_16_0__ap_done(krnl_partialKnn_wrapper_16_0__ap_done),
    .krnl_partialKnn_wrapper_16_0__ap_idle(krnl_partialKnn_wrapper_16_0__ap_idle),
    .krnl_partialKnn_wrapper_17_0___in_17__q0(krnl_partialKnn_wrapper_17_0___in_17__q0),
    .krnl_partialKnn_wrapper_17_0__ap_start(krnl_partialKnn_wrapper_17_0__ap_start),
    .krnl_partialKnn_wrapper_17_0__ap_ready(krnl_partialKnn_wrapper_17_0__ap_ready),
    .krnl_partialKnn_wrapper_17_0__ap_done(krnl_partialKnn_wrapper_17_0__ap_done),
    .krnl_partialKnn_wrapper_17_0__ap_idle(krnl_partialKnn_wrapper_17_0__ap_idle),
    .krnl_partialKnn_wrapper_18_0___in_18__q0(krnl_partialKnn_wrapper_18_0___in_18__q0),
    .krnl_partialKnn_wrapper_18_0__ap_start(krnl_partialKnn_wrapper_18_0__ap_start),
    .krnl_partialKnn_wrapper_18_0__ap_ready(krnl_partialKnn_wrapper_18_0__ap_ready),
    .krnl_partialKnn_wrapper_18_0__ap_done(krnl_partialKnn_wrapper_18_0__ap_done),
    .krnl_partialKnn_wrapper_18_0__ap_idle(krnl_partialKnn_wrapper_18_0__ap_idle),
    .krnl_partialKnn_wrapper_19_0___in_19__q0(krnl_partialKnn_wrapper_19_0___in_19__q0),
    .krnl_partialKnn_wrapper_19_0__ap_start(krnl_partialKnn_wrapper_19_0__ap_start),
    .krnl_partialKnn_wrapper_19_0__ap_ready(krnl_partialKnn_wrapper_19_0__ap_ready),
    .krnl_partialKnn_wrapper_19_0__ap_done(krnl_partialKnn_wrapper_19_0__ap_done),
    .krnl_partialKnn_wrapper_19_0__ap_idle(krnl_partialKnn_wrapper_19_0__ap_idle),
    .krnl_partialKnn_wrapper_2_0___in_2__q0(krnl_partialKnn_wrapper_2_0___in_2__q0),
    .krnl_partialKnn_wrapper_2_0__ap_start(krnl_partialKnn_wrapper_2_0__ap_start),
    .krnl_partialKnn_wrapper_2_0__ap_ready(krnl_partialKnn_wrapper_2_0__ap_ready),
    .krnl_partialKnn_wrapper_2_0__ap_done(krnl_partialKnn_wrapper_2_0__ap_done),
    .krnl_partialKnn_wrapper_2_0__ap_idle(krnl_partialKnn_wrapper_2_0__ap_idle),
    .krnl_partialKnn_wrapper_20_0___in_20__q0(krnl_partialKnn_wrapper_20_0___in_20__q0),
    .krnl_partialKnn_wrapper_20_0__ap_start(krnl_partialKnn_wrapper_20_0__ap_start),
    .krnl_partialKnn_wrapper_20_0__ap_ready(krnl_partialKnn_wrapper_20_0__ap_ready),
    .krnl_partialKnn_wrapper_20_0__ap_done(krnl_partialKnn_wrapper_20_0__ap_done),
    .krnl_partialKnn_wrapper_20_0__ap_idle(krnl_partialKnn_wrapper_20_0__ap_idle),
    .krnl_partialKnn_wrapper_21_0___in_21__q0(krnl_partialKnn_wrapper_21_0___in_21__q0),
    .krnl_partialKnn_wrapper_21_0__ap_start(krnl_partialKnn_wrapper_21_0__ap_start),
    .krnl_partialKnn_wrapper_21_0__ap_ready(krnl_partialKnn_wrapper_21_0__ap_ready),
    .krnl_partialKnn_wrapper_21_0__ap_done(krnl_partialKnn_wrapper_21_0__ap_done),
    .krnl_partialKnn_wrapper_21_0__ap_idle(krnl_partialKnn_wrapper_21_0__ap_idle),
    .krnl_partialKnn_wrapper_22_0___in_22__q0(krnl_partialKnn_wrapper_22_0___in_22__q0),
    .krnl_partialKnn_wrapper_22_0__ap_start(krnl_partialKnn_wrapper_22_0__ap_start),
    .krnl_partialKnn_wrapper_22_0__ap_ready(krnl_partialKnn_wrapper_22_0__ap_ready),
    .krnl_partialKnn_wrapper_22_0__ap_done(krnl_partialKnn_wrapper_22_0__ap_done),
    .krnl_partialKnn_wrapper_22_0__ap_idle(krnl_partialKnn_wrapper_22_0__ap_idle),
    .krnl_partialKnn_wrapper_23_0___in_23__q0(krnl_partialKnn_wrapper_23_0___in_23__q0),
    .krnl_partialKnn_wrapper_23_0__ap_start(krnl_partialKnn_wrapper_23_0__ap_start),
    .krnl_partialKnn_wrapper_23_0__ap_ready(krnl_partialKnn_wrapper_23_0__ap_ready),
    .krnl_partialKnn_wrapper_23_0__ap_done(krnl_partialKnn_wrapper_23_0__ap_done),
    .krnl_partialKnn_wrapper_23_0__ap_idle(krnl_partialKnn_wrapper_23_0__ap_idle),
    .krnl_partialKnn_wrapper_24_0___in_24__q0(krnl_partialKnn_wrapper_24_0___in_24__q0),
    .krnl_partialKnn_wrapper_24_0__ap_start(krnl_partialKnn_wrapper_24_0__ap_start),
    .krnl_partialKnn_wrapper_24_0__ap_ready(krnl_partialKnn_wrapper_24_0__ap_ready),
    .krnl_partialKnn_wrapper_24_0__ap_done(krnl_partialKnn_wrapper_24_0__ap_done),
    .krnl_partialKnn_wrapper_24_0__ap_idle(krnl_partialKnn_wrapper_24_0__ap_idle),
    .krnl_partialKnn_wrapper_25_0___in_25__q0(krnl_partialKnn_wrapper_25_0___in_25__q0),
    .krnl_partialKnn_wrapper_25_0__ap_start(krnl_partialKnn_wrapper_25_0__ap_start),
    .krnl_partialKnn_wrapper_25_0__ap_ready(krnl_partialKnn_wrapper_25_0__ap_ready),
    .krnl_partialKnn_wrapper_25_0__ap_done(krnl_partialKnn_wrapper_25_0__ap_done),
    .krnl_partialKnn_wrapper_25_0__ap_idle(krnl_partialKnn_wrapper_25_0__ap_idle),
    .krnl_partialKnn_wrapper_26_0___in_26__q0(krnl_partialKnn_wrapper_26_0___in_26__q0),
    .krnl_partialKnn_wrapper_26_0__ap_start(krnl_partialKnn_wrapper_26_0__ap_start),
    .krnl_partialKnn_wrapper_26_0__ap_ready(krnl_partialKnn_wrapper_26_0__ap_ready),
    .krnl_partialKnn_wrapper_26_0__ap_done(krnl_partialKnn_wrapper_26_0__ap_done),
    .krnl_partialKnn_wrapper_26_0__ap_idle(krnl_partialKnn_wrapper_26_0__ap_idle),
    .krnl_partialKnn_wrapper_3_0___in_3__q0(krnl_partialKnn_wrapper_3_0___in_3__q0),
    .krnl_partialKnn_wrapper_3_0__ap_start(krnl_partialKnn_wrapper_3_0__ap_start),
    .krnl_partialKnn_wrapper_3_0__ap_ready(krnl_partialKnn_wrapper_3_0__ap_ready),
    .krnl_partialKnn_wrapper_3_0__ap_done(krnl_partialKnn_wrapper_3_0__ap_done),
    .krnl_partialKnn_wrapper_3_0__ap_idle(krnl_partialKnn_wrapper_3_0__ap_idle),
    .krnl_partialKnn_wrapper_4_0___in_4__q0(krnl_partialKnn_wrapper_4_0___in_4__q0),
    .krnl_partialKnn_wrapper_4_0__ap_start(krnl_partialKnn_wrapper_4_0__ap_start),
    .krnl_partialKnn_wrapper_4_0__ap_ready(krnl_partialKnn_wrapper_4_0__ap_ready),
    .krnl_partialKnn_wrapper_4_0__ap_done(krnl_partialKnn_wrapper_4_0__ap_done),
    .krnl_partialKnn_wrapper_4_0__ap_idle(krnl_partialKnn_wrapper_4_0__ap_idle),
    .krnl_partialKnn_wrapper_5_0___in_5__q0(krnl_partialKnn_wrapper_5_0___in_5__q0),
    .krnl_partialKnn_wrapper_5_0__ap_start(krnl_partialKnn_wrapper_5_0__ap_start),
    .krnl_partialKnn_wrapper_5_0__ap_ready(krnl_partialKnn_wrapper_5_0__ap_ready),
    .krnl_partialKnn_wrapper_5_0__ap_done(krnl_partialKnn_wrapper_5_0__ap_done),
    .krnl_partialKnn_wrapper_5_0__ap_idle(krnl_partialKnn_wrapper_5_0__ap_idle),
    .krnl_partialKnn_wrapper_6_0___in_6__q0(krnl_partialKnn_wrapper_6_0___in_6__q0),
    .krnl_partialKnn_wrapper_6_0__ap_start(krnl_partialKnn_wrapper_6_0__ap_start),
    .krnl_partialKnn_wrapper_6_0__ap_ready(krnl_partialKnn_wrapper_6_0__ap_ready),
    .krnl_partialKnn_wrapper_6_0__ap_done(krnl_partialKnn_wrapper_6_0__ap_done),
    .krnl_partialKnn_wrapper_6_0__ap_idle(krnl_partialKnn_wrapper_6_0__ap_idle),
    .krnl_partialKnn_wrapper_7_0___in_7__q0(krnl_partialKnn_wrapper_7_0___in_7__q0),
    .krnl_partialKnn_wrapper_7_0__ap_start(krnl_partialKnn_wrapper_7_0__ap_start),
    .krnl_partialKnn_wrapper_7_0__ap_ready(krnl_partialKnn_wrapper_7_0__ap_ready),
    .krnl_partialKnn_wrapper_7_0__ap_done(krnl_partialKnn_wrapper_7_0__ap_done),
    .krnl_partialKnn_wrapper_7_0__ap_idle(krnl_partialKnn_wrapper_7_0__ap_idle),
    .krnl_partialKnn_wrapper_8_0___in_8__q0(krnl_partialKnn_wrapper_8_0___in_8__q0),
    .krnl_partialKnn_wrapper_8_0__ap_start(krnl_partialKnn_wrapper_8_0__ap_start),
    .krnl_partialKnn_wrapper_8_0__ap_ready(krnl_partialKnn_wrapper_8_0__ap_ready),
    .krnl_partialKnn_wrapper_8_0__ap_done(krnl_partialKnn_wrapper_8_0__ap_done),
    .krnl_partialKnn_wrapper_8_0__ap_idle(krnl_partialKnn_wrapper_8_0__ap_idle),
    .krnl_partialKnn_wrapper_9_0___in_9__q0(krnl_partialKnn_wrapper_9_0___in_9__q0),
    .krnl_partialKnn_wrapper_9_0__ap_start(krnl_partialKnn_wrapper_9_0__ap_start),
    .krnl_partialKnn_wrapper_9_0__ap_ready(krnl_partialKnn_wrapper_9_0__ap_ready),
    .krnl_partialKnn_wrapper_9_0__ap_done(krnl_partialKnn_wrapper_9_0__ap_done),
    .krnl_partialKnn_wrapper_9_0__ap_idle(krnl_partialKnn_wrapper_9_0__ap_idle)
  );

  assign ap_rst_n_inv = (~ap_rst_n);

endmodule

