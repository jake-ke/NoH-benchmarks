`timescale 1 ns / 1 ps
 
(* CORE_GENERATION_INFO = "Serpens_Serpens,hls_ip_2023_2_2,{HLS_INPUT_TYPE=cxx,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=0,HLS_INPUT_PART=xcvh1582-vsva3697-2MP-e-S,HLS_INPUT_CLOCK=3.330000,HLS_INPUT_ARCH=others,HLS_SYN_CLOCK=1.000000,HLS_SYN_LAT=0,HLS_SYN_TPT=none,HLS_SYN_MEM=0,HLS_SYN_DSP=0,HLS_SYN_FF=3942,HLS_SYN_LUT=7144,HLS_VERSION=2023_2_2}" *)module __rs_Serpens_aux #(
    parameter C_S_AXI_CONTROL_DATA_WIDTH  = 32,
    parameter C_S_AXI_CONTROL_ADDR_WIDTH  = 10,
    parameter C_S_AXI_DATA_WIDTH          = 32,
    parameter C_S_AXI_CONTROL_WSTRB_WIDTH = 4,
    parameter C_S_AXI_WSTRB_WIDTH         = 4
) (
    input wire                                           s_axi_control_AWVALID,
    output wire                                          s_axi_control_AWREADY,
    input wire  [    (C_S_AXI_CONTROL_ADDR_WIDTH - 1):0] s_axi_control_AWADDR,
    input wire                                           s_axi_control_WVALID,
    output wire                                          s_axi_control_WREADY,
    input wire  [    (C_S_AXI_CONTROL_DATA_WIDTH - 1):0] s_axi_control_WDATA,
    input wire  [   (C_S_AXI_CONTROL_WSTRB_WIDTH - 1):0] s_axi_control_WSTRB,
    input wire                                           s_axi_control_ARVALID,
    output wire                                          s_axi_control_ARREADY,
    input wire  [    (C_S_AXI_CONTROL_ADDR_WIDTH - 1):0] s_axi_control_ARADDR,
    output wire                                          s_axi_control_RVALID,
    input wire                                           s_axi_control_RREADY,
    output wire [    (C_S_AXI_CONTROL_DATA_WIDTH - 1):0] s_axi_control_RDATA,
    output wire [                                   1:0] s_axi_control_RRESP,
    output wire                                          s_axi_control_BVALID,
    input wire                                           s_axi_control_BREADY,
    output wire [                                   1:0] s_axi_control_BRESP,
    input wire                                           ap_clk,
    input wire                                           ap_rst_n,
    output wire                                          interrupt,
    output wire [                                  63:0] m_axi_edge_list_ch_0_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_0_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_0_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_0_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_0_ARLEN,
    output wire                                          m_axi_edge_list_ch_0_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_0_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_0_ARQOS,
    input wire                                           m_axi_edge_list_ch_0_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_0_ARSIZE,
    output wire                                          m_axi_edge_list_ch_0_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_0_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_0_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_0_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_0_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_0_AWLEN,
    output wire                                          m_axi_edge_list_ch_0_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_0_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_0_AWQOS,
    input wire                                           m_axi_edge_list_ch_0_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_0_AWSIZE,
    output wire                                          m_axi_edge_list_ch_0_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_0_BID,
    output wire                                          m_axi_edge_list_ch_0_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_0_BRESP,
    input wire                                           m_axi_edge_list_ch_0_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_0_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_0_RID,
    input wire                                           m_axi_edge_list_ch_0_RLAST,
    output wire                                          m_axi_edge_list_ch_0_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_0_RRESP,
    input wire                                           m_axi_edge_list_ch_0_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_0_WDATA,
    output wire                                          m_axi_edge_list_ch_0_WLAST,
    input wire                                           m_axi_edge_list_ch_0_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_0_WSTRB,
    output wire                                          m_axi_edge_list_ch_0_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_1_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_1_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_1_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_1_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_1_ARLEN,
    output wire                                          m_axi_edge_list_ch_1_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_1_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_1_ARQOS,
    input wire                                           m_axi_edge_list_ch_1_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_1_ARSIZE,
    output wire                                          m_axi_edge_list_ch_1_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_1_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_1_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_1_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_1_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_1_AWLEN,
    output wire                                          m_axi_edge_list_ch_1_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_1_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_1_AWQOS,
    input wire                                           m_axi_edge_list_ch_1_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_1_AWSIZE,
    output wire                                          m_axi_edge_list_ch_1_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_1_BID,
    output wire                                          m_axi_edge_list_ch_1_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_1_BRESP,
    input wire                                           m_axi_edge_list_ch_1_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_1_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_1_RID,
    input wire                                           m_axi_edge_list_ch_1_RLAST,
    output wire                                          m_axi_edge_list_ch_1_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_1_RRESP,
    input wire                                           m_axi_edge_list_ch_1_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_1_WDATA,
    output wire                                          m_axi_edge_list_ch_1_WLAST,
    input wire                                           m_axi_edge_list_ch_1_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_1_WSTRB,
    output wire                                          m_axi_edge_list_ch_1_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_2_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_2_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_2_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_2_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_2_ARLEN,
    output wire                                          m_axi_edge_list_ch_2_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_2_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_2_ARQOS,
    input wire                                           m_axi_edge_list_ch_2_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_2_ARSIZE,
    output wire                                          m_axi_edge_list_ch_2_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_2_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_2_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_2_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_2_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_2_AWLEN,
    output wire                                          m_axi_edge_list_ch_2_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_2_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_2_AWQOS,
    input wire                                           m_axi_edge_list_ch_2_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_2_AWSIZE,
    output wire                                          m_axi_edge_list_ch_2_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_2_BID,
    output wire                                          m_axi_edge_list_ch_2_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_2_BRESP,
    input wire                                           m_axi_edge_list_ch_2_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_2_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_2_RID,
    input wire                                           m_axi_edge_list_ch_2_RLAST,
    output wire                                          m_axi_edge_list_ch_2_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_2_RRESP,
    input wire                                           m_axi_edge_list_ch_2_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_2_WDATA,
    output wire                                          m_axi_edge_list_ch_2_WLAST,
    input wire                                           m_axi_edge_list_ch_2_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_2_WSTRB,
    output wire                                          m_axi_edge_list_ch_2_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_3_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_3_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_3_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_3_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_3_ARLEN,
    output wire                                          m_axi_edge_list_ch_3_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_3_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_3_ARQOS,
    input wire                                           m_axi_edge_list_ch_3_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_3_ARSIZE,
    output wire                                          m_axi_edge_list_ch_3_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_3_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_3_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_3_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_3_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_3_AWLEN,
    output wire                                          m_axi_edge_list_ch_3_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_3_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_3_AWQOS,
    input wire                                           m_axi_edge_list_ch_3_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_3_AWSIZE,
    output wire                                          m_axi_edge_list_ch_3_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_3_BID,
    output wire                                          m_axi_edge_list_ch_3_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_3_BRESP,
    input wire                                           m_axi_edge_list_ch_3_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_3_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_3_RID,
    input wire                                           m_axi_edge_list_ch_3_RLAST,
    output wire                                          m_axi_edge_list_ch_3_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_3_RRESP,
    input wire                                           m_axi_edge_list_ch_3_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_3_WDATA,
    output wire                                          m_axi_edge_list_ch_3_WLAST,
    input wire                                           m_axi_edge_list_ch_3_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_3_WSTRB,
    output wire                                          m_axi_edge_list_ch_3_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_4_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_4_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_4_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_4_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_4_ARLEN,
    output wire                                          m_axi_edge_list_ch_4_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_4_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_4_ARQOS,
    input wire                                           m_axi_edge_list_ch_4_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_4_ARSIZE,
    output wire                                          m_axi_edge_list_ch_4_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_4_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_4_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_4_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_4_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_4_AWLEN,
    output wire                                          m_axi_edge_list_ch_4_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_4_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_4_AWQOS,
    input wire                                           m_axi_edge_list_ch_4_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_4_AWSIZE,
    output wire                                          m_axi_edge_list_ch_4_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_4_BID,
    output wire                                          m_axi_edge_list_ch_4_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_4_BRESP,
    input wire                                           m_axi_edge_list_ch_4_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_4_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_4_RID,
    input wire                                           m_axi_edge_list_ch_4_RLAST,
    output wire                                          m_axi_edge_list_ch_4_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_4_RRESP,
    input wire                                           m_axi_edge_list_ch_4_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_4_WDATA,
    output wire                                          m_axi_edge_list_ch_4_WLAST,
    input wire                                           m_axi_edge_list_ch_4_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_4_WSTRB,
    output wire                                          m_axi_edge_list_ch_4_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_5_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_5_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_5_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_5_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_5_ARLEN,
    output wire                                          m_axi_edge_list_ch_5_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_5_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_5_ARQOS,
    input wire                                           m_axi_edge_list_ch_5_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_5_ARSIZE,
    output wire                                          m_axi_edge_list_ch_5_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_5_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_5_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_5_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_5_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_5_AWLEN,
    output wire                                          m_axi_edge_list_ch_5_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_5_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_5_AWQOS,
    input wire                                           m_axi_edge_list_ch_5_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_5_AWSIZE,
    output wire                                          m_axi_edge_list_ch_5_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_5_BID,
    output wire                                          m_axi_edge_list_ch_5_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_5_BRESP,
    input wire                                           m_axi_edge_list_ch_5_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_5_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_5_RID,
    input wire                                           m_axi_edge_list_ch_5_RLAST,
    output wire                                          m_axi_edge_list_ch_5_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_5_RRESP,
    input wire                                           m_axi_edge_list_ch_5_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_5_WDATA,
    output wire                                          m_axi_edge_list_ch_5_WLAST,
    input wire                                           m_axi_edge_list_ch_5_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_5_WSTRB,
    output wire                                          m_axi_edge_list_ch_5_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_6_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_6_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_6_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_6_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_6_ARLEN,
    output wire                                          m_axi_edge_list_ch_6_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_6_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_6_ARQOS,
    input wire                                           m_axi_edge_list_ch_6_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_6_ARSIZE,
    output wire                                          m_axi_edge_list_ch_6_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_6_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_6_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_6_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_6_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_6_AWLEN,
    output wire                                          m_axi_edge_list_ch_6_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_6_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_6_AWQOS,
    input wire                                           m_axi_edge_list_ch_6_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_6_AWSIZE,
    output wire                                          m_axi_edge_list_ch_6_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_6_BID,
    output wire                                          m_axi_edge_list_ch_6_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_6_BRESP,
    input wire                                           m_axi_edge_list_ch_6_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_6_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_6_RID,
    input wire                                           m_axi_edge_list_ch_6_RLAST,
    output wire                                          m_axi_edge_list_ch_6_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_6_RRESP,
    input wire                                           m_axi_edge_list_ch_6_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_6_WDATA,
    output wire                                          m_axi_edge_list_ch_6_WLAST,
    input wire                                           m_axi_edge_list_ch_6_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_6_WSTRB,
    output wire                                          m_axi_edge_list_ch_6_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_7_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_7_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_7_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_7_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_7_ARLEN,
    output wire                                          m_axi_edge_list_ch_7_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_7_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_7_ARQOS,
    input wire                                           m_axi_edge_list_ch_7_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_7_ARSIZE,
    output wire                                          m_axi_edge_list_ch_7_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_7_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_7_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_7_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_7_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_7_AWLEN,
    output wire                                          m_axi_edge_list_ch_7_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_7_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_7_AWQOS,
    input wire                                           m_axi_edge_list_ch_7_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_7_AWSIZE,
    output wire                                          m_axi_edge_list_ch_7_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_7_BID,
    output wire                                          m_axi_edge_list_ch_7_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_7_BRESP,
    input wire                                           m_axi_edge_list_ch_7_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_7_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_7_RID,
    input wire                                           m_axi_edge_list_ch_7_RLAST,
    output wire                                          m_axi_edge_list_ch_7_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_7_RRESP,
    input wire                                           m_axi_edge_list_ch_7_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_7_WDATA,
    output wire                                          m_axi_edge_list_ch_7_WLAST,
    input wire                                           m_axi_edge_list_ch_7_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_7_WSTRB,
    output wire                                          m_axi_edge_list_ch_7_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_8_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_8_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_8_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_8_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_8_ARLEN,
    output wire                                          m_axi_edge_list_ch_8_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_8_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_8_ARQOS,
    input wire                                           m_axi_edge_list_ch_8_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_8_ARSIZE,
    output wire                                          m_axi_edge_list_ch_8_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_8_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_8_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_8_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_8_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_8_AWLEN,
    output wire                                          m_axi_edge_list_ch_8_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_8_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_8_AWQOS,
    input wire                                           m_axi_edge_list_ch_8_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_8_AWSIZE,
    output wire                                          m_axi_edge_list_ch_8_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_8_BID,
    output wire                                          m_axi_edge_list_ch_8_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_8_BRESP,
    input wire                                           m_axi_edge_list_ch_8_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_8_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_8_RID,
    input wire                                           m_axi_edge_list_ch_8_RLAST,
    output wire                                          m_axi_edge_list_ch_8_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_8_RRESP,
    input wire                                           m_axi_edge_list_ch_8_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_8_WDATA,
    output wire                                          m_axi_edge_list_ch_8_WLAST,
    input wire                                           m_axi_edge_list_ch_8_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_8_WSTRB,
    output wire                                          m_axi_edge_list_ch_8_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_9_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_9_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_9_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_9_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_9_ARLEN,
    output wire                                          m_axi_edge_list_ch_9_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_9_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_9_ARQOS,
    input wire                                           m_axi_edge_list_ch_9_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_9_ARSIZE,
    output wire                                          m_axi_edge_list_ch_9_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_9_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_9_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_9_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_9_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_9_AWLEN,
    output wire                                          m_axi_edge_list_ch_9_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_9_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_9_AWQOS,
    input wire                                           m_axi_edge_list_ch_9_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_9_AWSIZE,
    output wire                                          m_axi_edge_list_ch_9_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_9_BID,
    output wire                                          m_axi_edge_list_ch_9_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_9_BRESP,
    input wire                                           m_axi_edge_list_ch_9_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_9_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_9_RID,
    input wire                                           m_axi_edge_list_ch_9_RLAST,
    output wire                                          m_axi_edge_list_ch_9_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_9_RRESP,
    input wire                                           m_axi_edge_list_ch_9_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_9_WDATA,
    output wire                                          m_axi_edge_list_ch_9_WLAST,
    input wire                                           m_axi_edge_list_ch_9_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_9_WSTRB,
    output wire                                          m_axi_edge_list_ch_9_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_10_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_10_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_10_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_10_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_10_ARLEN,
    output wire                                          m_axi_edge_list_ch_10_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_10_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_10_ARQOS,
    input wire                                           m_axi_edge_list_ch_10_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_10_ARSIZE,
    output wire                                          m_axi_edge_list_ch_10_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_10_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_10_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_10_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_10_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_10_AWLEN,
    output wire                                          m_axi_edge_list_ch_10_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_10_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_10_AWQOS,
    input wire                                           m_axi_edge_list_ch_10_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_10_AWSIZE,
    output wire                                          m_axi_edge_list_ch_10_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_10_BID,
    output wire                                          m_axi_edge_list_ch_10_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_10_BRESP,
    input wire                                           m_axi_edge_list_ch_10_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_10_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_10_RID,
    input wire                                           m_axi_edge_list_ch_10_RLAST,
    output wire                                          m_axi_edge_list_ch_10_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_10_RRESP,
    input wire                                           m_axi_edge_list_ch_10_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_10_WDATA,
    output wire                                          m_axi_edge_list_ch_10_WLAST,
    input wire                                           m_axi_edge_list_ch_10_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_10_WSTRB,
    output wire                                          m_axi_edge_list_ch_10_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_11_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_11_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_11_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_11_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_11_ARLEN,
    output wire                                          m_axi_edge_list_ch_11_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_11_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_11_ARQOS,
    input wire                                           m_axi_edge_list_ch_11_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_11_ARSIZE,
    output wire                                          m_axi_edge_list_ch_11_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_11_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_11_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_11_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_11_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_11_AWLEN,
    output wire                                          m_axi_edge_list_ch_11_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_11_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_11_AWQOS,
    input wire                                           m_axi_edge_list_ch_11_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_11_AWSIZE,
    output wire                                          m_axi_edge_list_ch_11_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_11_BID,
    output wire                                          m_axi_edge_list_ch_11_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_11_BRESP,
    input wire                                           m_axi_edge_list_ch_11_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_11_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_11_RID,
    input wire                                           m_axi_edge_list_ch_11_RLAST,
    output wire                                          m_axi_edge_list_ch_11_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_11_RRESP,
    input wire                                           m_axi_edge_list_ch_11_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_11_WDATA,
    output wire                                          m_axi_edge_list_ch_11_WLAST,
    input wire                                           m_axi_edge_list_ch_11_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_11_WSTRB,
    output wire                                          m_axi_edge_list_ch_11_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_12_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_12_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_12_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_12_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_12_ARLEN,
    output wire                                          m_axi_edge_list_ch_12_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_12_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_12_ARQOS,
    input wire                                           m_axi_edge_list_ch_12_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_12_ARSIZE,
    output wire                                          m_axi_edge_list_ch_12_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_12_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_12_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_12_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_12_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_12_AWLEN,
    output wire                                          m_axi_edge_list_ch_12_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_12_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_12_AWQOS,
    input wire                                           m_axi_edge_list_ch_12_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_12_AWSIZE,
    output wire                                          m_axi_edge_list_ch_12_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_12_BID,
    output wire                                          m_axi_edge_list_ch_12_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_12_BRESP,
    input wire                                           m_axi_edge_list_ch_12_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_12_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_12_RID,
    input wire                                           m_axi_edge_list_ch_12_RLAST,
    output wire                                          m_axi_edge_list_ch_12_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_12_RRESP,
    input wire                                           m_axi_edge_list_ch_12_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_12_WDATA,
    output wire                                          m_axi_edge_list_ch_12_WLAST,
    input wire                                           m_axi_edge_list_ch_12_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_12_WSTRB,
    output wire                                          m_axi_edge_list_ch_12_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_13_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_13_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_13_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_13_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_13_ARLEN,
    output wire                                          m_axi_edge_list_ch_13_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_13_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_13_ARQOS,
    input wire                                           m_axi_edge_list_ch_13_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_13_ARSIZE,
    output wire                                          m_axi_edge_list_ch_13_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_13_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_13_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_13_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_13_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_13_AWLEN,
    output wire                                          m_axi_edge_list_ch_13_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_13_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_13_AWQOS,
    input wire                                           m_axi_edge_list_ch_13_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_13_AWSIZE,
    output wire                                          m_axi_edge_list_ch_13_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_13_BID,
    output wire                                          m_axi_edge_list_ch_13_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_13_BRESP,
    input wire                                           m_axi_edge_list_ch_13_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_13_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_13_RID,
    input wire                                           m_axi_edge_list_ch_13_RLAST,
    output wire                                          m_axi_edge_list_ch_13_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_13_RRESP,
    input wire                                           m_axi_edge_list_ch_13_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_13_WDATA,
    output wire                                          m_axi_edge_list_ch_13_WLAST,
    input wire                                           m_axi_edge_list_ch_13_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_13_WSTRB,
    output wire                                          m_axi_edge_list_ch_13_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_14_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_14_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_14_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_14_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_14_ARLEN,
    output wire                                          m_axi_edge_list_ch_14_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_14_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_14_ARQOS,
    input wire                                           m_axi_edge_list_ch_14_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_14_ARSIZE,
    output wire                                          m_axi_edge_list_ch_14_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_14_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_14_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_14_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_14_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_14_AWLEN,
    output wire                                          m_axi_edge_list_ch_14_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_14_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_14_AWQOS,
    input wire                                           m_axi_edge_list_ch_14_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_14_AWSIZE,
    output wire                                          m_axi_edge_list_ch_14_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_14_BID,
    output wire                                          m_axi_edge_list_ch_14_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_14_BRESP,
    input wire                                           m_axi_edge_list_ch_14_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_14_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_14_RID,
    input wire                                           m_axi_edge_list_ch_14_RLAST,
    output wire                                          m_axi_edge_list_ch_14_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_14_RRESP,
    input wire                                           m_axi_edge_list_ch_14_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_14_WDATA,
    output wire                                          m_axi_edge_list_ch_14_WLAST,
    input wire                                           m_axi_edge_list_ch_14_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_14_WSTRB,
    output wire                                          m_axi_edge_list_ch_14_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_15_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_15_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_15_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_15_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_15_ARLEN,
    output wire                                          m_axi_edge_list_ch_15_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_15_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_15_ARQOS,
    input wire                                           m_axi_edge_list_ch_15_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_15_ARSIZE,
    output wire                                          m_axi_edge_list_ch_15_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_15_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_15_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_15_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_15_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_15_AWLEN,
    output wire                                          m_axi_edge_list_ch_15_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_15_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_15_AWQOS,
    input wire                                           m_axi_edge_list_ch_15_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_15_AWSIZE,
    output wire                                          m_axi_edge_list_ch_15_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_15_BID,
    output wire                                          m_axi_edge_list_ch_15_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_15_BRESP,
    input wire                                           m_axi_edge_list_ch_15_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_15_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_15_RID,
    input wire                                           m_axi_edge_list_ch_15_RLAST,
    output wire                                          m_axi_edge_list_ch_15_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_15_RRESP,
    input wire                                           m_axi_edge_list_ch_15_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_15_WDATA,
    output wire                                          m_axi_edge_list_ch_15_WLAST,
    input wire                                           m_axi_edge_list_ch_15_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_15_WSTRB,
    output wire                                          m_axi_edge_list_ch_15_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_16_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_16_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_16_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_16_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_16_ARLEN,
    output wire                                          m_axi_edge_list_ch_16_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_16_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_16_ARQOS,
    input wire                                           m_axi_edge_list_ch_16_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_16_ARSIZE,
    output wire                                          m_axi_edge_list_ch_16_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_16_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_16_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_16_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_16_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_16_AWLEN,
    output wire                                          m_axi_edge_list_ch_16_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_16_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_16_AWQOS,
    input wire                                           m_axi_edge_list_ch_16_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_16_AWSIZE,
    output wire                                          m_axi_edge_list_ch_16_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_16_BID,
    output wire                                          m_axi_edge_list_ch_16_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_16_BRESP,
    input wire                                           m_axi_edge_list_ch_16_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_16_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_16_RID,
    input wire                                           m_axi_edge_list_ch_16_RLAST,
    output wire                                          m_axi_edge_list_ch_16_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_16_RRESP,
    input wire                                           m_axi_edge_list_ch_16_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_16_WDATA,
    output wire                                          m_axi_edge_list_ch_16_WLAST,
    input wire                                           m_axi_edge_list_ch_16_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_16_WSTRB,
    output wire                                          m_axi_edge_list_ch_16_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_17_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_17_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_17_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_17_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_17_ARLEN,
    output wire                                          m_axi_edge_list_ch_17_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_17_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_17_ARQOS,
    input wire                                           m_axi_edge_list_ch_17_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_17_ARSIZE,
    output wire                                          m_axi_edge_list_ch_17_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_17_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_17_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_17_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_17_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_17_AWLEN,
    output wire                                          m_axi_edge_list_ch_17_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_17_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_17_AWQOS,
    input wire                                           m_axi_edge_list_ch_17_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_17_AWSIZE,
    output wire                                          m_axi_edge_list_ch_17_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_17_BID,
    output wire                                          m_axi_edge_list_ch_17_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_17_BRESP,
    input wire                                           m_axi_edge_list_ch_17_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_17_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_17_RID,
    input wire                                           m_axi_edge_list_ch_17_RLAST,
    output wire                                          m_axi_edge_list_ch_17_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_17_RRESP,
    input wire                                           m_axi_edge_list_ch_17_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_17_WDATA,
    output wire                                          m_axi_edge_list_ch_17_WLAST,
    input wire                                           m_axi_edge_list_ch_17_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_17_WSTRB,
    output wire                                          m_axi_edge_list_ch_17_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_18_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_18_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_18_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_18_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_18_ARLEN,
    output wire                                          m_axi_edge_list_ch_18_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_18_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_18_ARQOS,
    input wire                                           m_axi_edge_list_ch_18_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_18_ARSIZE,
    output wire                                          m_axi_edge_list_ch_18_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_18_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_18_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_18_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_18_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_18_AWLEN,
    output wire                                          m_axi_edge_list_ch_18_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_18_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_18_AWQOS,
    input wire                                           m_axi_edge_list_ch_18_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_18_AWSIZE,
    output wire                                          m_axi_edge_list_ch_18_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_18_BID,
    output wire                                          m_axi_edge_list_ch_18_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_18_BRESP,
    input wire                                           m_axi_edge_list_ch_18_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_18_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_18_RID,
    input wire                                           m_axi_edge_list_ch_18_RLAST,
    output wire                                          m_axi_edge_list_ch_18_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_18_RRESP,
    input wire                                           m_axi_edge_list_ch_18_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_18_WDATA,
    output wire                                          m_axi_edge_list_ch_18_WLAST,
    input wire                                           m_axi_edge_list_ch_18_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_18_WSTRB,
    output wire                                          m_axi_edge_list_ch_18_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_19_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_19_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_19_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_19_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_19_ARLEN,
    output wire                                          m_axi_edge_list_ch_19_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_19_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_19_ARQOS,
    input wire                                           m_axi_edge_list_ch_19_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_19_ARSIZE,
    output wire                                          m_axi_edge_list_ch_19_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_19_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_19_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_19_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_19_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_19_AWLEN,
    output wire                                          m_axi_edge_list_ch_19_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_19_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_19_AWQOS,
    input wire                                           m_axi_edge_list_ch_19_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_19_AWSIZE,
    output wire                                          m_axi_edge_list_ch_19_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_19_BID,
    output wire                                          m_axi_edge_list_ch_19_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_19_BRESP,
    input wire                                           m_axi_edge_list_ch_19_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_19_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_19_RID,
    input wire                                           m_axi_edge_list_ch_19_RLAST,
    output wire                                          m_axi_edge_list_ch_19_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_19_RRESP,
    input wire                                           m_axi_edge_list_ch_19_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_19_WDATA,
    output wire                                          m_axi_edge_list_ch_19_WLAST,
    input wire                                           m_axi_edge_list_ch_19_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_19_WSTRB,
    output wire                                          m_axi_edge_list_ch_19_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_20_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_20_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_20_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_20_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_20_ARLEN,
    output wire                                          m_axi_edge_list_ch_20_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_20_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_20_ARQOS,
    input wire                                           m_axi_edge_list_ch_20_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_20_ARSIZE,
    output wire                                          m_axi_edge_list_ch_20_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_20_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_20_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_20_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_20_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_20_AWLEN,
    output wire                                          m_axi_edge_list_ch_20_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_20_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_20_AWQOS,
    input wire                                           m_axi_edge_list_ch_20_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_20_AWSIZE,
    output wire                                          m_axi_edge_list_ch_20_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_20_BID,
    output wire                                          m_axi_edge_list_ch_20_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_20_BRESP,
    input wire                                           m_axi_edge_list_ch_20_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_20_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_20_RID,
    input wire                                           m_axi_edge_list_ch_20_RLAST,
    output wire                                          m_axi_edge_list_ch_20_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_20_RRESP,
    input wire                                           m_axi_edge_list_ch_20_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_20_WDATA,
    output wire                                          m_axi_edge_list_ch_20_WLAST,
    input wire                                           m_axi_edge_list_ch_20_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_20_WSTRB,
    output wire                                          m_axi_edge_list_ch_20_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_21_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_21_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_21_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_21_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_21_ARLEN,
    output wire                                          m_axi_edge_list_ch_21_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_21_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_21_ARQOS,
    input wire                                           m_axi_edge_list_ch_21_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_21_ARSIZE,
    output wire                                          m_axi_edge_list_ch_21_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_21_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_21_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_21_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_21_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_21_AWLEN,
    output wire                                          m_axi_edge_list_ch_21_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_21_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_21_AWQOS,
    input wire                                           m_axi_edge_list_ch_21_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_21_AWSIZE,
    output wire                                          m_axi_edge_list_ch_21_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_21_BID,
    output wire                                          m_axi_edge_list_ch_21_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_21_BRESP,
    input wire                                           m_axi_edge_list_ch_21_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_21_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_21_RID,
    input wire                                           m_axi_edge_list_ch_21_RLAST,
    output wire                                          m_axi_edge_list_ch_21_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_21_RRESP,
    input wire                                           m_axi_edge_list_ch_21_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_21_WDATA,
    output wire                                          m_axi_edge_list_ch_21_WLAST,
    input wire                                           m_axi_edge_list_ch_21_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_21_WSTRB,
    output wire                                          m_axi_edge_list_ch_21_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_22_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_22_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_22_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_22_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_22_ARLEN,
    output wire                                          m_axi_edge_list_ch_22_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_22_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_22_ARQOS,
    input wire                                           m_axi_edge_list_ch_22_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_22_ARSIZE,
    output wire                                          m_axi_edge_list_ch_22_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_22_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_22_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_22_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_22_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_22_AWLEN,
    output wire                                          m_axi_edge_list_ch_22_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_22_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_22_AWQOS,
    input wire                                           m_axi_edge_list_ch_22_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_22_AWSIZE,
    output wire                                          m_axi_edge_list_ch_22_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_22_BID,
    output wire                                          m_axi_edge_list_ch_22_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_22_BRESP,
    input wire                                           m_axi_edge_list_ch_22_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_22_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_22_RID,
    input wire                                           m_axi_edge_list_ch_22_RLAST,
    output wire                                          m_axi_edge_list_ch_22_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_22_RRESP,
    input wire                                           m_axi_edge_list_ch_22_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_22_WDATA,
    output wire                                          m_axi_edge_list_ch_22_WLAST,
    input wire                                           m_axi_edge_list_ch_22_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_22_WSTRB,
    output wire                                          m_axi_edge_list_ch_22_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_23_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_23_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_23_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_23_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_23_ARLEN,
    output wire                                          m_axi_edge_list_ch_23_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_23_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_23_ARQOS,
    input wire                                           m_axi_edge_list_ch_23_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_23_ARSIZE,
    output wire                                          m_axi_edge_list_ch_23_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_23_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_23_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_23_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_23_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_23_AWLEN,
    output wire                                          m_axi_edge_list_ch_23_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_23_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_23_AWQOS,
    input wire                                           m_axi_edge_list_ch_23_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_23_AWSIZE,
    output wire                                          m_axi_edge_list_ch_23_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_23_BID,
    output wire                                          m_axi_edge_list_ch_23_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_23_BRESP,
    input wire                                           m_axi_edge_list_ch_23_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_23_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_23_RID,
    input wire                                           m_axi_edge_list_ch_23_RLAST,
    output wire                                          m_axi_edge_list_ch_23_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_23_RRESP,
    input wire                                           m_axi_edge_list_ch_23_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_23_WDATA,
    output wire                                          m_axi_edge_list_ch_23_WLAST,
    input wire                                           m_axi_edge_list_ch_23_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_23_WSTRB,
    output wire                                          m_axi_edge_list_ch_23_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_24_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_24_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_24_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_24_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_24_ARLEN,
    output wire                                          m_axi_edge_list_ch_24_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_24_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_24_ARQOS,
    input wire                                           m_axi_edge_list_ch_24_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_24_ARSIZE,
    output wire                                          m_axi_edge_list_ch_24_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_24_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_24_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_24_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_24_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_24_AWLEN,
    output wire                                          m_axi_edge_list_ch_24_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_24_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_24_AWQOS,
    input wire                                           m_axi_edge_list_ch_24_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_24_AWSIZE,
    output wire                                          m_axi_edge_list_ch_24_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_24_BID,
    output wire                                          m_axi_edge_list_ch_24_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_24_BRESP,
    input wire                                           m_axi_edge_list_ch_24_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_24_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_24_RID,
    input wire                                           m_axi_edge_list_ch_24_RLAST,
    output wire                                          m_axi_edge_list_ch_24_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_24_RRESP,
    input wire                                           m_axi_edge_list_ch_24_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_24_WDATA,
    output wire                                          m_axi_edge_list_ch_24_WLAST,
    input wire                                           m_axi_edge_list_ch_24_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_24_WSTRB,
    output wire                                          m_axi_edge_list_ch_24_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_25_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_25_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_25_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_25_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_25_ARLEN,
    output wire                                          m_axi_edge_list_ch_25_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_25_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_25_ARQOS,
    input wire                                           m_axi_edge_list_ch_25_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_25_ARSIZE,
    output wire                                          m_axi_edge_list_ch_25_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_25_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_25_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_25_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_25_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_25_AWLEN,
    output wire                                          m_axi_edge_list_ch_25_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_25_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_25_AWQOS,
    input wire                                           m_axi_edge_list_ch_25_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_25_AWSIZE,
    output wire                                          m_axi_edge_list_ch_25_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_25_BID,
    output wire                                          m_axi_edge_list_ch_25_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_25_BRESP,
    input wire                                           m_axi_edge_list_ch_25_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_25_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_25_RID,
    input wire                                           m_axi_edge_list_ch_25_RLAST,
    output wire                                          m_axi_edge_list_ch_25_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_25_RRESP,
    input wire                                           m_axi_edge_list_ch_25_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_25_WDATA,
    output wire                                          m_axi_edge_list_ch_25_WLAST,
    input wire                                           m_axi_edge_list_ch_25_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_25_WSTRB,
    output wire                                          m_axi_edge_list_ch_25_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_26_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_26_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_26_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_26_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_26_ARLEN,
    output wire                                          m_axi_edge_list_ch_26_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_26_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_26_ARQOS,
    input wire                                           m_axi_edge_list_ch_26_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_26_ARSIZE,
    output wire                                          m_axi_edge_list_ch_26_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_26_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_26_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_26_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_26_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_26_AWLEN,
    output wire                                          m_axi_edge_list_ch_26_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_26_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_26_AWQOS,
    input wire                                           m_axi_edge_list_ch_26_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_26_AWSIZE,
    output wire                                          m_axi_edge_list_ch_26_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_26_BID,
    output wire                                          m_axi_edge_list_ch_26_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_26_BRESP,
    input wire                                           m_axi_edge_list_ch_26_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_26_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_26_RID,
    input wire                                           m_axi_edge_list_ch_26_RLAST,
    output wire                                          m_axi_edge_list_ch_26_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_26_RRESP,
    input wire                                           m_axi_edge_list_ch_26_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_26_WDATA,
    output wire                                          m_axi_edge_list_ch_26_WLAST,
    input wire                                           m_axi_edge_list_ch_26_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_26_WSTRB,
    output wire                                          m_axi_edge_list_ch_26_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_27_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_27_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_27_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_27_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_27_ARLEN,
    output wire                                          m_axi_edge_list_ch_27_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_27_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_27_ARQOS,
    input wire                                           m_axi_edge_list_ch_27_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_27_ARSIZE,
    output wire                                          m_axi_edge_list_ch_27_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_27_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_27_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_27_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_27_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_27_AWLEN,
    output wire                                          m_axi_edge_list_ch_27_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_27_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_27_AWQOS,
    input wire                                           m_axi_edge_list_ch_27_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_27_AWSIZE,
    output wire                                          m_axi_edge_list_ch_27_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_27_BID,
    output wire                                          m_axi_edge_list_ch_27_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_27_BRESP,
    input wire                                           m_axi_edge_list_ch_27_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_27_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_27_RID,
    input wire                                           m_axi_edge_list_ch_27_RLAST,
    output wire                                          m_axi_edge_list_ch_27_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_27_RRESP,
    input wire                                           m_axi_edge_list_ch_27_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_27_WDATA,
    output wire                                          m_axi_edge_list_ch_27_WLAST,
    input wire                                           m_axi_edge_list_ch_27_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_27_WSTRB,
    output wire                                          m_axi_edge_list_ch_27_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_28_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_28_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_28_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_28_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_28_ARLEN,
    output wire                                          m_axi_edge_list_ch_28_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_28_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_28_ARQOS,
    input wire                                           m_axi_edge_list_ch_28_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_28_ARSIZE,
    output wire                                          m_axi_edge_list_ch_28_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_28_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_28_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_28_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_28_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_28_AWLEN,
    output wire                                          m_axi_edge_list_ch_28_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_28_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_28_AWQOS,
    input wire                                           m_axi_edge_list_ch_28_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_28_AWSIZE,
    output wire                                          m_axi_edge_list_ch_28_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_28_BID,
    output wire                                          m_axi_edge_list_ch_28_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_28_BRESP,
    input wire                                           m_axi_edge_list_ch_28_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_28_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_28_RID,
    input wire                                           m_axi_edge_list_ch_28_RLAST,
    output wire                                          m_axi_edge_list_ch_28_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_28_RRESP,
    input wire                                           m_axi_edge_list_ch_28_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_28_WDATA,
    output wire                                          m_axi_edge_list_ch_28_WLAST,
    input wire                                           m_axi_edge_list_ch_28_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_28_WSTRB,
    output wire                                          m_axi_edge_list_ch_28_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_29_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_29_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_29_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_29_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_29_ARLEN,
    output wire                                          m_axi_edge_list_ch_29_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_29_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_29_ARQOS,
    input wire                                           m_axi_edge_list_ch_29_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_29_ARSIZE,
    output wire                                          m_axi_edge_list_ch_29_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_29_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_29_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_29_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_29_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_29_AWLEN,
    output wire                                          m_axi_edge_list_ch_29_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_29_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_29_AWQOS,
    input wire                                           m_axi_edge_list_ch_29_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_29_AWSIZE,
    output wire                                          m_axi_edge_list_ch_29_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_29_BID,
    output wire                                          m_axi_edge_list_ch_29_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_29_BRESP,
    input wire                                           m_axi_edge_list_ch_29_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_29_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_29_RID,
    input wire                                           m_axi_edge_list_ch_29_RLAST,
    output wire                                          m_axi_edge_list_ch_29_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_29_RRESP,
    input wire                                           m_axi_edge_list_ch_29_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_29_WDATA,
    output wire                                          m_axi_edge_list_ch_29_WLAST,
    input wire                                           m_axi_edge_list_ch_29_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_29_WSTRB,
    output wire                                          m_axi_edge_list_ch_29_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_30_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_30_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_30_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_30_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_30_ARLEN,
    output wire                                          m_axi_edge_list_ch_30_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_30_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_30_ARQOS,
    input wire                                           m_axi_edge_list_ch_30_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_30_ARSIZE,
    output wire                                          m_axi_edge_list_ch_30_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_30_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_30_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_30_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_30_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_30_AWLEN,
    output wire                                          m_axi_edge_list_ch_30_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_30_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_30_AWQOS,
    input wire                                           m_axi_edge_list_ch_30_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_30_AWSIZE,
    output wire                                          m_axi_edge_list_ch_30_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_30_BID,
    output wire                                          m_axi_edge_list_ch_30_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_30_BRESP,
    input wire                                           m_axi_edge_list_ch_30_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_30_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_30_RID,
    input wire                                           m_axi_edge_list_ch_30_RLAST,
    output wire                                          m_axi_edge_list_ch_30_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_30_RRESP,
    input wire                                           m_axi_edge_list_ch_30_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_30_WDATA,
    output wire                                          m_axi_edge_list_ch_30_WLAST,
    input wire                                           m_axi_edge_list_ch_30_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_30_WSTRB,
    output wire                                          m_axi_edge_list_ch_30_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_31_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_31_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_31_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_31_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_31_ARLEN,
    output wire                                          m_axi_edge_list_ch_31_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_31_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_31_ARQOS,
    input wire                                           m_axi_edge_list_ch_31_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_31_ARSIZE,
    output wire                                          m_axi_edge_list_ch_31_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_31_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_31_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_31_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_31_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_31_AWLEN,
    output wire                                          m_axi_edge_list_ch_31_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_31_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_31_AWQOS,
    input wire                                           m_axi_edge_list_ch_31_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_31_AWSIZE,
    output wire                                          m_axi_edge_list_ch_31_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_31_BID,
    output wire                                          m_axi_edge_list_ch_31_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_31_BRESP,
    input wire                                           m_axi_edge_list_ch_31_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_31_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_31_RID,
    input wire                                           m_axi_edge_list_ch_31_RLAST,
    output wire                                          m_axi_edge_list_ch_31_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_31_RRESP,
    input wire                                           m_axi_edge_list_ch_31_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_31_WDATA,
    output wire                                          m_axi_edge_list_ch_31_WLAST,
    input wire                                           m_axi_edge_list_ch_31_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_31_WSTRB,
    output wire                                          m_axi_edge_list_ch_31_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_32_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_32_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_32_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_32_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_32_ARLEN,
    output wire                                          m_axi_edge_list_ch_32_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_32_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_32_ARQOS,
    input wire                                           m_axi_edge_list_ch_32_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_32_ARSIZE,
    output wire                                          m_axi_edge_list_ch_32_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_32_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_32_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_32_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_32_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_32_AWLEN,
    output wire                                          m_axi_edge_list_ch_32_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_32_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_32_AWQOS,
    input wire                                           m_axi_edge_list_ch_32_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_32_AWSIZE,
    output wire                                          m_axi_edge_list_ch_32_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_32_BID,
    output wire                                          m_axi_edge_list_ch_32_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_32_BRESP,
    input wire                                           m_axi_edge_list_ch_32_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_32_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_32_RID,
    input wire                                           m_axi_edge_list_ch_32_RLAST,
    output wire                                          m_axi_edge_list_ch_32_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_32_RRESP,
    input wire                                           m_axi_edge_list_ch_32_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_32_WDATA,
    output wire                                          m_axi_edge_list_ch_32_WLAST,
    input wire                                           m_axi_edge_list_ch_32_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_32_WSTRB,
    output wire                                          m_axi_edge_list_ch_32_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_33_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_33_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_33_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_33_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_33_ARLEN,
    output wire                                          m_axi_edge_list_ch_33_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_33_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_33_ARQOS,
    input wire                                           m_axi_edge_list_ch_33_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_33_ARSIZE,
    output wire                                          m_axi_edge_list_ch_33_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_33_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_33_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_33_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_33_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_33_AWLEN,
    output wire                                          m_axi_edge_list_ch_33_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_33_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_33_AWQOS,
    input wire                                           m_axi_edge_list_ch_33_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_33_AWSIZE,
    output wire                                          m_axi_edge_list_ch_33_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_33_BID,
    output wire                                          m_axi_edge_list_ch_33_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_33_BRESP,
    input wire                                           m_axi_edge_list_ch_33_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_33_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_33_RID,
    input wire                                           m_axi_edge_list_ch_33_RLAST,
    output wire                                          m_axi_edge_list_ch_33_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_33_RRESP,
    input wire                                           m_axi_edge_list_ch_33_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_33_WDATA,
    output wire                                          m_axi_edge_list_ch_33_WLAST,
    input wire                                           m_axi_edge_list_ch_33_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_33_WSTRB,
    output wire                                          m_axi_edge_list_ch_33_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_34_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_34_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_34_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_34_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_34_ARLEN,
    output wire                                          m_axi_edge_list_ch_34_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_34_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_34_ARQOS,
    input wire                                           m_axi_edge_list_ch_34_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_34_ARSIZE,
    output wire                                          m_axi_edge_list_ch_34_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_34_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_34_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_34_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_34_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_34_AWLEN,
    output wire                                          m_axi_edge_list_ch_34_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_34_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_34_AWQOS,
    input wire                                           m_axi_edge_list_ch_34_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_34_AWSIZE,
    output wire                                          m_axi_edge_list_ch_34_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_34_BID,
    output wire                                          m_axi_edge_list_ch_34_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_34_BRESP,
    input wire                                           m_axi_edge_list_ch_34_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_34_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_34_RID,
    input wire                                           m_axi_edge_list_ch_34_RLAST,
    output wire                                          m_axi_edge_list_ch_34_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_34_RRESP,
    input wire                                           m_axi_edge_list_ch_34_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_34_WDATA,
    output wire                                          m_axi_edge_list_ch_34_WLAST,
    input wire                                           m_axi_edge_list_ch_34_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_34_WSTRB,
    output wire                                          m_axi_edge_list_ch_34_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_35_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_35_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_35_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_35_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_35_ARLEN,
    output wire                                          m_axi_edge_list_ch_35_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_35_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_35_ARQOS,
    input wire                                           m_axi_edge_list_ch_35_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_35_ARSIZE,
    output wire                                          m_axi_edge_list_ch_35_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_35_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_35_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_35_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_35_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_35_AWLEN,
    output wire                                          m_axi_edge_list_ch_35_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_35_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_35_AWQOS,
    input wire                                           m_axi_edge_list_ch_35_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_35_AWSIZE,
    output wire                                          m_axi_edge_list_ch_35_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_35_BID,
    output wire                                          m_axi_edge_list_ch_35_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_35_BRESP,
    input wire                                           m_axi_edge_list_ch_35_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_35_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_35_RID,
    input wire                                           m_axi_edge_list_ch_35_RLAST,
    output wire                                          m_axi_edge_list_ch_35_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_35_RRESP,
    input wire                                           m_axi_edge_list_ch_35_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_35_WDATA,
    output wire                                          m_axi_edge_list_ch_35_WLAST,
    input wire                                           m_axi_edge_list_ch_35_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_35_WSTRB,
    output wire                                          m_axi_edge_list_ch_35_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_36_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_36_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_36_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_36_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_36_ARLEN,
    output wire                                          m_axi_edge_list_ch_36_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_36_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_36_ARQOS,
    input wire                                           m_axi_edge_list_ch_36_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_36_ARSIZE,
    output wire                                          m_axi_edge_list_ch_36_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_36_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_36_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_36_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_36_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_36_AWLEN,
    output wire                                          m_axi_edge_list_ch_36_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_36_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_36_AWQOS,
    input wire                                           m_axi_edge_list_ch_36_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_36_AWSIZE,
    output wire                                          m_axi_edge_list_ch_36_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_36_BID,
    output wire                                          m_axi_edge_list_ch_36_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_36_BRESP,
    input wire                                           m_axi_edge_list_ch_36_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_36_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_36_RID,
    input wire                                           m_axi_edge_list_ch_36_RLAST,
    output wire                                          m_axi_edge_list_ch_36_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_36_RRESP,
    input wire                                           m_axi_edge_list_ch_36_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_36_WDATA,
    output wire                                          m_axi_edge_list_ch_36_WLAST,
    input wire                                           m_axi_edge_list_ch_36_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_36_WSTRB,
    output wire                                          m_axi_edge_list_ch_36_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_37_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_37_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_37_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_37_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_37_ARLEN,
    output wire                                          m_axi_edge_list_ch_37_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_37_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_37_ARQOS,
    input wire                                           m_axi_edge_list_ch_37_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_37_ARSIZE,
    output wire                                          m_axi_edge_list_ch_37_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_37_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_37_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_37_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_37_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_37_AWLEN,
    output wire                                          m_axi_edge_list_ch_37_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_37_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_37_AWQOS,
    input wire                                           m_axi_edge_list_ch_37_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_37_AWSIZE,
    output wire                                          m_axi_edge_list_ch_37_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_37_BID,
    output wire                                          m_axi_edge_list_ch_37_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_37_BRESP,
    input wire                                           m_axi_edge_list_ch_37_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_37_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_37_RID,
    input wire                                           m_axi_edge_list_ch_37_RLAST,
    output wire                                          m_axi_edge_list_ch_37_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_37_RRESP,
    input wire                                           m_axi_edge_list_ch_37_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_37_WDATA,
    output wire                                          m_axi_edge_list_ch_37_WLAST,
    input wire                                           m_axi_edge_list_ch_37_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_37_WSTRB,
    output wire                                          m_axi_edge_list_ch_37_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_38_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_38_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_38_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_38_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_38_ARLEN,
    output wire                                          m_axi_edge_list_ch_38_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_38_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_38_ARQOS,
    input wire                                           m_axi_edge_list_ch_38_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_38_ARSIZE,
    output wire                                          m_axi_edge_list_ch_38_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_38_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_38_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_38_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_38_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_38_AWLEN,
    output wire                                          m_axi_edge_list_ch_38_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_38_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_38_AWQOS,
    input wire                                           m_axi_edge_list_ch_38_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_38_AWSIZE,
    output wire                                          m_axi_edge_list_ch_38_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_38_BID,
    output wire                                          m_axi_edge_list_ch_38_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_38_BRESP,
    input wire                                           m_axi_edge_list_ch_38_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_38_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_38_RID,
    input wire                                           m_axi_edge_list_ch_38_RLAST,
    output wire                                          m_axi_edge_list_ch_38_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_38_RRESP,
    input wire                                           m_axi_edge_list_ch_38_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_38_WDATA,
    output wire                                          m_axi_edge_list_ch_38_WLAST,
    input wire                                           m_axi_edge_list_ch_38_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_38_WSTRB,
    output wire                                          m_axi_edge_list_ch_38_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_39_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_39_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_39_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_39_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_39_ARLEN,
    output wire                                          m_axi_edge_list_ch_39_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_39_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_39_ARQOS,
    input wire                                           m_axi_edge_list_ch_39_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_39_ARSIZE,
    output wire                                          m_axi_edge_list_ch_39_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_39_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_39_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_39_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_39_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_39_AWLEN,
    output wire                                          m_axi_edge_list_ch_39_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_39_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_39_AWQOS,
    input wire                                           m_axi_edge_list_ch_39_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_39_AWSIZE,
    output wire                                          m_axi_edge_list_ch_39_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_39_BID,
    output wire                                          m_axi_edge_list_ch_39_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_39_BRESP,
    input wire                                           m_axi_edge_list_ch_39_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_39_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_39_RID,
    input wire                                           m_axi_edge_list_ch_39_RLAST,
    output wire                                          m_axi_edge_list_ch_39_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_39_RRESP,
    input wire                                           m_axi_edge_list_ch_39_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_39_WDATA,
    output wire                                          m_axi_edge_list_ch_39_WLAST,
    input wire                                           m_axi_edge_list_ch_39_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_39_WSTRB,
    output wire                                          m_axi_edge_list_ch_39_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_40_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_40_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_40_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_40_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_40_ARLEN,
    output wire                                          m_axi_edge_list_ch_40_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_40_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_40_ARQOS,
    input wire                                           m_axi_edge_list_ch_40_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_40_ARSIZE,
    output wire                                          m_axi_edge_list_ch_40_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_40_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_40_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_40_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_40_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_40_AWLEN,
    output wire                                          m_axi_edge_list_ch_40_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_40_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_40_AWQOS,
    input wire                                           m_axi_edge_list_ch_40_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_40_AWSIZE,
    output wire                                          m_axi_edge_list_ch_40_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_40_BID,
    output wire                                          m_axi_edge_list_ch_40_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_40_BRESP,
    input wire                                           m_axi_edge_list_ch_40_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_40_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_40_RID,
    input wire                                           m_axi_edge_list_ch_40_RLAST,
    output wire                                          m_axi_edge_list_ch_40_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_40_RRESP,
    input wire                                           m_axi_edge_list_ch_40_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_40_WDATA,
    output wire                                          m_axi_edge_list_ch_40_WLAST,
    input wire                                           m_axi_edge_list_ch_40_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_40_WSTRB,
    output wire                                          m_axi_edge_list_ch_40_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_41_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_41_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_41_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_41_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_41_ARLEN,
    output wire                                          m_axi_edge_list_ch_41_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_41_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_41_ARQOS,
    input wire                                           m_axi_edge_list_ch_41_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_41_ARSIZE,
    output wire                                          m_axi_edge_list_ch_41_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_41_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_41_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_41_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_41_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_41_AWLEN,
    output wire                                          m_axi_edge_list_ch_41_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_41_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_41_AWQOS,
    input wire                                           m_axi_edge_list_ch_41_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_41_AWSIZE,
    output wire                                          m_axi_edge_list_ch_41_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_41_BID,
    output wire                                          m_axi_edge_list_ch_41_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_41_BRESP,
    input wire                                           m_axi_edge_list_ch_41_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_41_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_41_RID,
    input wire                                           m_axi_edge_list_ch_41_RLAST,
    output wire                                          m_axi_edge_list_ch_41_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_41_RRESP,
    input wire                                           m_axi_edge_list_ch_41_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_41_WDATA,
    output wire                                          m_axi_edge_list_ch_41_WLAST,
    input wire                                           m_axi_edge_list_ch_41_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_41_WSTRB,
    output wire                                          m_axi_edge_list_ch_41_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_42_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_42_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_42_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_42_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_42_ARLEN,
    output wire                                          m_axi_edge_list_ch_42_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_42_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_42_ARQOS,
    input wire                                           m_axi_edge_list_ch_42_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_42_ARSIZE,
    output wire                                          m_axi_edge_list_ch_42_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_42_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_42_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_42_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_42_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_42_AWLEN,
    output wire                                          m_axi_edge_list_ch_42_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_42_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_42_AWQOS,
    input wire                                           m_axi_edge_list_ch_42_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_42_AWSIZE,
    output wire                                          m_axi_edge_list_ch_42_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_42_BID,
    output wire                                          m_axi_edge_list_ch_42_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_42_BRESP,
    input wire                                           m_axi_edge_list_ch_42_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_42_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_42_RID,
    input wire                                           m_axi_edge_list_ch_42_RLAST,
    output wire                                          m_axi_edge_list_ch_42_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_42_RRESP,
    input wire                                           m_axi_edge_list_ch_42_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_42_WDATA,
    output wire                                          m_axi_edge_list_ch_42_WLAST,
    input wire                                           m_axi_edge_list_ch_42_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_42_WSTRB,
    output wire                                          m_axi_edge_list_ch_42_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_43_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_43_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_43_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_43_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_43_ARLEN,
    output wire                                          m_axi_edge_list_ch_43_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_43_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_43_ARQOS,
    input wire                                           m_axi_edge_list_ch_43_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_43_ARSIZE,
    output wire                                          m_axi_edge_list_ch_43_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_43_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_43_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_43_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_43_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_43_AWLEN,
    output wire                                          m_axi_edge_list_ch_43_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_43_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_43_AWQOS,
    input wire                                           m_axi_edge_list_ch_43_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_43_AWSIZE,
    output wire                                          m_axi_edge_list_ch_43_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_43_BID,
    output wire                                          m_axi_edge_list_ch_43_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_43_BRESP,
    input wire                                           m_axi_edge_list_ch_43_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_43_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_43_RID,
    input wire                                           m_axi_edge_list_ch_43_RLAST,
    output wire                                          m_axi_edge_list_ch_43_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_43_RRESP,
    input wire                                           m_axi_edge_list_ch_43_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_43_WDATA,
    output wire                                          m_axi_edge_list_ch_43_WLAST,
    input wire                                           m_axi_edge_list_ch_43_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_43_WSTRB,
    output wire                                          m_axi_edge_list_ch_43_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_44_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_44_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_44_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_44_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_44_ARLEN,
    output wire                                          m_axi_edge_list_ch_44_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_44_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_44_ARQOS,
    input wire                                           m_axi_edge_list_ch_44_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_44_ARSIZE,
    output wire                                          m_axi_edge_list_ch_44_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_44_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_44_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_44_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_44_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_44_AWLEN,
    output wire                                          m_axi_edge_list_ch_44_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_44_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_44_AWQOS,
    input wire                                           m_axi_edge_list_ch_44_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_44_AWSIZE,
    output wire                                          m_axi_edge_list_ch_44_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_44_BID,
    output wire                                          m_axi_edge_list_ch_44_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_44_BRESP,
    input wire                                           m_axi_edge_list_ch_44_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_44_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_44_RID,
    input wire                                           m_axi_edge_list_ch_44_RLAST,
    output wire                                          m_axi_edge_list_ch_44_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_44_RRESP,
    input wire                                           m_axi_edge_list_ch_44_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_44_WDATA,
    output wire                                          m_axi_edge_list_ch_44_WLAST,
    input wire                                           m_axi_edge_list_ch_44_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_44_WSTRB,
    output wire                                          m_axi_edge_list_ch_44_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_45_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_45_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_45_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_45_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_45_ARLEN,
    output wire                                          m_axi_edge_list_ch_45_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_45_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_45_ARQOS,
    input wire                                           m_axi_edge_list_ch_45_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_45_ARSIZE,
    output wire                                          m_axi_edge_list_ch_45_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_45_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_45_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_45_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_45_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_45_AWLEN,
    output wire                                          m_axi_edge_list_ch_45_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_45_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_45_AWQOS,
    input wire                                           m_axi_edge_list_ch_45_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_45_AWSIZE,
    output wire                                          m_axi_edge_list_ch_45_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_45_BID,
    output wire                                          m_axi_edge_list_ch_45_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_45_BRESP,
    input wire                                           m_axi_edge_list_ch_45_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_45_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_45_RID,
    input wire                                           m_axi_edge_list_ch_45_RLAST,
    output wire                                          m_axi_edge_list_ch_45_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_45_RRESP,
    input wire                                           m_axi_edge_list_ch_45_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_45_WDATA,
    output wire                                          m_axi_edge_list_ch_45_WLAST,
    input wire                                           m_axi_edge_list_ch_45_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_45_WSTRB,
    output wire                                          m_axi_edge_list_ch_45_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_46_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_46_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_46_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_46_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_46_ARLEN,
    output wire                                          m_axi_edge_list_ch_46_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_46_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_46_ARQOS,
    input wire                                           m_axi_edge_list_ch_46_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_46_ARSIZE,
    output wire                                          m_axi_edge_list_ch_46_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_46_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_46_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_46_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_46_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_46_AWLEN,
    output wire                                          m_axi_edge_list_ch_46_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_46_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_46_AWQOS,
    input wire                                           m_axi_edge_list_ch_46_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_46_AWSIZE,
    output wire                                          m_axi_edge_list_ch_46_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_46_BID,
    output wire                                          m_axi_edge_list_ch_46_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_46_BRESP,
    input wire                                           m_axi_edge_list_ch_46_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_46_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_46_RID,
    input wire                                           m_axi_edge_list_ch_46_RLAST,
    output wire                                          m_axi_edge_list_ch_46_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_46_RRESP,
    input wire                                           m_axi_edge_list_ch_46_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_46_WDATA,
    output wire                                          m_axi_edge_list_ch_46_WLAST,
    input wire                                           m_axi_edge_list_ch_46_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_46_WSTRB,
    output wire                                          m_axi_edge_list_ch_46_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_47_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_47_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_47_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_47_ARID,
    output wire [                                   7:0] m_axi_edge_list_ch_47_ARLEN,
    output wire                                          m_axi_edge_list_ch_47_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_47_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_47_ARQOS,
    input wire                                           m_axi_edge_list_ch_47_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_47_ARSIZE,
    output wire                                          m_axi_edge_list_ch_47_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ch_47_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ch_47_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ch_47_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ch_47_AWID,
    output wire [                                   7:0] m_axi_edge_list_ch_47_AWLEN,
    output wire                                          m_axi_edge_list_ch_47_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ch_47_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ch_47_AWQOS,
    input wire                                           m_axi_edge_list_ch_47_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ch_47_AWSIZE,
    output wire                                          m_axi_edge_list_ch_47_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ch_47_BID,
    output wire                                          m_axi_edge_list_ch_47_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_47_BRESP,
    input wire                                           m_axi_edge_list_ch_47_BVALID,
    input wire  [                                 255:0] m_axi_edge_list_ch_47_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ch_47_RID,
    input wire                                           m_axi_edge_list_ch_47_RLAST,
    output wire                                          m_axi_edge_list_ch_47_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ch_47_RRESP,
    input wire                                           m_axi_edge_list_ch_47_RVALID,
    output wire [                                 255:0] m_axi_edge_list_ch_47_WDATA,
    output wire                                          m_axi_edge_list_ch_47_WLAST,
    input wire                                           m_axi_edge_list_ch_47_WREADY,
    output wire [                                  31:0] m_axi_edge_list_ch_47_WSTRB,
    output wire                                          m_axi_edge_list_ch_47_WVALID,
    output wire [                                  63:0] m_axi_vec_X_ARADDR,
    output wire [                                   1:0] m_axi_vec_X_ARBURST,
    output wire [                                   3:0] m_axi_vec_X_ARCACHE,
    output wire [                                   0:0] m_axi_vec_X_ARID,
    output wire [                                   7:0] m_axi_vec_X_ARLEN,
    output wire                                          m_axi_vec_X_ARLOCK,
    output wire [                                   2:0] m_axi_vec_X_ARPROT,
    output wire [                                   3:0] m_axi_vec_X_ARQOS,
    input wire                                           m_axi_vec_X_ARREADY,
    output wire [                                   2:0] m_axi_vec_X_ARSIZE,
    output wire                                          m_axi_vec_X_ARVALID,
    output wire [                                  63:0] m_axi_vec_X_AWADDR,
    output wire [                                   1:0] m_axi_vec_X_AWBURST,
    output wire [                                   3:0] m_axi_vec_X_AWCACHE,
    output wire [                                   0:0] m_axi_vec_X_AWID,
    output wire [                                   7:0] m_axi_vec_X_AWLEN,
    output wire                                          m_axi_vec_X_AWLOCK,
    output wire [                                   2:0] m_axi_vec_X_AWPROT,
    output wire [                                   3:0] m_axi_vec_X_AWQOS,
    input wire                                           m_axi_vec_X_AWREADY,
    output wire [                                   2:0] m_axi_vec_X_AWSIZE,
    output wire                                          m_axi_vec_X_AWVALID,
    input wire  [                                   0:0] m_axi_vec_X_BID,
    output wire                                          m_axi_vec_X_BREADY,
    input wire  [                                   1:0] m_axi_vec_X_BRESP,
    input wire                                           m_axi_vec_X_BVALID,
    input wire  [                                 255:0] m_axi_vec_X_RDATA,
    input wire  [                                   0:0] m_axi_vec_X_RID,
    input wire                                           m_axi_vec_X_RLAST,
    output wire                                          m_axi_vec_X_RREADY,
    input wire  [                                   1:0] m_axi_vec_X_RRESP,
    input wire                                           m_axi_vec_X_RVALID,
    output wire [                                 255:0] m_axi_vec_X_WDATA,
    output wire                                          m_axi_vec_X_WLAST,
    input wire                                           m_axi_vec_X_WREADY,
    output wire [                                  31:0] m_axi_vec_X_WSTRB,
    output wire                                          m_axi_vec_X_WVALID,
    output wire [                                  63:0] m_axi_vec_Y_ARADDR,
    output wire [                                   1:0] m_axi_vec_Y_ARBURST,
    output wire [                                   3:0] m_axi_vec_Y_ARCACHE,
    output wire [                                   0:0] m_axi_vec_Y_ARID,
    output wire [                                   7:0] m_axi_vec_Y_ARLEN,
    output wire                                          m_axi_vec_Y_ARLOCK,
    output wire [                                   2:0] m_axi_vec_Y_ARPROT,
    output wire [                                   3:0] m_axi_vec_Y_ARQOS,
    input wire                                           m_axi_vec_Y_ARREADY,
    output wire [                                   2:0] m_axi_vec_Y_ARSIZE,
    output wire                                          m_axi_vec_Y_ARVALID,
    output wire [                                  63:0] m_axi_vec_Y_AWADDR,
    output wire [                                   1:0] m_axi_vec_Y_AWBURST,
    output wire [                                   3:0] m_axi_vec_Y_AWCACHE,
    output wire [                                   0:0] m_axi_vec_Y_AWID,
    output wire [                                   7:0] m_axi_vec_Y_AWLEN,
    output wire                                          m_axi_vec_Y_AWLOCK,
    output wire [                                   2:0] m_axi_vec_Y_AWPROT,
    output wire [                                   3:0] m_axi_vec_Y_AWQOS,
    input wire                                           m_axi_vec_Y_AWREADY,
    output wire [                                   2:0] m_axi_vec_Y_AWSIZE,
    output wire                                          m_axi_vec_Y_AWVALID,
    input wire  [                                   0:0] m_axi_vec_Y_BID,
    output wire                                          m_axi_vec_Y_BREADY,
    input wire  [                                   1:0] m_axi_vec_Y_BRESP,
    input wire                                           m_axi_vec_Y_BVALID,
    input wire  [                                 255:0] m_axi_vec_Y_RDATA,
    input wire  [                                   0:0] m_axi_vec_Y_RID,
    input wire                                           m_axi_vec_Y_RLAST,
    output wire                                          m_axi_vec_Y_RREADY,
    input wire  [                                   1:0] m_axi_vec_Y_RRESP,
    input wire                                           m_axi_vec_Y_RVALID,
    output wire [                                 255:0] m_axi_vec_Y_WDATA,
    output wire                                          m_axi_vec_Y_WLAST,
    input wire                                           m_axi_vec_Y_WREADY,
    output wire [                                  31:0] m_axi_vec_Y_WSTRB,
    output wire                                          m_axi_vec_Y_WVALID,
    output wire [                                  63:0] m_axi_edge_list_ptr_ARADDR,
    output wire [                                   1:0] m_axi_edge_list_ptr_ARBURST,
    output wire [                                   3:0] m_axi_edge_list_ptr_ARCACHE,
    output wire [                                   0:0] m_axi_edge_list_ptr_ARID,
    output wire [                                   7:0] m_axi_edge_list_ptr_ARLEN,
    output wire                                          m_axi_edge_list_ptr_ARLOCK,
    output wire [                                   2:0] m_axi_edge_list_ptr_ARPROT,
    output wire [                                   3:0] m_axi_edge_list_ptr_ARQOS,
    input wire                                           m_axi_edge_list_ptr_ARREADY,
    output wire [                                   2:0] m_axi_edge_list_ptr_ARSIZE,
    output wire                                          m_axi_edge_list_ptr_ARVALID,
    output wire [                                  63:0] m_axi_edge_list_ptr_AWADDR,
    output wire [                                   1:0] m_axi_edge_list_ptr_AWBURST,
    output wire [                                   3:0] m_axi_edge_list_ptr_AWCACHE,
    output wire [                                   0:0] m_axi_edge_list_ptr_AWID,
    output wire [                                   7:0] m_axi_edge_list_ptr_AWLEN,
    output wire                                          m_axi_edge_list_ptr_AWLOCK,
    output wire [                                   2:0] m_axi_edge_list_ptr_AWPROT,
    output wire [                                   3:0] m_axi_edge_list_ptr_AWQOS,
    input wire                                           m_axi_edge_list_ptr_AWREADY,
    output wire [                                   2:0] m_axi_edge_list_ptr_AWSIZE,
    output wire                                          m_axi_edge_list_ptr_AWVALID,
    input wire  [                                   0:0] m_axi_edge_list_ptr_BID,
    output wire                                          m_axi_edge_list_ptr_BREADY,
    input wire  [                                   1:0] m_axi_edge_list_ptr_BRESP,
    input wire                                           m_axi_edge_list_ptr_BVALID,
    input wire  [                                  31:0] m_axi_edge_list_ptr_RDATA,
    input wire  [                                   0:0] m_axi_edge_list_ptr_RID,
    input wire                                           m_axi_edge_list_ptr_RLAST,
    output wire                                          m_axi_edge_list_ptr_RREADY,
    input wire  [                                   1:0] m_axi_edge_list_ptr_RRESP,
    input wire                                           m_axi_edge_list_ptr_RVALID,
    output wire [                                  31:0] m_axi_edge_list_ptr_WDATA,
    output wire                                          m_axi_edge_list_ptr_WLAST,
    input wire                                           m_axi_edge_list_ptr_WREADY,
    output wire [                                   3:0] m_axi_edge_list_ptr_WSTRB,
    output wire                                          m_axi_edge_list_ptr_WVALID,
    output wire [                                  63:0] m_axi_vec_Y_out_ARADDR,
    output wire [                                   1:0] m_axi_vec_Y_out_ARBURST,
    output wire [                                   3:0] m_axi_vec_Y_out_ARCACHE,
    output wire [                                   0:0] m_axi_vec_Y_out_ARID,
    output wire [                                   7:0] m_axi_vec_Y_out_ARLEN,
    output wire                                          m_axi_vec_Y_out_ARLOCK,
    output wire [                                   2:0] m_axi_vec_Y_out_ARPROT,
    output wire [                                   3:0] m_axi_vec_Y_out_ARQOS,
    input wire                                           m_axi_vec_Y_out_ARREADY,
    output wire [                                   2:0] m_axi_vec_Y_out_ARSIZE,
    output wire                                          m_axi_vec_Y_out_ARVALID,
    output wire [                                  63:0] m_axi_vec_Y_out_AWADDR,
    output wire [                                   1:0] m_axi_vec_Y_out_AWBURST,
    output wire [                                   3:0] m_axi_vec_Y_out_AWCACHE,
    output wire [                                   0:0] m_axi_vec_Y_out_AWID,
    output wire [                                   7:0] m_axi_vec_Y_out_AWLEN,
    output wire                                          m_axi_vec_Y_out_AWLOCK,
    output wire [                                   2:0] m_axi_vec_Y_out_AWPROT,
    output wire [                                   3:0] m_axi_vec_Y_out_AWQOS,
    input wire                                           m_axi_vec_Y_out_AWREADY,
    output wire [                                   2:0] m_axi_vec_Y_out_AWSIZE,
    output wire                                          m_axi_vec_Y_out_AWVALID,
    input wire  [                                   0:0] m_axi_vec_Y_out_BID,
    output wire                                          m_axi_vec_Y_out_BREADY,
    input wire  [                                   1:0] m_axi_vec_Y_out_BRESP,
    input wire                                           m_axi_vec_Y_out_BVALID,
    input wire  [                                 255:0] m_axi_vec_Y_out_RDATA,
    input wire  [                                   0:0] m_axi_vec_Y_out_RID,
    input wire                                           m_axi_vec_Y_out_RLAST,
    output wire                                          m_axi_vec_Y_out_RREADY,
    input wire  [                                   1:0] m_axi_vec_Y_out_RRESP,
    input wire                                           m_axi_vec_Y_out_RVALID,
    output wire [                                 255:0] m_axi_vec_Y_out_WDATA,
    output wire                                          m_axi_vec_Y_out_WLAST,
    input wire                                           m_axi_vec_Y_out_WREADY,
    output wire [                                  31:0] m_axi_vec_Y_out_WSTRB,
    output wire                                          m_axi_vec_Y_out_WVALID,
    output wire                                          control_s_axi_U_ACLK,
    output wire                                          control_s_axi_U_ACLK_EN,
    output wire [    (C_S_AXI_CONTROL_ADDR_WIDTH - 1):0] control_s_axi_U_ARADDR,
    output wire                                          control_s_axi_U_ARESET,
    input wire                                           control_s_axi_U_ARREADY,
    output wire                                          control_s_axi_U_ARVALID,
    output wire [    (C_S_AXI_CONTROL_ADDR_WIDTH - 1):0] control_s_axi_U_AWADDR,
    input wire                                           control_s_axi_U_AWREADY,
    output wire                                          control_s_axi_U_AWVALID,
    output wire                                          control_s_axi_U_BREADY,
    input wire  [                                   1:0] control_s_axi_U_BRESP,
    input wire                                           control_s_axi_U_BVALID,
    input wire  [                                  31:0] control_s_axi_U_K,
    input wire  [                                  31:0] control_s_axi_U_M,
    input wire  [                                  31:0] control_s_axi_U_NUM_A_LEN,
    input wire  [                                  31:0] control_s_axi_U_NUM_ITE,
    input wire  [                                  31:0] control_s_axi_U_P_N,
    input wire  [    (C_S_AXI_CONTROL_DATA_WIDTH - 1):0] control_s_axi_U_RDATA,
    output wire                                          control_s_axi_U_RREADY,
    input wire  [                                   1:0] control_s_axi_U_RRESP,
    input wire                                           control_s_axi_U_RVALID,
    output wire [    (C_S_AXI_CONTROL_DATA_WIDTH - 1):0] control_s_axi_U_WDATA,
    input wire                                           control_s_axi_U_WREADY,
    output wire [(C_S_AXI_CONTROL_DATA_WIDTH / 8 - 1):0] control_s_axi_U_WSTRB,
    output wire                                          control_s_axi_U_WVALID,
    input wire  [                                  31:0] control_s_axi_U_alpha_u,
    output wire                                          control_s_axi_U_ap_done,
    output wire                                          control_s_axi_U_ap_idle,
    output wire                                          control_s_axi_U_ap_ready,
    input wire                                           control_s_axi_U_ap_start,
    input wire  [                                  31:0] control_s_axi_U_beta_u,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_0,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_1,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_10,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_11,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_12,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_13,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_14,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_15,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_16,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_17,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_18,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_19,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_2,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_20,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_21,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_22,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_23,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_24,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_25,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_26,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_27,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_28,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_29,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_3,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_30,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_31,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_32,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_33,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_34,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_35,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_36,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_37,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_38,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_39,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_4,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_40,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_41,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_42,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_43,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_44,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_45,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_46,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_47,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_5,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_6,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_7,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_8,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ch_9,
    input wire  [                                  63:0] control_s_axi_U_edge_list_ptr,
    input wire                                           control_s_axi_U_interrupt,
    input wire  [                                  63:0] control_s_axi_U_vec_X,
    input wire  [                                  63:0] control_s_axi_U_vec_Y,
    input wire  [                                  63:0] control_s_axi_U_vec_Y_out,
    output wire                                          PE_inst_0_clk,
    output wire [                                  32:0] PE_inst_0_if_din,
    input wire  [                                  32:0] PE_inst_0_if_dout,
    input wire                                           PE_inst_0_if_empty_n,
    input wire                                           PE_inst_0_if_full_n,
    output wire                                          PE_inst_0_if_read,
    output wire                                          PE_inst_0_if_read_ce,
    output wire                                          PE_inst_0_if_write,
    output wire                                          PE_inst_0_if_write_ce,
    output wire                                          PE_inst_0_reset,
    output wire                                          PE_inst_10_clk,
    output wire [                                  32:0] PE_inst_10_if_din,
    input wire  [                                  32:0] PE_inst_10_if_dout,
    input wire                                           PE_inst_10_if_empty_n,
    input wire                                           PE_inst_10_if_full_n,
    output wire                                          PE_inst_10_if_read,
    output wire                                          PE_inst_10_if_read_ce,
    output wire                                          PE_inst_10_if_write,
    output wire                                          PE_inst_10_if_write_ce,
    output wire                                          PE_inst_10_reset,
    output wire                                          PE_inst_11_clk,
    output wire [                                  32:0] PE_inst_11_if_din,
    input wire  [                                  32:0] PE_inst_11_if_dout,
    input wire                                           PE_inst_11_if_empty_n,
    input wire                                           PE_inst_11_if_full_n,
    output wire                                          PE_inst_11_if_read,
    output wire                                          PE_inst_11_if_read_ce,
    output wire                                          PE_inst_11_if_write,
    output wire                                          PE_inst_11_if_write_ce,
    output wire                                          PE_inst_11_reset,
    output wire                                          PE_inst_12_clk,
    output wire [                                  32:0] PE_inst_12_if_din,
    input wire  [                                  32:0] PE_inst_12_if_dout,
    input wire                                           PE_inst_12_if_empty_n,
    input wire                                           PE_inst_12_if_full_n,
    output wire                                          PE_inst_12_if_read,
    output wire                                          PE_inst_12_if_read_ce,
    output wire                                          PE_inst_12_if_write,
    output wire                                          PE_inst_12_if_write_ce,
    output wire                                          PE_inst_12_reset,
    output wire                                          PE_inst_13_clk,
    output wire [                                  32:0] PE_inst_13_if_din,
    input wire  [                                  32:0] PE_inst_13_if_dout,
    input wire                                           PE_inst_13_if_empty_n,
    input wire                                           PE_inst_13_if_full_n,
    output wire                                          PE_inst_13_if_read,
    output wire                                          PE_inst_13_if_read_ce,
    output wire                                          PE_inst_13_if_write,
    output wire                                          PE_inst_13_if_write_ce,
    output wire                                          PE_inst_13_reset,
    output wire                                          PE_inst_14_clk,
    output wire [                                  32:0] PE_inst_14_if_din,
    input wire  [                                  32:0] PE_inst_14_if_dout,
    input wire                                           PE_inst_14_if_empty_n,
    input wire                                           PE_inst_14_if_full_n,
    output wire                                          PE_inst_14_if_read,
    output wire                                          PE_inst_14_if_read_ce,
    output wire                                          PE_inst_14_if_write,
    output wire                                          PE_inst_14_if_write_ce,
    output wire                                          PE_inst_14_reset,
    output wire                                          PE_inst_15_clk,
    output wire [                                  32:0] PE_inst_15_if_din,
    input wire  [                                  32:0] PE_inst_15_if_dout,
    input wire                                           PE_inst_15_if_empty_n,
    input wire                                           PE_inst_15_if_full_n,
    output wire                                          PE_inst_15_if_read,
    output wire                                          PE_inst_15_if_read_ce,
    output wire                                          PE_inst_15_if_write,
    output wire                                          PE_inst_15_if_write_ce,
    output wire                                          PE_inst_15_reset,
    output wire                                          PE_inst_16_clk,
    output wire [                                  32:0] PE_inst_16_if_din,
    input wire  [                                  32:0] PE_inst_16_if_dout,
    input wire                                           PE_inst_16_if_empty_n,
    input wire                                           PE_inst_16_if_full_n,
    output wire                                          PE_inst_16_if_read,
    output wire                                          PE_inst_16_if_read_ce,
    output wire                                          PE_inst_16_if_write,
    output wire                                          PE_inst_16_if_write_ce,
    output wire                                          PE_inst_16_reset,
    output wire                                          PE_inst_17_clk,
    output wire [                                  32:0] PE_inst_17_if_din,
    input wire  [                                  32:0] PE_inst_17_if_dout,
    input wire                                           PE_inst_17_if_empty_n,
    input wire                                           PE_inst_17_if_full_n,
    output wire                                          PE_inst_17_if_read,
    output wire                                          PE_inst_17_if_read_ce,
    output wire                                          PE_inst_17_if_write,
    output wire                                          PE_inst_17_if_write_ce,
    output wire                                          PE_inst_17_reset,
    output wire                                          PE_inst_18_clk,
    output wire [                                  32:0] PE_inst_18_if_din,
    input wire  [                                  32:0] PE_inst_18_if_dout,
    input wire                                           PE_inst_18_if_empty_n,
    input wire                                           PE_inst_18_if_full_n,
    output wire                                          PE_inst_18_if_read,
    output wire                                          PE_inst_18_if_read_ce,
    output wire                                          PE_inst_18_if_write,
    output wire                                          PE_inst_18_if_write_ce,
    output wire                                          PE_inst_18_reset,
    output wire                                          PE_inst_19_clk,
    output wire [                                  32:0] PE_inst_19_if_din,
    input wire  [                                  32:0] PE_inst_19_if_dout,
    input wire                                           PE_inst_19_if_empty_n,
    input wire                                           PE_inst_19_if_full_n,
    output wire                                          PE_inst_19_if_read,
    output wire                                          PE_inst_19_if_read_ce,
    output wire                                          PE_inst_19_if_write,
    output wire                                          PE_inst_19_if_write_ce,
    output wire                                          PE_inst_19_reset,
    output wire                                          PE_inst_1_clk,
    output wire [                                  32:0] PE_inst_1_if_din,
    input wire  [                                  32:0] PE_inst_1_if_dout,
    input wire                                           PE_inst_1_if_empty_n,
    input wire                                           PE_inst_1_if_full_n,
    output wire                                          PE_inst_1_if_read,
    output wire                                          PE_inst_1_if_read_ce,
    output wire                                          PE_inst_1_if_write,
    output wire                                          PE_inst_1_if_write_ce,
    output wire                                          PE_inst_1_reset,
    output wire                                          PE_inst_20_clk,
    output wire [                                  32:0] PE_inst_20_if_din,
    input wire  [                                  32:0] PE_inst_20_if_dout,
    input wire                                           PE_inst_20_if_empty_n,
    input wire                                           PE_inst_20_if_full_n,
    output wire                                          PE_inst_20_if_read,
    output wire                                          PE_inst_20_if_read_ce,
    output wire                                          PE_inst_20_if_write,
    output wire                                          PE_inst_20_if_write_ce,
    output wire                                          PE_inst_20_reset,
    output wire                                          PE_inst_21_clk,
    output wire [                                  32:0] PE_inst_21_if_din,
    input wire  [                                  32:0] PE_inst_21_if_dout,
    input wire                                           PE_inst_21_if_empty_n,
    input wire                                           PE_inst_21_if_full_n,
    output wire                                          PE_inst_21_if_read,
    output wire                                          PE_inst_21_if_read_ce,
    output wire                                          PE_inst_21_if_write,
    output wire                                          PE_inst_21_if_write_ce,
    output wire                                          PE_inst_21_reset,
    output wire                                          PE_inst_22_clk,
    output wire [                                  32:0] PE_inst_22_if_din,
    input wire  [                                  32:0] PE_inst_22_if_dout,
    input wire                                           PE_inst_22_if_empty_n,
    input wire                                           PE_inst_22_if_full_n,
    output wire                                          PE_inst_22_if_read,
    output wire                                          PE_inst_22_if_read_ce,
    output wire                                          PE_inst_22_if_write,
    output wire                                          PE_inst_22_if_write_ce,
    output wire                                          PE_inst_22_reset,
    output wire                                          PE_inst_23_clk,
    output wire [                                  32:0] PE_inst_23_if_din,
    input wire  [                                  32:0] PE_inst_23_if_dout,
    input wire                                           PE_inst_23_if_empty_n,
    input wire                                           PE_inst_23_if_full_n,
    output wire                                          PE_inst_23_if_read,
    output wire                                          PE_inst_23_if_read_ce,
    output wire                                          PE_inst_23_if_write,
    output wire                                          PE_inst_23_if_write_ce,
    output wire                                          PE_inst_23_reset,
    output wire                                          PE_inst_24_clk,
    output wire [                                  32:0] PE_inst_24_if_din,
    input wire  [                                  32:0] PE_inst_24_if_dout,
    input wire                                           PE_inst_24_if_empty_n,
    input wire                                           PE_inst_24_if_full_n,
    output wire                                          PE_inst_24_if_read,
    output wire                                          PE_inst_24_if_read_ce,
    output wire                                          PE_inst_24_if_write,
    output wire                                          PE_inst_24_if_write_ce,
    output wire                                          PE_inst_24_reset,
    output wire                                          PE_inst_25_clk,
    output wire [                                  32:0] PE_inst_25_if_din,
    input wire  [                                  32:0] PE_inst_25_if_dout,
    input wire                                           PE_inst_25_if_empty_n,
    input wire                                           PE_inst_25_if_full_n,
    output wire                                          PE_inst_25_if_read,
    output wire                                          PE_inst_25_if_read_ce,
    output wire                                          PE_inst_25_if_write,
    output wire                                          PE_inst_25_if_write_ce,
    output wire                                          PE_inst_25_reset,
    output wire                                          PE_inst_26_clk,
    output wire [                                  32:0] PE_inst_26_if_din,
    input wire  [                                  32:0] PE_inst_26_if_dout,
    input wire                                           PE_inst_26_if_empty_n,
    input wire                                           PE_inst_26_if_full_n,
    output wire                                          PE_inst_26_if_read,
    output wire                                          PE_inst_26_if_read_ce,
    output wire                                          PE_inst_26_if_write,
    output wire                                          PE_inst_26_if_write_ce,
    output wire                                          PE_inst_26_reset,
    output wire                                          PE_inst_27_clk,
    output wire [                                  32:0] PE_inst_27_if_din,
    input wire  [                                  32:0] PE_inst_27_if_dout,
    input wire                                           PE_inst_27_if_empty_n,
    input wire                                           PE_inst_27_if_full_n,
    output wire                                          PE_inst_27_if_read,
    output wire                                          PE_inst_27_if_read_ce,
    output wire                                          PE_inst_27_if_write,
    output wire                                          PE_inst_27_if_write_ce,
    output wire                                          PE_inst_27_reset,
    output wire                                          PE_inst_28_clk,
    output wire [                                  32:0] PE_inst_28_if_din,
    input wire  [                                  32:0] PE_inst_28_if_dout,
    input wire                                           PE_inst_28_if_empty_n,
    input wire                                           PE_inst_28_if_full_n,
    output wire                                          PE_inst_28_if_read,
    output wire                                          PE_inst_28_if_read_ce,
    output wire                                          PE_inst_28_if_write,
    output wire                                          PE_inst_28_if_write_ce,
    output wire                                          PE_inst_28_reset,
    output wire                                          PE_inst_29_clk,
    output wire [                                  32:0] PE_inst_29_if_din,
    input wire  [                                  32:0] PE_inst_29_if_dout,
    input wire                                           PE_inst_29_if_empty_n,
    input wire                                           PE_inst_29_if_full_n,
    output wire                                          PE_inst_29_if_read,
    output wire                                          PE_inst_29_if_read_ce,
    output wire                                          PE_inst_29_if_write,
    output wire                                          PE_inst_29_if_write_ce,
    output wire                                          PE_inst_29_reset,
    output wire                                          PE_inst_2_clk,
    output wire [                                  32:0] PE_inst_2_if_din,
    input wire  [                                  32:0] PE_inst_2_if_dout,
    input wire                                           PE_inst_2_if_empty_n,
    input wire                                           PE_inst_2_if_full_n,
    output wire                                          PE_inst_2_if_read,
    output wire                                          PE_inst_2_if_read_ce,
    output wire                                          PE_inst_2_if_write,
    output wire                                          PE_inst_2_if_write_ce,
    output wire                                          PE_inst_2_reset,
    output wire                                          PE_inst_30_clk,
    output wire [                                  32:0] PE_inst_30_if_din,
    input wire  [                                  32:0] PE_inst_30_if_dout,
    input wire                                           PE_inst_30_if_empty_n,
    input wire                                           PE_inst_30_if_full_n,
    output wire                                          PE_inst_30_if_read,
    output wire                                          PE_inst_30_if_read_ce,
    output wire                                          PE_inst_30_if_write,
    output wire                                          PE_inst_30_if_write_ce,
    output wire                                          PE_inst_30_reset,
    output wire                                          PE_inst_31_clk,
    output wire [                                  32:0] PE_inst_31_if_din,
    input wire  [                                  32:0] PE_inst_31_if_dout,
    input wire                                           PE_inst_31_if_empty_n,
    input wire                                           PE_inst_31_if_full_n,
    output wire                                          PE_inst_31_if_read,
    output wire                                          PE_inst_31_if_read_ce,
    output wire                                          PE_inst_31_if_write,
    output wire                                          PE_inst_31_if_write_ce,
    output wire                                          PE_inst_31_reset,
    output wire                                          PE_inst_32_clk,
    output wire [                                  32:0] PE_inst_32_if_din,
    input wire  [                                  32:0] PE_inst_32_if_dout,
    input wire                                           PE_inst_32_if_empty_n,
    input wire                                           PE_inst_32_if_full_n,
    output wire                                          PE_inst_32_if_read,
    output wire                                          PE_inst_32_if_read_ce,
    output wire                                          PE_inst_32_if_write,
    output wire                                          PE_inst_32_if_write_ce,
    output wire                                          PE_inst_32_reset,
    output wire                                          PE_inst_33_clk,
    output wire [                                  32:0] PE_inst_33_if_din,
    input wire  [                                  32:0] PE_inst_33_if_dout,
    input wire                                           PE_inst_33_if_empty_n,
    input wire                                           PE_inst_33_if_full_n,
    output wire                                          PE_inst_33_if_read,
    output wire                                          PE_inst_33_if_read_ce,
    output wire                                          PE_inst_33_if_write,
    output wire                                          PE_inst_33_if_write_ce,
    output wire                                          PE_inst_33_reset,
    output wire                                          PE_inst_34_clk,
    output wire [                                  32:0] PE_inst_34_if_din,
    input wire  [                                  32:0] PE_inst_34_if_dout,
    input wire                                           PE_inst_34_if_empty_n,
    input wire                                           PE_inst_34_if_full_n,
    output wire                                          PE_inst_34_if_read,
    output wire                                          PE_inst_34_if_read_ce,
    output wire                                          PE_inst_34_if_write,
    output wire                                          PE_inst_34_if_write_ce,
    output wire                                          PE_inst_34_reset,
    output wire                                          PE_inst_35_clk,
    output wire [                                  32:0] PE_inst_35_if_din,
    input wire  [                                  32:0] PE_inst_35_if_dout,
    input wire                                           PE_inst_35_if_empty_n,
    input wire                                           PE_inst_35_if_full_n,
    output wire                                          PE_inst_35_if_read,
    output wire                                          PE_inst_35_if_read_ce,
    output wire                                          PE_inst_35_if_write,
    output wire                                          PE_inst_35_if_write_ce,
    output wire                                          PE_inst_35_reset,
    output wire                                          PE_inst_36_clk,
    output wire [                                  32:0] PE_inst_36_if_din,
    input wire  [                                  32:0] PE_inst_36_if_dout,
    input wire                                           PE_inst_36_if_empty_n,
    input wire                                           PE_inst_36_if_full_n,
    output wire                                          PE_inst_36_if_read,
    output wire                                          PE_inst_36_if_read_ce,
    output wire                                          PE_inst_36_if_write,
    output wire                                          PE_inst_36_if_write_ce,
    output wire                                          PE_inst_36_reset,
    output wire                                          PE_inst_37_clk,
    output wire [                                  32:0] PE_inst_37_if_din,
    input wire  [                                  32:0] PE_inst_37_if_dout,
    input wire                                           PE_inst_37_if_empty_n,
    input wire                                           PE_inst_37_if_full_n,
    output wire                                          PE_inst_37_if_read,
    output wire                                          PE_inst_37_if_read_ce,
    output wire                                          PE_inst_37_if_write,
    output wire                                          PE_inst_37_if_write_ce,
    output wire                                          PE_inst_37_reset,
    output wire                                          PE_inst_38_clk,
    output wire [                                  32:0] PE_inst_38_if_din,
    input wire  [                                  32:0] PE_inst_38_if_dout,
    input wire                                           PE_inst_38_if_empty_n,
    input wire                                           PE_inst_38_if_full_n,
    output wire                                          PE_inst_38_if_read,
    output wire                                          PE_inst_38_if_read_ce,
    output wire                                          PE_inst_38_if_write,
    output wire                                          PE_inst_38_if_write_ce,
    output wire                                          PE_inst_38_reset,
    output wire                                          PE_inst_39_clk,
    output wire [                                  32:0] PE_inst_39_if_din,
    input wire  [                                  32:0] PE_inst_39_if_dout,
    input wire                                           PE_inst_39_if_empty_n,
    input wire                                           PE_inst_39_if_full_n,
    output wire                                          PE_inst_39_if_read,
    output wire                                          PE_inst_39_if_read_ce,
    output wire                                          PE_inst_39_if_write,
    output wire                                          PE_inst_39_if_write_ce,
    output wire                                          PE_inst_39_reset,
    output wire                                          PE_inst_3_clk,
    output wire [                                  32:0] PE_inst_3_if_din,
    input wire  [                                  32:0] PE_inst_3_if_dout,
    input wire                                           PE_inst_3_if_empty_n,
    input wire                                           PE_inst_3_if_full_n,
    output wire                                          PE_inst_3_if_read,
    output wire                                          PE_inst_3_if_read_ce,
    output wire                                          PE_inst_3_if_write,
    output wire                                          PE_inst_3_if_write_ce,
    output wire                                          PE_inst_3_reset,
    output wire                                          PE_inst_40_clk,
    output wire [                                  32:0] PE_inst_40_if_din,
    input wire  [                                  32:0] PE_inst_40_if_dout,
    input wire                                           PE_inst_40_if_empty_n,
    input wire                                           PE_inst_40_if_full_n,
    output wire                                          PE_inst_40_if_read,
    output wire                                          PE_inst_40_if_read_ce,
    output wire                                          PE_inst_40_if_write,
    output wire                                          PE_inst_40_if_write_ce,
    output wire                                          PE_inst_40_reset,
    output wire                                          PE_inst_41_clk,
    output wire [                                  32:0] PE_inst_41_if_din,
    input wire  [                                  32:0] PE_inst_41_if_dout,
    input wire                                           PE_inst_41_if_empty_n,
    input wire                                           PE_inst_41_if_full_n,
    output wire                                          PE_inst_41_if_read,
    output wire                                          PE_inst_41_if_read_ce,
    output wire                                          PE_inst_41_if_write,
    output wire                                          PE_inst_41_if_write_ce,
    output wire                                          PE_inst_41_reset,
    output wire                                          PE_inst_42_clk,
    output wire [                                  32:0] PE_inst_42_if_din,
    input wire  [                                  32:0] PE_inst_42_if_dout,
    input wire                                           PE_inst_42_if_empty_n,
    input wire                                           PE_inst_42_if_full_n,
    output wire                                          PE_inst_42_if_read,
    output wire                                          PE_inst_42_if_read_ce,
    output wire                                          PE_inst_42_if_write,
    output wire                                          PE_inst_42_if_write_ce,
    output wire                                          PE_inst_42_reset,
    output wire                                          PE_inst_43_clk,
    output wire [                                  32:0] PE_inst_43_if_din,
    input wire  [                                  32:0] PE_inst_43_if_dout,
    input wire                                           PE_inst_43_if_empty_n,
    input wire                                           PE_inst_43_if_full_n,
    output wire                                          PE_inst_43_if_read,
    output wire                                          PE_inst_43_if_read_ce,
    output wire                                          PE_inst_43_if_write,
    output wire                                          PE_inst_43_if_write_ce,
    output wire                                          PE_inst_43_reset,
    output wire                                          PE_inst_44_clk,
    output wire [                                  32:0] PE_inst_44_if_din,
    input wire  [                                  32:0] PE_inst_44_if_dout,
    input wire                                           PE_inst_44_if_empty_n,
    input wire                                           PE_inst_44_if_full_n,
    output wire                                          PE_inst_44_if_read,
    output wire                                          PE_inst_44_if_read_ce,
    output wire                                          PE_inst_44_if_write,
    output wire                                          PE_inst_44_if_write_ce,
    output wire                                          PE_inst_44_reset,
    output wire                                          PE_inst_45_clk,
    output wire [                                  32:0] PE_inst_45_if_din,
    input wire  [                                  32:0] PE_inst_45_if_dout,
    input wire                                           PE_inst_45_if_empty_n,
    input wire                                           PE_inst_45_if_full_n,
    output wire                                          PE_inst_45_if_read,
    output wire                                          PE_inst_45_if_read_ce,
    output wire                                          PE_inst_45_if_write,
    output wire                                          PE_inst_45_if_write_ce,
    output wire                                          PE_inst_45_reset,
    output wire                                          PE_inst_46_clk,
    output wire [                                  32:0] PE_inst_46_if_din,
    input wire  [                                  32:0] PE_inst_46_if_dout,
    input wire                                           PE_inst_46_if_empty_n,
    input wire                                           PE_inst_46_if_full_n,
    output wire                                          PE_inst_46_if_read,
    output wire                                          PE_inst_46_if_read_ce,
    output wire                                          PE_inst_46_if_write,
    output wire                                          PE_inst_46_if_write_ce,
    output wire                                          PE_inst_46_reset,
    output wire                                          PE_inst_47_clk,
    output wire [                                  32:0] PE_inst_47_if_din,
    input wire  [                                  32:0] PE_inst_47_if_dout,
    input wire                                           PE_inst_47_if_empty_n,
    input wire                                           PE_inst_47_if_full_n,
    output wire                                          PE_inst_47_if_read,
    output wire                                          PE_inst_47_if_read_ce,
    output wire                                          PE_inst_47_if_write,
    output wire                                          PE_inst_47_if_write_ce,
    output wire                                          PE_inst_47_reset,
    output wire                                          PE_inst_48_clk,
    output wire [                                  32:0] PE_inst_48_if_din,
    input wire  [                                  32:0] PE_inst_48_if_dout,
    input wire                                           PE_inst_48_if_empty_n,
    input wire                                           PE_inst_48_if_full_n,
    output wire                                          PE_inst_48_if_read,
    output wire                                          PE_inst_48_if_read_ce,
    output wire                                          PE_inst_48_if_write,
    output wire                                          PE_inst_48_if_write_ce,
    output wire                                          PE_inst_48_reset,
    output wire                                          PE_inst_4_clk,
    output wire [                                  32:0] PE_inst_4_if_din,
    input wire  [                                  32:0] PE_inst_4_if_dout,
    input wire                                           PE_inst_4_if_empty_n,
    input wire                                           PE_inst_4_if_full_n,
    output wire                                          PE_inst_4_if_read,
    output wire                                          PE_inst_4_if_read_ce,
    output wire                                          PE_inst_4_if_write,
    output wire                                          PE_inst_4_if_write_ce,
    output wire                                          PE_inst_4_reset,
    output wire                                          PE_inst_5_clk,
    output wire [                                  32:0] PE_inst_5_if_din,
    input wire  [                                  32:0] PE_inst_5_if_dout,
    input wire                                           PE_inst_5_if_empty_n,
    input wire                                           PE_inst_5_if_full_n,
    output wire                                          PE_inst_5_if_read,
    output wire                                          PE_inst_5_if_read_ce,
    output wire                                          PE_inst_5_if_write,
    output wire                                          PE_inst_5_if_write_ce,
    output wire                                          PE_inst_5_reset,
    output wire                                          PE_inst_6_clk,
    output wire [                                  32:0] PE_inst_6_if_din,
    input wire  [                                  32:0] PE_inst_6_if_dout,
    input wire                                           PE_inst_6_if_empty_n,
    input wire                                           PE_inst_6_if_full_n,
    output wire                                          PE_inst_6_if_read,
    output wire                                          PE_inst_6_if_read_ce,
    output wire                                          PE_inst_6_if_write,
    output wire                                          PE_inst_6_if_write_ce,
    output wire                                          PE_inst_6_reset,
    output wire                                          PE_inst_7_clk,
    output wire [                                  32:0] PE_inst_7_if_din,
    input wire  [                                  32:0] PE_inst_7_if_dout,
    input wire                                           PE_inst_7_if_empty_n,
    input wire                                           PE_inst_7_if_full_n,
    output wire                                          PE_inst_7_if_read,
    output wire                                          PE_inst_7_if_read_ce,
    output wire                                          PE_inst_7_if_write,
    output wire                                          PE_inst_7_if_write_ce,
    output wire                                          PE_inst_7_reset,
    output wire                                          PE_inst_8_clk,
    output wire [                                  32:0] PE_inst_8_if_din,
    input wire  [                                  32:0] PE_inst_8_if_dout,
    input wire                                           PE_inst_8_if_empty_n,
    input wire                                           PE_inst_8_if_full_n,
    output wire                                          PE_inst_8_if_read,
    output wire                                          PE_inst_8_if_read_ce,
    output wire                                          PE_inst_8_if_write,
    output wire                                          PE_inst_8_if_write_ce,
    output wire                                          PE_inst_8_reset,
    output wire                                          PE_inst_9_clk,
    output wire [                                  32:0] PE_inst_9_if_din,
    input wire  [                                  32:0] PE_inst_9_if_dout,
    input wire                                           PE_inst_9_if_empty_n,
    input wire                                           PE_inst_9_if_full_n,
    output wire                                          PE_inst_9_if_read,
    output wire                                          PE_inst_9_if_read_ce,
    output wire                                          PE_inst_9_if_write,
    output wire                                          PE_inst_9_if_write_ce,
    output wire                                          PE_inst_9_reset,
    output wire                                          Yvec_inst_0_clk,
    output wire [                                  32:0] Yvec_inst_0_if_din,
    input wire  [                                  32:0] Yvec_inst_0_if_dout,
    input wire                                           Yvec_inst_0_if_empty_n,
    input wire                                           Yvec_inst_0_if_full_n,
    output wire                                          Yvec_inst_0_if_read,
    output wire                                          Yvec_inst_0_if_read_ce,
    output wire                                          Yvec_inst_0_if_write,
    output wire                                          Yvec_inst_0_if_write_ce,
    output wire                                          Yvec_inst_0_reset,
    output wire                                          Yvec_inst_10_clk,
    output wire [                                  32:0] Yvec_inst_10_if_din,
    input wire  [                                  32:0] Yvec_inst_10_if_dout,
    input wire                                           Yvec_inst_10_if_empty_n,
    input wire                                           Yvec_inst_10_if_full_n,
    output wire                                          Yvec_inst_10_if_read,
    output wire                                          Yvec_inst_10_if_read_ce,
    output wire                                          Yvec_inst_10_if_write,
    output wire                                          Yvec_inst_10_if_write_ce,
    output wire                                          Yvec_inst_10_reset,
    output wire                                          Yvec_inst_11_clk,
    output wire [                                  32:0] Yvec_inst_11_if_din,
    input wire  [                                  32:0] Yvec_inst_11_if_dout,
    input wire                                           Yvec_inst_11_if_empty_n,
    input wire                                           Yvec_inst_11_if_full_n,
    output wire                                          Yvec_inst_11_if_read,
    output wire                                          Yvec_inst_11_if_read_ce,
    output wire                                          Yvec_inst_11_if_write,
    output wire                                          Yvec_inst_11_if_write_ce,
    output wire                                          Yvec_inst_11_reset,
    output wire                                          Yvec_inst_12_clk,
    output wire [                                  32:0] Yvec_inst_12_if_din,
    input wire  [                                  32:0] Yvec_inst_12_if_dout,
    input wire                                           Yvec_inst_12_if_empty_n,
    input wire                                           Yvec_inst_12_if_full_n,
    output wire                                          Yvec_inst_12_if_read,
    output wire                                          Yvec_inst_12_if_read_ce,
    output wire                                          Yvec_inst_12_if_write,
    output wire                                          Yvec_inst_12_if_write_ce,
    output wire                                          Yvec_inst_12_reset,
    output wire                                          Yvec_inst_13_clk,
    output wire [                                  32:0] Yvec_inst_13_if_din,
    input wire  [                                  32:0] Yvec_inst_13_if_dout,
    input wire                                           Yvec_inst_13_if_empty_n,
    input wire                                           Yvec_inst_13_if_full_n,
    output wire                                          Yvec_inst_13_if_read,
    output wire                                          Yvec_inst_13_if_read_ce,
    output wire                                          Yvec_inst_13_if_write,
    output wire                                          Yvec_inst_13_if_write_ce,
    output wire                                          Yvec_inst_13_reset,
    output wire                                          Yvec_inst_14_clk,
    output wire [                                  32:0] Yvec_inst_14_if_din,
    input wire  [                                  32:0] Yvec_inst_14_if_dout,
    input wire                                           Yvec_inst_14_if_empty_n,
    input wire                                           Yvec_inst_14_if_full_n,
    output wire                                          Yvec_inst_14_if_read,
    output wire                                          Yvec_inst_14_if_read_ce,
    output wire                                          Yvec_inst_14_if_write,
    output wire                                          Yvec_inst_14_if_write_ce,
    output wire                                          Yvec_inst_14_reset,
    output wire                                          Yvec_inst_15_clk,
    output wire [                                  32:0] Yvec_inst_15_if_din,
    input wire  [                                  32:0] Yvec_inst_15_if_dout,
    input wire                                           Yvec_inst_15_if_empty_n,
    input wire                                           Yvec_inst_15_if_full_n,
    output wire                                          Yvec_inst_15_if_read,
    output wire                                          Yvec_inst_15_if_read_ce,
    output wire                                          Yvec_inst_15_if_write,
    output wire                                          Yvec_inst_15_if_write_ce,
    output wire                                          Yvec_inst_15_reset,
    output wire                                          Yvec_inst_16_clk,
    output wire [                                  32:0] Yvec_inst_16_if_din,
    input wire  [                                  32:0] Yvec_inst_16_if_dout,
    input wire                                           Yvec_inst_16_if_empty_n,
    input wire                                           Yvec_inst_16_if_full_n,
    output wire                                          Yvec_inst_16_if_read,
    output wire                                          Yvec_inst_16_if_read_ce,
    output wire                                          Yvec_inst_16_if_write,
    output wire                                          Yvec_inst_16_if_write_ce,
    output wire                                          Yvec_inst_16_reset,
    output wire                                          Yvec_inst_17_clk,
    output wire [                                  32:0] Yvec_inst_17_if_din,
    input wire  [                                  32:0] Yvec_inst_17_if_dout,
    input wire                                           Yvec_inst_17_if_empty_n,
    input wire                                           Yvec_inst_17_if_full_n,
    output wire                                          Yvec_inst_17_if_read,
    output wire                                          Yvec_inst_17_if_read_ce,
    output wire                                          Yvec_inst_17_if_write,
    output wire                                          Yvec_inst_17_if_write_ce,
    output wire                                          Yvec_inst_17_reset,
    output wire                                          Yvec_inst_18_clk,
    output wire [                                  32:0] Yvec_inst_18_if_din,
    input wire  [                                  32:0] Yvec_inst_18_if_dout,
    input wire                                           Yvec_inst_18_if_empty_n,
    input wire                                           Yvec_inst_18_if_full_n,
    output wire                                          Yvec_inst_18_if_read,
    output wire                                          Yvec_inst_18_if_read_ce,
    output wire                                          Yvec_inst_18_if_write,
    output wire                                          Yvec_inst_18_if_write_ce,
    output wire                                          Yvec_inst_18_reset,
    output wire                                          Yvec_inst_19_clk,
    output wire [                                  32:0] Yvec_inst_19_if_din,
    input wire  [                                  32:0] Yvec_inst_19_if_dout,
    input wire                                           Yvec_inst_19_if_empty_n,
    input wire                                           Yvec_inst_19_if_full_n,
    output wire                                          Yvec_inst_19_if_read,
    output wire                                          Yvec_inst_19_if_read_ce,
    output wire                                          Yvec_inst_19_if_write,
    output wire                                          Yvec_inst_19_if_write_ce,
    output wire                                          Yvec_inst_19_reset,
    output wire                                          Yvec_inst_1_clk,
    output wire [                                  32:0] Yvec_inst_1_if_din,
    input wire  [                                  32:0] Yvec_inst_1_if_dout,
    input wire                                           Yvec_inst_1_if_empty_n,
    input wire                                           Yvec_inst_1_if_full_n,
    output wire                                          Yvec_inst_1_if_read,
    output wire                                          Yvec_inst_1_if_read_ce,
    output wire                                          Yvec_inst_1_if_write,
    output wire                                          Yvec_inst_1_if_write_ce,
    output wire                                          Yvec_inst_1_reset,
    output wire                                          Yvec_inst_20_clk,
    output wire [                                  32:0] Yvec_inst_20_if_din,
    input wire  [                                  32:0] Yvec_inst_20_if_dout,
    input wire                                           Yvec_inst_20_if_empty_n,
    input wire                                           Yvec_inst_20_if_full_n,
    output wire                                          Yvec_inst_20_if_read,
    output wire                                          Yvec_inst_20_if_read_ce,
    output wire                                          Yvec_inst_20_if_write,
    output wire                                          Yvec_inst_20_if_write_ce,
    output wire                                          Yvec_inst_20_reset,
    output wire                                          Yvec_inst_21_clk,
    output wire [                                  32:0] Yvec_inst_21_if_din,
    input wire  [                                  32:0] Yvec_inst_21_if_dout,
    input wire                                           Yvec_inst_21_if_empty_n,
    input wire                                           Yvec_inst_21_if_full_n,
    output wire                                          Yvec_inst_21_if_read,
    output wire                                          Yvec_inst_21_if_read_ce,
    output wire                                          Yvec_inst_21_if_write,
    output wire                                          Yvec_inst_21_if_write_ce,
    output wire                                          Yvec_inst_21_reset,
    output wire                                          Yvec_inst_22_clk,
    output wire [                                  32:0] Yvec_inst_22_if_din,
    input wire  [                                  32:0] Yvec_inst_22_if_dout,
    input wire                                           Yvec_inst_22_if_empty_n,
    input wire                                           Yvec_inst_22_if_full_n,
    output wire                                          Yvec_inst_22_if_read,
    output wire                                          Yvec_inst_22_if_read_ce,
    output wire                                          Yvec_inst_22_if_write,
    output wire                                          Yvec_inst_22_if_write_ce,
    output wire                                          Yvec_inst_22_reset,
    output wire                                          Yvec_inst_23_clk,
    output wire [                                  32:0] Yvec_inst_23_if_din,
    input wire  [                                  32:0] Yvec_inst_23_if_dout,
    input wire                                           Yvec_inst_23_if_empty_n,
    input wire                                           Yvec_inst_23_if_full_n,
    output wire                                          Yvec_inst_23_if_read,
    output wire                                          Yvec_inst_23_if_read_ce,
    output wire                                          Yvec_inst_23_if_write,
    output wire                                          Yvec_inst_23_if_write_ce,
    output wire                                          Yvec_inst_23_reset,
    output wire                                          Yvec_inst_24_clk,
    output wire [                                  32:0] Yvec_inst_24_if_din,
    input wire  [                                  32:0] Yvec_inst_24_if_dout,
    input wire                                           Yvec_inst_24_if_empty_n,
    input wire                                           Yvec_inst_24_if_full_n,
    output wire                                          Yvec_inst_24_if_read,
    output wire                                          Yvec_inst_24_if_read_ce,
    output wire                                          Yvec_inst_24_if_write,
    output wire                                          Yvec_inst_24_if_write_ce,
    output wire                                          Yvec_inst_24_reset,
    output wire                                          Yvec_inst_25_clk,
    output wire [                                  32:0] Yvec_inst_25_if_din,
    input wire  [                                  32:0] Yvec_inst_25_if_dout,
    input wire                                           Yvec_inst_25_if_empty_n,
    input wire                                           Yvec_inst_25_if_full_n,
    output wire                                          Yvec_inst_25_if_read,
    output wire                                          Yvec_inst_25_if_read_ce,
    output wire                                          Yvec_inst_25_if_write,
    output wire                                          Yvec_inst_25_if_write_ce,
    output wire                                          Yvec_inst_25_reset,
    output wire                                          Yvec_inst_26_clk,
    output wire [                                  32:0] Yvec_inst_26_if_din,
    input wire  [                                  32:0] Yvec_inst_26_if_dout,
    input wire                                           Yvec_inst_26_if_empty_n,
    input wire                                           Yvec_inst_26_if_full_n,
    output wire                                          Yvec_inst_26_if_read,
    output wire                                          Yvec_inst_26_if_read_ce,
    output wire                                          Yvec_inst_26_if_write,
    output wire                                          Yvec_inst_26_if_write_ce,
    output wire                                          Yvec_inst_26_reset,
    output wire                                          Yvec_inst_27_clk,
    output wire [                                  32:0] Yvec_inst_27_if_din,
    input wire  [                                  32:0] Yvec_inst_27_if_dout,
    input wire                                           Yvec_inst_27_if_empty_n,
    input wire                                           Yvec_inst_27_if_full_n,
    output wire                                          Yvec_inst_27_if_read,
    output wire                                          Yvec_inst_27_if_read_ce,
    output wire                                          Yvec_inst_27_if_write,
    output wire                                          Yvec_inst_27_if_write_ce,
    output wire                                          Yvec_inst_27_reset,
    output wire                                          Yvec_inst_28_clk,
    output wire [                                  32:0] Yvec_inst_28_if_din,
    input wire  [                                  32:0] Yvec_inst_28_if_dout,
    input wire                                           Yvec_inst_28_if_empty_n,
    input wire                                           Yvec_inst_28_if_full_n,
    output wire                                          Yvec_inst_28_if_read,
    output wire                                          Yvec_inst_28_if_read_ce,
    output wire                                          Yvec_inst_28_if_write,
    output wire                                          Yvec_inst_28_if_write_ce,
    output wire                                          Yvec_inst_28_reset,
    output wire                                          Yvec_inst_29_clk,
    output wire [                                  32:0] Yvec_inst_29_if_din,
    input wire  [                                  32:0] Yvec_inst_29_if_dout,
    input wire                                           Yvec_inst_29_if_empty_n,
    input wire                                           Yvec_inst_29_if_full_n,
    output wire                                          Yvec_inst_29_if_read,
    output wire                                          Yvec_inst_29_if_read_ce,
    output wire                                          Yvec_inst_29_if_write,
    output wire                                          Yvec_inst_29_if_write_ce,
    output wire                                          Yvec_inst_29_reset,
    output wire                                          Yvec_inst_2_clk,
    output wire [                                  32:0] Yvec_inst_2_if_din,
    input wire  [                                  32:0] Yvec_inst_2_if_dout,
    input wire                                           Yvec_inst_2_if_empty_n,
    input wire                                           Yvec_inst_2_if_full_n,
    output wire                                          Yvec_inst_2_if_read,
    output wire                                          Yvec_inst_2_if_read_ce,
    output wire                                          Yvec_inst_2_if_write,
    output wire                                          Yvec_inst_2_if_write_ce,
    output wire                                          Yvec_inst_2_reset,
    output wire                                          Yvec_inst_30_clk,
    output wire [                                  32:0] Yvec_inst_30_if_din,
    input wire  [                                  32:0] Yvec_inst_30_if_dout,
    input wire                                           Yvec_inst_30_if_empty_n,
    input wire                                           Yvec_inst_30_if_full_n,
    output wire                                          Yvec_inst_30_if_read,
    output wire                                          Yvec_inst_30_if_read_ce,
    output wire                                          Yvec_inst_30_if_write,
    output wire                                          Yvec_inst_30_if_write_ce,
    output wire                                          Yvec_inst_30_reset,
    output wire                                          Yvec_inst_31_clk,
    output wire [                                  32:0] Yvec_inst_31_if_din,
    input wire  [                                  32:0] Yvec_inst_31_if_dout,
    input wire                                           Yvec_inst_31_if_empty_n,
    input wire                                           Yvec_inst_31_if_full_n,
    output wire                                          Yvec_inst_31_if_read,
    output wire                                          Yvec_inst_31_if_read_ce,
    output wire                                          Yvec_inst_31_if_write,
    output wire                                          Yvec_inst_31_if_write_ce,
    output wire                                          Yvec_inst_31_reset,
    output wire                                          Yvec_inst_32_clk,
    output wire [                                  32:0] Yvec_inst_32_if_din,
    input wire  [                                  32:0] Yvec_inst_32_if_dout,
    input wire                                           Yvec_inst_32_if_empty_n,
    input wire                                           Yvec_inst_32_if_full_n,
    output wire                                          Yvec_inst_32_if_read,
    output wire                                          Yvec_inst_32_if_read_ce,
    output wire                                          Yvec_inst_32_if_write,
    output wire                                          Yvec_inst_32_if_write_ce,
    output wire                                          Yvec_inst_32_reset,
    output wire                                          Yvec_inst_33_clk,
    output wire [                                  32:0] Yvec_inst_33_if_din,
    input wire  [                                  32:0] Yvec_inst_33_if_dout,
    input wire                                           Yvec_inst_33_if_empty_n,
    input wire                                           Yvec_inst_33_if_full_n,
    output wire                                          Yvec_inst_33_if_read,
    output wire                                          Yvec_inst_33_if_read_ce,
    output wire                                          Yvec_inst_33_if_write,
    output wire                                          Yvec_inst_33_if_write_ce,
    output wire                                          Yvec_inst_33_reset,
    output wire                                          Yvec_inst_34_clk,
    output wire [                                  32:0] Yvec_inst_34_if_din,
    input wire  [                                  32:0] Yvec_inst_34_if_dout,
    input wire                                           Yvec_inst_34_if_empty_n,
    input wire                                           Yvec_inst_34_if_full_n,
    output wire                                          Yvec_inst_34_if_read,
    output wire                                          Yvec_inst_34_if_read_ce,
    output wire                                          Yvec_inst_34_if_write,
    output wire                                          Yvec_inst_34_if_write_ce,
    output wire                                          Yvec_inst_34_reset,
    output wire                                          Yvec_inst_35_clk,
    output wire [                                  32:0] Yvec_inst_35_if_din,
    input wire  [                                  32:0] Yvec_inst_35_if_dout,
    input wire                                           Yvec_inst_35_if_empty_n,
    input wire                                           Yvec_inst_35_if_full_n,
    output wire                                          Yvec_inst_35_if_read,
    output wire                                          Yvec_inst_35_if_read_ce,
    output wire                                          Yvec_inst_35_if_write,
    output wire                                          Yvec_inst_35_if_write_ce,
    output wire                                          Yvec_inst_35_reset,
    output wire                                          Yvec_inst_36_clk,
    output wire [                                  32:0] Yvec_inst_36_if_din,
    input wire  [                                  32:0] Yvec_inst_36_if_dout,
    input wire                                           Yvec_inst_36_if_empty_n,
    input wire                                           Yvec_inst_36_if_full_n,
    output wire                                          Yvec_inst_36_if_read,
    output wire                                          Yvec_inst_36_if_read_ce,
    output wire                                          Yvec_inst_36_if_write,
    output wire                                          Yvec_inst_36_if_write_ce,
    output wire                                          Yvec_inst_36_reset,
    output wire                                          Yvec_inst_37_clk,
    output wire [                                  32:0] Yvec_inst_37_if_din,
    input wire  [                                  32:0] Yvec_inst_37_if_dout,
    input wire                                           Yvec_inst_37_if_empty_n,
    input wire                                           Yvec_inst_37_if_full_n,
    output wire                                          Yvec_inst_37_if_read,
    output wire                                          Yvec_inst_37_if_read_ce,
    output wire                                          Yvec_inst_37_if_write,
    output wire                                          Yvec_inst_37_if_write_ce,
    output wire                                          Yvec_inst_37_reset,
    output wire                                          Yvec_inst_38_clk,
    output wire [                                  32:0] Yvec_inst_38_if_din,
    input wire  [                                  32:0] Yvec_inst_38_if_dout,
    input wire                                           Yvec_inst_38_if_empty_n,
    input wire                                           Yvec_inst_38_if_full_n,
    output wire                                          Yvec_inst_38_if_read,
    output wire                                          Yvec_inst_38_if_read_ce,
    output wire                                          Yvec_inst_38_if_write,
    output wire                                          Yvec_inst_38_if_write_ce,
    output wire                                          Yvec_inst_38_reset,
    output wire                                          Yvec_inst_39_clk,
    output wire [                                  32:0] Yvec_inst_39_if_din,
    input wire  [                                  32:0] Yvec_inst_39_if_dout,
    input wire                                           Yvec_inst_39_if_empty_n,
    input wire                                           Yvec_inst_39_if_full_n,
    output wire                                          Yvec_inst_39_if_read,
    output wire                                          Yvec_inst_39_if_read_ce,
    output wire                                          Yvec_inst_39_if_write,
    output wire                                          Yvec_inst_39_if_write_ce,
    output wire                                          Yvec_inst_39_reset,
    output wire                                          Yvec_inst_3_clk,
    output wire [                                  32:0] Yvec_inst_3_if_din,
    input wire  [                                  32:0] Yvec_inst_3_if_dout,
    input wire                                           Yvec_inst_3_if_empty_n,
    input wire                                           Yvec_inst_3_if_full_n,
    output wire                                          Yvec_inst_3_if_read,
    output wire                                          Yvec_inst_3_if_read_ce,
    output wire                                          Yvec_inst_3_if_write,
    output wire                                          Yvec_inst_3_if_write_ce,
    output wire                                          Yvec_inst_3_reset,
    output wire                                          Yvec_inst_40_clk,
    output wire [                                  32:0] Yvec_inst_40_if_din,
    input wire  [                                  32:0] Yvec_inst_40_if_dout,
    input wire                                           Yvec_inst_40_if_empty_n,
    input wire                                           Yvec_inst_40_if_full_n,
    output wire                                          Yvec_inst_40_if_read,
    output wire                                          Yvec_inst_40_if_read_ce,
    output wire                                          Yvec_inst_40_if_write,
    output wire                                          Yvec_inst_40_if_write_ce,
    output wire                                          Yvec_inst_40_reset,
    output wire                                          Yvec_inst_41_clk,
    output wire [                                  32:0] Yvec_inst_41_if_din,
    input wire  [                                  32:0] Yvec_inst_41_if_dout,
    input wire                                           Yvec_inst_41_if_empty_n,
    input wire                                           Yvec_inst_41_if_full_n,
    output wire                                          Yvec_inst_41_if_read,
    output wire                                          Yvec_inst_41_if_read_ce,
    output wire                                          Yvec_inst_41_if_write,
    output wire                                          Yvec_inst_41_if_write_ce,
    output wire                                          Yvec_inst_41_reset,
    output wire                                          Yvec_inst_42_clk,
    output wire [                                  32:0] Yvec_inst_42_if_din,
    input wire  [                                  32:0] Yvec_inst_42_if_dout,
    input wire                                           Yvec_inst_42_if_empty_n,
    input wire                                           Yvec_inst_42_if_full_n,
    output wire                                          Yvec_inst_42_if_read,
    output wire                                          Yvec_inst_42_if_read_ce,
    output wire                                          Yvec_inst_42_if_write,
    output wire                                          Yvec_inst_42_if_write_ce,
    output wire                                          Yvec_inst_42_reset,
    output wire                                          Yvec_inst_43_clk,
    output wire [                                  32:0] Yvec_inst_43_if_din,
    input wire  [                                  32:0] Yvec_inst_43_if_dout,
    input wire                                           Yvec_inst_43_if_empty_n,
    input wire                                           Yvec_inst_43_if_full_n,
    output wire                                          Yvec_inst_43_if_read,
    output wire                                          Yvec_inst_43_if_read_ce,
    output wire                                          Yvec_inst_43_if_write,
    output wire                                          Yvec_inst_43_if_write_ce,
    output wire                                          Yvec_inst_43_reset,
    output wire                                          Yvec_inst_44_clk,
    output wire [                                  32:0] Yvec_inst_44_if_din,
    input wire  [                                  32:0] Yvec_inst_44_if_dout,
    input wire                                           Yvec_inst_44_if_empty_n,
    input wire                                           Yvec_inst_44_if_full_n,
    output wire                                          Yvec_inst_44_if_read,
    output wire                                          Yvec_inst_44_if_read_ce,
    output wire                                          Yvec_inst_44_if_write,
    output wire                                          Yvec_inst_44_if_write_ce,
    output wire                                          Yvec_inst_44_reset,
    output wire                                          Yvec_inst_45_clk,
    output wire [                                  32:0] Yvec_inst_45_if_din,
    input wire  [                                  32:0] Yvec_inst_45_if_dout,
    input wire                                           Yvec_inst_45_if_empty_n,
    input wire                                           Yvec_inst_45_if_full_n,
    output wire                                          Yvec_inst_45_if_read,
    output wire                                          Yvec_inst_45_if_read_ce,
    output wire                                          Yvec_inst_45_if_write,
    output wire                                          Yvec_inst_45_if_write_ce,
    output wire                                          Yvec_inst_45_reset,
    output wire                                          Yvec_inst_46_clk,
    output wire [                                  32:0] Yvec_inst_46_if_din,
    input wire  [                                  32:0] Yvec_inst_46_if_dout,
    input wire                                           Yvec_inst_46_if_empty_n,
    input wire                                           Yvec_inst_46_if_full_n,
    output wire                                          Yvec_inst_46_if_read,
    output wire                                          Yvec_inst_46_if_read_ce,
    output wire                                          Yvec_inst_46_if_write,
    output wire                                          Yvec_inst_46_if_write_ce,
    output wire                                          Yvec_inst_46_reset,
    output wire                                          Yvec_inst_47_clk,
    output wire [                                  32:0] Yvec_inst_47_if_din,
    input wire  [                                  32:0] Yvec_inst_47_if_dout,
    input wire                                           Yvec_inst_47_if_empty_n,
    input wire                                           Yvec_inst_47_if_full_n,
    output wire                                          Yvec_inst_47_if_read,
    output wire                                          Yvec_inst_47_if_read_ce,
    output wire                                          Yvec_inst_47_if_write,
    output wire                                          Yvec_inst_47_if_write_ce,
    output wire                                          Yvec_inst_47_reset,
    output wire                                          Yvec_inst_4_clk,
    output wire [                                  32:0] Yvec_inst_4_if_din,
    input wire  [                                  32:0] Yvec_inst_4_if_dout,
    input wire                                           Yvec_inst_4_if_empty_n,
    input wire                                           Yvec_inst_4_if_full_n,
    output wire                                          Yvec_inst_4_if_read,
    output wire                                          Yvec_inst_4_if_read_ce,
    output wire                                          Yvec_inst_4_if_write,
    output wire                                          Yvec_inst_4_if_write_ce,
    output wire                                          Yvec_inst_4_reset,
    output wire                                          Yvec_inst_5_clk,
    output wire [                                  32:0] Yvec_inst_5_if_din,
    input wire  [                                  32:0] Yvec_inst_5_if_dout,
    input wire                                           Yvec_inst_5_if_empty_n,
    input wire                                           Yvec_inst_5_if_full_n,
    output wire                                          Yvec_inst_5_if_read,
    output wire                                          Yvec_inst_5_if_read_ce,
    output wire                                          Yvec_inst_5_if_write,
    output wire                                          Yvec_inst_5_if_write_ce,
    output wire                                          Yvec_inst_5_reset,
    output wire                                          Yvec_inst_6_clk,
    output wire [                                  32:0] Yvec_inst_6_if_din,
    input wire  [                                  32:0] Yvec_inst_6_if_dout,
    input wire                                           Yvec_inst_6_if_empty_n,
    input wire                                           Yvec_inst_6_if_full_n,
    output wire                                          Yvec_inst_6_if_read,
    output wire                                          Yvec_inst_6_if_read_ce,
    output wire                                          Yvec_inst_6_if_write,
    output wire                                          Yvec_inst_6_if_write_ce,
    output wire                                          Yvec_inst_6_reset,
    output wire                                          Yvec_inst_7_clk,
    output wire [                                  32:0] Yvec_inst_7_if_din,
    input wire  [                                  32:0] Yvec_inst_7_if_dout,
    input wire                                           Yvec_inst_7_if_empty_n,
    input wire                                           Yvec_inst_7_if_full_n,
    output wire                                          Yvec_inst_7_if_read,
    output wire                                          Yvec_inst_7_if_read_ce,
    output wire                                          Yvec_inst_7_if_write,
    output wire                                          Yvec_inst_7_if_write_ce,
    output wire                                          Yvec_inst_7_reset,
    output wire                                          Yvec_inst_8_clk,
    output wire [                                  32:0] Yvec_inst_8_if_din,
    input wire  [                                  32:0] Yvec_inst_8_if_dout,
    input wire                                           Yvec_inst_8_if_empty_n,
    input wire                                           Yvec_inst_8_if_full_n,
    output wire                                          Yvec_inst_8_if_read,
    output wire                                          Yvec_inst_8_if_read_ce,
    output wire                                          Yvec_inst_8_if_write,
    output wire                                          Yvec_inst_8_if_write_ce,
    output wire                                          Yvec_inst_8_reset,
    output wire                                          Yvec_inst_9_clk,
    output wire [                                  32:0] Yvec_inst_9_if_din,
    input wire  [                                  32:0] Yvec_inst_9_if_dout,
    input wire                                           Yvec_inst_9_if_empty_n,
    input wire                                           Yvec_inst_9_if_full_n,
    output wire                                          Yvec_inst_9_if_read,
    output wire                                          Yvec_inst_9_if_read_ce,
    output wire                                          Yvec_inst_9_if_write,
    output wire                                          Yvec_inst_9_if_write_ce,
    output wire                                          Yvec_inst_9_reset,
    output wire                                          fifo_A_0_clk,
    output wire [                                 512:0] fifo_A_0_if_din,
    input wire  [                                 512:0] fifo_A_0_if_dout,
    input wire                                           fifo_A_0_if_empty_n,
    input wire                                           fifo_A_0_if_full_n,
    output wire                                          fifo_A_0_if_read,
    output wire                                          fifo_A_0_if_read_ce,
    output wire                                          fifo_A_0_if_write,
    output wire                                          fifo_A_0_if_write_ce,
    output wire                                          fifo_A_0_reset,
    output wire                                          fifo_A_10_clk,
    output wire [                                 512:0] fifo_A_10_if_din,
    input wire  [                                 512:0] fifo_A_10_if_dout,
    input wire                                           fifo_A_10_if_empty_n,
    input wire                                           fifo_A_10_if_full_n,
    output wire                                          fifo_A_10_if_read,
    output wire                                          fifo_A_10_if_read_ce,
    output wire                                          fifo_A_10_if_write,
    output wire                                          fifo_A_10_if_write_ce,
    output wire                                          fifo_A_10_reset,
    output wire                                          fifo_A_11_clk,
    output wire [                                 512:0] fifo_A_11_if_din,
    input wire  [                                 512:0] fifo_A_11_if_dout,
    input wire                                           fifo_A_11_if_empty_n,
    input wire                                           fifo_A_11_if_full_n,
    output wire                                          fifo_A_11_if_read,
    output wire                                          fifo_A_11_if_read_ce,
    output wire                                          fifo_A_11_if_write,
    output wire                                          fifo_A_11_if_write_ce,
    output wire                                          fifo_A_11_reset,
    output wire                                          fifo_A_12_clk,
    output wire [                                 512:0] fifo_A_12_if_din,
    input wire  [                                 512:0] fifo_A_12_if_dout,
    input wire                                           fifo_A_12_if_empty_n,
    input wire                                           fifo_A_12_if_full_n,
    output wire                                          fifo_A_12_if_read,
    output wire                                          fifo_A_12_if_read_ce,
    output wire                                          fifo_A_12_if_write,
    output wire                                          fifo_A_12_if_write_ce,
    output wire                                          fifo_A_12_reset,
    output wire                                          fifo_A_13_clk,
    output wire [                                 512:0] fifo_A_13_if_din,
    input wire  [                                 512:0] fifo_A_13_if_dout,
    input wire                                           fifo_A_13_if_empty_n,
    input wire                                           fifo_A_13_if_full_n,
    output wire                                          fifo_A_13_if_read,
    output wire                                          fifo_A_13_if_read_ce,
    output wire                                          fifo_A_13_if_write,
    output wire                                          fifo_A_13_if_write_ce,
    output wire                                          fifo_A_13_reset,
    output wire                                          fifo_A_14_clk,
    output wire [                                 512:0] fifo_A_14_if_din,
    input wire  [                                 512:0] fifo_A_14_if_dout,
    input wire                                           fifo_A_14_if_empty_n,
    input wire                                           fifo_A_14_if_full_n,
    output wire                                          fifo_A_14_if_read,
    output wire                                          fifo_A_14_if_read_ce,
    output wire                                          fifo_A_14_if_write,
    output wire                                          fifo_A_14_if_write_ce,
    output wire                                          fifo_A_14_reset,
    output wire                                          fifo_A_15_clk,
    output wire [                                 512:0] fifo_A_15_if_din,
    input wire  [                                 512:0] fifo_A_15_if_dout,
    input wire                                           fifo_A_15_if_empty_n,
    input wire                                           fifo_A_15_if_full_n,
    output wire                                          fifo_A_15_if_read,
    output wire                                          fifo_A_15_if_read_ce,
    output wire                                          fifo_A_15_if_write,
    output wire                                          fifo_A_15_if_write_ce,
    output wire                                          fifo_A_15_reset,
    output wire                                          fifo_A_16_clk,
    output wire [                                 512:0] fifo_A_16_if_din,
    input wire  [                                 512:0] fifo_A_16_if_dout,
    input wire                                           fifo_A_16_if_empty_n,
    input wire                                           fifo_A_16_if_full_n,
    output wire                                          fifo_A_16_if_read,
    output wire                                          fifo_A_16_if_read_ce,
    output wire                                          fifo_A_16_if_write,
    output wire                                          fifo_A_16_if_write_ce,
    output wire                                          fifo_A_16_reset,
    output wire                                          fifo_A_17_clk,
    output wire [                                 512:0] fifo_A_17_if_din,
    input wire  [                                 512:0] fifo_A_17_if_dout,
    input wire                                           fifo_A_17_if_empty_n,
    input wire                                           fifo_A_17_if_full_n,
    output wire                                          fifo_A_17_if_read,
    output wire                                          fifo_A_17_if_read_ce,
    output wire                                          fifo_A_17_if_write,
    output wire                                          fifo_A_17_if_write_ce,
    output wire                                          fifo_A_17_reset,
    output wire                                          fifo_A_18_clk,
    output wire [                                 512:0] fifo_A_18_if_din,
    input wire  [                                 512:0] fifo_A_18_if_dout,
    input wire                                           fifo_A_18_if_empty_n,
    input wire                                           fifo_A_18_if_full_n,
    output wire                                          fifo_A_18_if_read,
    output wire                                          fifo_A_18_if_read_ce,
    output wire                                          fifo_A_18_if_write,
    output wire                                          fifo_A_18_if_write_ce,
    output wire                                          fifo_A_18_reset,
    output wire                                          fifo_A_19_clk,
    output wire [                                 512:0] fifo_A_19_if_din,
    input wire  [                                 512:0] fifo_A_19_if_dout,
    input wire                                           fifo_A_19_if_empty_n,
    input wire                                           fifo_A_19_if_full_n,
    output wire                                          fifo_A_19_if_read,
    output wire                                          fifo_A_19_if_read_ce,
    output wire                                          fifo_A_19_if_write,
    output wire                                          fifo_A_19_if_write_ce,
    output wire                                          fifo_A_19_reset,
    output wire                                          fifo_A_1_clk,
    output wire [                                 512:0] fifo_A_1_if_din,
    input wire  [                                 512:0] fifo_A_1_if_dout,
    input wire                                           fifo_A_1_if_empty_n,
    input wire                                           fifo_A_1_if_full_n,
    output wire                                          fifo_A_1_if_read,
    output wire                                          fifo_A_1_if_read_ce,
    output wire                                          fifo_A_1_if_write,
    output wire                                          fifo_A_1_if_write_ce,
    output wire                                          fifo_A_1_reset,
    output wire                                          fifo_A_20_clk,
    output wire [                                 512:0] fifo_A_20_if_din,
    input wire  [                                 512:0] fifo_A_20_if_dout,
    input wire                                           fifo_A_20_if_empty_n,
    input wire                                           fifo_A_20_if_full_n,
    output wire                                          fifo_A_20_if_read,
    output wire                                          fifo_A_20_if_read_ce,
    output wire                                          fifo_A_20_if_write,
    output wire                                          fifo_A_20_if_write_ce,
    output wire                                          fifo_A_20_reset,
    output wire                                          fifo_A_21_clk,
    output wire [                                 512:0] fifo_A_21_if_din,
    input wire  [                                 512:0] fifo_A_21_if_dout,
    input wire                                           fifo_A_21_if_empty_n,
    input wire                                           fifo_A_21_if_full_n,
    output wire                                          fifo_A_21_if_read,
    output wire                                          fifo_A_21_if_read_ce,
    output wire                                          fifo_A_21_if_write,
    output wire                                          fifo_A_21_if_write_ce,
    output wire                                          fifo_A_21_reset,
    output wire                                          fifo_A_22_clk,
    output wire [                                 512:0] fifo_A_22_if_din,
    input wire  [                                 512:0] fifo_A_22_if_dout,
    input wire                                           fifo_A_22_if_empty_n,
    input wire                                           fifo_A_22_if_full_n,
    output wire                                          fifo_A_22_if_read,
    output wire                                          fifo_A_22_if_read_ce,
    output wire                                          fifo_A_22_if_write,
    output wire                                          fifo_A_22_if_write_ce,
    output wire                                          fifo_A_22_reset,
    output wire                                          fifo_A_23_clk,
    output wire [                                 512:0] fifo_A_23_if_din,
    input wire  [                                 512:0] fifo_A_23_if_dout,
    input wire                                           fifo_A_23_if_empty_n,
    input wire                                           fifo_A_23_if_full_n,
    output wire                                          fifo_A_23_if_read,
    output wire                                          fifo_A_23_if_read_ce,
    output wire                                          fifo_A_23_if_write,
    output wire                                          fifo_A_23_if_write_ce,
    output wire                                          fifo_A_23_reset,
    output wire                                          fifo_A_24_clk,
    output wire [                                 512:0] fifo_A_24_if_din,
    input wire  [                                 512:0] fifo_A_24_if_dout,
    input wire                                           fifo_A_24_if_empty_n,
    input wire                                           fifo_A_24_if_full_n,
    output wire                                          fifo_A_24_if_read,
    output wire                                          fifo_A_24_if_read_ce,
    output wire                                          fifo_A_24_if_write,
    output wire                                          fifo_A_24_if_write_ce,
    output wire                                          fifo_A_24_reset,
    output wire                                          fifo_A_25_clk,
    output wire [                                 512:0] fifo_A_25_if_din,
    input wire  [                                 512:0] fifo_A_25_if_dout,
    input wire                                           fifo_A_25_if_empty_n,
    input wire                                           fifo_A_25_if_full_n,
    output wire                                          fifo_A_25_if_read,
    output wire                                          fifo_A_25_if_read_ce,
    output wire                                          fifo_A_25_if_write,
    output wire                                          fifo_A_25_if_write_ce,
    output wire                                          fifo_A_25_reset,
    output wire                                          fifo_A_26_clk,
    output wire [                                 512:0] fifo_A_26_if_din,
    input wire  [                                 512:0] fifo_A_26_if_dout,
    input wire                                           fifo_A_26_if_empty_n,
    input wire                                           fifo_A_26_if_full_n,
    output wire                                          fifo_A_26_if_read,
    output wire                                          fifo_A_26_if_read_ce,
    output wire                                          fifo_A_26_if_write,
    output wire                                          fifo_A_26_if_write_ce,
    output wire                                          fifo_A_26_reset,
    output wire                                          fifo_A_27_clk,
    output wire [                                 512:0] fifo_A_27_if_din,
    input wire  [                                 512:0] fifo_A_27_if_dout,
    input wire                                           fifo_A_27_if_empty_n,
    input wire                                           fifo_A_27_if_full_n,
    output wire                                          fifo_A_27_if_read,
    output wire                                          fifo_A_27_if_read_ce,
    output wire                                          fifo_A_27_if_write,
    output wire                                          fifo_A_27_if_write_ce,
    output wire                                          fifo_A_27_reset,
    output wire                                          fifo_A_28_clk,
    output wire [                                 512:0] fifo_A_28_if_din,
    input wire  [                                 512:0] fifo_A_28_if_dout,
    input wire                                           fifo_A_28_if_empty_n,
    input wire                                           fifo_A_28_if_full_n,
    output wire                                          fifo_A_28_if_read,
    output wire                                          fifo_A_28_if_read_ce,
    output wire                                          fifo_A_28_if_write,
    output wire                                          fifo_A_28_if_write_ce,
    output wire                                          fifo_A_28_reset,
    output wire                                          fifo_A_29_clk,
    output wire [                                 512:0] fifo_A_29_if_din,
    input wire  [                                 512:0] fifo_A_29_if_dout,
    input wire                                           fifo_A_29_if_empty_n,
    input wire                                           fifo_A_29_if_full_n,
    output wire                                          fifo_A_29_if_read,
    output wire                                          fifo_A_29_if_read_ce,
    output wire                                          fifo_A_29_if_write,
    output wire                                          fifo_A_29_if_write_ce,
    output wire                                          fifo_A_29_reset,
    output wire                                          fifo_A_2_clk,
    output wire [                                 512:0] fifo_A_2_if_din,
    input wire  [                                 512:0] fifo_A_2_if_dout,
    input wire                                           fifo_A_2_if_empty_n,
    input wire                                           fifo_A_2_if_full_n,
    output wire                                          fifo_A_2_if_read,
    output wire                                          fifo_A_2_if_read_ce,
    output wire                                          fifo_A_2_if_write,
    output wire                                          fifo_A_2_if_write_ce,
    output wire                                          fifo_A_2_reset,
    output wire                                          fifo_A_30_clk,
    output wire [                                 512:0] fifo_A_30_if_din,
    input wire  [                                 512:0] fifo_A_30_if_dout,
    input wire                                           fifo_A_30_if_empty_n,
    input wire                                           fifo_A_30_if_full_n,
    output wire                                          fifo_A_30_if_read,
    output wire                                          fifo_A_30_if_read_ce,
    output wire                                          fifo_A_30_if_write,
    output wire                                          fifo_A_30_if_write_ce,
    output wire                                          fifo_A_30_reset,
    output wire                                          fifo_A_31_clk,
    output wire [                                 512:0] fifo_A_31_if_din,
    input wire  [                                 512:0] fifo_A_31_if_dout,
    input wire                                           fifo_A_31_if_empty_n,
    input wire                                           fifo_A_31_if_full_n,
    output wire                                          fifo_A_31_if_read,
    output wire                                          fifo_A_31_if_read_ce,
    output wire                                          fifo_A_31_if_write,
    output wire                                          fifo_A_31_if_write_ce,
    output wire                                          fifo_A_31_reset,
    output wire                                          fifo_A_32_clk,
    output wire [                                 512:0] fifo_A_32_if_din,
    input wire  [                                 512:0] fifo_A_32_if_dout,
    input wire                                           fifo_A_32_if_empty_n,
    input wire                                           fifo_A_32_if_full_n,
    output wire                                          fifo_A_32_if_read,
    output wire                                          fifo_A_32_if_read_ce,
    output wire                                          fifo_A_32_if_write,
    output wire                                          fifo_A_32_if_write_ce,
    output wire                                          fifo_A_32_reset,
    output wire                                          fifo_A_33_clk,
    output wire [                                 512:0] fifo_A_33_if_din,
    input wire  [                                 512:0] fifo_A_33_if_dout,
    input wire                                           fifo_A_33_if_empty_n,
    input wire                                           fifo_A_33_if_full_n,
    output wire                                          fifo_A_33_if_read,
    output wire                                          fifo_A_33_if_read_ce,
    output wire                                          fifo_A_33_if_write,
    output wire                                          fifo_A_33_if_write_ce,
    output wire                                          fifo_A_33_reset,
    output wire                                          fifo_A_34_clk,
    output wire [                                 512:0] fifo_A_34_if_din,
    input wire  [                                 512:0] fifo_A_34_if_dout,
    input wire                                           fifo_A_34_if_empty_n,
    input wire                                           fifo_A_34_if_full_n,
    output wire                                          fifo_A_34_if_read,
    output wire                                          fifo_A_34_if_read_ce,
    output wire                                          fifo_A_34_if_write,
    output wire                                          fifo_A_34_if_write_ce,
    output wire                                          fifo_A_34_reset,
    output wire                                          fifo_A_35_clk,
    output wire [                                 512:0] fifo_A_35_if_din,
    input wire  [                                 512:0] fifo_A_35_if_dout,
    input wire                                           fifo_A_35_if_empty_n,
    input wire                                           fifo_A_35_if_full_n,
    output wire                                          fifo_A_35_if_read,
    output wire                                          fifo_A_35_if_read_ce,
    output wire                                          fifo_A_35_if_write,
    output wire                                          fifo_A_35_if_write_ce,
    output wire                                          fifo_A_35_reset,
    output wire                                          fifo_A_36_clk,
    output wire [                                 512:0] fifo_A_36_if_din,
    input wire  [                                 512:0] fifo_A_36_if_dout,
    input wire                                           fifo_A_36_if_empty_n,
    input wire                                           fifo_A_36_if_full_n,
    output wire                                          fifo_A_36_if_read,
    output wire                                          fifo_A_36_if_read_ce,
    output wire                                          fifo_A_36_if_write,
    output wire                                          fifo_A_36_if_write_ce,
    output wire                                          fifo_A_36_reset,
    output wire                                          fifo_A_37_clk,
    output wire [                                 512:0] fifo_A_37_if_din,
    input wire  [                                 512:0] fifo_A_37_if_dout,
    input wire                                           fifo_A_37_if_empty_n,
    input wire                                           fifo_A_37_if_full_n,
    output wire                                          fifo_A_37_if_read,
    output wire                                          fifo_A_37_if_read_ce,
    output wire                                          fifo_A_37_if_write,
    output wire                                          fifo_A_37_if_write_ce,
    output wire                                          fifo_A_37_reset,
    output wire                                          fifo_A_38_clk,
    output wire [                                 512:0] fifo_A_38_if_din,
    input wire  [                                 512:0] fifo_A_38_if_dout,
    input wire                                           fifo_A_38_if_empty_n,
    input wire                                           fifo_A_38_if_full_n,
    output wire                                          fifo_A_38_if_read,
    output wire                                          fifo_A_38_if_read_ce,
    output wire                                          fifo_A_38_if_write,
    output wire                                          fifo_A_38_if_write_ce,
    output wire                                          fifo_A_38_reset,
    output wire                                          fifo_A_39_clk,
    output wire [                                 512:0] fifo_A_39_if_din,
    input wire  [                                 512:0] fifo_A_39_if_dout,
    input wire                                           fifo_A_39_if_empty_n,
    input wire                                           fifo_A_39_if_full_n,
    output wire                                          fifo_A_39_if_read,
    output wire                                          fifo_A_39_if_read_ce,
    output wire                                          fifo_A_39_if_write,
    output wire                                          fifo_A_39_if_write_ce,
    output wire                                          fifo_A_39_reset,
    output wire                                          fifo_A_3_clk,
    output wire [                                 512:0] fifo_A_3_if_din,
    input wire  [                                 512:0] fifo_A_3_if_dout,
    input wire                                           fifo_A_3_if_empty_n,
    input wire                                           fifo_A_3_if_full_n,
    output wire                                          fifo_A_3_if_read,
    output wire                                          fifo_A_3_if_read_ce,
    output wire                                          fifo_A_3_if_write,
    output wire                                          fifo_A_3_if_write_ce,
    output wire                                          fifo_A_3_reset,
    output wire                                          fifo_A_40_clk,
    output wire [                                 512:0] fifo_A_40_if_din,
    input wire  [                                 512:0] fifo_A_40_if_dout,
    input wire                                           fifo_A_40_if_empty_n,
    input wire                                           fifo_A_40_if_full_n,
    output wire                                          fifo_A_40_if_read,
    output wire                                          fifo_A_40_if_read_ce,
    output wire                                          fifo_A_40_if_write,
    output wire                                          fifo_A_40_if_write_ce,
    output wire                                          fifo_A_40_reset,
    output wire                                          fifo_A_41_clk,
    output wire [                                 512:0] fifo_A_41_if_din,
    input wire  [                                 512:0] fifo_A_41_if_dout,
    input wire                                           fifo_A_41_if_empty_n,
    input wire                                           fifo_A_41_if_full_n,
    output wire                                          fifo_A_41_if_read,
    output wire                                          fifo_A_41_if_read_ce,
    output wire                                          fifo_A_41_if_write,
    output wire                                          fifo_A_41_if_write_ce,
    output wire                                          fifo_A_41_reset,
    output wire                                          fifo_A_42_clk,
    output wire [                                 512:0] fifo_A_42_if_din,
    input wire  [                                 512:0] fifo_A_42_if_dout,
    input wire                                           fifo_A_42_if_empty_n,
    input wire                                           fifo_A_42_if_full_n,
    output wire                                          fifo_A_42_if_read,
    output wire                                          fifo_A_42_if_read_ce,
    output wire                                          fifo_A_42_if_write,
    output wire                                          fifo_A_42_if_write_ce,
    output wire                                          fifo_A_42_reset,
    output wire                                          fifo_A_43_clk,
    output wire [                                 512:0] fifo_A_43_if_din,
    input wire  [                                 512:0] fifo_A_43_if_dout,
    input wire                                           fifo_A_43_if_empty_n,
    input wire                                           fifo_A_43_if_full_n,
    output wire                                          fifo_A_43_if_read,
    output wire                                          fifo_A_43_if_read_ce,
    output wire                                          fifo_A_43_if_write,
    output wire                                          fifo_A_43_if_write_ce,
    output wire                                          fifo_A_43_reset,
    output wire                                          fifo_A_44_clk,
    output wire [                                 512:0] fifo_A_44_if_din,
    input wire  [                                 512:0] fifo_A_44_if_dout,
    input wire                                           fifo_A_44_if_empty_n,
    input wire                                           fifo_A_44_if_full_n,
    output wire                                          fifo_A_44_if_read,
    output wire                                          fifo_A_44_if_read_ce,
    output wire                                          fifo_A_44_if_write,
    output wire                                          fifo_A_44_if_write_ce,
    output wire                                          fifo_A_44_reset,
    output wire                                          fifo_A_45_clk,
    output wire [                                 512:0] fifo_A_45_if_din,
    input wire  [                                 512:0] fifo_A_45_if_dout,
    input wire                                           fifo_A_45_if_empty_n,
    input wire                                           fifo_A_45_if_full_n,
    output wire                                          fifo_A_45_if_read,
    output wire                                          fifo_A_45_if_read_ce,
    output wire                                          fifo_A_45_if_write,
    output wire                                          fifo_A_45_if_write_ce,
    output wire                                          fifo_A_45_reset,
    output wire                                          fifo_A_46_clk,
    output wire [                                 512:0] fifo_A_46_if_din,
    input wire  [                                 512:0] fifo_A_46_if_dout,
    input wire                                           fifo_A_46_if_empty_n,
    input wire                                           fifo_A_46_if_full_n,
    output wire                                          fifo_A_46_if_read,
    output wire                                          fifo_A_46_if_read_ce,
    output wire                                          fifo_A_46_if_write,
    output wire                                          fifo_A_46_if_write_ce,
    output wire                                          fifo_A_46_reset,
    output wire                                          fifo_A_47_clk,
    output wire [                                 512:0] fifo_A_47_if_din,
    input wire  [                                 512:0] fifo_A_47_if_dout,
    input wire                                           fifo_A_47_if_empty_n,
    input wire                                           fifo_A_47_if_full_n,
    output wire                                          fifo_A_47_if_read,
    output wire                                          fifo_A_47_if_read_ce,
    output wire                                          fifo_A_47_if_write,
    output wire                                          fifo_A_47_if_write_ce,
    output wire                                          fifo_A_47_reset,
    output wire                                          fifo_A_4_clk,
    output wire [                                 512:0] fifo_A_4_if_din,
    input wire  [                                 512:0] fifo_A_4_if_dout,
    input wire                                           fifo_A_4_if_empty_n,
    input wire                                           fifo_A_4_if_full_n,
    output wire                                          fifo_A_4_if_read,
    output wire                                          fifo_A_4_if_read_ce,
    output wire                                          fifo_A_4_if_write,
    output wire                                          fifo_A_4_if_write_ce,
    output wire                                          fifo_A_4_reset,
    output wire                                          fifo_A_5_clk,
    output wire [                                 512:0] fifo_A_5_if_din,
    input wire  [                                 512:0] fifo_A_5_if_dout,
    input wire                                           fifo_A_5_if_empty_n,
    input wire                                           fifo_A_5_if_full_n,
    output wire                                          fifo_A_5_if_read,
    output wire                                          fifo_A_5_if_read_ce,
    output wire                                          fifo_A_5_if_write,
    output wire                                          fifo_A_5_if_write_ce,
    output wire                                          fifo_A_5_reset,
    output wire                                          fifo_A_6_clk,
    output wire [                                 512:0] fifo_A_6_if_din,
    input wire  [                                 512:0] fifo_A_6_if_dout,
    input wire                                           fifo_A_6_if_empty_n,
    input wire                                           fifo_A_6_if_full_n,
    output wire                                          fifo_A_6_if_read,
    output wire                                          fifo_A_6_if_read_ce,
    output wire                                          fifo_A_6_if_write,
    output wire                                          fifo_A_6_if_write_ce,
    output wire                                          fifo_A_6_reset,
    output wire                                          fifo_A_7_clk,
    output wire [                                 512:0] fifo_A_7_if_din,
    input wire  [                                 512:0] fifo_A_7_if_dout,
    input wire                                           fifo_A_7_if_empty_n,
    input wire                                           fifo_A_7_if_full_n,
    output wire                                          fifo_A_7_if_read,
    output wire                                          fifo_A_7_if_read_ce,
    output wire                                          fifo_A_7_if_write,
    output wire                                          fifo_A_7_if_write_ce,
    output wire                                          fifo_A_7_reset,
    output wire                                          fifo_A_8_clk,
    output wire [                                 512:0] fifo_A_8_if_din,
    input wire  [                                 512:0] fifo_A_8_if_dout,
    input wire                                           fifo_A_8_if_empty_n,
    input wire                                           fifo_A_8_if_full_n,
    output wire                                          fifo_A_8_if_read,
    output wire                                          fifo_A_8_if_read_ce,
    output wire                                          fifo_A_8_if_write,
    output wire                                          fifo_A_8_if_write_ce,
    output wire                                          fifo_A_8_reset,
    output wire                                          fifo_A_9_clk,
    output wire [                                 512:0] fifo_A_9_if_din,
    input wire  [                                 512:0] fifo_A_9_if_dout,
    input wire                                           fifo_A_9_if_empty_n,
    input wire                                           fifo_A_9_if_full_n,
    output wire                                          fifo_A_9_if_read,
    output wire                                          fifo_A_9_if_read_ce,
    output wire                                          fifo_A_9_if_write,
    output wire                                          fifo_A_9_if_write_ce,
    output wire                                          fifo_A_9_reset,
    output wire                                          fifo_X_pe_0_clk,
    output wire [                                 512:0] fifo_X_pe_0_if_din,
    input wire  [                                 512:0] fifo_X_pe_0_if_dout,
    input wire                                           fifo_X_pe_0_if_empty_n,
    input wire                                           fifo_X_pe_0_if_full_n,
    output wire                                          fifo_X_pe_0_if_read,
    output wire                                          fifo_X_pe_0_if_read_ce,
    output wire                                          fifo_X_pe_0_if_write,
    output wire                                          fifo_X_pe_0_if_write_ce,
    output wire                                          fifo_X_pe_0_reset,
    output wire                                          fifo_X_pe_10_clk,
    output wire [                                 512:0] fifo_X_pe_10_if_din,
    input wire  [                                 512:0] fifo_X_pe_10_if_dout,
    input wire                                           fifo_X_pe_10_if_empty_n,
    input wire                                           fifo_X_pe_10_if_full_n,
    output wire                                          fifo_X_pe_10_if_read,
    output wire                                          fifo_X_pe_10_if_read_ce,
    output wire                                          fifo_X_pe_10_if_write,
    output wire                                          fifo_X_pe_10_if_write_ce,
    output wire                                          fifo_X_pe_10_reset,
    output wire                                          fifo_X_pe_11_clk,
    output wire [                                 512:0] fifo_X_pe_11_if_din,
    input wire  [                                 512:0] fifo_X_pe_11_if_dout,
    input wire                                           fifo_X_pe_11_if_empty_n,
    input wire                                           fifo_X_pe_11_if_full_n,
    output wire                                          fifo_X_pe_11_if_read,
    output wire                                          fifo_X_pe_11_if_read_ce,
    output wire                                          fifo_X_pe_11_if_write,
    output wire                                          fifo_X_pe_11_if_write_ce,
    output wire                                          fifo_X_pe_11_reset,
    output wire                                          fifo_X_pe_12_clk,
    output wire [                                 512:0] fifo_X_pe_12_if_din,
    input wire  [                                 512:0] fifo_X_pe_12_if_dout,
    input wire                                           fifo_X_pe_12_if_empty_n,
    input wire                                           fifo_X_pe_12_if_full_n,
    output wire                                          fifo_X_pe_12_if_read,
    output wire                                          fifo_X_pe_12_if_read_ce,
    output wire                                          fifo_X_pe_12_if_write,
    output wire                                          fifo_X_pe_12_if_write_ce,
    output wire                                          fifo_X_pe_12_reset,
    output wire                                          fifo_X_pe_13_clk,
    output wire [                                 512:0] fifo_X_pe_13_if_din,
    input wire  [                                 512:0] fifo_X_pe_13_if_dout,
    input wire                                           fifo_X_pe_13_if_empty_n,
    input wire                                           fifo_X_pe_13_if_full_n,
    output wire                                          fifo_X_pe_13_if_read,
    output wire                                          fifo_X_pe_13_if_read_ce,
    output wire                                          fifo_X_pe_13_if_write,
    output wire                                          fifo_X_pe_13_if_write_ce,
    output wire                                          fifo_X_pe_13_reset,
    output wire                                          fifo_X_pe_14_clk,
    output wire [                                 512:0] fifo_X_pe_14_if_din,
    input wire  [                                 512:0] fifo_X_pe_14_if_dout,
    input wire                                           fifo_X_pe_14_if_empty_n,
    input wire                                           fifo_X_pe_14_if_full_n,
    output wire                                          fifo_X_pe_14_if_read,
    output wire                                          fifo_X_pe_14_if_read_ce,
    output wire                                          fifo_X_pe_14_if_write,
    output wire                                          fifo_X_pe_14_if_write_ce,
    output wire                                          fifo_X_pe_14_reset,
    output wire                                          fifo_X_pe_15_clk,
    output wire [                                 512:0] fifo_X_pe_15_if_din,
    input wire  [                                 512:0] fifo_X_pe_15_if_dout,
    input wire                                           fifo_X_pe_15_if_empty_n,
    input wire                                           fifo_X_pe_15_if_full_n,
    output wire                                          fifo_X_pe_15_if_read,
    output wire                                          fifo_X_pe_15_if_read_ce,
    output wire                                          fifo_X_pe_15_if_write,
    output wire                                          fifo_X_pe_15_if_write_ce,
    output wire                                          fifo_X_pe_15_reset,
    output wire                                          fifo_X_pe_16_clk,
    output wire [                                 512:0] fifo_X_pe_16_if_din,
    input wire  [                                 512:0] fifo_X_pe_16_if_dout,
    input wire                                           fifo_X_pe_16_if_empty_n,
    input wire                                           fifo_X_pe_16_if_full_n,
    output wire                                          fifo_X_pe_16_if_read,
    output wire                                          fifo_X_pe_16_if_read_ce,
    output wire                                          fifo_X_pe_16_if_write,
    output wire                                          fifo_X_pe_16_if_write_ce,
    output wire                                          fifo_X_pe_16_reset,
    output wire                                          fifo_X_pe_17_clk,
    output wire [                                 512:0] fifo_X_pe_17_if_din,
    input wire  [                                 512:0] fifo_X_pe_17_if_dout,
    input wire                                           fifo_X_pe_17_if_empty_n,
    input wire                                           fifo_X_pe_17_if_full_n,
    output wire                                          fifo_X_pe_17_if_read,
    output wire                                          fifo_X_pe_17_if_read_ce,
    output wire                                          fifo_X_pe_17_if_write,
    output wire                                          fifo_X_pe_17_if_write_ce,
    output wire                                          fifo_X_pe_17_reset,
    output wire                                          fifo_X_pe_18_clk,
    output wire [                                 512:0] fifo_X_pe_18_if_din,
    input wire  [                                 512:0] fifo_X_pe_18_if_dout,
    input wire                                           fifo_X_pe_18_if_empty_n,
    input wire                                           fifo_X_pe_18_if_full_n,
    output wire                                          fifo_X_pe_18_if_read,
    output wire                                          fifo_X_pe_18_if_read_ce,
    output wire                                          fifo_X_pe_18_if_write,
    output wire                                          fifo_X_pe_18_if_write_ce,
    output wire                                          fifo_X_pe_18_reset,
    output wire                                          fifo_X_pe_19_clk,
    output wire [                                 512:0] fifo_X_pe_19_if_din,
    input wire  [                                 512:0] fifo_X_pe_19_if_dout,
    input wire                                           fifo_X_pe_19_if_empty_n,
    input wire                                           fifo_X_pe_19_if_full_n,
    output wire                                          fifo_X_pe_19_if_read,
    output wire                                          fifo_X_pe_19_if_read_ce,
    output wire                                          fifo_X_pe_19_if_write,
    output wire                                          fifo_X_pe_19_if_write_ce,
    output wire                                          fifo_X_pe_19_reset,
    output wire                                          fifo_X_pe_1_clk,
    output wire [                                 512:0] fifo_X_pe_1_if_din,
    input wire  [                                 512:0] fifo_X_pe_1_if_dout,
    input wire                                           fifo_X_pe_1_if_empty_n,
    input wire                                           fifo_X_pe_1_if_full_n,
    output wire                                          fifo_X_pe_1_if_read,
    output wire                                          fifo_X_pe_1_if_read_ce,
    output wire                                          fifo_X_pe_1_if_write,
    output wire                                          fifo_X_pe_1_if_write_ce,
    output wire                                          fifo_X_pe_1_reset,
    output wire                                          fifo_X_pe_20_clk,
    output wire [                                 512:0] fifo_X_pe_20_if_din,
    input wire  [                                 512:0] fifo_X_pe_20_if_dout,
    input wire                                           fifo_X_pe_20_if_empty_n,
    input wire                                           fifo_X_pe_20_if_full_n,
    output wire                                          fifo_X_pe_20_if_read,
    output wire                                          fifo_X_pe_20_if_read_ce,
    output wire                                          fifo_X_pe_20_if_write,
    output wire                                          fifo_X_pe_20_if_write_ce,
    output wire                                          fifo_X_pe_20_reset,
    output wire                                          fifo_X_pe_21_clk,
    output wire [                                 512:0] fifo_X_pe_21_if_din,
    input wire  [                                 512:0] fifo_X_pe_21_if_dout,
    input wire                                           fifo_X_pe_21_if_empty_n,
    input wire                                           fifo_X_pe_21_if_full_n,
    output wire                                          fifo_X_pe_21_if_read,
    output wire                                          fifo_X_pe_21_if_read_ce,
    output wire                                          fifo_X_pe_21_if_write,
    output wire                                          fifo_X_pe_21_if_write_ce,
    output wire                                          fifo_X_pe_21_reset,
    output wire                                          fifo_X_pe_22_clk,
    output wire [                                 512:0] fifo_X_pe_22_if_din,
    input wire  [                                 512:0] fifo_X_pe_22_if_dout,
    input wire                                           fifo_X_pe_22_if_empty_n,
    input wire                                           fifo_X_pe_22_if_full_n,
    output wire                                          fifo_X_pe_22_if_read,
    output wire                                          fifo_X_pe_22_if_read_ce,
    output wire                                          fifo_X_pe_22_if_write,
    output wire                                          fifo_X_pe_22_if_write_ce,
    output wire                                          fifo_X_pe_22_reset,
    output wire                                          fifo_X_pe_23_clk,
    output wire [                                 512:0] fifo_X_pe_23_if_din,
    input wire  [                                 512:0] fifo_X_pe_23_if_dout,
    input wire                                           fifo_X_pe_23_if_empty_n,
    input wire                                           fifo_X_pe_23_if_full_n,
    output wire                                          fifo_X_pe_23_if_read,
    output wire                                          fifo_X_pe_23_if_read_ce,
    output wire                                          fifo_X_pe_23_if_write,
    output wire                                          fifo_X_pe_23_if_write_ce,
    output wire                                          fifo_X_pe_23_reset,
    output wire                                          fifo_X_pe_24_clk,
    output wire [                                 512:0] fifo_X_pe_24_if_din,
    input wire  [                                 512:0] fifo_X_pe_24_if_dout,
    input wire                                           fifo_X_pe_24_if_empty_n,
    input wire                                           fifo_X_pe_24_if_full_n,
    output wire                                          fifo_X_pe_24_if_read,
    output wire                                          fifo_X_pe_24_if_read_ce,
    output wire                                          fifo_X_pe_24_if_write,
    output wire                                          fifo_X_pe_24_if_write_ce,
    output wire                                          fifo_X_pe_24_reset,
    output wire                                          fifo_X_pe_25_clk,
    output wire [                                 512:0] fifo_X_pe_25_if_din,
    input wire  [                                 512:0] fifo_X_pe_25_if_dout,
    input wire                                           fifo_X_pe_25_if_empty_n,
    input wire                                           fifo_X_pe_25_if_full_n,
    output wire                                          fifo_X_pe_25_if_read,
    output wire                                          fifo_X_pe_25_if_read_ce,
    output wire                                          fifo_X_pe_25_if_write,
    output wire                                          fifo_X_pe_25_if_write_ce,
    output wire                                          fifo_X_pe_25_reset,
    output wire                                          fifo_X_pe_26_clk,
    output wire [                                 512:0] fifo_X_pe_26_if_din,
    input wire  [                                 512:0] fifo_X_pe_26_if_dout,
    input wire                                           fifo_X_pe_26_if_empty_n,
    input wire                                           fifo_X_pe_26_if_full_n,
    output wire                                          fifo_X_pe_26_if_read,
    output wire                                          fifo_X_pe_26_if_read_ce,
    output wire                                          fifo_X_pe_26_if_write,
    output wire                                          fifo_X_pe_26_if_write_ce,
    output wire                                          fifo_X_pe_26_reset,
    output wire                                          fifo_X_pe_27_clk,
    output wire [                                 512:0] fifo_X_pe_27_if_din,
    input wire  [                                 512:0] fifo_X_pe_27_if_dout,
    input wire                                           fifo_X_pe_27_if_empty_n,
    input wire                                           fifo_X_pe_27_if_full_n,
    output wire                                          fifo_X_pe_27_if_read,
    output wire                                          fifo_X_pe_27_if_read_ce,
    output wire                                          fifo_X_pe_27_if_write,
    output wire                                          fifo_X_pe_27_if_write_ce,
    output wire                                          fifo_X_pe_27_reset,
    output wire                                          fifo_X_pe_28_clk,
    output wire [                                 512:0] fifo_X_pe_28_if_din,
    input wire  [                                 512:0] fifo_X_pe_28_if_dout,
    input wire                                           fifo_X_pe_28_if_empty_n,
    input wire                                           fifo_X_pe_28_if_full_n,
    output wire                                          fifo_X_pe_28_if_read,
    output wire                                          fifo_X_pe_28_if_read_ce,
    output wire                                          fifo_X_pe_28_if_write,
    output wire                                          fifo_X_pe_28_if_write_ce,
    output wire                                          fifo_X_pe_28_reset,
    output wire                                          fifo_X_pe_29_clk,
    output wire [                                 512:0] fifo_X_pe_29_if_din,
    input wire  [                                 512:0] fifo_X_pe_29_if_dout,
    input wire                                           fifo_X_pe_29_if_empty_n,
    input wire                                           fifo_X_pe_29_if_full_n,
    output wire                                          fifo_X_pe_29_if_read,
    output wire                                          fifo_X_pe_29_if_read_ce,
    output wire                                          fifo_X_pe_29_if_write,
    output wire                                          fifo_X_pe_29_if_write_ce,
    output wire                                          fifo_X_pe_29_reset,
    output wire                                          fifo_X_pe_2_clk,
    output wire [                                 512:0] fifo_X_pe_2_if_din,
    input wire  [                                 512:0] fifo_X_pe_2_if_dout,
    input wire                                           fifo_X_pe_2_if_empty_n,
    input wire                                           fifo_X_pe_2_if_full_n,
    output wire                                          fifo_X_pe_2_if_read,
    output wire                                          fifo_X_pe_2_if_read_ce,
    output wire                                          fifo_X_pe_2_if_write,
    output wire                                          fifo_X_pe_2_if_write_ce,
    output wire                                          fifo_X_pe_2_reset,
    output wire                                          fifo_X_pe_30_clk,
    output wire [                                 512:0] fifo_X_pe_30_if_din,
    input wire  [                                 512:0] fifo_X_pe_30_if_dout,
    input wire                                           fifo_X_pe_30_if_empty_n,
    input wire                                           fifo_X_pe_30_if_full_n,
    output wire                                          fifo_X_pe_30_if_read,
    output wire                                          fifo_X_pe_30_if_read_ce,
    output wire                                          fifo_X_pe_30_if_write,
    output wire                                          fifo_X_pe_30_if_write_ce,
    output wire                                          fifo_X_pe_30_reset,
    output wire                                          fifo_X_pe_31_clk,
    output wire [                                 512:0] fifo_X_pe_31_if_din,
    input wire  [                                 512:0] fifo_X_pe_31_if_dout,
    input wire                                           fifo_X_pe_31_if_empty_n,
    input wire                                           fifo_X_pe_31_if_full_n,
    output wire                                          fifo_X_pe_31_if_read,
    output wire                                          fifo_X_pe_31_if_read_ce,
    output wire                                          fifo_X_pe_31_if_write,
    output wire                                          fifo_X_pe_31_if_write_ce,
    output wire                                          fifo_X_pe_31_reset,
    output wire                                          fifo_X_pe_32_clk,
    output wire [                                 512:0] fifo_X_pe_32_if_din,
    input wire  [                                 512:0] fifo_X_pe_32_if_dout,
    input wire                                           fifo_X_pe_32_if_empty_n,
    input wire                                           fifo_X_pe_32_if_full_n,
    output wire                                          fifo_X_pe_32_if_read,
    output wire                                          fifo_X_pe_32_if_read_ce,
    output wire                                          fifo_X_pe_32_if_write,
    output wire                                          fifo_X_pe_32_if_write_ce,
    output wire                                          fifo_X_pe_32_reset,
    output wire                                          fifo_X_pe_33_clk,
    output wire [                                 512:0] fifo_X_pe_33_if_din,
    input wire  [                                 512:0] fifo_X_pe_33_if_dout,
    input wire                                           fifo_X_pe_33_if_empty_n,
    input wire                                           fifo_X_pe_33_if_full_n,
    output wire                                          fifo_X_pe_33_if_read,
    output wire                                          fifo_X_pe_33_if_read_ce,
    output wire                                          fifo_X_pe_33_if_write,
    output wire                                          fifo_X_pe_33_if_write_ce,
    output wire                                          fifo_X_pe_33_reset,
    output wire                                          fifo_X_pe_34_clk,
    output wire [                                 512:0] fifo_X_pe_34_if_din,
    input wire  [                                 512:0] fifo_X_pe_34_if_dout,
    input wire                                           fifo_X_pe_34_if_empty_n,
    input wire                                           fifo_X_pe_34_if_full_n,
    output wire                                          fifo_X_pe_34_if_read,
    output wire                                          fifo_X_pe_34_if_read_ce,
    output wire                                          fifo_X_pe_34_if_write,
    output wire                                          fifo_X_pe_34_if_write_ce,
    output wire                                          fifo_X_pe_34_reset,
    output wire                                          fifo_X_pe_35_clk,
    output wire [                                 512:0] fifo_X_pe_35_if_din,
    input wire  [                                 512:0] fifo_X_pe_35_if_dout,
    input wire                                           fifo_X_pe_35_if_empty_n,
    input wire                                           fifo_X_pe_35_if_full_n,
    output wire                                          fifo_X_pe_35_if_read,
    output wire                                          fifo_X_pe_35_if_read_ce,
    output wire                                          fifo_X_pe_35_if_write,
    output wire                                          fifo_X_pe_35_if_write_ce,
    output wire                                          fifo_X_pe_35_reset,
    output wire                                          fifo_X_pe_36_clk,
    output wire [                                 512:0] fifo_X_pe_36_if_din,
    input wire  [                                 512:0] fifo_X_pe_36_if_dout,
    input wire                                           fifo_X_pe_36_if_empty_n,
    input wire                                           fifo_X_pe_36_if_full_n,
    output wire                                          fifo_X_pe_36_if_read,
    output wire                                          fifo_X_pe_36_if_read_ce,
    output wire                                          fifo_X_pe_36_if_write,
    output wire                                          fifo_X_pe_36_if_write_ce,
    output wire                                          fifo_X_pe_36_reset,
    output wire                                          fifo_X_pe_37_clk,
    output wire [                                 512:0] fifo_X_pe_37_if_din,
    input wire  [                                 512:0] fifo_X_pe_37_if_dout,
    input wire                                           fifo_X_pe_37_if_empty_n,
    input wire                                           fifo_X_pe_37_if_full_n,
    output wire                                          fifo_X_pe_37_if_read,
    output wire                                          fifo_X_pe_37_if_read_ce,
    output wire                                          fifo_X_pe_37_if_write,
    output wire                                          fifo_X_pe_37_if_write_ce,
    output wire                                          fifo_X_pe_37_reset,
    output wire                                          fifo_X_pe_38_clk,
    output wire [                                 512:0] fifo_X_pe_38_if_din,
    input wire  [                                 512:0] fifo_X_pe_38_if_dout,
    input wire                                           fifo_X_pe_38_if_empty_n,
    input wire                                           fifo_X_pe_38_if_full_n,
    output wire                                          fifo_X_pe_38_if_read,
    output wire                                          fifo_X_pe_38_if_read_ce,
    output wire                                          fifo_X_pe_38_if_write,
    output wire                                          fifo_X_pe_38_if_write_ce,
    output wire                                          fifo_X_pe_38_reset,
    output wire                                          fifo_X_pe_39_clk,
    output wire [                                 512:0] fifo_X_pe_39_if_din,
    input wire  [                                 512:0] fifo_X_pe_39_if_dout,
    input wire                                           fifo_X_pe_39_if_empty_n,
    input wire                                           fifo_X_pe_39_if_full_n,
    output wire                                          fifo_X_pe_39_if_read,
    output wire                                          fifo_X_pe_39_if_read_ce,
    output wire                                          fifo_X_pe_39_if_write,
    output wire                                          fifo_X_pe_39_if_write_ce,
    output wire                                          fifo_X_pe_39_reset,
    output wire                                          fifo_X_pe_3_clk,
    output wire [                                 512:0] fifo_X_pe_3_if_din,
    input wire  [                                 512:0] fifo_X_pe_3_if_dout,
    input wire                                           fifo_X_pe_3_if_empty_n,
    input wire                                           fifo_X_pe_3_if_full_n,
    output wire                                          fifo_X_pe_3_if_read,
    output wire                                          fifo_X_pe_3_if_read_ce,
    output wire                                          fifo_X_pe_3_if_write,
    output wire                                          fifo_X_pe_3_if_write_ce,
    output wire                                          fifo_X_pe_3_reset,
    output wire                                          fifo_X_pe_40_clk,
    output wire [                                 512:0] fifo_X_pe_40_if_din,
    input wire  [                                 512:0] fifo_X_pe_40_if_dout,
    input wire                                           fifo_X_pe_40_if_empty_n,
    input wire                                           fifo_X_pe_40_if_full_n,
    output wire                                          fifo_X_pe_40_if_read,
    output wire                                          fifo_X_pe_40_if_read_ce,
    output wire                                          fifo_X_pe_40_if_write,
    output wire                                          fifo_X_pe_40_if_write_ce,
    output wire                                          fifo_X_pe_40_reset,
    output wire                                          fifo_X_pe_41_clk,
    output wire [                                 512:0] fifo_X_pe_41_if_din,
    input wire  [                                 512:0] fifo_X_pe_41_if_dout,
    input wire                                           fifo_X_pe_41_if_empty_n,
    input wire                                           fifo_X_pe_41_if_full_n,
    output wire                                          fifo_X_pe_41_if_read,
    output wire                                          fifo_X_pe_41_if_read_ce,
    output wire                                          fifo_X_pe_41_if_write,
    output wire                                          fifo_X_pe_41_if_write_ce,
    output wire                                          fifo_X_pe_41_reset,
    output wire                                          fifo_X_pe_42_clk,
    output wire [                                 512:0] fifo_X_pe_42_if_din,
    input wire  [                                 512:0] fifo_X_pe_42_if_dout,
    input wire                                           fifo_X_pe_42_if_empty_n,
    input wire                                           fifo_X_pe_42_if_full_n,
    output wire                                          fifo_X_pe_42_if_read,
    output wire                                          fifo_X_pe_42_if_read_ce,
    output wire                                          fifo_X_pe_42_if_write,
    output wire                                          fifo_X_pe_42_if_write_ce,
    output wire                                          fifo_X_pe_42_reset,
    output wire                                          fifo_X_pe_43_clk,
    output wire [                                 512:0] fifo_X_pe_43_if_din,
    input wire  [                                 512:0] fifo_X_pe_43_if_dout,
    input wire                                           fifo_X_pe_43_if_empty_n,
    input wire                                           fifo_X_pe_43_if_full_n,
    output wire                                          fifo_X_pe_43_if_read,
    output wire                                          fifo_X_pe_43_if_read_ce,
    output wire                                          fifo_X_pe_43_if_write,
    output wire                                          fifo_X_pe_43_if_write_ce,
    output wire                                          fifo_X_pe_43_reset,
    output wire                                          fifo_X_pe_44_clk,
    output wire [                                 512:0] fifo_X_pe_44_if_din,
    input wire  [                                 512:0] fifo_X_pe_44_if_dout,
    input wire                                           fifo_X_pe_44_if_empty_n,
    input wire                                           fifo_X_pe_44_if_full_n,
    output wire                                          fifo_X_pe_44_if_read,
    output wire                                          fifo_X_pe_44_if_read_ce,
    output wire                                          fifo_X_pe_44_if_write,
    output wire                                          fifo_X_pe_44_if_write_ce,
    output wire                                          fifo_X_pe_44_reset,
    output wire                                          fifo_X_pe_45_clk,
    output wire [                                 512:0] fifo_X_pe_45_if_din,
    input wire  [                                 512:0] fifo_X_pe_45_if_dout,
    input wire                                           fifo_X_pe_45_if_empty_n,
    input wire                                           fifo_X_pe_45_if_full_n,
    output wire                                          fifo_X_pe_45_if_read,
    output wire                                          fifo_X_pe_45_if_read_ce,
    output wire                                          fifo_X_pe_45_if_write,
    output wire                                          fifo_X_pe_45_if_write_ce,
    output wire                                          fifo_X_pe_45_reset,
    output wire                                          fifo_X_pe_46_clk,
    output wire [                                 512:0] fifo_X_pe_46_if_din,
    input wire  [                                 512:0] fifo_X_pe_46_if_dout,
    input wire                                           fifo_X_pe_46_if_empty_n,
    input wire                                           fifo_X_pe_46_if_full_n,
    output wire                                          fifo_X_pe_46_if_read,
    output wire                                          fifo_X_pe_46_if_read_ce,
    output wire                                          fifo_X_pe_46_if_write,
    output wire                                          fifo_X_pe_46_if_write_ce,
    output wire                                          fifo_X_pe_46_reset,
    output wire                                          fifo_X_pe_47_clk,
    output wire [                                 512:0] fifo_X_pe_47_if_din,
    input wire  [                                 512:0] fifo_X_pe_47_if_dout,
    input wire                                           fifo_X_pe_47_if_empty_n,
    input wire                                           fifo_X_pe_47_if_full_n,
    output wire                                          fifo_X_pe_47_if_read,
    output wire                                          fifo_X_pe_47_if_read_ce,
    output wire                                          fifo_X_pe_47_if_write,
    output wire                                          fifo_X_pe_47_if_write_ce,
    output wire                                          fifo_X_pe_47_reset,
    output wire                                          fifo_X_pe_48_clk,
    output wire [                                 512:0] fifo_X_pe_48_if_din,
    input wire  [                                 512:0] fifo_X_pe_48_if_dout,
    input wire                                           fifo_X_pe_48_if_empty_n,
    input wire                                           fifo_X_pe_48_if_full_n,
    output wire                                          fifo_X_pe_48_if_read,
    output wire                                          fifo_X_pe_48_if_read_ce,
    output wire                                          fifo_X_pe_48_if_write,
    output wire                                          fifo_X_pe_48_if_write_ce,
    output wire                                          fifo_X_pe_48_reset,
    output wire                                          fifo_X_pe_4_clk,
    output wire [                                 512:0] fifo_X_pe_4_if_din,
    input wire  [                                 512:0] fifo_X_pe_4_if_dout,
    input wire                                           fifo_X_pe_4_if_empty_n,
    input wire                                           fifo_X_pe_4_if_full_n,
    output wire                                          fifo_X_pe_4_if_read,
    output wire                                          fifo_X_pe_4_if_read_ce,
    output wire                                          fifo_X_pe_4_if_write,
    output wire                                          fifo_X_pe_4_if_write_ce,
    output wire                                          fifo_X_pe_4_reset,
    output wire                                          fifo_X_pe_5_clk,
    output wire [                                 512:0] fifo_X_pe_5_if_din,
    input wire  [                                 512:0] fifo_X_pe_5_if_dout,
    input wire                                           fifo_X_pe_5_if_empty_n,
    input wire                                           fifo_X_pe_5_if_full_n,
    output wire                                          fifo_X_pe_5_if_read,
    output wire                                          fifo_X_pe_5_if_read_ce,
    output wire                                          fifo_X_pe_5_if_write,
    output wire                                          fifo_X_pe_5_if_write_ce,
    output wire                                          fifo_X_pe_5_reset,
    output wire                                          fifo_X_pe_6_clk,
    output wire [                                 512:0] fifo_X_pe_6_if_din,
    input wire  [                                 512:0] fifo_X_pe_6_if_dout,
    input wire                                           fifo_X_pe_6_if_empty_n,
    input wire                                           fifo_X_pe_6_if_full_n,
    output wire                                          fifo_X_pe_6_if_read,
    output wire                                          fifo_X_pe_6_if_read_ce,
    output wire                                          fifo_X_pe_6_if_write,
    output wire                                          fifo_X_pe_6_if_write_ce,
    output wire                                          fifo_X_pe_6_reset,
    output wire                                          fifo_X_pe_7_clk,
    output wire [                                 512:0] fifo_X_pe_7_if_din,
    input wire  [                                 512:0] fifo_X_pe_7_if_dout,
    input wire                                           fifo_X_pe_7_if_empty_n,
    input wire                                           fifo_X_pe_7_if_full_n,
    output wire                                          fifo_X_pe_7_if_read,
    output wire                                          fifo_X_pe_7_if_read_ce,
    output wire                                          fifo_X_pe_7_if_write,
    output wire                                          fifo_X_pe_7_if_write_ce,
    output wire                                          fifo_X_pe_7_reset,
    output wire                                          fifo_X_pe_8_clk,
    output wire [                                 512:0] fifo_X_pe_8_if_din,
    input wire  [                                 512:0] fifo_X_pe_8_if_dout,
    input wire                                           fifo_X_pe_8_if_empty_n,
    input wire                                           fifo_X_pe_8_if_full_n,
    output wire                                          fifo_X_pe_8_if_read,
    output wire                                          fifo_X_pe_8_if_read_ce,
    output wire                                          fifo_X_pe_8_if_write,
    output wire                                          fifo_X_pe_8_if_write_ce,
    output wire                                          fifo_X_pe_8_reset,
    output wire                                          fifo_X_pe_9_clk,
    output wire [                                 512:0] fifo_X_pe_9_if_din,
    input wire  [                                 512:0] fifo_X_pe_9_if_dout,
    input wire                                           fifo_X_pe_9_if_empty_n,
    input wire                                           fifo_X_pe_9_if_full_n,
    output wire                                          fifo_X_pe_9_if_read,
    output wire                                          fifo_X_pe_9_if_read_ce,
    output wire                                          fifo_X_pe_9_if_write,
    output wire                                          fifo_X_pe_9_if_write_ce,
    output wire                                          fifo_X_pe_9_reset,
    output wire                                          fifo_Y_AX_clk,
    output wire [                                 512:0] fifo_Y_AX_if_din,
    input wire  [                                 512:0] fifo_Y_AX_if_dout,
    input wire                                           fifo_Y_AX_if_empty_n,
    input wire                                           fifo_Y_AX_if_full_n,
    output wire                                          fifo_Y_AX_if_read,
    output wire                                          fifo_Y_AX_if_read_ce,
    output wire                                          fifo_Y_AX_if_write,
    output wire                                          fifo_Y_AX_if_write_ce,
    output wire                                          fifo_Y_AX_reset,
    output wire                                          fifo_Y_alpha_AX_clk,
    output wire [                                 512:0] fifo_Y_alpha_AX_if_din,
    input wire  [                                 512:0] fifo_Y_alpha_AX_if_dout,
    input wire                                           fifo_Y_alpha_AX_if_empty_n,
    input wire                                           fifo_Y_alpha_AX_if_full_n,
    output wire                                          fifo_Y_alpha_AX_if_read,
    output wire                                          fifo_Y_alpha_AX_if_read_ce,
    output wire                                          fifo_Y_alpha_AX_if_write,
    output wire                                          fifo_Y_alpha_AX_if_write_ce,
    output wire                                          fifo_Y_alpha_AX_reset,
    output wire                                          fifo_Y_in_clk,
    output wire [                                 512:0] fifo_Y_in_if_din,
    input wire  [                                 512:0] fifo_Y_in_if_dout,
    input wire                                           fifo_Y_in_if_empty_n,
    input wire                                           fifo_Y_in_if_full_n,
    output wire                                          fifo_Y_in_if_read,
    output wire                                          fifo_Y_in_if_read_ce,
    output wire                                          fifo_Y_in_if_write,
    output wire                                          fifo_Y_in_if_write_ce,
    output wire                                          fifo_Y_in_reset,
    output wire                                          fifo_Y_in_beta_clk,
    output wire [                                 512:0] fifo_Y_in_beta_if_din,
    input wire  [                                 512:0] fifo_Y_in_beta_if_dout,
    input wire                                           fifo_Y_in_beta_if_empty_n,
    input wire                                           fifo_Y_in_beta_if_full_n,
    output wire                                          fifo_Y_in_beta_if_read,
    output wire                                          fifo_Y_in_beta_if_read_ce,
    output wire                                          fifo_Y_in_beta_if_write,
    output wire                                          fifo_Y_in_beta_if_write_ce,
    output wire                                          fifo_Y_in_beta_reset,
    output wire                                          fifo_Y_out_clk,
    output wire [                                 512:0] fifo_Y_out_if_din,
    input wire  [                                 512:0] fifo_Y_out_if_dout,
    input wire                                           fifo_Y_out_if_empty_n,
    input wire                                           fifo_Y_out_if_full_n,
    output wire                                          fifo_Y_out_if_read,
    output wire                                          fifo_Y_out_if_read_ce,
    output wire                                          fifo_Y_out_if_write,
    output wire                                          fifo_Y_out_if_write_ce,
    output wire                                          fifo_Y_out_reset,
    output wire                                          fifo_Y_pe_0_clk,
    output wire [                                  64:0] fifo_Y_pe_0_if_din,
    input wire  [                                  64:0] fifo_Y_pe_0_if_dout,
    input wire                                           fifo_Y_pe_0_if_empty_n,
    input wire                                           fifo_Y_pe_0_if_full_n,
    output wire                                          fifo_Y_pe_0_if_read,
    output wire                                          fifo_Y_pe_0_if_read_ce,
    output wire                                          fifo_Y_pe_0_if_write,
    output wire                                          fifo_Y_pe_0_if_write_ce,
    output wire                                          fifo_Y_pe_0_reset,
    output wire                                          fifo_Y_pe_10_clk,
    output wire [                                  64:0] fifo_Y_pe_10_if_din,
    input wire  [                                  64:0] fifo_Y_pe_10_if_dout,
    input wire                                           fifo_Y_pe_10_if_empty_n,
    input wire                                           fifo_Y_pe_10_if_full_n,
    output wire                                          fifo_Y_pe_10_if_read,
    output wire                                          fifo_Y_pe_10_if_read_ce,
    output wire                                          fifo_Y_pe_10_if_write,
    output wire                                          fifo_Y_pe_10_if_write_ce,
    output wire                                          fifo_Y_pe_10_reset,
    output wire                                          fifo_Y_pe_11_clk,
    output wire [                                  64:0] fifo_Y_pe_11_if_din,
    input wire  [                                  64:0] fifo_Y_pe_11_if_dout,
    input wire                                           fifo_Y_pe_11_if_empty_n,
    input wire                                           fifo_Y_pe_11_if_full_n,
    output wire                                          fifo_Y_pe_11_if_read,
    output wire                                          fifo_Y_pe_11_if_read_ce,
    output wire                                          fifo_Y_pe_11_if_write,
    output wire                                          fifo_Y_pe_11_if_write_ce,
    output wire                                          fifo_Y_pe_11_reset,
    output wire                                          fifo_Y_pe_12_clk,
    output wire [                                  64:0] fifo_Y_pe_12_if_din,
    input wire  [                                  64:0] fifo_Y_pe_12_if_dout,
    input wire                                           fifo_Y_pe_12_if_empty_n,
    input wire                                           fifo_Y_pe_12_if_full_n,
    output wire                                          fifo_Y_pe_12_if_read,
    output wire                                          fifo_Y_pe_12_if_read_ce,
    output wire                                          fifo_Y_pe_12_if_write,
    output wire                                          fifo_Y_pe_12_if_write_ce,
    output wire                                          fifo_Y_pe_12_reset,
    output wire                                          fifo_Y_pe_13_clk,
    output wire [                                  64:0] fifo_Y_pe_13_if_din,
    input wire  [                                  64:0] fifo_Y_pe_13_if_dout,
    input wire                                           fifo_Y_pe_13_if_empty_n,
    input wire                                           fifo_Y_pe_13_if_full_n,
    output wire                                          fifo_Y_pe_13_if_read,
    output wire                                          fifo_Y_pe_13_if_read_ce,
    output wire                                          fifo_Y_pe_13_if_write,
    output wire                                          fifo_Y_pe_13_if_write_ce,
    output wire                                          fifo_Y_pe_13_reset,
    output wire                                          fifo_Y_pe_14_clk,
    output wire [                                  64:0] fifo_Y_pe_14_if_din,
    input wire  [                                  64:0] fifo_Y_pe_14_if_dout,
    input wire                                           fifo_Y_pe_14_if_empty_n,
    input wire                                           fifo_Y_pe_14_if_full_n,
    output wire                                          fifo_Y_pe_14_if_read,
    output wire                                          fifo_Y_pe_14_if_read_ce,
    output wire                                          fifo_Y_pe_14_if_write,
    output wire                                          fifo_Y_pe_14_if_write_ce,
    output wire                                          fifo_Y_pe_14_reset,
    output wire                                          fifo_Y_pe_15_clk,
    output wire [                                  64:0] fifo_Y_pe_15_if_din,
    input wire  [                                  64:0] fifo_Y_pe_15_if_dout,
    input wire                                           fifo_Y_pe_15_if_empty_n,
    input wire                                           fifo_Y_pe_15_if_full_n,
    output wire                                          fifo_Y_pe_15_if_read,
    output wire                                          fifo_Y_pe_15_if_read_ce,
    output wire                                          fifo_Y_pe_15_if_write,
    output wire                                          fifo_Y_pe_15_if_write_ce,
    output wire                                          fifo_Y_pe_15_reset,
    output wire                                          fifo_Y_pe_16_clk,
    output wire [                                  64:0] fifo_Y_pe_16_if_din,
    input wire  [                                  64:0] fifo_Y_pe_16_if_dout,
    input wire                                           fifo_Y_pe_16_if_empty_n,
    input wire                                           fifo_Y_pe_16_if_full_n,
    output wire                                          fifo_Y_pe_16_if_read,
    output wire                                          fifo_Y_pe_16_if_read_ce,
    output wire                                          fifo_Y_pe_16_if_write,
    output wire                                          fifo_Y_pe_16_if_write_ce,
    output wire                                          fifo_Y_pe_16_reset,
    output wire                                          fifo_Y_pe_17_clk,
    output wire [                                  64:0] fifo_Y_pe_17_if_din,
    input wire  [                                  64:0] fifo_Y_pe_17_if_dout,
    input wire                                           fifo_Y_pe_17_if_empty_n,
    input wire                                           fifo_Y_pe_17_if_full_n,
    output wire                                          fifo_Y_pe_17_if_read,
    output wire                                          fifo_Y_pe_17_if_read_ce,
    output wire                                          fifo_Y_pe_17_if_write,
    output wire                                          fifo_Y_pe_17_if_write_ce,
    output wire                                          fifo_Y_pe_17_reset,
    output wire                                          fifo_Y_pe_18_clk,
    output wire [                                  64:0] fifo_Y_pe_18_if_din,
    input wire  [                                  64:0] fifo_Y_pe_18_if_dout,
    input wire                                           fifo_Y_pe_18_if_empty_n,
    input wire                                           fifo_Y_pe_18_if_full_n,
    output wire                                          fifo_Y_pe_18_if_read,
    output wire                                          fifo_Y_pe_18_if_read_ce,
    output wire                                          fifo_Y_pe_18_if_write,
    output wire                                          fifo_Y_pe_18_if_write_ce,
    output wire                                          fifo_Y_pe_18_reset,
    output wire                                          fifo_Y_pe_19_clk,
    output wire [                                  64:0] fifo_Y_pe_19_if_din,
    input wire  [                                  64:0] fifo_Y_pe_19_if_dout,
    input wire                                           fifo_Y_pe_19_if_empty_n,
    input wire                                           fifo_Y_pe_19_if_full_n,
    output wire                                          fifo_Y_pe_19_if_read,
    output wire                                          fifo_Y_pe_19_if_read_ce,
    output wire                                          fifo_Y_pe_19_if_write,
    output wire                                          fifo_Y_pe_19_if_write_ce,
    output wire                                          fifo_Y_pe_19_reset,
    output wire                                          fifo_Y_pe_1_clk,
    output wire [                                  64:0] fifo_Y_pe_1_if_din,
    input wire  [                                  64:0] fifo_Y_pe_1_if_dout,
    input wire                                           fifo_Y_pe_1_if_empty_n,
    input wire                                           fifo_Y_pe_1_if_full_n,
    output wire                                          fifo_Y_pe_1_if_read,
    output wire                                          fifo_Y_pe_1_if_read_ce,
    output wire                                          fifo_Y_pe_1_if_write,
    output wire                                          fifo_Y_pe_1_if_write_ce,
    output wire                                          fifo_Y_pe_1_reset,
    output wire                                          fifo_Y_pe_20_clk,
    output wire [                                  64:0] fifo_Y_pe_20_if_din,
    input wire  [                                  64:0] fifo_Y_pe_20_if_dout,
    input wire                                           fifo_Y_pe_20_if_empty_n,
    input wire                                           fifo_Y_pe_20_if_full_n,
    output wire                                          fifo_Y_pe_20_if_read,
    output wire                                          fifo_Y_pe_20_if_read_ce,
    output wire                                          fifo_Y_pe_20_if_write,
    output wire                                          fifo_Y_pe_20_if_write_ce,
    output wire                                          fifo_Y_pe_20_reset,
    output wire                                          fifo_Y_pe_21_clk,
    output wire [                                  64:0] fifo_Y_pe_21_if_din,
    input wire  [                                  64:0] fifo_Y_pe_21_if_dout,
    input wire                                           fifo_Y_pe_21_if_empty_n,
    input wire                                           fifo_Y_pe_21_if_full_n,
    output wire                                          fifo_Y_pe_21_if_read,
    output wire                                          fifo_Y_pe_21_if_read_ce,
    output wire                                          fifo_Y_pe_21_if_write,
    output wire                                          fifo_Y_pe_21_if_write_ce,
    output wire                                          fifo_Y_pe_21_reset,
    output wire                                          fifo_Y_pe_22_clk,
    output wire [                                  64:0] fifo_Y_pe_22_if_din,
    input wire  [                                  64:0] fifo_Y_pe_22_if_dout,
    input wire                                           fifo_Y_pe_22_if_empty_n,
    input wire                                           fifo_Y_pe_22_if_full_n,
    output wire                                          fifo_Y_pe_22_if_read,
    output wire                                          fifo_Y_pe_22_if_read_ce,
    output wire                                          fifo_Y_pe_22_if_write,
    output wire                                          fifo_Y_pe_22_if_write_ce,
    output wire                                          fifo_Y_pe_22_reset,
    output wire                                          fifo_Y_pe_23_clk,
    output wire [                                  64:0] fifo_Y_pe_23_if_din,
    input wire  [                                  64:0] fifo_Y_pe_23_if_dout,
    input wire                                           fifo_Y_pe_23_if_empty_n,
    input wire                                           fifo_Y_pe_23_if_full_n,
    output wire                                          fifo_Y_pe_23_if_read,
    output wire                                          fifo_Y_pe_23_if_read_ce,
    output wire                                          fifo_Y_pe_23_if_write,
    output wire                                          fifo_Y_pe_23_if_write_ce,
    output wire                                          fifo_Y_pe_23_reset,
    output wire                                          fifo_Y_pe_24_clk,
    output wire [                                  64:0] fifo_Y_pe_24_if_din,
    input wire  [                                  64:0] fifo_Y_pe_24_if_dout,
    input wire                                           fifo_Y_pe_24_if_empty_n,
    input wire                                           fifo_Y_pe_24_if_full_n,
    output wire                                          fifo_Y_pe_24_if_read,
    output wire                                          fifo_Y_pe_24_if_read_ce,
    output wire                                          fifo_Y_pe_24_if_write,
    output wire                                          fifo_Y_pe_24_if_write_ce,
    output wire                                          fifo_Y_pe_24_reset,
    output wire                                          fifo_Y_pe_25_clk,
    output wire [                                  64:0] fifo_Y_pe_25_if_din,
    input wire  [                                  64:0] fifo_Y_pe_25_if_dout,
    input wire                                           fifo_Y_pe_25_if_empty_n,
    input wire                                           fifo_Y_pe_25_if_full_n,
    output wire                                          fifo_Y_pe_25_if_read,
    output wire                                          fifo_Y_pe_25_if_read_ce,
    output wire                                          fifo_Y_pe_25_if_write,
    output wire                                          fifo_Y_pe_25_if_write_ce,
    output wire                                          fifo_Y_pe_25_reset,
    output wire                                          fifo_Y_pe_26_clk,
    output wire [                                  64:0] fifo_Y_pe_26_if_din,
    input wire  [                                  64:0] fifo_Y_pe_26_if_dout,
    input wire                                           fifo_Y_pe_26_if_empty_n,
    input wire                                           fifo_Y_pe_26_if_full_n,
    output wire                                          fifo_Y_pe_26_if_read,
    output wire                                          fifo_Y_pe_26_if_read_ce,
    output wire                                          fifo_Y_pe_26_if_write,
    output wire                                          fifo_Y_pe_26_if_write_ce,
    output wire                                          fifo_Y_pe_26_reset,
    output wire                                          fifo_Y_pe_27_clk,
    output wire [                                  64:0] fifo_Y_pe_27_if_din,
    input wire  [                                  64:0] fifo_Y_pe_27_if_dout,
    input wire                                           fifo_Y_pe_27_if_empty_n,
    input wire                                           fifo_Y_pe_27_if_full_n,
    output wire                                          fifo_Y_pe_27_if_read,
    output wire                                          fifo_Y_pe_27_if_read_ce,
    output wire                                          fifo_Y_pe_27_if_write,
    output wire                                          fifo_Y_pe_27_if_write_ce,
    output wire                                          fifo_Y_pe_27_reset,
    output wire                                          fifo_Y_pe_28_clk,
    output wire [                                  64:0] fifo_Y_pe_28_if_din,
    input wire  [                                  64:0] fifo_Y_pe_28_if_dout,
    input wire                                           fifo_Y_pe_28_if_empty_n,
    input wire                                           fifo_Y_pe_28_if_full_n,
    output wire                                          fifo_Y_pe_28_if_read,
    output wire                                          fifo_Y_pe_28_if_read_ce,
    output wire                                          fifo_Y_pe_28_if_write,
    output wire                                          fifo_Y_pe_28_if_write_ce,
    output wire                                          fifo_Y_pe_28_reset,
    output wire                                          fifo_Y_pe_29_clk,
    output wire [                                  64:0] fifo_Y_pe_29_if_din,
    input wire  [                                  64:0] fifo_Y_pe_29_if_dout,
    input wire                                           fifo_Y_pe_29_if_empty_n,
    input wire                                           fifo_Y_pe_29_if_full_n,
    output wire                                          fifo_Y_pe_29_if_read,
    output wire                                          fifo_Y_pe_29_if_read_ce,
    output wire                                          fifo_Y_pe_29_if_write,
    output wire                                          fifo_Y_pe_29_if_write_ce,
    output wire                                          fifo_Y_pe_29_reset,
    output wire                                          fifo_Y_pe_2_clk,
    output wire [                                  64:0] fifo_Y_pe_2_if_din,
    input wire  [                                  64:0] fifo_Y_pe_2_if_dout,
    input wire                                           fifo_Y_pe_2_if_empty_n,
    input wire                                           fifo_Y_pe_2_if_full_n,
    output wire                                          fifo_Y_pe_2_if_read,
    output wire                                          fifo_Y_pe_2_if_read_ce,
    output wire                                          fifo_Y_pe_2_if_write,
    output wire                                          fifo_Y_pe_2_if_write_ce,
    output wire                                          fifo_Y_pe_2_reset,
    output wire                                          fifo_Y_pe_30_clk,
    output wire [                                  64:0] fifo_Y_pe_30_if_din,
    input wire  [                                  64:0] fifo_Y_pe_30_if_dout,
    input wire                                           fifo_Y_pe_30_if_empty_n,
    input wire                                           fifo_Y_pe_30_if_full_n,
    output wire                                          fifo_Y_pe_30_if_read,
    output wire                                          fifo_Y_pe_30_if_read_ce,
    output wire                                          fifo_Y_pe_30_if_write,
    output wire                                          fifo_Y_pe_30_if_write_ce,
    output wire                                          fifo_Y_pe_30_reset,
    output wire                                          fifo_Y_pe_31_clk,
    output wire [                                  64:0] fifo_Y_pe_31_if_din,
    input wire  [                                  64:0] fifo_Y_pe_31_if_dout,
    input wire                                           fifo_Y_pe_31_if_empty_n,
    input wire                                           fifo_Y_pe_31_if_full_n,
    output wire                                          fifo_Y_pe_31_if_read,
    output wire                                          fifo_Y_pe_31_if_read_ce,
    output wire                                          fifo_Y_pe_31_if_write,
    output wire                                          fifo_Y_pe_31_if_write_ce,
    output wire                                          fifo_Y_pe_31_reset,
    output wire                                          fifo_Y_pe_32_clk,
    output wire [                                  64:0] fifo_Y_pe_32_if_din,
    input wire  [                                  64:0] fifo_Y_pe_32_if_dout,
    input wire                                           fifo_Y_pe_32_if_empty_n,
    input wire                                           fifo_Y_pe_32_if_full_n,
    output wire                                          fifo_Y_pe_32_if_read,
    output wire                                          fifo_Y_pe_32_if_read_ce,
    output wire                                          fifo_Y_pe_32_if_write,
    output wire                                          fifo_Y_pe_32_if_write_ce,
    output wire                                          fifo_Y_pe_32_reset,
    output wire                                          fifo_Y_pe_33_clk,
    output wire [                                  64:0] fifo_Y_pe_33_if_din,
    input wire  [                                  64:0] fifo_Y_pe_33_if_dout,
    input wire                                           fifo_Y_pe_33_if_empty_n,
    input wire                                           fifo_Y_pe_33_if_full_n,
    output wire                                          fifo_Y_pe_33_if_read,
    output wire                                          fifo_Y_pe_33_if_read_ce,
    output wire                                          fifo_Y_pe_33_if_write,
    output wire                                          fifo_Y_pe_33_if_write_ce,
    output wire                                          fifo_Y_pe_33_reset,
    output wire                                          fifo_Y_pe_34_clk,
    output wire [                                  64:0] fifo_Y_pe_34_if_din,
    input wire  [                                  64:0] fifo_Y_pe_34_if_dout,
    input wire                                           fifo_Y_pe_34_if_empty_n,
    input wire                                           fifo_Y_pe_34_if_full_n,
    output wire                                          fifo_Y_pe_34_if_read,
    output wire                                          fifo_Y_pe_34_if_read_ce,
    output wire                                          fifo_Y_pe_34_if_write,
    output wire                                          fifo_Y_pe_34_if_write_ce,
    output wire                                          fifo_Y_pe_34_reset,
    output wire                                          fifo_Y_pe_35_clk,
    output wire [                                  64:0] fifo_Y_pe_35_if_din,
    input wire  [                                  64:0] fifo_Y_pe_35_if_dout,
    input wire                                           fifo_Y_pe_35_if_empty_n,
    input wire                                           fifo_Y_pe_35_if_full_n,
    output wire                                          fifo_Y_pe_35_if_read,
    output wire                                          fifo_Y_pe_35_if_read_ce,
    output wire                                          fifo_Y_pe_35_if_write,
    output wire                                          fifo_Y_pe_35_if_write_ce,
    output wire                                          fifo_Y_pe_35_reset,
    output wire                                          fifo_Y_pe_36_clk,
    output wire [                                  64:0] fifo_Y_pe_36_if_din,
    input wire  [                                  64:0] fifo_Y_pe_36_if_dout,
    input wire                                           fifo_Y_pe_36_if_empty_n,
    input wire                                           fifo_Y_pe_36_if_full_n,
    output wire                                          fifo_Y_pe_36_if_read,
    output wire                                          fifo_Y_pe_36_if_read_ce,
    output wire                                          fifo_Y_pe_36_if_write,
    output wire                                          fifo_Y_pe_36_if_write_ce,
    output wire                                          fifo_Y_pe_36_reset,
    output wire                                          fifo_Y_pe_37_clk,
    output wire [                                  64:0] fifo_Y_pe_37_if_din,
    input wire  [                                  64:0] fifo_Y_pe_37_if_dout,
    input wire                                           fifo_Y_pe_37_if_empty_n,
    input wire                                           fifo_Y_pe_37_if_full_n,
    output wire                                          fifo_Y_pe_37_if_read,
    output wire                                          fifo_Y_pe_37_if_read_ce,
    output wire                                          fifo_Y_pe_37_if_write,
    output wire                                          fifo_Y_pe_37_if_write_ce,
    output wire                                          fifo_Y_pe_37_reset,
    output wire                                          fifo_Y_pe_38_clk,
    output wire [                                  64:0] fifo_Y_pe_38_if_din,
    input wire  [                                  64:0] fifo_Y_pe_38_if_dout,
    input wire                                           fifo_Y_pe_38_if_empty_n,
    input wire                                           fifo_Y_pe_38_if_full_n,
    output wire                                          fifo_Y_pe_38_if_read,
    output wire                                          fifo_Y_pe_38_if_read_ce,
    output wire                                          fifo_Y_pe_38_if_write,
    output wire                                          fifo_Y_pe_38_if_write_ce,
    output wire                                          fifo_Y_pe_38_reset,
    output wire                                          fifo_Y_pe_39_clk,
    output wire [                                  64:0] fifo_Y_pe_39_if_din,
    input wire  [                                  64:0] fifo_Y_pe_39_if_dout,
    input wire                                           fifo_Y_pe_39_if_empty_n,
    input wire                                           fifo_Y_pe_39_if_full_n,
    output wire                                          fifo_Y_pe_39_if_read,
    output wire                                          fifo_Y_pe_39_if_read_ce,
    output wire                                          fifo_Y_pe_39_if_write,
    output wire                                          fifo_Y_pe_39_if_write_ce,
    output wire                                          fifo_Y_pe_39_reset,
    output wire                                          fifo_Y_pe_3_clk,
    output wire [                                  64:0] fifo_Y_pe_3_if_din,
    input wire  [                                  64:0] fifo_Y_pe_3_if_dout,
    input wire                                           fifo_Y_pe_3_if_empty_n,
    input wire                                           fifo_Y_pe_3_if_full_n,
    output wire                                          fifo_Y_pe_3_if_read,
    output wire                                          fifo_Y_pe_3_if_read_ce,
    output wire                                          fifo_Y_pe_3_if_write,
    output wire                                          fifo_Y_pe_3_if_write_ce,
    output wire                                          fifo_Y_pe_3_reset,
    output wire                                          fifo_Y_pe_40_clk,
    output wire [                                  64:0] fifo_Y_pe_40_if_din,
    input wire  [                                  64:0] fifo_Y_pe_40_if_dout,
    input wire                                           fifo_Y_pe_40_if_empty_n,
    input wire                                           fifo_Y_pe_40_if_full_n,
    output wire                                          fifo_Y_pe_40_if_read,
    output wire                                          fifo_Y_pe_40_if_read_ce,
    output wire                                          fifo_Y_pe_40_if_write,
    output wire                                          fifo_Y_pe_40_if_write_ce,
    output wire                                          fifo_Y_pe_40_reset,
    output wire                                          fifo_Y_pe_41_clk,
    output wire [                                  64:0] fifo_Y_pe_41_if_din,
    input wire  [                                  64:0] fifo_Y_pe_41_if_dout,
    input wire                                           fifo_Y_pe_41_if_empty_n,
    input wire                                           fifo_Y_pe_41_if_full_n,
    output wire                                          fifo_Y_pe_41_if_read,
    output wire                                          fifo_Y_pe_41_if_read_ce,
    output wire                                          fifo_Y_pe_41_if_write,
    output wire                                          fifo_Y_pe_41_if_write_ce,
    output wire                                          fifo_Y_pe_41_reset,
    output wire                                          fifo_Y_pe_42_clk,
    output wire [                                  64:0] fifo_Y_pe_42_if_din,
    input wire  [                                  64:0] fifo_Y_pe_42_if_dout,
    input wire                                           fifo_Y_pe_42_if_empty_n,
    input wire                                           fifo_Y_pe_42_if_full_n,
    output wire                                          fifo_Y_pe_42_if_read,
    output wire                                          fifo_Y_pe_42_if_read_ce,
    output wire                                          fifo_Y_pe_42_if_write,
    output wire                                          fifo_Y_pe_42_if_write_ce,
    output wire                                          fifo_Y_pe_42_reset,
    output wire                                          fifo_Y_pe_43_clk,
    output wire [                                  64:0] fifo_Y_pe_43_if_din,
    input wire  [                                  64:0] fifo_Y_pe_43_if_dout,
    input wire                                           fifo_Y_pe_43_if_empty_n,
    input wire                                           fifo_Y_pe_43_if_full_n,
    output wire                                          fifo_Y_pe_43_if_read,
    output wire                                          fifo_Y_pe_43_if_read_ce,
    output wire                                          fifo_Y_pe_43_if_write,
    output wire                                          fifo_Y_pe_43_if_write_ce,
    output wire                                          fifo_Y_pe_43_reset,
    output wire                                          fifo_Y_pe_44_clk,
    output wire [                                  64:0] fifo_Y_pe_44_if_din,
    input wire  [                                  64:0] fifo_Y_pe_44_if_dout,
    input wire                                           fifo_Y_pe_44_if_empty_n,
    input wire                                           fifo_Y_pe_44_if_full_n,
    output wire                                          fifo_Y_pe_44_if_read,
    output wire                                          fifo_Y_pe_44_if_read_ce,
    output wire                                          fifo_Y_pe_44_if_write,
    output wire                                          fifo_Y_pe_44_if_write_ce,
    output wire                                          fifo_Y_pe_44_reset,
    output wire                                          fifo_Y_pe_45_clk,
    output wire [                                  64:0] fifo_Y_pe_45_if_din,
    input wire  [                                  64:0] fifo_Y_pe_45_if_dout,
    input wire                                           fifo_Y_pe_45_if_empty_n,
    input wire                                           fifo_Y_pe_45_if_full_n,
    output wire                                          fifo_Y_pe_45_if_read,
    output wire                                          fifo_Y_pe_45_if_read_ce,
    output wire                                          fifo_Y_pe_45_if_write,
    output wire                                          fifo_Y_pe_45_if_write_ce,
    output wire                                          fifo_Y_pe_45_reset,
    output wire                                          fifo_Y_pe_46_clk,
    output wire [                                  64:0] fifo_Y_pe_46_if_din,
    input wire  [                                  64:0] fifo_Y_pe_46_if_dout,
    input wire                                           fifo_Y_pe_46_if_empty_n,
    input wire                                           fifo_Y_pe_46_if_full_n,
    output wire                                          fifo_Y_pe_46_if_read,
    output wire                                          fifo_Y_pe_46_if_read_ce,
    output wire                                          fifo_Y_pe_46_if_write,
    output wire                                          fifo_Y_pe_46_if_write_ce,
    output wire                                          fifo_Y_pe_46_reset,
    output wire                                          fifo_Y_pe_47_clk,
    output wire [                                  64:0] fifo_Y_pe_47_if_din,
    input wire  [                                  64:0] fifo_Y_pe_47_if_dout,
    input wire                                           fifo_Y_pe_47_if_empty_n,
    input wire                                           fifo_Y_pe_47_if_full_n,
    output wire                                          fifo_Y_pe_47_if_read,
    output wire                                          fifo_Y_pe_47_if_read_ce,
    output wire                                          fifo_Y_pe_47_if_write,
    output wire                                          fifo_Y_pe_47_if_write_ce,
    output wire                                          fifo_Y_pe_47_reset,
    output wire                                          fifo_Y_pe_4_clk,
    output wire [                                  64:0] fifo_Y_pe_4_if_din,
    input wire  [                                  64:0] fifo_Y_pe_4_if_dout,
    input wire                                           fifo_Y_pe_4_if_empty_n,
    input wire                                           fifo_Y_pe_4_if_full_n,
    output wire                                          fifo_Y_pe_4_if_read,
    output wire                                          fifo_Y_pe_4_if_read_ce,
    output wire                                          fifo_Y_pe_4_if_write,
    output wire                                          fifo_Y_pe_4_if_write_ce,
    output wire                                          fifo_Y_pe_4_reset,
    output wire                                          fifo_Y_pe_5_clk,
    output wire [                                  64:0] fifo_Y_pe_5_if_din,
    input wire  [                                  64:0] fifo_Y_pe_5_if_dout,
    input wire                                           fifo_Y_pe_5_if_empty_n,
    input wire                                           fifo_Y_pe_5_if_full_n,
    output wire                                          fifo_Y_pe_5_if_read,
    output wire                                          fifo_Y_pe_5_if_read_ce,
    output wire                                          fifo_Y_pe_5_if_write,
    output wire                                          fifo_Y_pe_5_if_write_ce,
    output wire                                          fifo_Y_pe_5_reset,
    output wire                                          fifo_Y_pe_6_clk,
    output wire [                                  64:0] fifo_Y_pe_6_if_din,
    input wire  [                                  64:0] fifo_Y_pe_6_if_dout,
    input wire                                           fifo_Y_pe_6_if_empty_n,
    input wire                                           fifo_Y_pe_6_if_full_n,
    output wire                                          fifo_Y_pe_6_if_read,
    output wire                                          fifo_Y_pe_6_if_read_ce,
    output wire                                          fifo_Y_pe_6_if_write,
    output wire                                          fifo_Y_pe_6_if_write_ce,
    output wire                                          fifo_Y_pe_6_reset,
    output wire                                          fifo_Y_pe_7_clk,
    output wire [                                  64:0] fifo_Y_pe_7_if_din,
    input wire  [                                  64:0] fifo_Y_pe_7_if_dout,
    input wire                                           fifo_Y_pe_7_if_empty_n,
    input wire                                           fifo_Y_pe_7_if_full_n,
    output wire                                          fifo_Y_pe_7_if_read,
    output wire                                          fifo_Y_pe_7_if_read_ce,
    output wire                                          fifo_Y_pe_7_if_write,
    output wire                                          fifo_Y_pe_7_if_write_ce,
    output wire                                          fifo_Y_pe_7_reset,
    output wire                                          fifo_Y_pe_8_clk,
    output wire [                                  64:0] fifo_Y_pe_8_if_din,
    input wire  [                                  64:0] fifo_Y_pe_8_if_dout,
    input wire                                           fifo_Y_pe_8_if_empty_n,
    input wire                                           fifo_Y_pe_8_if_full_n,
    output wire                                          fifo_Y_pe_8_if_read,
    output wire                                          fifo_Y_pe_8_if_read_ce,
    output wire                                          fifo_Y_pe_8_if_write,
    output wire                                          fifo_Y_pe_8_if_write_ce,
    output wire                                          fifo_Y_pe_8_reset,
    output wire                                          fifo_Y_pe_9_clk,
    output wire [                                  64:0] fifo_Y_pe_9_if_din,
    input wire  [                                  64:0] fifo_Y_pe_9_if_dout,
    input wire                                           fifo_Y_pe_9_if_empty_n,
    input wire                                           fifo_Y_pe_9_if_full_n,
    output wire                                          fifo_Y_pe_9_if_read,
    output wire                                          fifo_Y_pe_9_if_read_ce,
    output wire                                          fifo_Y_pe_9_if_write,
    output wire                                          fifo_Y_pe_9_if_write_ce,
    output wire                                          fifo_Y_pe_9_reset,
    output wire                                          fifo_Y_pe_abd_0_clk,
    output wire [                                  64:0] fifo_Y_pe_abd_0_if_din,
    input wire  [                                  64:0] fifo_Y_pe_abd_0_if_dout,
    input wire                                           fifo_Y_pe_abd_0_if_empty_n,
    input wire                                           fifo_Y_pe_abd_0_if_full_n,
    output wire                                          fifo_Y_pe_abd_0_if_read,
    output wire                                          fifo_Y_pe_abd_0_if_read_ce,
    output wire                                          fifo_Y_pe_abd_0_if_write,
    output wire                                          fifo_Y_pe_abd_0_if_write_ce,
    output wire                                          fifo_Y_pe_abd_0_reset,
    output wire                                          fifo_Y_pe_abd_1_clk,
    output wire [                                  64:0] fifo_Y_pe_abd_1_if_din,
    input wire  [                                  64:0] fifo_Y_pe_abd_1_if_dout,
    input wire                                           fifo_Y_pe_abd_1_if_empty_n,
    input wire                                           fifo_Y_pe_abd_1_if_full_n,
    output wire                                          fifo_Y_pe_abd_1_if_read,
    output wire                                          fifo_Y_pe_abd_1_if_read_ce,
    output wire                                          fifo_Y_pe_abd_1_if_write,
    output wire                                          fifo_Y_pe_abd_1_if_write_ce,
    output wire                                          fifo_Y_pe_abd_1_reset,
    output wire                                          fifo_Y_pe_abd_2_clk,
    output wire [                                  64:0] fifo_Y_pe_abd_2_if_din,
    input wire  [                                  64:0] fifo_Y_pe_abd_2_if_dout,
    input wire                                           fifo_Y_pe_abd_2_if_empty_n,
    input wire                                           fifo_Y_pe_abd_2_if_full_n,
    output wire                                          fifo_Y_pe_abd_2_if_read,
    output wire                                          fifo_Y_pe_abd_2_if_read_ce,
    output wire                                          fifo_Y_pe_abd_2_if_write,
    output wire                                          fifo_Y_pe_abd_2_if_write_ce,
    output wire                                          fifo_Y_pe_abd_2_reset,
    output wire                                          fifo_Y_pe_abd_3_clk,
    output wire [                                  64:0] fifo_Y_pe_abd_3_if_din,
    input wire  [                                  64:0] fifo_Y_pe_abd_3_if_dout,
    input wire                                           fifo_Y_pe_abd_3_if_empty_n,
    input wire                                           fifo_Y_pe_abd_3_if_full_n,
    output wire                                          fifo_Y_pe_abd_3_if_read,
    output wire                                          fifo_Y_pe_abd_3_if_read_ce,
    output wire                                          fifo_Y_pe_abd_3_if_write,
    output wire                                          fifo_Y_pe_abd_3_if_write_ce,
    output wire                                          fifo_Y_pe_abd_3_reset,
    output wire                                          fifo_Y_pe_abd_4_clk,
    output wire [                                  64:0] fifo_Y_pe_abd_4_if_din,
    input wire  [                                  64:0] fifo_Y_pe_abd_4_if_dout,
    input wire                                           fifo_Y_pe_abd_4_if_empty_n,
    input wire                                           fifo_Y_pe_abd_4_if_full_n,
    output wire                                          fifo_Y_pe_abd_4_if_read,
    output wire                                          fifo_Y_pe_abd_4_if_read_ce,
    output wire                                          fifo_Y_pe_abd_4_if_write,
    output wire                                          fifo_Y_pe_abd_4_if_write_ce,
    output wire                                          fifo_Y_pe_abd_4_reset,
    output wire                                          fifo_Y_pe_abd_5_clk,
    output wire [                                  64:0] fifo_Y_pe_abd_5_if_din,
    input wire  [                                  64:0] fifo_Y_pe_abd_5_if_dout,
    input wire                                           fifo_Y_pe_abd_5_if_empty_n,
    input wire                                           fifo_Y_pe_abd_5_if_full_n,
    output wire                                          fifo_Y_pe_abd_5_if_read,
    output wire                                          fifo_Y_pe_abd_5_if_read_ce,
    output wire                                          fifo_Y_pe_abd_5_if_write,
    output wire                                          fifo_Y_pe_abd_5_if_write_ce,
    output wire                                          fifo_Y_pe_abd_5_reset,
    output wire                                          fifo_Y_pe_abd_6_clk,
    output wire [                                  64:0] fifo_Y_pe_abd_6_if_din,
    input wire  [                                  64:0] fifo_Y_pe_abd_6_if_dout,
    input wire                                           fifo_Y_pe_abd_6_if_empty_n,
    input wire                                           fifo_Y_pe_abd_6_if_full_n,
    output wire                                          fifo_Y_pe_abd_6_if_read,
    output wire                                          fifo_Y_pe_abd_6_if_read_ce,
    output wire                                          fifo_Y_pe_abd_6_if_write,
    output wire                                          fifo_Y_pe_abd_6_if_write_ce,
    output wire                                          fifo_Y_pe_abd_6_reset,
    output wire                                          fifo_Y_pe_abd_7_clk,
    output wire [                                  64:0] fifo_Y_pe_abd_7_if_din,
    input wire  [                                  64:0] fifo_Y_pe_abd_7_if_dout,
    input wire                                           fifo_Y_pe_abd_7_if_empty_n,
    input wire                                           fifo_Y_pe_abd_7_if_full_n,
    output wire                                          fifo_Y_pe_abd_7_if_read,
    output wire                                          fifo_Y_pe_abd_7_if_read_ce,
    output wire                                          fifo_Y_pe_abd_7_if_write,
    output wire                                          fifo_Y_pe_abd_7_if_write_ce,
    output wire                                          fifo_Y_pe_abd_7_reset,
    output wire                                          fifo_aXvec_0_clk,
    output wire [                                 400:0] fifo_aXvec_0_if_din,
    input wire  [                                 400:0] fifo_aXvec_0_if_dout,
    input wire                                           fifo_aXvec_0_if_empty_n,
    input wire                                           fifo_aXvec_0_if_full_n,
    output wire                                          fifo_aXvec_0_if_read,
    output wire                                          fifo_aXvec_0_if_read_ce,
    output wire                                          fifo_aXvec_0_if_write,
    output wire                                          fifo_aXvec_0_if_write_ce,
    output wire                                          fifo_aXvec_0_reset,
    output wire                                          fifo_aXvec_10_clk,
    output wire [                                 400:0] fifo_aXvec_10_if_din,
    input wire  [                                 400:0] fifo_aXvec_10_if_dout,
    input wire                                           fifo_aXvec_10_if_empty_n,
    input wire                                           fifo_aXvec_10_if_full_n,
    output wire                                          fifo_aXvec_10_if_read,
    output wire                                          fifo_aXvec_10_if_read_ce,
    output wire                                          fifo_aXvec_10_if_write,
    output wire                                          fifo_aXvec_10_if_write_ce,
    output wire                                          fifo_aXvec_10_reset,
    output wire                                          fifo_aXvec_11_clk,
    output wire [                                 400:0] fifo_aXvec_11_if_din,
    input wire  [                                 400:0] fifo_aXvec_11_if_dout,
    input wire                                           fifo_aXvec_11_if_empty_n,
    input wire                                           fifo_aXvec_11_if_full_n,
    output wire                                          fifo_aXvec_11_if_read,
    output wire                                          fifo_aXvec_11_if_read_ce,
    output wire                                          fifo_aXvec_11_if_write,
    output wire                                          fifo_aXvec_11_if_write_ce,
    output wire                                          fifo_aXvec_11_reset,
    output wire                                          fifo_aXvec_12_clk,
    output wire [                                 400:0] fifo_aXvec_12_if_din,
    input wire  [                                 400:0] fifo_aXvec_12_if_dout,
    input wire                                           fifo_aXvec_12_if_empty_n,
    input wire                                           fifo_aXvec_12_if_full_n,
    output wire                                          fifo_aXvec_12_if_read,
    output wire                                          fifo_aXvec_12_if_read_ce,
    output wire                                          fifo_aXvec_12_if_write,
    output wire                                          fifo_aXvec_12_if_write_ce,
    output wire                                          fifo_aXvec_12_reset,
    output wire                                          fifo_aXvec_13_clk,
    output wire [                                 400:0] fifo_aXvec_13_if_din,
    input wire  [                                 400:0] fifo_aXvec_13_if_dout,
    input wire                                           fifo_aXvec_13_if_empty_n,
    input wire                                           fifo_aXvec_13_if_full_n,
    output wire                                          fifo_aXvec_13_if_read,
    output wire                                          fifo_aXvec_13_if_read_ce,
    output wire                                          fifo_aXvec_13_if_write,
    output wire                                          fifo_aXvec_13_if_write_ce,
    output wire                                          fifo_aXvec_13_reset,
    output wire                                          fifo_aXvec_14_clk,
    output wire [                                 400:0] fifo_aXvec_14_if_din,
    input wire  [                                 400:0] fifo_aXvec_14_if_dout,
    input wire                                           fifo_aXvec_14_if_empty_n,
    input wire                                           fifo_aXvec_14_if_full_n,
    output wire                                          fifo_aXvec_14_if_read,
    output wire                                          fifo_aXvec_14_if_read_ce,
    output wire                                          fifo_aXvec_14_if_write,
    output wire                                          fifo_aXvec_14_if_write_ce,
    output wire                                          fifo_aXvec_14_reset,
    output wire                                          fifo_aXvec_15_clk,
    output wire [                                 400:0] fifo_aXvec_15_if_din,
    input wire  [                                 400:0] fifo_aXvec_15_if_dout,
    input wire                                           fifo_aXvec_15_if_empty_n,
    input wire                                           fifo_aXvec_15_if_full_n,
    output wire                                          fifo_aXvec_15_if_read,
    output wire                                          fifo_aXvec_15_if_read_ce,
    output wire                                          fifo_aXvec_15_if_write,
    output wire                                          fifo_aXvec_15_if_write_ce,
    output wire                                          fifo_aXvec_15_reset,
    output wire                                          fifo_aXvec_16_clk,
    output wire [                                 400:0] fifo_aXvec_16_if_din,
    input wire  [                                 400:0] fifo_aXvec_16_if_dout,
    input wire                                           fifo_aXvec_16_if_empty_n,
    input wire                                           fifo_aXvec_16_if_full_n,
    output wire                                          fifo_aXvec_16_if_read,
    output wire                                          fifo_aXvec_16_if_read_ce,
    output wire                                          fifo_aXvec_16_if_write,
    output wire                                          fifo_aXvec_16_if_write_ce,
    output wire                                          fifo_aXvec_16_reset,
    output wire                                          fifo_aXvec_17_clk,
    output wire [                                 400:0] fifo_aXvec_17_if_din,
    input wire  [                                 400:0] fifo_aXvec_17_if_dout,
    input wire                                           fifo_aXvec_17_if_empty_n,
    input wire                                           fifo_aXvec_17_if_full_n,
    output wire                                          fifo_aXvec_17_if_read,
    output wire                                          fifo_aXvec_17_if_read_ce,
    output wire                                          fifo_aXvec_17_if_write,
    output wire                                          fifo_aXvec_17_if_write_ce,
    output wire                                          fifo_aXvec_17_reset,
    output wire                                          fifo_aXvec_18_clk,
    output wire [                                 400:0] fifo_aXvec_18_if_din,
    input wire  [                                 400:0] fifo_aXvec_18_if_dout,
    input wire                                           fifo_aXvec_18_if_empty_n,
    input wire                                           fifo_aXvec_18_if_full_n,
    output wire                                          fifo_aXvec_18_if_read,
    output wire                                          fifo_aXvec_18_if_read_ce,
    output wire                                          fifo_aXvec_18_if_write,
    output wire                                          fifo_aXvec_18_if_write_ce,
    output wire                                          fifo_aXvec_18_reset,
    output wire                                          fifo_aXvec_19_clk,
    output wire [                                 400:0] fifo_aXvec_19_if_din,
    input wire  [                                 400:0] fifo_aXvec_19_if_dout,
    input wire                                           fifo_aXvec_19_if_empty_n,
    input wire                                           fifo_aXvec_19_if_full_n,
    output wire                                          fifo_aXvec_19_if_read,
    output wire                                          fifo_aXvec_19_if_read_ce,
    output wire                                          fifo_aXvec_19_if_write,
    output wire                                          fifo_aXvec_19_if_write_ce,
    output wire                                          fifo_aXvec_19_reset,
    output wire                                          fifo_aXvec_1_clk,
    output wire [                                 400:0] fifo_aXvec_1_if_din,
    input wire  [                                 400:0] fifo_aXvec_1_if_dout,
    input wire                                           fifo_aXvec_1_if_empty_n,
    input wire                                           fifo_aXvec_1_if_full_n,
    output wire                                          fifo_aXvec_1_if_read,
    output wire                                          fifo_aXvec_1_if_read_ce,
    output wire                                          fifo_aXvec_1_if_write,
    output wire                                          fifo_aXvec_1_if_write_ce,
    output wire                                          fifo_aXvec_1_reset,
    output wire                                          fifo_aXvec_20_clk,
    output wire [                                 400:0] fifo_aXvec_20_if_din,
    input wire  [                                 400:0] fifo_aXvec_20_if_dout,
    input wire                                           fifo_aXvec_20_if_empty_n,
    input wire                                           fifo_aXvec_20_if_full_n,
    output wire                                          fifo_aXvec_20_if_read,
    output wire                                          fifo_aXvec_20_if_read_ce,
    output wire                                          fifo_aXvec_20_if_write,
    output wire                                          fifo_aXvec_20_if_write_ce,
    output wire                                          fifo_aXvec_20_reset,
    output wire                                          fifo_aXvec_21_clk,
    output wire [                                 400:0] fifo_aXvec_21_if_din,
    input wire  [                                 400:0] fifo_aXvec_21_if_dout,
    input wire                                           fifo_aXvec_21_if_empty_n,
    input wire                                           fifo_aXvec_21_if_full_n,
    output wire                                          fifo_aXvec_21_if_read,
    output wire                                          fifo_aXvec_21_if_read_ce,
    output wire                                          fifo_aXvec_21_if_write,
    output wire                                          fifo_aXvec_21_if_write_ce,
    output wire                                          fifo_aXvec_21_reset,
    output wire                                          fifo_aXvec_22_clk,
    output wire [                                 400:0] fifo_aXvec_22_if_din,
    input wire  [                                 400:0] fifo_aXvec_22_if_dout,
    input wire                                           fifo_aXvec_22_if_empty_n,
    input wire                                           fifo_aXvec_22_if_full_n,
    output wire                                          fifo_aXvec_22_if_read,
    output wire                                          fifo_aXvec_22_if_read_ce,
    output wire                                          fifo_aXvec_22_if_write,
    output wire                                          fifo_aXvec_22_if_write_ce,
    output wire                                          fifo_aXvec_22_reset,
    output wire                                          fifo_aXvec_23_clk,
    output wire [                                 400:0] fifo_aXvec_23_if_din,
    input wire  [                                 400:0] fifo_aXvec_23_if_dout,
    input wire                                           fifo_aXvec_23_if_empty_n,
    input wire                                           fifo_aXvec_23_if_full_n,
    output wire                                          fifo_aXvec_23_if_read,
    output wire                                          fifo_aXvec_23_if_read_ce,
    output wire                                          fifo_aXvec_23_if_write,
    output wire                                          fifo_aXvec_23_if_write_ce,
    output wire                                          fifo_aXvec_23_reset,
    output wire                                          fifo_aXvec_24_clk,
    output wire [                                 400:0] fifo_aXvec_24_if_din,
    input wire  [                                 400:0] fifo_aXvec_24_if_dout,
    input wire                                           fifo_aXvec_24_if_empty_n,
    input wire                                           fifo_aXvec_24_if_full_n,
    output wire                                          fifo_aXvec_24_if_read,
    output wire                                          fifo_aXvec_24_if_read_ce,
    output wire                                          fifo_aXvec_24_if_write,
    output wire                                          fifo_aXvec_24_if_write_ce,
    output wire                                          fifo_aXvec_24_reset,
    output wire                                          fifo_aXvec_25_clk,
    output wire [                                 400:0] fifo_aXvec_25_if_din,
    input wire  [                                 400:0] fifo_aXvec_25_if_dout,
    input wire                                           fifo_aXvec_25_if_empty_n,
    input wire                                           fifo_aXvec_25_if_full_n,
    output wire                                          fifo_aXvec_25_if_read,
    output wire                                          fifo_aXvec_25_if_read_ce,
    output wire                                          fifo_aXvec_25_if_write,
    output wire                                          fifo_aXvec_25_if_write_ce,
    output wire                                          fifo_aXvec_25_reset,
    output wire                                          fifo_aXvec_26_clk,
    output wire [                                 400:0] fifo_aXvec_26_if_din,
    input wire  [                                 400:0] fifo_aXvec_26_if_dout,
    input wire                                           fifo_aXvec_26_if_empty_n,
    input wire                                           fifo_aXvec_26_if_full_n,
    output wire                                          fifo_aXvec_26_if_read,
    output wire                                          fifo_aXvec_26_if_read_ce,
    output wire                                          fifo_aXvec_26_if_write,
    output wire                                          fifo_aXvec_26_if_write_ce,
    output wire                                          fifo_aXvec_26_reset,
    output wire                                          fifo_aXvec_27_clk,
    output wire [                                 400:0] fifo_aXvec_27_if_din,
    input wire  [                                 400:0] fifo_aXvec_27_if_dout,
    input wire                                           fifo_aXvec_27_if_empty_n,
    input wire                                           fifo_aXvec_27_if_full_n,
    output wire                                          fifo_aXvec_27_if_read,
    output wire                                          fifo_aXvec_27_if_read_ce,
    output wire                                          fifo_aXvec_27_if_write,
    output wire                                          fifo_aXvec_27_if_write_ce,
    output wire                                          fifo_aXvec_27_reset,
    output wire                                          fifo_aXvec_28_clk,
    output wire [                                 400:0] fifo_aXvec_28_if_din,
    input wire  [                                 400:0] fifo_aXvec_28_if_dout,
    input wire                                           fifo_aXvec_28_if_empty_n,
    input wire                                           fifo_aXvec_28_if_full_n,
    output wire                                          fifo_aXvec_28_if_read,
    output wire                                          fifo_aXvec_28_if_read_ce,
    output wire                                          fifo_aXvec_28_if_write,
    output wire                                          fifo_aXvec_28_if_write_ce,
    output wire                                          fifo_aXvec_28_reset,
    output wire                                          fifo_aXvec_29_clk,
    output wire [                                 400:0] fifo_aXvec_29_if_din,
    input wire  [                                 400:0] fifo_aXvec_29_if_dout,
    input wire                                           fifo_aXvec_29_if_empty_n,
    input wire                                           fifo_aXvec_29_if_full_n,
    output wire                                          fifo_aXvec_29_if_read,
    output wire                                          fifo_aXvec_29_if_read_ce,
    output wire                                          fifo_aXvec_29_if_write,
    output wire                                          fifo_aXvec_29_if_write_ce,
    output wire                                          fifo_aXvec_29_reset,
    output wire                                          fifo_aXvec_2_clk,
    output wire [                                 400:0] fifo_aXvec_2_if_din,
    input wire  [                                 400:0] fifo_aXvec_2_if_dout,
    input wire                                           fifo_aXvec_2_if_empty_n,
    input wire                                           fifo_aXvec_2_if_full_n,
    output wire                                          fifo_aXvec_2_if_read,
    output wire                                          fifo_aXvec_2_if_read_ce,
    output wire                                          fifo_aXvec_2_if_write,
    output wire                                          fifo_aXvec_2_if_write_ce,
    output wire                                          fifo_aXvec_2_reset,
    output wire                                          fifo_aXvec_30_clk,
    output wire [                                 400:0] fifo_aXvec_30_if_din,
    input wire  [                                 400:0] fifo_aXvec_30_if_dout,
    input wire                                           fifo_aXvec_30_if_empty_n,
    input wire                                           fifo_aXvec_30_if_full_n,
    output wire                                          fifo_aXvec_30_if_read,
    output wire                                          fifo_aXvec_30_if_read_ce,
    output wire                                          fifo_aXvec_30_if_write,
    output wire                                          fifo_aXvec_30_if_write_ce,
    output wire                                          fifo_aXvec_30_reset,
    output wire                                          fifo_aXvec_31_clk,
    output wire [                                 400:0] fifo_aXvec_31_if_din,
    input wire  [                                 400:0] fifo_aXvec_31_if_dout,
    input wire                                           fifo_aXvec_31_if_empty_n,
    input wire                                           fifo_aXvec_31_if_full_n,
    output wire                                          fifo_aXvec_31_if_read,
    output wire                                          fifo_aXvec_31_if_read_ce,
    output wire                                          fifo_aXvec_31_if_write,
    output wire                                          fifo_aXvec_31_if_write_ce,
    output wire                                          fifo_aXvec_31_reset,
    output wire                                          fifo_aXvec_32_clk,
    output wire [                                 400:0] fifo_aXvec_32_if_din,
    input wire  [                                 400:0] fifo_aXvec_32_if_dout,
    input wire                                           fifo_aXvec_32_if_empty_n,
    input wire                                           fifo_aXvec_32_if_full_n,
    output wire                                          fifo_aXvec_32_if_read,
    output wire                                          fifo_aXvec_32_if_read_ce,
    output wire                                          fifo_aXvec_32_if_write,
    output wire                                          fifo_aXvec_32_if_write_ce,
    output wire                                          fifo_aXvec_32_reset,
    output wire                                          fifo_aXvec_33_clk,
    output wire [                                 400:0] fifo_aXvec_33_if_din,
    input wire  [                                 400:0] fifo_aXvec_33_if_dout,
    input wire                                           fifo_aXvec_33_if_empty_n,
    input wire                                           fifo_aXvec_33_if_full_n,
    output wire                                          fifo_aXvec_33_if_read,
    output wire                                          fifo_aXvec_33_if_read_ce,
    output wire                                          fifo_aXvec_33_if_write,
    output wire                                          fifo_aXvec_33_if_write_ce,
    output wire                                          fifo_aXvec_33_reset,
    output wire                                          fifo_aXvec_34_clk,
    output wire [                                 400:0] fifo_aXvec_34_if_din,
    input wire  [                                 400:0] fifo_aXvec_34_if_dout,
    input wire                                           fifo_aXvec_34_if_empty_n,
    input wire                                           fifo_aXvec_34_if_full_n,
    output wire                                          fifo_aXvec_34_if_read,
    output wire                                          fifo_aXvec_34_if_read_ce,
    output wire                                          fifo_aXvec_34_if_write,
    output wire                                          fifo_aXvec_34_if_write_ce,
    output wire                                          fifo_aXvec_34_reset,
    output wire                                          fifo_aXvec_35_clk,
    output wire [                                 400:0] fifo_aXvec_35_if_din,
    input wire  [                                 400:0] fifo_aXvec_35_if_dout,
    input wire                                           fifo_aXvec_35_if_empty_n,
    input wire                                           fifo_aXvec_35_if_full_n,
    output wire                                          fifo_aXvec_35_if_read,
    output wire                                          fifo_aXvec_35_if_read_ce,
    output wire                                          fifo_aXvec_35_if_write,
    output wire                                          fifo_aXvec_35_if_write_ce,
    output wire                                          fifo_aXvec_35_reset,
    output wire                                          fifo_aXvec_36_clk,
    output wire [                                 400:0] fifo_aXvec_36_if_din,
    input wire  [                                 400:0] fifo_aXvec_36_if_dout,
    input wire                                           fifo_aXvec_36_if_empty_n,
    input wire                                           fifo_aXvec_36_if_full_n,
    output wire                                          fifo_aXvec_36_if_read,
    output wire                                          fifo_aXvec_36_if_read_ce,
    output wire                                          fifo_aXvec_36_if_write,
    output wire                                          fifo_aXvec_36_if_write_ce,
    output wire                                          fifo_aXvec_36_reset,
    output wire                                          fifo_aXvec_37_clk,
    output wire [                                 400:0] fifo_aXvec_37_if_din,
    input wire  [                                 400:0] fifo_aXvec_37_if_dout,
    input wire                                           fifo_aXvec_37_if_empty_n,
    input wire                                           fifo_aXvec_37_if_full_n,
    output wire                                          fifo_aXvec_37_if_read,
    output wire                                          fifo_aXvec_37_if_read_ce,
    output wire                                          fifo_aXvec_37_if_write,
    output wire                                          fifo_aXvec_37_if_write_ce,
    output wire                                          fifo_aXvec_37_reset,
    output wire                                          fifo_aXvec_38_clk,
    output wire [                                 400:0] fifo_aXvec_38_if_din,
    input wire  [                                 400:0] fifo_aXvec_38_if_dout,
    input wire                                           fifo_aXvec_38_if_empty_n,
    input wire                                           fifo_aXvec_38_if_full_n,
    output wire                                          fifo_aXvec_38_if_read,
    output wire                                          fifo_aXvec_38_if_read_ce,
    output wire                                          fifo_aXvec_38_if_write,
    output wire                                          fifo_aXvec_38_if_write_ce,
    output wire                                          fifo_aXvec_38_reset,
    output wire                                          fifo_aXvec_39_clk,
    output wire [                                 400:0] fifo_aXvec_39_if_din,
    input wire  [                                 400:0] fifo_aXvec_39_if_dout,
    input wire                                           fifo_aXvec_39_if_empty_n,
    input wire                                           fifo_aXvec_39_if_full_n,
    output wire                                          fifo_aXvec_39_if_read,
    output wire                                          fifo_aXvec_39_if_read_ce,
    output wire                                          fifo_aXvec_39_if_write,
    output wire                                          fifo_aXvec_39_if_write_ce,
    output wire                                          fifo_aXvec_39_reset,
    output wire                                          fifo_aXvec_3_clk,
    output wire [                                 400:0] fifo_aXvec_3_if_din,
    input wire  [                                 400:0] fifo_aXvec_3_if_dout,
    input wire                                           fifo_aXvec_3_if_empty_n,
    input wire                                           fifo_aXvec_3_if_full_n,
    output wire                                          fifo_aXvec_3_if_read,
    output wire                                          fifo_aXvec_3_if_read_ce,
    output wire                                          fifo_aXvec_3_if_write,
    output wire                                          fifo_aXvec_3_if_write_ce,
    output wire                                          fifo_aXvec_3_reset,
    output wire                                          fifo_aXvec_40_clk,
    output wire [                                 400:0] fifo_aXvec_40_if_din,
    input wire  [                                 400:0] fifo_aXvec_40_if_dout,
    input wire                                           fifo_aXvec_40_if_empty_n,
    input wire                                           fifo_aXvec_40_if_full_n,
    output wire                                          fifo_aXvec_40_if_read,
    output wire                                          fifo_aXvec_40_if_read_ce,
    output wire                                          fifo_aXvec_40_if_write,
    output wire                                          fifo_aXvec_40_if_write_ce,
    output wire                                          fifo_aXvec_40_reset,
    output wire                                          fifo_aXvec_41_clk,
    output wire [                                 400:0] fifo_aXvec_41_if_din,
    input wire  [                                 400:0] fifo_aXvec_41_if_dout,
    input wire                                           fifo_aXvec_41_if_empty_n,
    input wire                                           fifo_aXvec_41_if_full_n,
    output wire                                          fifo_aXvec_41_if_read,
    output wire                                          fifo_aXvec_41_if_read_ce,
    output wire                                          fifo_aXvec_41_if_write,
    output wire                                          fifo_aXvec_41_if_write_ce,
    output wire                                          fifo_aXvec_41_reset,
    output wire                                          fifo_aXvec_42_clk,
    output wire [                                 400:0] fifo_aXvec_42_if_din,
    input wire  [                                 400:0] fifo_aXvec_42_if_dout,
    input wire                                           fifo_aXvec_42_if_empty_n,
    input wire                                           fifo_aXvec_42_if_full_n,
    output wire                                          fifo_aXvec_42_if_read,
    output wire                                          fifo_aXvec_42_if_read_ce,
    output wire                                          fifo_aXvec_42_if_write,
    output wire                                          fifo_aXvec_42_if_write_ce,
    output wire                                          fifo_aXvec_42_reset,
    output wire                                          fifo_aXvec_43_clk,
    output wire [                                 400:0] fifo_aXvec_43_if_din,
    input wire  [                                 400:0] fifo_aXvec_43_if_dout,
    input wire                                           fifo_aXvec_43_if_empty_n,
    input wire                                           fifo_aXvec_43_if_full_n,
    output wire                                          fifo_aXvec_43_if_read,
    output wire                                          fifo_aXvec_43_if_read_ce,
    output wire                                          fifo_aXvec_43_if_write,
    output wire                                          fifo_aXvec_43_if_write_ce,
    output wire                                          fifo_aXvec_43_reset,
    output wire                                          fifo_aXvec_44_clk,
    output wire [                                 400:0] fifo_aXvec_44_if_din,
    input wire  [                                 400:0] fifo_aXvec_44_if_dout,
    input wire                                           fifo_aXvec_44_if_empty_n,
    input wire                                           fifo_aXvec_44_if_full_n,
    output wire                                          fifo_aXvec_44_if_read,
    output wire                                          fifo_aXvec_44_if_read_ce,
    output wire                                          fifo_aXvec_44_if_write,
    output wire                                          fifo_aXvec_44_if_write_ce,
    output wire                                          fifo_aXvec_44_reset,
    output wire                                          fifo_aXvec_45_clk,
    output wire [                                 400:0] fifo_aXvec_45_if_din,
    input wire  [                                 400:0] fifo_aXvec_45_if_dout,
    input wire                                           fifo_aXvec_45_if_empty_n,
    input wire                                           fifo_aXvec_45_if_full_n,
    output wire                                          fifo_aXvec_45_if_read,
    output wire                                          fifo_aXvec_45_if_read_ce,
    output wire                                          fifo_aXvec_45_if_write,
    output wire                                          fifo_aXvec_45_if_write_ce,
    output wire                                          fifo_aXvec_45_reset,
    output wire                                          fifo_aXvec_46_clk,
    output wire [                                 400:0] fifo_aXvec_46_if_din,
    input wire  [                                 400:0] fifo_aXvec_46_if_dout,
    input wire                                           fifo_aXvec_46_if_empty_n,
    input wire                                           fifo_aXvec_46_if_full_n,
    output wire                                          fifo_aXvec_46_if_read,
    output wire                                          fifo_aXvec_46_if_read_ce,
    output wire                                          fifo_aXvec_46_if_write,
    output wire                                          fifo_aXvec_46_if_write_ce,
    output wire                                          fifo_aXvec_46_reset,
    output wire                                          fifo_aXvec_47_clk,
    output wire [                                 400:0] fifo_aXvec_47_if_din,
    input wire  [                                 400:0] fifo_aXvec_47_if_dout,
    input wire                                           fifo_aXvec_47_if_empty_n,
    input wire                                           fifo_aXvec_47_if_full_n,
    output wire                                          fifo_aXvec_47_if_read,
    output wire                                          fifo_aXvec_47_if_read_ce,
    output wire                                          fifo_aXvec_47_if_write,
    output wire                                          fifo_aXvec_47_if_write_ce,
    output wire                                          fifo_aXvec_47_reset,
    output wire                                          fifo_aXvec_4_clk,
    output wire [                                 400:0] fifo_aXvec_4_if_din,
    input wire  [                                 400:0] fifo_aXvec_4_if_dout,
    input wire                                           fifo_aXvec_4_if_empty_n,
    input wire                                           fifo_aXvec_4_if_full_n,
    output wire                                          fifo_aXvec_4_if_read,
    output wire                                          fifo_aXvec_4_if_read_ce,
    output wire                                          fifo_aXvec_4_if_write,
    output wire                                          fifo_aXvec_4_if_write_ce,
    output wire                                          fifo_aXvec_4_reset,
    output wire                                          fifo_aXvec_5_clk,
    output wire [                                 400:0] fifo_aXvec_5_if_din,
    input wire  [                                 400:0] fifo_aXvec_5_if_dout,
    input wire                                           fifo_aXvec_5_if_empty_n,
    input wire                                           fifo_aXvec_5_if_full_n,
    output wire                                          fifo_aXvec_5_if_read,
    output wire                                          fifo_aXvec_5_if_read_ce,
    output wire                                          fifo_aXvec_5_if_write,
    output wire                                          fifo_aXvec_5_if_write_ce,
    output wire                                          fifo_aXvec_5_reset,
    output wire                                          fifo_aXvec_6_clk,
    output wire [                                 400:0] fifo_aXvec_6_if_din,
    input wire  [                                 400:0] fifo_aXvec_6_if_dout,
    input wire                                           fifo_aXvec_6_if_empty_n,
    input wire                                           fifo_aXvec_6_if_full_n,
    output wire                                          fifo_aXvec_6_if_read,
    output wire                                          fifo_aXvec_6_if_read_ce,
    output wire                                          fifo_aXvec_6_if_write,
    output wire                                          fifo_aXvec_6_if_write_ce,
    output wire                                          fifo_aXvec_6_reset,
    output wire                                          fifo_aXvec_7_clk,
    output wire [                                 400:0] fifo_aXvec_7_if_din,
    input wire  [                                 400:0] fifo_aXvec_7_if_dout,
    input wire                                           fifo_aXvec_7_if_empty_n,
    input wire                                           fifo_aXvec_7_if_full_n,
    output wire                                          fifo_aXvec_7_if_read,
    output wire                                          fifo_aXvec_7_if_read_ce,
    output wire                                          fifo_aXvec_7_if_write,
    output wire                                          fifo_aXvec_7_if_write_ce,
    output wire                                          fifo_aXvec_7_reset,
    output wire                                          fifo_aXvec_8_clk,
    output wire [                                 400:0] fifo_aXvec_8_if_din,
    input wire  [                                 400:0] fifo_aXvec_8_if_dout,
    input wire                                           fifo_aXvec_8_if_empty_n,
    input wire                                           fifo_aXvec_8_if_full_n,
    output wire                                          fifo_aXvec_8_if_read,
    output wire                                          fifo_aXvec_8_if_read_ce,
    output wire                                          fifo_aXvec_8_if_write,
    output wire                                          fifo_aXvec_8_if_write_ce,
    output wire                                          fifo_aXvec_8_reset,
    output wire                                          fifo_aXvec_9_clk,
    output wire [                                 400:0] fifo_aXvec_9_if_din,
    input wire  [                                 400:0] fifo_aXvec_9_if_dout,
    input wire                                           fifo_aXvec_9_if_empty_n,
    input wire                                           fifo_aXvec_9_if_full_n,
    output wire                                          fifo_aXvec_9_if_read,
    output wire                                          fifo_aXvec_9_if_read_ce,
    output wire                                          fifo_aXvec_9_if_write,
    output wire                                          fifo_aXvec_9_if_write_ce,
    output wire                                          fifo_aXvec_9_reset,
    output wire [                                  31:0] Arbiter_Y_0_M,
    output wire [                                  31:0] Arbiter_Y_0_P_N,
    output wire                                          Arbiter_Y_0_ap_clk,
    input wire                                           Arbiter_Y_0_ap_done,
    input wire                                           Arbiter_Y_0_ap_idle,
    input wire                                           Arbiter_Y_0_ap_ready,
    output wire                                          Arbiter_Y_0_ap_rst_n,
    output wire                                          Arbiter_Y_0_ap_start,
    output wire [                                  64:0] Arbiter_Y_0_fifo_in_0_dout,
    output wire                                          Arbiter_Y_0_fifo_in_0_empty_n,
    input wire                                           Arbiter_Y_0_fifo_in_0_read,
    output wire [                                  64:0] Arbiter_Y_0_fifo_in_1_dout,
    output wire                                          Arbiter_Y_0_fifo_in_1_empty_n,
    input wire                                           Arbiter_Y_0_fifo_in_1_read,
    output wire [                                  64:0] Arbiter_Y_0_fifo_in_2_dout,
    output wire                                          Arbiter_Y_0_fifo_in_2_empty_n,
    input wire                                           Arbiter_Y_0_fifo_in_2_read,
    output wire [                                  64:0] Arbiter_Y_0_fifo_in_3_dout,
    output wire                                          Arbiter_Y_0_fifo_in_3_empty_n,
    input wire                                           Arbiter_Y_0_fifo_in_3_read,
    output wire [                                  64:0] Arbiter_Y_0_fifo_in_4_dout,
    output wire                                          Arbiter_Y_0_fifo_in_4_empty_n,
    input wire                                           Arbiter_Y_0_fifo_in_4_read,
    output wire [                                  64:0] Arbiter_Y_0_fifo_in_5_dout,
    output wire                                          Arbiter_Y_0_fifo_in_5_empty_n,
    input wire                                           Arbiter_Y_0_fifo_in_5_read,
    output wire [                                  64:0] Arbiter_Y_0_fifo_in_peek_0_dout,
    output wire                                          Arbiter_Y_0_fifo_in_peek_0_empty_n,
    input wire                                           Arbiter_Y_0_fifo_in_peek_0_read,
    output wire [                                  64:0] Arbiter_Y_0_fifo_in_peek_1_dout,
    output wire                                          Arbiter_Y_0_fifo_in_peek_1_empty_n,
    input wire                                           Arbiter_Y_0_fifo_in_peek_1_read,
    output wire [                                  64:0] Arbiter_Y_0_fifo_in_peek_2_dout,
    output wire                                          Arbiter_Y_0_fifo_in_peek_2_empty_n,
    input wire                                           Arbiter_Y_0_fifo_in_peek_2_read,
    output wire [                                  64:0] Arbiter_Y_0_fifo_in_peek_3_dout,
    output wire                                          Arbiter_Y_0_fifo_in_peek_3_empty_n,
    input wire                                           Arbiter_Y_0_fifo_in_peek_3_read,
    output wire [                                  64:0] Arbiter_Y_0_fifo_in_peek_4_dout,
    output wire                                          Arbiter_Y_0_fifo_in_peek_4_empty_n,
    input wire                                           Arbiter_Y_0_fifo_in_peek_4_read,
    output wire [                                  64:0] Arbiter_Y_0_fifo_in_peek_5_dout,
    output wire                                          Arbiter_Y_0_fifo_in_peek_5_empty_n,
    input wire                                           Arbiter_Y_0_fifo_in_peek_5_read,
    input wire  [                                  64:0] Arbiter_Y_0_fifo_out_din,
    output wire                                          Arbiter_Y_0_fifo_out_full_n,
    input wire                                           Arbiter_Y_0_fifo_out_write,
    output wire [                                  31:0] Arbiter_Y_1_M,
    output wire [                                  31:0] Arbiter_Y_1_P_N,
    output wire                                          Arbiter_Y_1_ap_clk,
    input wire                                           Arbiter_Y_1_ap_done,
    input wire                                           Arbiter_Y_1_ap_idle,
    input wire                                           Arbiter_Y_1_ap_ready,
    output wire                                          Arbiter_Y_1_ap_rst_n,
    output wire                                          Arbiter_Y_1_ap_start,
    output wire [                                  64:0] Arbiter_Y_1_fifo_in_0_dout,
    output wire                                          Arbiter_Y_1_fifo_in_0_empty_n,
    input wire                                           Arbiter_Y_1_fifo_in_0_read,
    output wire [                                  64:0] Arbiter_Y_1_fifo_in_1_dout,
    output wire                                          Arbiter_Y_1_fifo_in_1_empty_n,
    input wire                                           Arbiter_Y_1_fifo_in_1_read,
    output wire [                                  64:0] Arbiter_Y_1_fifo_in_2_dout,
    output wire                                          Arbiter_Y_1_fifo_in_2_empty_n,
    input wire                                           Arbiter_Y_1_fifo_in_2_read,
    output wire [                                  64:0] Arbiter_Y_1_fifo_in_3_dout,
    output wire                                          Arbiter_Y_1_fifo_in_3_empty_n,
    input wire                                           Arbiter_Y_1_fifo_in_3_read,
    output wire [                                  64:0] Arbiter_Y_1_fifo_in_4_dout,
    output wire                                          Arbiter_Y_1_fifo_in_4_empty_n,
    input wire                                           Arbiter_Y_1_fifo_in_4_read,
    output wire [                                  64:0] Arbiter_Y_1_fifo_in_5_dout,
    output wire                                          Arbiter_Y_1_fifo_in_5_empty_n,
    input wire                                           Arbiter_Y_1_fifo_in_5_read,
    output wire [                                  64:0] Arbiter_Y_1_fifo_in_peek_0_dout,
    output wire                                          Arbiter_Y_1_fifo_in_peek_0_empty_n,
    input wire                                           Arbiter_Y_1_fifo_in_peek_0_read,
    output wire [                                  64:0] Arbiter_Y_1_fifo_in_peek_1_dout,
    output wire                                          Arbiter_Y_1_fifo_in_peek_1_empty_n,
    input wire                                           Arbiter_Y_1_fifo_in_peek_1_read,
    output wire [                                  64:0] Arbiter_Y_1_fifo_in_peek_2_dout,
    output wire                                          Arbiter_Y_1_fifo_in_peek_2_empty_n,
    input wire                                           Arbiter_Y_1_fifo_in_peek_2_read,
    output wire [                                  64:0] Arbiter_Y_1_fifo_in_peek_3_dout,
    output wire                                          Arbiter_Y_1_fifo_in_peek_3_empty_n,
    input wire                                           Arbiter_Y_1_fifo_in_peek_3_read,
    output wire [                                  64:0] Arbiter_Y_1_fifo_in_peek_4_dout,
    output wire                                          Arbiter_Y_1_fifo_in_peek_4_empty_n,
    input wire                                           Arbiter_Y_1_fifo_in_peek_4_read,
    output wire [                                  64:0] Arbiter_Y_1_fifo_in_peek_5_dout,
    output wire                                          Arbiter_Y_1_fifo_in_peek_5_empty_n,
    input wire                                           Arbiter_Y_1_fifo_in_peek_5_read,
    input wire  [                                  64:0] Arbiter_Y_1_fifo_out_din,
    output wire                                          Arbiter_Y_1_fifo_out_full_n,
    input wire                                           Arbiter_Y_1_fifo_out_write,
    output wire [                                  31:0] Arbiter_Y_2_M,
    output wire [                                  31:0] Arbiter_Y_2_P_N,
    output wire                                          Arbiter_Y_2_ap_clk,
    input wire                                           Arbiter_Y_2_ap_done,
    input wire                                           Arbiter_Y_2_ap_idle,
    input wire                                           Arbiter_Y_2_ap_ready,
    output wire                                          Arbiter_Y_2_ap_rst_n,
    output wire                                          Arbiter_Y_2_ap_start,
    output wire [                                  64:0] Arbiter_Y_2_fifo_in_0_dout,
    output wire                                          Arbiter_Y_2_fifo_in_0_empty_n,
    input wire                                           Arbiter_Y_2_fifo_in_0_read,
    output wire [                                  64:0] Arbiter_Y_2_fifo_in_1_dout,
    output wire                                          Arbiter_Y_2_fifo_in_1_empty_n,
    input wire                                           Arbiter_Y_2_fifo_in_1_read,
    output wire [                                  64:0] Arbiter_Y_2_fifo_in_2_dout,
    output wire                                          Arbiter_Y_2_fifo_in_2_empty_n,
    input wire                                           Arbiter_Y_2_fifo_in_2_read,
    output wire [                                  64:0] Arbiter_Y_2_fifo_in_3_dout,
    output wire                                          Arbiter_Y_2_fifo_in_3_empty_n,
    input wire                                           Arbiter_Y_2_fifo_in_3_read,
    output wire [                                  64:0] Arbiter_Y_2_fifo_in_4_dout,
    output wire                                          Arbiter_Y_2_fifo_in_4_empty_n,
    input wire                                           Arbiter_Y_2_fifo_in_4_read,
    output wire [                                  64:0] Arbiter_Y_2_fifo_in_5_dout,
    output wire                                          Arbiter_Y_2_fifo_in_5_empty_n,
    input wire                                           Arbiter_Y_2_fifo_in_5_read,
    output wire [                                  64:0] Arbiter_Y_2_fifo_in_peek_0_dout,
    output wire                                          Arbiter_Y_2_fifo_in_peek_0_empty_n,
    input wire                                           Arbiter_Y_2_fifo_in_peek_0_read,
    output wire [                                  64:0] Arbiter_Y_2_fifo_in_peek_1_dout,
    output wire                                          Arbiter_Y_2_fifo_in_peek_1_empty_n,
    input wire                                           Arbiter_Y_2_fifo_in_peek_1_read,
    output wire [                                  64:0] Arbiter_Y_2_fifo_in_peek_2_dout,
    output wire                                          Arbiter_Y_2_fifo_in_peek_2_empty_n,
    input wire                                           Arbiter_Y_2_fifo_in_peek_2_read,
    output wire [                                  64:0] Arbiter_Y_2_fifo_in_peek_3_dout,
    output wire                                          Arbiter_Y_2_fifo_in_peek_3_empty_n,
    input wire                                           Arbiter_Y_2_fifo_in_peek_3_read,
    output wire [                                  64:0] Arbiter_Y_2_fifo_in_peek_4_dout,
    output wire                                          Arbiter_Y_2_fifo_in_peek_4_empty_n,
    input wire                                           Arbiter_Y_2_fifo_in_peek_4_read,
    output wire [                                  64:0] Arbiter_Y_2_fifo_in_peek_5_dout,
    output wire                                          Arbiter_Y_2_fifo_in_peek_5_empty_n,
    input wire                                           Arbiter_Y_2_fifo_in_peek_5_read,
    input wire  [                                  64:0] Arbiter_Y_2_fifo_out_din,
    output wire                                          Arbiter_Y_2_fifo_out_full_n,
    input wire                                           Arbiter_Y_2_fifo_out_write,
    output wire [                                  31:0] Arbiter_Y_3_M,
    output wire [                                  31:0] Arbiter_Y_3_P_N,
    output wire                                          Arbiter_Y_3_ap_clk,
    input wire                                           Arbiter_Y_3_ap_done,
    input wire                                           Arbiter_Y_3_ap_idle,
    input wire                                           Arbiter_Y_3_ap_ready,
    output wire                                          Arbiter_Y_3_ap_rst_n,
    output wire                                          Arbiter_Y_3_ap_start,
    output wire [                                  64:0] Arbiter_Y_3_fifo_in_0_dout,
    output wire                                          Arbiter_Y_3_fifo_in_0_empty_n,
    input wire                                           Arbiter_Y_3_fifo_in_0_read,
    output wire [                                  64:0] Arbiter_Y_3_fifo_in_1_dout,
    output wire                                          Arbiter_Y_3_fifo_in_1_empty_n,
    input wire                                           Arbiter_Y_3_fifo_in_1_read,
    output wire [                                  64:0] Arbiter_Y_3_fifo_in_2_dout,
    output wire                                          Arbiter_Y_3_fifo_in_2_empty_n,
    input wire                                           Arbiter_Y_3_fifo_in_2_read,
    output wire [                                  64:0] Arbiter_Y_3_fifo_in_3_dout,
    output wire                                          Arbiter_Y_3_fifo_in_3_empty_n,
    input wire                                           Arbiter_Y_3_fifo_in_3_read,
    output wire [                                  64:0] Arbiter_Y_3_fifo_in_4_dout,
    output wire                                          Arbiter_Y_3_fifo_in_4_empty_n,
    input wire                                           Arbiter_Y_3_fifo_in_4_read,
    output wire [                                  64:0] Arbiter_Y_3_fifo_in_5_dout,
    output wire                                          Arbiter_Y_3_fifo_in_5_empty_n,
    input wire                                           Arbiter_Y_3_fifo_in_5_read,
    output wire [                                  64:0] Arbiter_Y_3_fifo_in_peek_0_dout,
    output wire                                          Arbiter_Y_3_fifo_in_peek_0_empty_n,
    input wire                                           Arbiter_Y_3_fifo_in_peek_0_read,
    output wire [                                  64:0] Arbiter_Y_3_fifo_in_peek_1_dout,
    output wire                                          Arbiter_Y_3_fifo_in_peek_1_empty_n,
    input wire                                           Arbiter_Y_3_fifo_in_peek_1_read,
    output wire [                                  64:0] Arbiter_Y_3_fifo_in_peek_2_dout,
    output wire                                          Arbiter_Y_3_fifo_in_peek_2_empty_n,
    input wire                                           Arbiter_Y_3_fifo_in_peek_2_read,
    output wire [                                  64:0] Arbiter_Y_3_fifo_in_peek_3_dout,
    output wire                                          Arbiter_Y_3_fifo_in_peek_3_empty_n,
    input wire                                           Arbiter_Y_3_fifo_in_peek_3_read,
    output wire [                                  64:0] Arbiter_Y_3_fifo_in_peek_4_dout,
    output wire                                          Arbiter_Y_3_fifo_in_peek_4_empty_n,
    input wire                                           Arbiter_Y_3_fifo_in_peek_4_read,
    output wire [                                  64:0] Arbiter_Y_3_fifo_in_peek_5_dout,
    output wire                                          Arbiter_Y_3_fifo_in_peek_5_empty_n,
    input wire                                           Arbiter_Y_3_fifo_in_peek_5_read,
    input wire  [                                  64:0] Arbiter_Y_3_fifo_out_din,
    output wire                                          Arbiter_Y_3_fifo_out_full_n,
    input wire                                           Arbiter_Y_3_fifo_out_write,
    output wire [                                  31:0] Arbiter_Y_4_M,
    output wire [                                  31:0] Arbiter_Y_4_P_N,
    output wire                                          Arbiter_Y_4_ap_clk,
    input wire                                           Arbiter_Y_4_ap_done,
    input wire                                           Arbiter_Y_4_ap_idle,
    input wire                                           Arbiter_Y_4_ap_ready,
    output wire                                          Arbiter_Y_4_ap_rst_n,
    output wire                                          Arbiter_Y_4_ap_start,
    output wire [                                  64:0] Arbiter_Y_4_fifo_in_0_dout,
    output wire                                          Arbiter_Y_4_fifo_in_0_empty_n,
    input wire                                           Arbiter_Y_4_fifo_in_0_read,
    output wire [                                  64:0] Arbiter_Y_4_fifo_in_1_dout,
    output wire                                          Arbiter_Y_4_fifo_in_1_empty_n,
    input wire                                           Arbiter_Y_4_fifo_in_1_read,
    output wire [                                  64:0] Arbiter_Y_4_fifo_in_2_dout,
    output wire                                          Arbiter_Y_4_fifo_in_2_empty_n,
    input wire                                           Arbiter_Y_4_fifo_in_2_read,
    output wire [                                  64:0] Arbiter_Y_4_fifo_in_3_dout,
    output wire                                          Arbiter_Y_4_fifo_in_3_empty_n,
    input wire                                           Arbiter_Y_4_fifo_in_3_read,
    output wire [                                  64:0] Arbiter_Y_4_fifo_in_4_dout,
    output wire                                          Arbiter_Y_4_fifo_in_4_empty_n,
    input wire                                           Arbiter_Y_4_fifo_in_4_read,
    output wire [                                  64:0] Arbiter_Y_4_fifo_in_5_dout,
    output wire                                          Arbiter_Y_4_fifo_in_5_empty_n,
    input wire                                           Arbiter_Y_4_fifo_in_5_read,
    output wire [                                  64:0] Arbiter_Y_4_fifo_in_peek_0_dout,
    output wire                                          Arbiter_Y_4_fifo_in_peek_0_empty_n,
    input wire                                           Arbiter_Y_4_fifo_in_peek_0_read,
    output wire [                                  64:0] Arbiter_Y_4_fifo_in_peek_1_dout,
    output wire                                          Arbiter_Y_4_fifo_in_peek_1_empty_n,
    input wire                                           Arbiter_Y_4_fifo_in_peek_1_read,
    output wire [                                  64:0] Arbiter_Y_4_fifo_in_peek_2_dout,
    output wire                                          Arbiter_Y_4_fifo_in_peek_2_empty_n,
    input wire                                           Arbiter_Y_4_fifo_in_peek_2_read,
    output wire [                                  64:0] Arbiter_Y_4_fifo_in_peek_3_dout,
    output wire                                          Arbiter_Y_4_fifo_in_peek_3_empty_n,
    input wire                                           Arbiter_Y_4_fifo_in_peek_3_read,
    output wire [                                  64:0] Arbiter_Y_4_fifo_in_peek_4_dout,
    output wire                                          Arbiter_Y_4_fifo_in_peek_4_empty_n,
    input wire                                           Arbiter_Y_4_fifo_in_peek_4_read,
    output wire [                                  64:0] Arbiter_Y_4_fifo_in_peek_5_dout,
    output wire                                          Arbiter_Y_4_fifo_in_peek_5_empty_n,
    input wire                                           Arbiter_Y_4_fifo_in_peek_5_read,
    input wire  [                                  64:0] Arbiter_Y_4_fifo_out_din,
    output wire                                          Arbiter_Y_4_fifo_out_full_n,
    input wire                                           Arbiter_Y_4_fifo_out_write,
    output wire [                                  31:0] Arbiter_Y_5_M,
    output wire [                                  31:0] Arbiter_Y_5_P_N,
    output wire                                          Arbiter_Y_5_ap_clk,
    input wire                                           Arbiter_Y_5_ap_done,
    input wire                                           Arbiter_Y_5_ap_idle,
    input wire                                           Arbiter_Y_5_ap_ready,
    output wire                                          Arbiter_Y_5_ap_rst_n,
    output wire                                          Arbiter_Y_5_ap_start,
    output wire [                                  64:0] Arbiter_Y_5_fifo_in_0_dout,
    output wire                                          Arbiter_Y_5_fifo_in_0_empty_n,
    input wire                                           Arbiter_Y_5_fifo_in_0_read,
    output wire [                                  64:0] Arbiter_Y_5_fifo_in_1_dout,
    output wire                                          Arbiter_Y_5_fifo_in_1_empty_n,
    input wire                                           Arbiter_Y_5_fifo_in_1_read,
    output wire [                                  64:0] Arbiter_Y_5_fifo_in_2_dout,
    output wire                                          Arbiter_Y_5_fifo_in_2_empty_n,
    input wire                                           Arbiter_Y_5_fifo_in_2_read,
    output wire [                                  64:0] Arbiter_Y_5_fifo_in_3_dout,
    output wire                                          Arbiter_Y_5_fifo_in_3_empty_n,
    input wire                                           Arbiter_Y_5_fifo_in_3_read,
    output wire [                                  64:0] Arbiter_Y_5_fifo_in_4_dout,
    output wire                                          Arbiter_Y_5_fifo_in_4_empty_n,
    input wire                                           Arbiter_Y_5_fifo_in_4_read,
    output wire [                                  64:0] Arbiter_Y_5_fifo_in_5_dout,
    output wire                                          Arbiter_Y_5_fifo_in_5_empty_n,
    input wire                                           Arbiter_Y_5_fifo_in_5_read,
    output wire [                                  64:0] Arbiter_Y_5_fifo_in_peek_0_dout,
    output wire                                          Arbiter_Y_5_fifo_in_peek_0_empty_n,
    input wire                                           Arbiter_Y_5_fifo_in_peek_0_read,
    output wire [                                  64:0] Arbiter_Y_5_fifo_in_peek_1_dout,
    output wire                                          Arbiter_Y_5_fifo_in_peek_1_empty_n,
    input wire                                           Arbiter_Y_5_fifo_in_peek_1_read,
    output wire [                                  64:0] Arbiter_Y_5_fifo_in_peek_2_dout,
    output wire                                          Arbiter_Y_5_fifo_in_peek_2_empty_n,
    input wire                                           Arbiter_Y_5_fifo_in_peek_2_read,
    output wire [                                  64:0] Arbiter_Y_5_fifo_in_peek_3_dout,
    output wire                                          Arbiter_Y_5_fifo_in_peek_3_empty_n,
    input wire                                           Arbiter_Y_5_fifo_in_peek_3_read,
    output wire [                                  64:0] Arbiter_Y_5_fifo_in_peek_4_dout,
    output wire                                          Arbiter_Y_5_fifo_in_peek_4_empty_n,
    input wire                                           Arbiter_Y_5_fifo_in_peek_4_read,
    output wire [                                  64:0] Arbiter_Y_5_fifo_in_peek_5_dout,
    output wire                                          Arbiter_Y_5_fifo_in_peek_5_empty_n,
    input wire                                           Arbiter_Y_5_fifo_in_peek_5_read,
    input wire  [                                  64:0] Arbiter_Y_5_fifo_out_din,
    output wire                                          Arbiter_Y_5_fifo_out_full_n,
    input wire                                           Arbiter_Y_5_fifo_out_write,
    output wire [                                  31:0] Arbiter_Y_6_M,
    output wire [                                  31:0] Arbiter_Y_6_P_N,
    output wire                                          Arbiter_Y_6_ap_clk,
    input wire                                           Arbiter_Y_6_ap_done,
    input wire                                           Arbiter_Y_6_ap_idle,
    input wire                                           Arbiter_Y_6_ap_ready,
    output wire                                          Arbiter_Y_6_ap_rst_n,
    output wire                                          Arbiter_Y_6_ap_start,
    output wire [                                  64:0] Arbiter_Y_6_fifo_in_0_dout,
    output wire                                          Arbiter_Y_6_fifo_in_0_empty_n,
    input wire                                           Arbiter_Y_6_fifo_in_0_read,
    output wire [                                  64:0] Arbiter_Y_6_fifo_in_1_dout,
    output wire                                          Arbiter_Y_6_fifo_in_1_empty_n,
    input wire                                           Arbiter_Y_6_fifo_in_1_read,
    output wire [                                  64:0] Arbiter_Y_6_fifo_in_2_dout,
    output wire                                          Arbiter_Y_6_fifo_in_2_empty_n,
    input wire                                           Arbiter_Y_6_fifo_in_2_read,
    output wire [                                  64:0] Arbiter_Y_6_fifo_in_3_dout,
    output wire                                          Arbiter_Y_6_fifo_in_3_empty_n,
    input wire                                           Arbiter_Y_6_fifo_in_3_read,
    output wire [                                  64:0] Arbiter_Y_6_fifo_in_4_dout,
    output wire                                          Arbiter_Y_6_fifo_in_4_empty_n,
    input wire                                           Arbiter_Y_6_fifo_in_4_read,
    output wire [                                  64:0] Arbiter_Y_6_fifo_in_5_dout,
    output wire                                          Arbiter_Y_6_fifo_in_5_empty_n,
    input wire                                           Arbiter_Y_6_fifo_in_5_read,
    output wire [                                  64:0] Arbiter_Y_6_fifo_in_peek_0_dout,
    output wire                                          Arbiter_Y_6_fifo_in_peek_0_empty_n,
    input wire                                           Arbiter_Y_6_fifo_in_peek_0_read,
    output wire [                                  64:0] Arbiter_Y_6_fifo_in_peek_1_dout,
    output wire                                          Arbiter_Y_6_fifo_in_peek_1_empty_n,
    input wire                                           Arbiter_Y_6_fifo_in_peek_1_read,
    output wire [                                  64:0] Arbiter_Y_6_fifo_in_peek_2_dout,
    output wire                                          Arbiter_Y_6_fifo_in_peek_2_empty_n,
    input wire                                           Arbiter_Y_6_fifo_in_peek_2_read,
    output wire [                                  64:0] Arbiter_Y_6_fifo_in_peek_3_dout,
    output wire                                          Arbiter_Y_6_fifo_in_peek_3_empty_n,
    input wire                                           Arbiter_Y_6_fifo_in_peek_3_read,
    output wire [                                  64:0] Arbiter_Y_6_fifo_in_peek_4_dout,
    output wire                                          Arbiter_Y_6_fifo_in_peek_4_empty_n,
    input wire                                           Arbiter_Y_6_fifo_in_peek_4_read,
    output wire [                                  64:0] Arbiter_Y_6_fifo_in_peek_5_dout,
    output wire                                          Arbiter_Y_6_fifo_in_peek_5_empty_n,
    input wire                                           Arbiter_Y_6_fifo_in_peek_5_read,
    input wire  [                                  64:0] Arbiter_Y_6_fifo_out_din,
    output wire                                          Arbiter_Y_6_fifo_out_full_n,
    input wire                                           Arbiter_Y_6_fifo_out_write,
    output wire [                                  31:0] Arbiter_Y_7_M,
    output wire [                                  31:0] Arbiter_Y_7_P_N,
    output wire                                          Arbiter_Y_7_ap_clk,
    input wire                                           Arbiter_Y_7_ap_done,
    input wire                                           Arbiter_Y_7_ap_idle,
    input wire                                           Arbiter_Y_7_ap_ready,
    output wire                                          Arbiter_Y_7_ap_rst_n,
    output wire                                          Arbiter_Y_7_ap_start,
    output wire [                                  64:0] Arbiter_Y_7_fifo_in_0_dout,
    output wire                                          Arbiter_Y_7_fifo_in_0_empty_n,
    input wire                                           Arbiter_Y_7_fifo_in_0_read,
    output wire [                                  64:0] Arbiter_Y_7_fifo_in_1_dout,
    output wire                                          Arbiter_Y_7_fifo_in_1_empty_n,
    input wire                                           Arbiter_Y_7_fifo_in_1_read,
    output wire [                                  64:0] Arbiter_Y_7_fifo_in_2_dout,
    output wire                                          Arbiter_Y_7_fifo_in_2_empty_n,
    input wire                                           Arbiter_Y_7_fifo_in_2_read,
    output wire [                                  64:0] Arbiter_Y_7_fifo_in_3_dout,
    output wire                                          Arbiter_Y_7_fifo_in_3_empty_n,
    input wire                                           Arbiter_Y_7_fifo_in_3_read,
    output wire [                                  64:0] Arbiter_Y_7_fifo_in_4_dout,
    output wire                                          Arbiter_Y_7_fifo_in_4_empty_n,
    input wire                                           Arbiter_Y_7_fifo_in_4_read,
    output wire [                                  64:0] Arbiter_Y_7_fifo_in_5_dout,
    output wire                                          Arbiter_Y_7_fifo_in_5_empty_n,
    input wire                                           Arbiter_Y_7_fifo_in_5_read,
    output wire [                                  64:0] Arbiter_Y_7_fifo_in_peek_0_dout,
    output wire                                          Arbiter_Y_7_fifo_in_peek_0_empty_n,
    input wire                                           Arbiter_Y_7_fifo_in_peek_0_read,
    output wire [                                  64:0] Arbiter_Y_7_fifo_in_peek_1_dout,
    output wire                                          Arbiter_Y_7_fifo_in_peek_1_empty_n,
    input wire                                           Arbiter_Y_7_fifo_in_peek_1_read,
    output wire [                                  64:0] Arbiter_Y_7_fifo_in_peek_2_dout,
    output wire                                          Arbiter_Y_7_fifo_in_peek_2_empty_n,
    input wire                                           Arbiter_Y_7_fifo_in_peek_2_read,
    output wire [                                  64:0] Arbiter_Y_7_fifo_in_peek_3_dout,
    output wire                                          Arbiter_Y_7_fifo_in_peek_3_empty_n,
    input wire                                           Arbiter_Y_7_fifo_in_peek_3_read,
    output wire [                                  64:0] Arbiter_Y_7_fifo_in_peek_4_dout,
    output wire                                          Arbiter_Y_7_fifo_in_peek_4_empty_n,
    input wire                                           Arbiter_Y_7_fifo_in_peek_4_read,
    output wire [                                  64:0] Arbiter_Y_7_fifo_in_peek_5_dout,
    output wire                                          Arbiter_Y_7_fifo_in_peek_5_empty_n,
    input wire                                           Arbiter_Y_7_fifo_in_peek_5_read,
    input wire  [                                  64:0] Arbiter_Y_7_fifo_out_din,
    output wire                                          Arbiter_Y_7_fifo_out_full_n,
    input wire                                           Arbiter_Y_7_fifo_out_write,
    output wire                                          FloatvAddFloatv_0_ap_clk,
    input wire                                           FloatvAddFloatv_0_ap_done,
    input wire                                           FloatvAddFloatv_0_ap_idle,
    input wire                                           FloatvAddFloatv_0_ap_ready,
    output wire                                          FloatvAddFloatv_0_ap_rst_n,
    output wire                                          FloatvAddFloatv_0_ap_start,
    output wire [                                 512:0] FloatvAddFloatv_0_fifo_in0_peek_dout,
    output wire                                          FloatvAddFloatv_0_fifo_in0_peek_empty_n,
    input wire                                           FloatvAddFloatv_0_fifo_in0_peek_read,
    output wire [                                 512:0] FloatvAddFloatv_0_fifo_in0_s_dout,
    output wire                                          FloatvAddFloatv_0_fifo_in0_s_empty_n,
    input wire                                           FloatvAddFloatv_0_fifo_in0_s_read,
    output wire [                                 512:0] FloatvAddFloatv_0_fifo_in1_peek_dout,
    output wire                                          FloatvAddFloatv_0_fifo_in1_peek_empty_n,
    input wire                                           FloatvAddFloatv_0_fifo_in1_peek_read,
    output wire [                                 512:0] FloatvAddFloatv_0_fifo_in1_s_dout,
    output wire                                          FloatvAddFloatv_0_fifo_in1_s_empty_n,
    input wire                                           FloatvAddFloatv_0_fifo_in1_s_read,
    input wire  [                                 512:0] FloatvAddFloatv_0_fifo_out_din,
    output wire                                          FloatvAddFloatv_0_fifo_out_full_n,
    input wire                                           FloatvAddFloatv_0_fifo_out_write,
    output wire [                                  31:0] FloatvMultConst_0_M,
    output wire [                                  31:0] FloatvMultConst_0_P_N,
    output wire [                                  31:0] FloatvMultConst_0_alpha_u,
    output wire                                          FloatvMultConst_0_ap_clk,
    input wire                                           FloatvMultConst_0_ap_done,
    input wire                                           FloatvMultConst_0_ap_idle,
    input wire                                           FloatvMultConst_0_ap_ready,
    output wire                                          FloatvMultConst_0_ap_rst_n,
    output wire                                          FloatvMultConst_0_ap_start,
    output wire [                                 512:0] FloatvMultConst_0_fifo_in_peek_dout,
    output wire                                          FloatvMultConst_0_fifo_in_peek_empty_n,
    input wire                                           FloatvMultConst_0_fifo_in_peek_read,
    output wire [                                 512:0] FloatvMultConst_0_fifo_in_s_dout,
    output wire                                          FloatvMultConst_0_fifo_in_s_empty_n,
    input wire                                           FloatvMultConst_0_fifo_in_s_read,
    input wire  [                                 512:0] FloatvMultConst_0_fifo_out_din,
    output wire                                          FloatvMultConst_0_fifo_out_full_n,
    input wire                                           FloatvMultConst_0_fifo_out_write,
    output wire [                                  31:0] FloatvMultConst_1_M,
    output wire [                                  31:0] FloatvMultConst_1_P_N,
    output wire [                                  31:0] FloatvMultConst_1_alpha_u,
    output wire                                          FloatvMultConst_1_ap_clk,
    input wire                                           FloatvMultConst_1_ap_done,
    input wire                                           FloatvMultConst_1_ap_idle,
    input wire                                           FloatvMultConst_1_ap_ready,
    output wire                                          FloatvMultConst_1_ap_rst_n,
    output wire                                          FloatvMultConst_1_ap_start,
    output wire [                                 512:0] FloatvMultConst_1_fifo_in_peek_dout,
    output wire                                          FloatvMultConst_1_fifo_in_peek_empty_n,
    input wire                                           FloatvMultConst_1_fifo_in_peek_read,
    output wire [                                 512:0] FloatvMultConst_1_fifo_in_s_dout,
    output wire                                          FloatvMultConst_1_fifo_in_s_empty_n,
    input wire                                           FloatvMultConst_1_fifo_in_s_read,
    input wire  [                                 512:0] FloatvMultConst_1_fifo_out_din,
    output wire                                          FloatvMultConst_1_fifo_out_full_n,
    input wire                                           FloatvMultConst_1_fifo_out_write,
    output wire                                          Merger_Y_0_ap_clk,
    input wire                                           Merger_Y_0_ap_done,
    input wire                                           Merger_Y_0_ap_idle,
    input wire                                           Merger_Y_0_ap_ready,
    output wire                                          Merger_Y_0_ap_rst_n,
    output wire                                          Merger_Y_0_ap_start,
    output wire [                                  64:0] Merger_Y_0_fifo_in_0_dout,
    output wire                                          Merger_Y_0_fifo_in_0_empty_n,
    input wire                                           Merger_Y_0_fifo_in_0_read,
    output wire [                                  64:0] Merger_Y_0_fifo_in_1_dout,
    output wire                                          Merger_Y_0_fifo_in_1_empty_n,
    input wire                                           Merger_Y_0_fifo_in_1_read,
    output wire [                                  64:0] Merger_Y_0_fifo_in_2_dout,
    output wire                                          Merger_Y_0_fifo_in_2_empty_n,
    input wire                                           Merger_Y_0_fifo_in_2_read,
    output wire [                                  64:0] Merger_Y_0_fifo_in_3_dout,
    output wire                                          Merger_Y_0_fifo_in_3_empty_n,
    input wire                                           Merger_Y_0_fifo_in_3_read,
    output wire [                                  64:0] Merger_Y_0_fifo_in_4_dout,
    output wire                                          Merger_Y_0_fifo_in_4_empty_n,
    input wire                                           Merger_Y_0_fifo_in_4_read,
    output wire [                                  64:0] Merger_Y_0_fifo_in_5_dout,
    output wire                                          Merger_Y_0_fifo_in_5_empty_n,
    input wire                                           Merger_Y_0_fifo_in_5_read,
    output wire [                                  64:0] Merger_Y_0_fifo_in_6_dout,
    output wire                                          Merger_Y_0_fifo_in_6_empty_n,
    input wire                                           Merger_Y_0_fifo_in_6_read,
    output wire [                                  64:0] Merger_Y_0_fifo_in_7_dout,
    output wire                                          Merger_Y_0_fifo_in_7_empty_n,
    input wire                                           Merger_Y_0_fifo_in_7_read,
    output wire [                                  64:0] Merger_Y_0_fifo_in_peek_0_dout,
    output wire                                          Merger_Y_0_fifo_in_peek_0_empty_n,
    input wire                                           Merger_Y_0_fifo_in_peek_0_read,
    output wire [                                  64:0] Merger_Y_0_fifo_in_peek_1_dout,
    output wire                                          Merger_Y_0_fifo_in_peek_1_empty_n,
    input wire                                           Merger_Y_0_fifo_in_peek_1_read,
    output wire [                                  64:0] Merger_Y_0_fifo_in_peek_2_dout,
    output wire                                          Merger_Y_0_fifo_in_peek_2_empty_n,
    input wire                                           Merger_Y_0_fifo_in_peek_2_read,
    output wire [                                  64:0] Merger_Y_0_fifo_in_peek_3_dout,
    output wire                                          Merger_Y_0_fifo_in_peek_3_empty_n,
    input wire                                           Merger_Y_0_fifo_in_peek_3_read,
    output wire [                                  64:0] Merger_Y_0_fifo_in_peek_4_dout,
    output wire                                          Merger_Y_0_fifo_in_peek_4_empty_n,
    input wire                                           Merger_Y_0_fifo_in_peek_4_read,
    output wire [                                  64:0] Merger_Y_0_fifo_in_peek_5_dout,
    output wire                                          Merger_Y_0_fifo_in_peek_5_empty_n,
    input wire                                           Merger_Y_0_fifo_in_peek_5_read,
    output wire [                                  64:0] Merger_Y_0_fifo_in_peek_6_dout,
    output wire                                          Merger_Y_0_fifo_in_peek_6_empty_n,
    input wire                                           Merger_Y_0_fifo_in_peek_6_read,
    output wire [                                  64:0] Merger_Y_0_fifo_in_peek_7_dout,
    output wire                                          Merger_Y_0_fifo_in_peek_7_empty_n,
    input wire                                           Merger_Y_0_fifo_in_peek_7_read,
    input wire  [                                 512:0] Merger_Y_0_fifo_out_din,
    output wire                                          Merger_Y_0_fifo_out_full_n,
    input wire                                           Merger_Y_0_fifo_out_write,
    output wire                                          PEG_Xvec_0_ap_clk,
    input wire                                           PEG_Xvec_0_ap_done,
    input wire                                           PEG_Xvec_0_ap_idle,
    input wire                                           PEG_Xvec_0_ap_ready,
    output wire                                          PEG_Xvec_0_ap_rst_n,
    output wire                                          PEG_Xvec_0_ap_start,
    output wire [                                 512:0] PEG_Xvec_0_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_0_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_0_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_0_fifo_A_s_dout,
    output wire                                          PEG_Xvec_0_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_0_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_0_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_0_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_0_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_0_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_0_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_0_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_0_fifo_X_out_din,
    output wire                                          PEG_Xvec_0_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_0_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_0_fifo_aXvec_din,
    output wire                                          PEG_Xvec_0_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_0_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_0_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_0_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_0_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_0_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_0_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_0_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_0_fifo_inst_out_din,
    output wire                                          PEG_Xvec_0_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_0_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_0_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_0_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_0_fifo_inst_out_write,
    output wire                                          PEG_Xvec_1_ap_clk,
    input wire                                           PEG_Xvec_1_ap_done,
    input wire                                           PEG_Xvec_1_ap_idle,
    input wire                                           PEG_Xvec_1_ap_ready,
    output wire                                          PEG_Xvec_1_ap_rst_n,
    output wire                                          PEG_Xvec_1_ap_start,
    output wire [                                 512:0] PEG_Xvec_1_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_1_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_1_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_1_fifo_A_s_dout,
    output wire                                          PEG_Xvec_1_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_1_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_1_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_1_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_1_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_1_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_1_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_1_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_1_fifo_X_out_din,
    output wire                                          PEG_Xvec_1_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_1_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_1_fifo_aXvec_din,
    output wire                                          PEG_Xvec_1_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_1_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_1_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_1_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_1_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_1_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_1_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_1_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_1_fifo_inst_out_din,
    output wire                                          PEG_Xvec_1_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_1_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_1_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_1_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_1_fifo_inst_out_write,
    output wire                                          PEG_Xvec_2_ap_clk,
    input wire                                           PEG_Xvec_2_ap_done,
    input wire                                           PEG_Xvec_2_ap_idle,
    input wire                                           PEG_Xvec_2_ap_ready,
    output wire                                          PEG_Xvec_2_ap_rst_n,
    output wire                                          PEG_Xvec_2_ap_start,
    output wire [                                 512:0] PEG_Xvec_2_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_2_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_2_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_2_fifo_A_s_dout,
    output wire                                          PEG_Xvec_2_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_2_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_2_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_2_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_2_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_2_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_2_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_2_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_2_fifo_X_out_din,
    output wire                                          PEG_Xvec_2_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_2_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_2_fifo_aXvec_din,
    output wire                                          PEG_Xvec_2_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_2_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_2_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_2_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_2_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_2_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_2_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_2_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_2_fifo_inst_out_din,
    output wire                                          PEG_Xvec_2_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_2_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_2_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_2_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_2_fifo_inst_out_write,
    output wire                                          PEG_Xvec_3_ap_clk,
    input wire                                           PEG_Xvec_3_ap_done,
    input wire                                           PEG_Xvec_3_ap_idle,
    input wire                                           PEG_Xvec_3_ap_ready,
    output wire                                          PEG_Xvec_3_ap_rst_n,
    output wire                                          PEG_Xvec_3_ap_start,
    output wire [                                 512:0] PEG_Xvec_3_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_3_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_3_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_3_fifo_A_s_dout,
    output wire                                          PEG_Xvec_3_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_3_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_3_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_3_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_3_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_3_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_3_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_3_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_3_fifo_X_out_din,
    output wire                                          PEG_Xvec_3_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_3_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_3_fifo_aXvec_din,
    output wire                                          PEG_Xvec_3_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_3_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_3_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_3_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_3_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_3_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_3_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_3_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_3_fifo_inst_out_din,
    output wire                                          PEG_Xvec_3_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_3_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_3_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_3_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_3_fifo_inst_out_write,
    output wire                                          PEG_Xvec_4_ap_clk,
    input wire                                           PEG_Xvec_4_ap_done,
    input wire                                           PEG_Xvec_4_ap_idle,
    input wire                                           PEG_Xvec_4_ap_ready,
    output wire                                          PEG_Xvec_4_ap_rst_n,
    output wire                                          PEG_Xvec_4_ap_start,
    output wire [                                 512:0] PEG_Xvec_4_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_4_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_4_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_4_fifo_A_s_dout,
    output wire                                          PEG_Xvec_4_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_4_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_4_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_4_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_4_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_4_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_4_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_4_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_4_fifo_X_out_din,
    output wire                                          PEG_Xvec_4_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_4_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_4_fifo_aXvec_din,
    output wire                                          PEG_Xvec_4_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_4_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_4_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_4_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_4_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_4_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_4_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_4_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_4_fifo_inst_out_din,
    output wire                                          PEG_Xvec_4_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_4_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_4_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_4_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_4_fifo_inst_out_write,
    output wire                                          PEG_Xvec_5_ap_clk,
    input wire                                           PEG_Xvec_5_ap_done,
    input wire                                           PEG_Xvec_5_ap_idle,
    input wire                                           PEG_Xvec_5_ap_ready,
    output wire                                          PEG_Xvec_5_ap_rst_n,
    output wire                                          PEG_Xvec_5_ap_start,
    output wire [                                 512:0] PEG_Xvec_5_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_5_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_5_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_5_fifo_A_s_dout,
    output wire                                          PEG_Xvec_5_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_5_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_5_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_5_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_5_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_5_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_5_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_5_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_5_fifo_X_out_din,
    output wire                                          PEG_Xvec_5_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_5_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_5_fifo_aXvec_din,
    output wire                                          PEG_Xvec_5_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_5_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_5_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_5_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_5_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_5_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_5_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_5_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_5_fifo_inst_out_din,
    output wire                                          PEG_Xvec_5_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_5_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_5_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_5_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_5_fifo_inst_out_write,
    output wire                                          PEG_Xvec_6_ap_clk,
    input wire                                           PEG_Xvec_6_ap_done,
    input wire                                           PEG_Xvec_6_ap_idle,
    input wire                                           PEG_Xvec_6_ap_ready,
    output wire                                          PEG_Xvec_6_ap_rst_n,
    output wire                                          PEG_Xvec_6_ap_start,
    output wire [                                 512:0] PEG_Xvec_6_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_6_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_6_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_6_fifo_A_s_dout,
    output wire                                          PEG_Xvec_6_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_6_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_6_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_6_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_6_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_6_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_6_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_6_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_6_fifo_X_out_din,
    output wire                                          PEG_Xvec_6_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_6_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_6_fifo_aXvec_din,
    output wire                                          PEG_Xvec_6_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_6_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_6_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_6_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_6_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_6_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_6_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_6_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_6_fifo_inst_out_din,
    output wire                                          PEG_Xvec_6_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_6_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_6_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_6_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_6_fifo_inst_out_write,
    output wire                                          PEG_Xvec_7_ap_clk,
    input wire                                           PEG_Xvec_7_ap_done,
    input wire                                           PEG_Xvec_7_ap_idle,
    input wire                                           PEG_Xvec_7_ap_ready,
    output wire                                          PEG_Xvec_7_ap_rst_n,
    output wire                                          PEG_Xvec_7_ap_start,
    output wire [                                 512:0] PEG_Xvec_7_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_7_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_7_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_7_fifo_A_s_dout,
    output wire                                          PEG_Xvec_7_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_7_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_7_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_7_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_7_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_7_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_7_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_7_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_7_fifo_X_out_din,
    output wire                                          PEG_Xvec_7_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_7_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_7_fifo_aXvec_din,
    output wire                                          PEG_Xvec_7_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_7_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_7_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_7_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_7_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_7_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_7_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_7_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_7_fifo_inst_out_din,
    output wire                                          PEG_Xvec_7_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_7_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_7_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_7_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_7_fifo_inst_out_write,
    output wire                                          PEG_Xvec_8_ap_clk,
    input wire                                           PEG_Xvec_8_ap_done,
    input wire                                           PEG_Xvec_8_ap_idle,
    input wire                                           PEG_Xvec_8_ap_ready,
    output wire                                          PEG_Xvec_8_ap_rst_n,
    output wire                                          PEG_Xvec_8_ap_start,
    output wire [                                 512:0] PEG_Xvec_8_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_8_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_8_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_8_fifo_A_s_dout,
    output wire                                          PEG_Xvec_8_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_8_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_8_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_8_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_8_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_8_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_8_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_8_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_8_fifo_X_out_din,
    output wire                                          PEG_Xvec_8_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_8_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_8_fifo_aXvec_din,
    output wire                                          PEG_Xvec_8_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_8_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_8_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_8_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_8_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_8_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_8_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_8_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_8_fifo_inst_out_din,
    output wire                                          PEG_Xvec_8_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_8_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_8_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_8_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_8_fifo_inst_out_write,
    output wire                                          PEG_Xvec_9_ap_clk,
    input wire                                           PEG_Xvec_9_ap_done,
    input wire                                           PEG_Xvec_9_ap_idle,
    input wire                                           PEG_Xvec_9_ap_ready,
    output wire                                          PEG_Xvec_9_ap_rst_n,
    output wire                                          PEG_Xvec_9_ap_start,
    output wire [                                 512:0] PEG_Xvec_9_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_9_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_9_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_9_fifo_A_s_dout,
    output wire                                          PEG_Xvec_9_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_9_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_9_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_9_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_9_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_9_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_9_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_9_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_9_fifo_X_out_din,
    output wire                                          PEG_Xvec_9_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_9_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_9_fifo_aXvec_din,
    output wire                                          PEG_Xvec_9_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_9_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_9_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_9_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_9_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_9_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_9_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_9_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_9_fifo_inst_out_din,
    output wire                                          PEG_Xvec_9_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_9_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_9_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_9_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_9_fifo_inst_out_write,
    output wire                                          PEG_Xvec_10_ap_clk,
    input wire                                           PEG_Xvec_10_ap_done,
    input wire                                           PEG_Xvec_10_ap_idle,
    input wire                                           PEG_Xvec_10_ap_ready,
    output wire                                          PEG_Xvec_10_ap_rst_n,
    output wire                                          PEG_Xvec_10_ap_start,
    output wire [                                 512:0] PEG_Xvec_10_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_10_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_10_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_10_fifo_A_s_dout,
    output wire                                          PEG_Xvec_10_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_10_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_10_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_10_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_10_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_10_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_10_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_10_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_10_fifo_X_out_din,
    output wire                                          PEG_Xvec_10_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_10_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_10_fifo_aXvec_din,
    output wire                                          PEG_Xvec_10_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_10_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_10_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_10_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_10_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_10_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_10_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_10_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_10_fifo_inst_out_din,
    output wire                                          PEG_Xvec_10_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_10_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_10_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_10_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_10_fifo_inst_out_write,
    output wire                                          PEG_Xvec_11_ap_clk,
    input wire                                           PEG_Xvec_11_ap_done,
    input wire                                           PEG_Xvec_11_ap_idle,
    input wire                                           PEG_Xvec_11_ap_ready,
    output wire                                          PEG_Xvec_11_ap_rst_n,
    output wire                                          PEG_Xvec_11_ap_start,
    output wire [                                 512:0] PEG_Xvec_11_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_11_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_11_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_11_fifo_A_s_dout,
    output wire                                          PEG_Xvec_11_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_11_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_11_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_11_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_11_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_11_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_11_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_11_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_11_fifo_X_out_din,
    output wire                                          PEG_Xvec_11_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_11_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_11_fifo_aXvec_din,
    output wire                                          PEG_Xvec_11_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_11_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_11_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_11_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_11_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_11_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_11_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_11_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_11_fifo_inst_out_din,
    output wire                                          PEG_Xvec_11_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_11_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_11_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_11_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_11_fifo_inst_out_write,
    output wire                                          PEG_Xvec_12_ap_clk,
    input wire                                           PEG_Xvec_12_ap_done,
    input wire                                           PEG_Xvec_12_ap_idle,
    input wire                                           PEG_Xvec_12_ap_ready,
    output wire                                          PEG_Xvec_12_ap_rst_n,
    output wire                                          PEG_Xvec_12_ap_start,
    output wire [                                 512:0] PEG_Xvec_12_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_12_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_12_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_12_fifo_A_s_dout,
    output wire                                          PEG_Xvec_12_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_12_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_12_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_12_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_12_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_12_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_12_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_12_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_12_fifo_X_out_din,
    output wire                                          PEG_Xvec_12_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_12_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_12_fifo_aXvec_din,
    output wire                                          PEG_Xvec_12_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_12_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_12_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_12_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_12_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_12_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_12_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_12_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_12_fifo_inst_out_din,
    output wire                                          PEG_Xvec_12_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_12_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_12_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_12_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_12_fifo_inst_out_write,
    output wire                                          PEG_Xvec_13_ap_clk,
    input wire                                           PEG_Xvec_13_ap_done,
    input wire                                           PEG_Xvec_13_ap_idle,
    input wire                                           PEG_Xvec_13_ap_ready,
    output wire                                          PEG_Xvec_13_ap_rst_n,
    output wire                                          PEG_Xvec_13_ap_start,
    output wire [                                 512:0] PEG_Xvec_13_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_13_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_13_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_13_fifo_A_s_dout,
    output wire                                          PEG_Xvec_13_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_13_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_13_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_13_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_13_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_13_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_13_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_13_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_13_fifo_X_out_din,
    output wire                                          PEG_Xvec_13_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_13_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_13_fifo_aXvec_din,
    output wire                                          PEG_Xvec_13_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_13_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_13_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_13_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_13_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_13_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_13_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_13_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_13_fifo_inst_out_din,
    output wire                                          PEG_Xvec_13_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_13_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_13_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_13_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_13_fifo_inst_out_write,
    output wire                                          PEG_Xvec_14_ap_clk,
    input wire                                           PEG_Xvec_14_ap_done,
    input wire                                           PEG_Xvec_14_ap_idle,
    input wire                                           PEG_Xvec_14_ap_ready,
    output wire                                          PEG_Xvec_14_ap_rst_n,
    output wire                                          PEG_Xvec_14_ap_start,
    output wire [                                 512:0] PEG_Xvec_14_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_14_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_14_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_14_fifo_A_s_dout,
    output wire                                          PEG_Xvec_14_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_14_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_14_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_14_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_14_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_14_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_14_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_14_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_14_fifo_X_out_din,
    output wire                                          PEG_Xvec_14_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_14_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_14_fifo_aXvec_din,
    output wire                                          PEG_Xvec_14_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_14_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_14_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_14_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_14_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_14_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_14_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_14_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_14_fifo_inst_out_din,
    output wire                                          PEG_Xvec_14_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_14_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_14_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_14_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_14_fifo_inst_out_write,
    output wire                                          PEG_Xvec_15_ap_clk,
    input wire                                           PEG_Xvec_15_ap_done,
    input wire                                           PEG_Xvec_15_ap_idle,
    input wire                                           PEG_Xvec_15_ap_ready,
    output wire                                          PEG_Xvec_15_ap_rst_n,
    output wire                                          PEG_Xvec_15_ap_start,
    output wire [                                 512:0] PEG_Xvec_15_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_15_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_15_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_15_fifo_A_s_dout,
    output wire                                          PEG_Xvec_15_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_15_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_15_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_15_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_15_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_15_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_15_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_15_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_15_fifo_X_out_din,
    output wire                                          PEG_Xvec_15_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_15_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_15_fifo_aXvec_din,
    output wire                                          PEG_Xvec_15_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_15_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_15_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_15_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_15_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_15_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_15_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_15_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_15_fifo_inst_out_din,
    output wire                                          PEG_Xvec_15_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_15_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_15_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_15_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_15_fifo_inst_out_write,
    output wire                                          PEG_Xvec_16_ap_clk,
    input wire                                           PEG_Xvec_16_ap_done,
    input wire                                           PEG_Xvec_16_ap_idle,
    input wire                                           PEG_Xvec_16_ap_ready,
    output wire                                          PEG_Xvec_16_ap_rst_n,
    output wire                                          PEG_Xvec_16_ap_start,
    output wire [                                 512:0] PEG_Xvec_16_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_16_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_16_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_16_fifo_A_s_dout,
    output wire                                          PEG_Xvec_16_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_16_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_16_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_16_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_16_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_16_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_16_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_16_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_16_fifo_X_out_din,
    output wire                                          PEG_Xvec_16_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_16_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_16_fifo_aXvec_din,
    output wire                                          PEG_Xvec_16_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_16_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_16_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_16_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_16_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_16_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_16_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_16_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_16_fifo_inst_out_din,
    output wire                                          PEG_Xvec_16_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_16_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_16_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_16_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_16_fifo_inst_out_write,
    output wire                                          PEG_Xvec_17_ap_clk,
    input wire                                           PEG_Xvec_17_ap_done,
    input wire                                           PEG_Xvec_17_ap_idle,
    input wire                                           PEG_Xvec_17_ap_ready,
    output wire                                          PEG_Xvec_17_ap_rst_n,
    output wire                                          PEG_Xvec_17_ap_start,
    output wire [                                 512:0] PEG_Xvec_17_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_17_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_17_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_17_fifo_A_s_dout,
    output wire                                          PEG_Xvec_17_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_17_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_17_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_17_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_17_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_17_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_17_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_17_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_17_fifo_X_out_din,
    output wire                                          PEG_Xvec_17_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_17_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_17_fifo_aXvec_din,
    output wire                                          PEG_Xvec_17_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_17_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_17_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_17_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_17_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_17_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_17_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_17_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_17_fifo_inst_out_din,
    output wire                                          PEG_Xvec_17_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_17_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_17_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_17_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_17_fifo_inst_out_write,
    output wire                                          PEG_Xvec_18_ap_clk,
    input wire                                           PEG_Xvec_18_ap_done,
    input wire                                           PEG_Xvec_18_ap_idle,
    input wire                                           PEG_Xvec_18_ap_ready,
    output wire                                          PEG_Xvec_18_ap_rst_n,
    output wire                                          PEG_Xvec_18_ap_start,
    output wire [                                 512:0] PEG_Xvec_18_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_18_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_18_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_18_fifo_A_s_dout,
    output wire                                          PEG_Xvec_18_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_18_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_18_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_18_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_18_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_18_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_18_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_18_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_18_fifo_X_out_din,
    output wire                                          PEG_Xvec_18_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_18_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_18_fifo_aXvec_din,
    output wire                                          PEG_Xvec_18_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_18_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_18_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_18_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_18_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_18_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_18_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_18_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_18_fifo_inst_out_din,
    output wire                                          PEG_Xvec_18_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_18_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_18_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_18_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_18_fifo_inst_out_write,
    output wire                                          PEG_Xvec_19_ap_clk,
    input wire                                           PEG_Xvec_19_ap_done,
    input wire                                           PEG_Xvec_19_ap_idle,
    input wire                                           PEG_Xvec_19_ap_ready,
    output wire                                          PEG_Xvec_19_ap_rst_n,
    output wire                                          PEG_Xvec_19_ap_start,
    output wire [                                 512:0] PEG_Xvec_19_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_19_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_19_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_19_fifo_A_s_dout,
    output wire                                          PEG_Xvec_19_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_19_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_19_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_19_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_19_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_19_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_19_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_19_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_19_fifo_X_out_din,
    output wire                                          PEG_Xvec_19_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_19_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_19_fifo_aXvec_din,
    output wire                                          PEG_Xvec_19_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_19_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_19_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_19_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_19_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_19_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_19_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_19_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_19_fifo_inst_out_din,
    output wire                                          PEG_Xvec_19_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_19_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_19_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_19_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_19_fifo_inst_out_write,
    output wire                                          PEG_Xvec_20_ap_clk,
    input wire                                           PEG_Xvec_20_ap_done,
    input wire                                           PEG_Xvec_20_ap_idle,
    input wire                                           PEG_Xvec_20_ap_ready,
    output wire                                          PEG_Xvec_20_ap_rst_n,
    output wire                                          PEG_Xvec_20_ap_start,
    output wire [                                 512:0] PEG_Xvec_20_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_20_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_20_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_20_fifo_A_s_dout,
    output wire                                          PEG_Xvec_20_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_20_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_20_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_20_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_20_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_20_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_20_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_20_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_20_fifo_X_out_din,
    output wire                                          PEG_Xvec_20_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_20_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_20_fifo_aXvec_din,
    output wire                                          PEG_Xvec_20_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_20_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_20_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_20_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_20_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_20_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_20_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_20_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_20_fifo_inst_out_din,
    output wire                                          PEG_Xvec_20_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_20_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_20_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_20_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_20_fifo_inst_out_write,
    output wire                                          PEG_Xvec_21_ap_clk,
    input wire                                           PEG_Xvec_21_ap_done,
    input wire                                           PEG_Xvec_21_ap_idle,
    input wire                                           PEG_Xvec_21_ap_ready,
    output wire                                          PEG_Xvec_21_ap_rst_n,
    output wire                                          PEG_Xvec_21_ap_start,
    output wire [                                 512:0] PEG_Xvec_21_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_21_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_21_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_21_fifo_A_s_dout,
    output wire                                          PEG_Xvec_21_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_21_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_21_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_21_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_21_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_21_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_21_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_21_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_21_fifo_X_out_din,
    output wire                                          PEG_Xvec_21_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_21_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_21_fifo_aXvec_din,
    output wire                                          PEG_Xvec_21_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_21_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_21_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_21_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_21_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_21_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_21_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_21_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_21_fifo_inst_out_din,
    output wire                                          PEG_Xvec_21_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_21_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_21_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_21_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_21_fifo_inst_out_write,
    output wire                                          PEG_Xvec_22_ap_clk,
    input wire                                           PEG_Xvec_22_ap_done,
    input wire                                           PEG_Xvec_22_ap_idle,
    input wire                                           PEG_Xvec_22_ap_ready,
    output wire                                          PEG_Xvec_22_ap_rst_n,
    output wire                                          PEG_Xvec_22_ap_start,
    output wire [                                 512:0] PEG_Xvec_22_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_22_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_22_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_22_fifo_A_s_dout,
    output wire                                          PEG_Xvec_22_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_22_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_22_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_22_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_22_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_22_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_22_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_22_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_22_fifo_X_out_din,
    output wire                                          PEG_Xvec_22_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_22_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_22_fifo_aXvec_din,
    output wire                                          PEG_Xvec_22_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_22_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_22_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_22_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_22_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_22_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_22_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_22_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_22_fifo_inst_out_din,
    output wire                                          PEG_Xvec_22_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_22_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_22_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_22_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_22_fifo_inst_out_write,
    output wire                                          PEG_Xvec_23_ap_clk,
    input wire                                           PEG_Xvec_23_ap_done,
    input wire                                           PEG_Xvec_23_ap_idle,
    input wire                                           PEG_Xvec_23_ap_ready,
    output wire                                          PEG_Xvec_23_ap_rst_n,
    output wire                                          PEG_Xvec_23_ap_start,
    output wire [                                 512:0] PEG_Xvec_23_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_23_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_23_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_23_fifo_A_s_dout,
    output wire                                          PEG_Xvec_23_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_23_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_23_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_23_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_23_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_23_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_23_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_23_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_23_fifo_X_out_din,
    output wire                                          PEG_Xvec_23_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_23_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_23_fifo_aXvec_din,
    output wire                                          PEG_Xvec_23_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_23_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_23_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_23_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_23_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_23_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_23_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_23_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_23_fifo_inst_out_din,
    output wire                                          PEG_Xvec_23_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_23_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_23_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_23_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_23_fifo_inst_out_write,
    output wire                                          PEG_Xvec_24_ap_clk,
    input wire                                           PEG_Xvec_24_ap_done,
    input wire                                           PEG_Xvec_24_ap_idle,
    input wire                                           PEG_Xvec_24_ap_ready,
    output wire                                          PEG_Xvec_24_ap_rst_n,
    output wire                                          PEG_Xvec_24_ap_start,
    output wire [                                 512:0] PEG_Xvec_24_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_24_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_24_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_24_fifo_A_s_dout,
    output wire                                          PEG_Xvec_24_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_24_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_24_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_24_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_24_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_24_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_24_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_24_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_24_fifo_X_out_din,
    output wire                                          PEG_Xvec_24_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_24_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_24_fifo_aXvec_din,
    output wire                                          PEG_Xvec_24_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_24_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_24_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_24_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_24_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_24_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_24_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_24_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_24_fifo_inst_out_din,
    output wire                                          PEG_Xvec_24_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_24_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_24_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_24_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_24_fifo_inst_out_write,
    output wire                                          PEG_Xvec_25_ap_clk,
    input wire                                           PEG_Xvec_25_ap_done,
    input wire                                           PEG_Xvec_25_ap_idle,
    input wire                                           PEG_Xvec_25_ap_ready,
    output wire                                          PEG_Xvec_25_ap_rst_n,
    output wire                                          PEG_Xvec_25_ap_start,
    output wire [                                 512:0] PEG_Xvec_25_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_25_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_25_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_25_fifo_A_s_dout,
    output wire                                          PEG_Xvec_25_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_25_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_25_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_25_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_25_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_25_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_25_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_25_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_25_fifo_X_out_din,
    output wire                                          PEG_Xvec_25_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_25_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_25_fifo_aXvec_din,
    output wire                                          PEG_Xvec_25_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_25_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_25_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_25_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_25_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_25_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_25_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_25_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_25_fifo_inst_out_din,
    output wire                                          PEG_Xvec_25_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_25_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_25_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_25_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_25_fifo_inst_out_write,
    output wire                                          PEG_Xvec_26_ap_clk,
    input wire                                           PEG_Xvec_26_ap_done,
    input wire                                           PEG_Xvec_26_ap_idle,
    input wire                                           PEG_Xvec_26_ap_ready,
    output wire                                          PEG_Xvec_26_ap_rst_n,
    output wire                                          PEG_Xvec_26_ap_start,
    output wire [                                 512:0] PEG_Xvec_26_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_26_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_26_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_26_fifo_A_s_dout,
    output wire                                          PEG_Xvec_26_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_26_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_26_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_26_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_26_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_26_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_26_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_26_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_26_fifo_X_out_din,
    output wire                                          PEG_Xvec_26_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_26_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_26_fifo_aXvec_din,
    output wire                                          PEG_Xvec_26_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_26_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_26_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_26_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_26_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_26_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_26_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_26_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_26_fifo_inst_out_din,
    output wire                                          PEG_Xvec_26_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_26_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_26_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_26_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_26_fifo_inst_out_write,
    output wire                                          PEG_Xvec_27_ap_clk,
    input wire                                           PEG_Xvec_27_ap_done,
    input wire                                           PEG_Xvec_27_ap_idle,
    input wire                                           PEG_Xvec_27_ap_ready,
    output wire                                          PEG_Xvec_27_ap_rst_n,
    output wire                                          PEG_Xvec_27_ap_start,
    output wire [                                 512:0] PEG_Xvec_27_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_27_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_27_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_27_fifo_A_s_dout,
    output wire                                          PEG_Xvec_27_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_27_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_27_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_27_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_27_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_27_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_27_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_27_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_27_fifo_X_out_din,
    output wire                                          PEG_Xvec_27_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_27_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_27_fifo_aXvec_din,
    output wire                                          PEG_Xvec_27_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_27_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_27_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_27_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_27_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_27_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_27_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_27_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_27_fifo_inst_out_din,
    output wire                                          PEG_Xvec_27_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_27_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_27_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_27_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_27_fifo_inst_out_write,
    output wire                                          PEG_Xvec_28_ap_clk,
    input wire                                           PEG_Xvec_28_ap_done,
    input wire                                           PEG_Xvec_28_ap_idle,
    input wire                                           PEG_Xvec_28_ap_ready,
    output wire                                          PEG_Xvec_28_ap_rst_n,
    output wire                                          PEG_Xvec_28_ap_start,
    output wire [                                 512:0] PEG_Xvec_28_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_28_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_28_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_28_fifo_A_s_dout,
    output wire                                          PEG_Xvec_28_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_28_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_28_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_28_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_28_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_28_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_28_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_28_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_28_fifo_X_out_din,
    output wire                                          PEG_Xvec_28_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_28_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_28_fifo_aXvec_din,
    output wire                                          PEG_Xvec_28_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_28_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_28_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_28_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_28_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_28_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_28_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_28_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_28_fifo_inst_out_din,
    output wire                                          PEG_Xvec_28_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_28_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_28_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_28_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_28_fifo_inst_out_write,
    output wire                                          PEG_Xvec_29_ap_clk,
    input wire                                           PEG_Xvec_29_ap_done,
    input wire                                           PEG_Xvec_29_ap_idle,
    input wire                                           PEG_Xvec_29_ap_ready,
    output wire                                          PEG_Xvec_29_ap_rst_n,
    output wire                                          PEG_Xvec_29_ap_start,
    output wire [                                 512:0] PEG_Xvec_29_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_29_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_29_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_29_fifo_A_s_dout,
    output wire                                          PEG_Xvec_29_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_29_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_29_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_29_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_29_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_29_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_29_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_29_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_29_fifo_X_out_din,
    output wire                                          PEG_Xvec_29_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_29_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_29_fifo_aXvec_din,
    output wire                                          PEG_Xvec_29_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_29_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_29_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_29_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_29_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_29_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_29_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_29_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_29_fifo_inst_out_din,
    output wire                                          PEG_Xvec_29_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_29_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_29_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_29_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_29_fifo_inst_out_write,
    output wire                                          PEG_Xvec_30_ap_clk,
    input wire                                           PEG_Xvec_30_ap_done,
    input wire                                           PEG_Xvec_30_ap_idle,
    input wire                                           PEG_Xvec_30_ap_ready,
    output wire                                          PEG_Xvec_30_ap_rst_n,
    output wire                                          PEG_Xvec_30_ap_start,
    output wire [                                 512:0] PEG_Xvec_30_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_30_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_30_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_30_fifo_A_s_dout,
    output wire                                          PEG_Xvec_30_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_30_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_30_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_30_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_30_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_30_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_30_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_30_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_30_fifo_X_out_din,
    output wire                                          PEG_Xvec_30_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_30_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_30_fifo_aXvec_din,
    output wire                                          PEG_Xvec_30_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_30_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_30_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_30_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_30_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_30_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_30_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_30_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_30_fifo_inst_out_din,
    output wire                                          PEG_Xvec_30_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_30_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_30_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_30_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_30_fifo_inst_out_write,
    output wire                                          PEG_Xvec_31_ap_clk,
    input wire                                           PEG_Xvec_31_ap_done,
    input wire                                           PEG_Xvec_31_ap_idle,
    input wire                                           PEG_Xvec_31_ap_ready,
    output wire                                          PEG_Xvec_31_ap_rst_n,
    output wire                                          PEG_Xvec_31_ap_start,
    output wire [                                 512:0] PEG_Xvec_31_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_31_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_31_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_31_fifo_A_s_dout,
    output wire                                          PEG_Xvec_31_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_31_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_31_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_31_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_31_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_31_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_31_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_31_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_31_fifo_X_out_din,
    output wire                                          PEG_Xvec_31_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_31_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_31_fifo_aXvec_din,
    output wire                                          PEG_Xvec_31_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_31_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_31_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_31_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_31_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_31_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_31_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_31_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_31_fifo_inst_out_din,
    output wire                                          PEG_Xvec_31_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_31_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_31_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_31_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_31_fifo_inst_out_write,
    output wire                                          PEG_Xvec_32_ap_clk,
    input wire                                           PEG_Xvec_32_ap_done,
    input wire                                           PEG_Xvec_32_ap_idle,
    input wire                                           PEG_Xvec_32_ap_ready,
    output wire                                          PEG_Xvec_32_ap_rst_n,
    output wire                                          PEG_Xvec_32_ap_start,
    output wire [                                 512:0] PEG_Xvec_32_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_32_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_32_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_32_fifo_A_s_dout,
    output wire                                          PEG_Xvec_32_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_32_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_32_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_32_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_32_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_32_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_32_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_32_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_32_fifo_X_out_din,
    output wire                                          PEG_Xvec_32_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_32_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_32_fifo_aXvec_din,
    output wire                                          PEG_Xvec_32_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_32_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_32_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_32_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_32_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_32_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_32_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_32_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_32_fifo_inst_out_din,
    output wire                                          PEG_Xvec_32_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_32_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_32_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_32_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_32_fifo_inst_out_write,
    output wire                                          PEG_Xvec_33_ap_clk,
    input wire                                           PEG_Xvec_33_ap_done,
    input wire                                           PEG_Xvec_33_ap_idle,
    input wire                                           PEG_Xvec_33_ap_ready,
    output wire                                          PEG_Xvec_33_ap_rst_n,
    output wire                                          PEG_Xvec_33_ap_start,
    output wire [                                 512:0] PEG_Xvec_33_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_33_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_33_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_33_fifo_A_s_dout,
    output wire                                          PEG_Xvec_33_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_33_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_33_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_33_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_33_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_33_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_33_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_33_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_33_fifo_X_out_din,
    output wire                                          PEG_Xvec_33_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_33_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_33_fifo_aXvec_din,
    output wire                                          PEG_Xvec_33_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_33_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_33_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_33_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_33_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_33_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_33_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_33_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_33_fifo_inst_out_din,
    output wire                                          PEG_Xvec_33_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_33_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_33_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_33_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_33_fifo_inst_out_write,
    output wire                                          PEG_Xvec_34_ap_clk,
    input wire                                           PEG_Xvec_34_ap_done,
    input wire                                           PEG_Xvec_34_ap_idle,
    input wire                                           PEG_Xvec_34_ap_ready,
    output wire                                          PEG_Xvec_34_ap_rst_n,
    output wire                                          PEG_Xvec_34_ap_start,
    output wire [                                 512:0] PEG_Xvec_34_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_34_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_34_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_34_fifo_A_s_dout,
    output wire                                          PEG_Xvec_34_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_34_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_34_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_34_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_34_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_34_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_34_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_34_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_34_fifo_X_out_din,
    output wire                                          PEG_Xvec_34_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_34_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_34_fifo_aXvec_din,
    output wire                                          PEG_Xvec_34_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_34_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_34_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_34_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_34_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_34_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_34_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_34_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_34_fifo_inst_out_din,
    output wire                                          PEG_Xvec_34_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_34_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_34_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_34_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_34_fifo_inst_out_write,
    output wire                                          PEG_Xvec_35_ap_clk,
    input wire                                           PEG_Xvec_35_ap_done,
    input wire                                           PEG_Xvec_35_ap_idle,
    input wire                                           PEG_Xvec_35_ap_ready,
    output wire                                          PEG_Xvec_35_ap_rst_n,
    output wire                                          PEG_Xvec_35_ap_start,
    output wire [                                 512:0] PEG_Xvec_35_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_35_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_35_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_35_fifo_A_s_dout,
    output wire                                          PEG_Xvec_35_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_35_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_35_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_35_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_35_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_35_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_35_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_35_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_35_fifo_X_out_din,
    output wire                                          PEG_Xvec_35_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_35_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_35_fifo_aXvec_din,
    output wire                                          PEG_Xvec_35_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_35_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_35_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_35_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_35_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_35_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_35_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_35_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_35_fifo_inst_out_din,
    output wire                                          PEG_Xvec_35_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_35_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_35_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_35_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_35_fifo_inst_out_write,
    output wire                                          PEG_Xvec_36_ap_clk,
    input wire                                           PEG_Xvec_36_ap_done,
    input wire                                           PEG_Xvec_36_ap_idle,
    input wire                                           PEG_Xvec_36_ap_ready,
    output wire                                          PEG_Xvec_36_ap_rst_n,
    output wire                                          PEG_Xvec_36_ap_start,
    output wire [                                 512:0] PEG_Xvec_36_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_36_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_36_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_36_fifo_A_s_dout,
    output wire                                          PEG_Xvec_36_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_36_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_36_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_36_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_36_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_36_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_36_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_36_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_36_fifo_X_out_din,
    output wire                                          PEG_Xvec_36_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_36_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_36_fifo_aXvec_din,
    output wire                                          PEG_Xvec_36_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_36_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_36_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_36_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_36_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_36_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_36_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_36_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_36_fifo_inst_out_din,
    output wire                                          PEG_Xvec_36_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_36_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_36_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_36_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_36_fifo_inst_out_write,
    output wire                                          PEG_Xvec_37_ap_clk,
    input wire                                           PEG_Xvec_37_ap_done,
    input wire                                           PEG_Xvec_37_ap_idle,
    input wire                                           PEG_Xvec_37_ap_ready,
    output wire                                          PEG_Xvec_37_ap_rst_n,
    output wire                                          PEG_Xvec_37_ap_start,
    output wire [                                 512:0] PEG_Xvec_37_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_37_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_37_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_37_fifo_A_s_dout,
    output wire                                          PEG_Xvec_37_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_37_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_37_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_37_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_37_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_37_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_37_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_37_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_37_fifo_X_out_din,
    output wire                                          PEG_Xvec_37_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_37_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_37_fifo_aXvec_din,
    output wire                                          PEG_Xvec_37_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_37_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_37_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_37_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_37_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_37_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_37_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_37_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_37_fifo_inst_out_din,
    output wire                                          PEG_Xvec_37_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_37_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_37_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_37_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_37_fifo_inst_out_write,
    output wire                                          PEG_Xvec_38_ap_clk,
    input wire                                           PEG_Xvec_38_ap_done,
    input wire                                           PEG_Xvec_38_ap_idle,
    input wire                                           PEG_Xvec_38_ap_ready,
    output wire                                          PEG_Xvec_38_ap_rst_n,
    output wire                                          PEG_Xvec_38_ap_start,
    output wire [                                 512:0] PEG_Xvec_38_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_38_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_38_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_38_fifo_A_s_dout,
    output wire                                          PEG_Xvec_38_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_38_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_38_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_38_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_38_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_38_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_38_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_38_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_38_fifo_X_out_din,
    output wire                                          PEG_Xvec_38_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_38_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_38_fifo_aXvec_din,
    output wire                                          PEG_Xvec_38_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_38_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_38_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_38_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_38_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_38_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_38_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_38_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_38_fifo_inst_out_din,
    output wire                                          PEG_Xvec_38_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_38_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_38_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_38_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_38_fifo_inst_out_write,
    output wire                                          PEG_Xvec_39_ap_clk,
    input wire                                           PEG_Xvec_39_ap_done,
    input wire                                           PEG_Xvec_39_ap_idle,
    input wire                                           PEG_Xvec_39_ap_ready,
    output wire                                          PEG_Xvec_39_ap_rst_n,
    output wire                                          PEG_Xvec_39_ap_start,
    output wire [                                 512:0] PEG_Xvec_39_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_39_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_39_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_39_fifo_A_s_dout,
    output wire                                          PEG_Xvec_39_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_39_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_39_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_39_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_39_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_39_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_39_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_39_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_39_fifo_X_out_din,
    output wire                                          PEG_Xvec_39_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_39_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_39_fifo_aXvec_din,
    output wire                                          PEG_Xvec_39_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_39_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_39_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_39_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_39_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_39_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_39_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_39_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_39_fifo_inst_out_din,
    output wire                                          PEG_Xvec_39_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_39_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_39_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_39_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_39_fifo_inst_out_write,
    output wire                                          PEG_Xvec_40_ap_clk,
    input wire                                           PEG_Xvec_40_ap_done,
    input wire                                           PEG_Xvec_40_ap_idle,
    input wire                                           PEG_Xvec_40_ap_ready,
    output wire                                          PEG_Xvec_40_ap_rst_n,
    output wire                                          PEG_Xvec_40_ap_start,
    output wire [                                 512:0] PEG_Xvec_40_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_40_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_40_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_40_fifo_A_s_dout,
    output wire                                          PEG_Xvec_40_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_40_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_40_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_40_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_40_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_40_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_40_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_40_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_40_fifo_X_out_din,
    output wire                                          PEG_Xvec_40_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_40_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_40_fifo_aXvec_din,
    output wire                                          PEG_Xvec_40_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_40_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_40_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_40_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_40_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_40_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_40_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_40_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_40_fifo_inst_out_din,
    output wire                                          PEG_Xvec_40_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_40_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_40_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_40_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_40_fifo_inst_out_write,
    output wire                                          PEG_Xvec_41_ap_clk,
    input wire                                           PEG_Xvec_41_ap_done,
    input wire                                           PEG_Xvec_41_ap_idle,
    input wire                                           PEG_Xvec_41_ap_ready,
    output wire                                          PEG_Xvec_41_ap_rst_n,
    output wire                                          PEG_Xvec_41_ap_start,
    output wire [                                 512:0] PEG_Xvec_41_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_41_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_41_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_41_fifo_A_s_dout,
    output wire                                          PEG_Xvec_41_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_41_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_41_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_41_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_41_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_41_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_41_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_41_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_41_fifo_X_out_din,
    output wire                                          PEG_Xvec_41_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_41_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_41_fifo_aXvec_din,
    output wire                                          PEG_Xvec_41_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_41_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_41_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_41_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_41_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_41_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_41_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_41_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_41_fifo_inst_out_din,
    output wire                                          PEG_Xvec_41_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_41_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_41_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_41_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_41_fifo_inst_out_write,
    output wire                                          PEG_Xvec_42_ap_clk,
    input wire                                           PEG_Xvec_42_ap_done,
    input wire                                           PEG_Xvec_42_ap_idle,
    input wire                                           PEG_Xvec_42_ap_ready,
    output wire                                          PEG_Xvec_42_ap_rst_n,
    output wire                                          PEG_Xvec_42_ap_start,
    output wire [                                 512:0] PEG_Xvec_42_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_42_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_42_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_42_fifo_A_s_dout,
    output wire                                          PEG_Xvec_42_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_42_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_42_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_42_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_42_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_42_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_42_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_42_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_42_fifo_X_out_din,
    output wire                                          PEG_Xvec_42_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_42_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_42_fifo_aXvec_din,
    output wire                                          PEG_Xvec_42_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_42_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_42_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_42_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_42_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_42_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_42_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_42_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_42_fifo_inst_out_din,
    output wire                                          PEG_Xvec_42_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_42_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_42_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_42_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_42_fifo_inst_out_write,
    output wire                                          PEG_Xvec_43_ap_clk,
    input wire                                           PEG_Xvec_43_ap_done,
    input wire                                           PEG_Xvec_43_ap_idle,
    input wire                                           PEG_Xvec_43_ap_ready,
    output wire                                          PEG_Xvec_43_ap_rst_n,
    output wire                                          PEG_Xvec_43_ap_start,
    output wire [                                 512:0] PEG_Xvec_43_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_43_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_43_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_43_fifo_A_s_dout,
    output wire                                          PEG_Xvec_43_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_43_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_43_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_43_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_43_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_43_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_43_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_43_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_43_fifo_X_out_din,
    output wire                                          PEG_Xvec_43_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_43_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_43_fifo_aXvec_din,
    output wire                                          PEG_Xvec_43_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_43_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_43_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_43_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_43_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_43_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_43_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_43_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_43_fifo_inst_out_din,
    output wire                                          PEG_Xvec_43_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_43_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_43_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_43_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_43_fifo_inst_out_write,
    output wire                                          PEG_Xvec_44_ap_clk,
    input wire                                           PEG_Xvec_44_ap_done,
    input wire                                           PEG_Xvec_44_ap_idle,
    input wire                                           PEG_Xvec_44_ap_ready,
    output wire                                          PEG_Xvec_44_ap_rst_n,
    output wire                                          PEG_Xvec_44_ap_start,
    output wire [                                 512:0] PEG_Xvec_44_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_44_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_44_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_44_fifo_A_s_dout,
    output wire                                          PEG_Xvec_44_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_44_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_44_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_44_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_44_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_44_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_44_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_44_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_44_fifo_X_out_din,
    output wire                                          PEG_Xvec_44_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_44_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_44_fifo_aXvec_din,
    output wire                                          PEG_Xvec_44_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_44_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_44_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_44_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_44_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_44_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_44_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_44_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_44_fifo_inst_out_din,
    output wire                                          PEG_Xvec_44_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_44_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_44_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_44_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_44_fifo_inst_out_write,
    output wire                                          PEG_Xvec_45_ap_clk,
    input wire                                           PEG_Xvec_45_ap_done,
    input wire                                           PEG_Xvec_45_ap_idle,
    input wire                                           PEG_Xvec_45_ap_ready,
    output wire                                          PEG_Xvec_45_ap_rst_n,
    output wire                                          PEG_Xvec_45_ap_start,
    output wire [                                 512:0] PEG_Xvec_45_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_45_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_45_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_45_fifo_A_s_dout,
    output wire                                          PEG_Xvec_45_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_45_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_45_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_45_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_45_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_45_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_45_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_45_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_45_fifo_X_out_din,
    output wire                                          PEG_Xvec_45_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_45_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_45_fifo_aXvec_din,
    output wire                                          PEG_Xvec_45_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_45_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_45_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_45_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_45_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_45_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_45_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_45_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_45_fifo_inst_out_din,
    output wire                                          PEG_Xvec_45_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_45_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_45_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_45_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_45_fifo_inst_out_write,
    output wire                                          PEG_Xvec_46_ap_clk,
    input wire                                           PEG_Xvec_46_ap_done,
    input wire                                           PEG_Xvec_46_ap_idle,
    input wire                                           PEG_Xvec_46_ap_ready,
    output wire                                          PEG_Xvec_46_ap_rst_n,
    output wire                                          PEG_Xvec_46_ap_start,
    output wire [                                 512:0] PEG_Xvec_46_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_46_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_46_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_46_fifo_A_s_dout,
    output wire                                          PEG_Xvec_46_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_46_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_46_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_46_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_46_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_46_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_46_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_46_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_46_fifo_X_out_din,
    output wire                                          PEG_Xvec_46_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_46_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_46_fifo_aXvec_din,
    output wire                                          PEG_Xvec_46_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_46_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_46_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_46_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_46_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_46_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_46_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_46_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_46_fifo_inst_out_din,
    output wire                                          PEG_Xvec_46_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_46_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_46_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_46_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_46_fifo_inst_out_write,
    output wire                                          PEG_Xvec_47_ap_clk,
    input wire                                           PEG_Xvec_47_ap_done,
    input wire                                           PEG_Xvec_47_ap_idle,
    input wire                                           PEG_Xvec_47_ap_ready,
    output wire                                          PEG_Xvec_47_ap_rst_n,
    output wire                                          PEG_Xvec_47_ap_start,
    output wire [                                 512:0] PEG_Xvec_47_fifo_A_peek_dout,
    output wire                                          PEG_Xvec_47_fifo_A_peek_empty_n,
    input wire                                           PEG_Xvec_47_fifo_A_peek_read,
    output wire [                                 512:0] PEG_Xvec_47_fifo_A_s_dout,
    output wire                                          PEG_Xvec_47_fifo_A_s_empty_n,
    input wire                                           PEG_Xvec_47_fifo_A_s_read,
    output wire [                                 512:0] PEG_Xvec_47_fifo_X_in_peek_dout,
    output wire                                          PEG_Xvec_47_fifo_X_in_peek_empty_n,
    input wire                                           PEG_Xvec_47_fifo_X_in_peek_read,
    output wire [                                 512:0] PEG_Xvec_47_fifo_X_in_s_dout,
    output wire                                          PEG_Xvec_47_fifo_X_in_s_empty_n,
    input wire                                           PEG_Xvec_47_fifo_X_in_s_read,
    input wire  [                                 512:0] PEG_Xvec_47_fifo_X_out_din,
    output wire                                          PEG_Xvec_47_fifo_X_out_full_n,
    input wire                                           PEG_Xvec_47_fifo_X_out_write,
    input wire  [                                 400:0] PEG_Xvec_47_fifo_aXvec_din,
    output wire                                          PEG_Xvec_47_fifo_aXvec_full_n,
    input wire                                           PEG_Xvec_47_fifo_aXvec_write,
    output wire [                                  32:0] PEG_Xvec_47_fifo_inst_in_peek_dout,
    output wire                                          PEG_Xvec_47_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Xvec_47_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Xvec_47_fifo_inst_in_s_dout,
    output wire                                          PEG_Xvec_47_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Xvec_47_fifo_inst_in_s_read,
    input wire  [                                  32:0] PEG_Xvec_47_fifo_inst_out_din,
    output wire                                          PEG_Xvec_47_fifo_inst_out_full_n,
    input wire  [                                  32:0] PEG_Xvec_47_fifo_inst_out_to_Yvec_din,
    output wire                                          PEG_Xvec_47_fifo_inst_out_to_Yvec_full_n,
    input wire                                           PEG_Xvec_47_fifo_inst_out_to_Yvec_write,
    input wire                                           PEG_Xvec_47_fifo_inst_out_write,
    output wire                                          PEG_Yvec_0_ap_clk,
    input wire                                           PEG_Yvec_0_ap_done,
    input wire                                           PEG_Yvec_0_ap_idle,
    input wire                                           PEG_Yvec_0_ap_ready,
    output wire                                          PEG_Yvec_0_ap_rst_n,
    output wire                                          PEG_Yvec_0_ap_start,
    input wire  [                                  64:0] PEG_Yvec_0_fifo_Y_out_din,
    output wire                                          PEG_Yvec_0_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_0_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_0_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_0_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_0_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_0_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_0_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_0_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_0_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_0_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_0_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_0_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_0_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_0_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_1_ap_clk,
    input wire                                           PEG_Yvec_1_ap_done,
    input wire                                           PEG_Yvec_1_ap_idle,
    input wire                                           PEG_Yvec_1_ap_ready,
    output wire                                          PEG_Yvec_1_ap_rst_n,
    output wire                                          PEG_Yvec_1_ap_start,
    input wire  [                                  64:0] PEG_Yvec_1_fifo_Y_out_din,
    output wire                                          PEG_Yvec_1_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_1_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_1_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_1_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_1_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_1_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_1_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_1_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_1_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_1_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_1_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_1_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_1_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_1_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_2_ap_clk,
    input wire                                           PEG_Yvec_2_ap_done,
    input wire                                           PEG_Yvec_2_ap_idle,
    input wire                                           PEG_Yvec_2_ap_ready,
    output wire                                          PEG_Yvec_2_ap_rst_n,
    output wire                                          PEG_Yvec_2_ap_start,
    input wire  [                                  64:0] PEG_Yvec_2_fifo_Y_out_din,
    output wire                                          PEG_Yvec_2_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_2_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_2_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_2_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_2_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_2_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_2_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_2_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_2_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_2_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_2_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_2_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_2_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_2_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_3_ap_clk,
    input wire                                           PEG_Yvec_3_ap_done,
    input wire                                           PEG_Yvec_3_ap_idle,
    input wire                                           PEG_Yvec_3_ap_ready,
    output wire                                          PEG_Yvec_3_ap_rst_n,
    output wire                                          PEG_Yvec_3_ap_start,
    input wire  [                                  64:0] PEG_Yvec_3_fifo_Y_out_din,
    output wire                                          PEG_Yvec_3_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_3_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_3_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_3_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_3_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_3_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_3_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_3_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_3_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_3_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_3_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_3_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_3_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_3_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_4_ap_clk,
    input wire                                           PEG_Yvec_4_ap_done,
    input wire                                           PEG_Yvec_4_ap_idle,
    input wire                                           PEG_Yvec_4_ap_ready,
    output wire                                          PEG_Yvec_4_ap_rst_n,
    output wire                                          PEG_Yvec_4_ap_start,
    input wire  [                                  64:0] PEG_Yvec_4_fifo_Y_out_din,
    output wire                                          PEG_Yvec_4_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_4_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_4_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_4_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_4_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_4_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_4_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_4_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_4_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_4_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_4_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_4_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_4_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_4_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_5_ap_clk,
    input wire                                           PEG_Yvec_5_ap_done,
    input wire                                           PEG_Yvec_5_ap_idle,
    input wire                                           PEG_Yvec_5_ap_ready,
    output wire                                          PEG_Yvec_5_ap_rst_n,
    output wire                                          PEG_Yvec_5_ap_start,
    input wire  [                                  64:0] PEG_Yvec_5_fifo_Y_out_din,
    output wire                                          PEG_Yvec_5_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_5_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_5_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_5_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_5_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_5_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_5_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_5_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_5_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_5_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_5_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_5_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_5_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_5_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_6_ap_clk,
    input wire                                           PEG_Yvec_6_ap_done,
    input wire                                           PEG_Yvec_6_ap_idle,
    input wire                                           PEG_Yvec_6_ap_ready,
    output wire                                          PEG_Yvec_6_ap_rst_n,
    output wire                                          PEG_Yvec_6_ap_start,
    input wire  [                                  64:0] PEG_Yvec_6_fifo_Y_out_din,
    output wire                                          PEG_Yvec_6_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_6_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_6_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_6_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_6_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_6_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_6_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_6_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_6_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_6_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_6_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_6_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_6_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_6_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_7_ap_clk,
    input wire                                           PEG_Yvec_7_ap_done,
    input wire                                           PEG_Yvec_7_ap_idle,
    input wire                                           PEG_Yvec_7_ap_ready,
    output wire                                          PEG_Yvec_7_ap_rst_n,
    output wire                                          PEG_Yvec_7_ap_start,
    input wire  [                                  64:0] PEG_Yvec_7_fifo_Y_out_din,
    output wire                                          PEG_Yvec_7_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_7_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_7_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_7_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_7_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_7_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_7_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_7_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_7_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_7_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_7_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_7_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_7_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_7_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_8_ap_clk,
    input wire                                           PEG_Yvec_8_ap_done,
    input wire                                           PEG_Yvec_8_ap_idle,
    input wire                                           PEG_Yvec_8_ap_ready,
    output wire                                          PEG_Yvec_8_ap_rst_n,
    output wire                                          PEG_Yvec_8_ap_start,
    input wire  [                                  64:0] PEG_Yvec_8_fifo_Y_out_din,
    output wire                                          PEG_Yvec_8_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_8_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_8_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_8_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_8_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_8_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_8_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_8_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_8_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_8_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_8_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_8_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_8_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_8_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_9_ap_clk,
    input wire                                           PEG_Yvec_9_ap_done,
    input wire                                           PEG_Yvec_9_ap_idle,
    input wire                                           PEG_Yvec_9_ap_ready,
    output wire                                          PEG_Yvec_9_ap_rst_n,
    output wire                                          PEG_Yvec_9_ap_start,
    input wire  [                                  64:0] PEG_Yvec_9_fifo_Y_out_din,
    output wire                                          PEG_Yvec_9_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_9_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_9_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_9_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_9_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_9_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_9_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_9_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_9_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_9_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_9_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_9_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_9_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_9_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_10_ap_clk,
    input wire                                           PEG_Yvec_10_ap_done,
    input wire                                           PEG_Yvec_10_ap_idle,
    input wire                                           PEG_Yvec_10_ap_ready,
    output wire                                          PEG_Yvec_10_ap_rst_n,
    output wire                                          PEG_Yvec_10_ap_start,
    input wire  [                                  64:0] PEG_Yvec_10_fifo_Y_out_din,
    output wire                                          PEG_Yvec_10_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_10_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_10_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_10_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_10_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_10_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_10_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_10_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_10_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_10_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_10_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_10_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_10_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_10_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_11_ap_clk,
    input wire                                           PEG_Yvec_11_ap_done,
    input wire                                           PEG_Yvec_11_ap_idle,
    input wire                                           PEG_Yvec_11_ap_ready,
    output wire                                          PEG_Yvec_11_ap_rst_n,
    output wire                                          PEG_Yvec_11_ap_start,
    input wire  [                                  64:0] PEG_Yvec_11_fifo_Y_out_din,
    output wire                                          PEG_Yvec_11_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_11_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_11_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_11_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_11_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_11_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_11_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_11_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_11_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_11_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_11_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_11_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_11_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_11_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_12_ap_clk,
    input wire                                           PEG_Yvec_12_ap_done,
    input wire                                           PEG_Yvec_12_ap_idle,
    input wire                                           PEG_Yvec_12_ap_ready,
    output wire                                          PEG_Yvec_12_ap_rst_n,
    output wire                                          PEG_Yvec_12_ap_start,
    input wire  [                                  64:0] PEG_Yvec_12_fifo_Y_out_din,
    output wire                                          PEG_Yvec_12_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_12_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_12_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_12_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_12_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_12_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_12_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_12_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_12_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_12_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_12_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_12_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_12_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_12_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_13_ap_clk,
    input wire                                           PEG_Yvec_13_ap_done,
    input wire                                           PEG_Yvec_13_ap_idle,
    input wire                                           PEG_Yvec_13_ap_ready,
    output wire                                          PEG_Yvec_13_ap_rst_n,
    output wire                                          PEG_Yvec_13_ap_start,
    input wire  [                                  64:0] PEG_Yvec_13_fifo_Y_out_din,
    output wire                                          PEG_Yvec_13_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_13_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_13_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_13_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_13_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_13_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_13_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_13_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_13_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_13_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_13_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_13_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_13_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_13_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_14_ap_clk,
    input wire                                           PEG_Yvec_14_ap_done,
    input wire                                           PEG_Yvec_14_ap_idle,
    input wire                                           PEG_Yvec_14_ap_ready,
    output wire                                          PEG_Yvec_14_ap_rst_n,
    output wire                                          PEG_Yvec_14_ap_start,
    input wire  [                                  64:0] PEG_Yvec_14_fifo_Y_out_din,
    output wire                                          PEG_Yvec_14_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_14_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_14_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_14_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_14_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_14_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_14_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_14_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_14_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_14_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_14_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_14_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_14_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_14_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_15_ap_clk,
    input wire                                           PEG_Yvec_15_ap_done,
    input wire                                           PEG_Yvec_15_ap_idle,
    input wire                                           PEG_Yvec_15_ap_ready,
    output wire                                          PEG_Yvec_15_ap_rst_n,
    output wire                                          PEG_Yvec_15_ap_start,
    input wire  [                                  64:0] PEG_Yvec_15_fifo_Y_out_din,
    output wire                                          PEG_Yvec_15_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_15_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_15_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_15_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_15_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_15_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_15_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_15_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_15_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_15_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_15_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_15_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_15_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_15_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_16_ap_clk,
    input wire                                           PEG_Yvec_16_ap_done,
    input wire                                           PEG_Yvec_16_ap_idle,
    input wire                                           PEG_Yvec_16_ap_ready,
    output wire                                          PEG_Yvec_16_ap_rst_n,
    output wire                                          PEG_Yvec_16_ap_start,
    input wire  [                                  64:0] PEG_Yvec_16_fifo_Y_out_din,
    output wire                                          PEG_Yvec_16_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_16_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_16_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_16_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_16_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_16_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_16_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_16_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_16_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_16_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_16_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_16_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_16_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_16_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_17_ap_clk,
    input wire                                           PEG_Yvec_17_ap_done,
    input wire                                           PEG_Yvec_17_ap_idle,
    input wire                                           PEG_Yvec_17_ap_ready,
    output wire                                          PEG_Yvec_17_ap_rst_n,
    output wire                                          PEG_Yvec_17_ap_start,
    input wire  [                                  64:0] PEG_Yvec_17_fifo_Y_out_din,
    output wire                                          PEG_Yvec_17_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_17_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_17_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_17_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_17_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_17_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_17_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_17_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_17_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_17_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_17_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_17_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_17_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_17_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_18_ap_clk,
    input wire                                           PEG_Yvec_18_ap_done,
    input wire                                           PEG_Yvec_18_ap_idle,
    input wire                                           PEG_Yvec_18_ap_ready,
    output wire                                          PEG_Yvec_18_ap_rst_n,
    output wire                                          PEG_Yvec_18_ap_start,
    input wire  [                                  64:0] PEG_Yvec_18_fifo_Y_out_din,
    output wire                                          PEG_Yvec_18_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_18_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_18_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_18_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_18_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_18_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_18_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_18_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_18_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_18_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_18_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_18_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_18_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_18_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_19_ap_clk,
    input wire                                           PEG_Yvec_19_ap_done,
    input wire                                           PEG_Yvec_19_ap_idle,
    input wire                                           PEG_Yvec_19_ap_ready,
    output wire                                          PEG_Yvec_19_ap_rst_n,
    output wire                                          PEG_Yvec_19_ap_start,
    input wire  [                                  64:0] PEG_Yvec_19_fifo_Y_out_din,
    output wire                                          PEG_Yvec_19_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_19_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_19_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_19_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_19_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_19_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_19_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_19_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_19_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_19_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_19_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_19_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_19_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_19_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_20_ap_clk,
    input wire                                           PEG_Yvec_20_ap_done,
    input wire                                           PEG_Yvec_20_ap_idle,
    input wire                                           PEG_Yvec_20_ap_ready,
    output wire                                          PEG_Yvec_20_ap_rst_n,
    output wire                                          PEG_Yvec_20_ap_start,
    input wire  [                                  64:0] PEG_Yvec_20_fifo_Y_out_din,
    output wire                                          PEG_Yvec_20_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_20_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_20_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_20_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_20_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_20_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_20_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_20_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_20_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_20_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_20_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_20_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_20_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_20_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_21_ap_clk,
    input wire                                           PEG_Yvec_21_ap_done,
    input wire                                           PEG_Yvec_21_ap_idle,
    input wire                                           PEG_Yvec_21_ap_ready,
    output wire                                          PEG_Yvec_21_ap_rst_n,
    output wire                                          PEG_Yvec_21_ap_start,
    input wire  [                                  64:0] PEG_Yvec_21_fifo_Y_out_din,
    output wire                                          PEG_Yvec_21_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_21_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_21_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_21_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_21_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_21_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_21_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_21_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_21_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_21_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_21_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_21_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_21_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_21_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_22_ap_clk,
    input wire                                           PEG_Yvec_22_ap_done,
    input wire                                           PEG_Yvec_22_ap_idle,
    input wire                                           PEG_Yvec_22_ap_ready,
    output wire                                          PEG_Yvec_22_ap_rst_n,
    output wire                                          PEG_Yvec_22_ap_start,
    input wire  [                                  64:0] PEG_Yvec_22_fifo_Y_out_din,
    output wire                                          PEG_Yvec_22_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_22_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_22_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_22_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_22_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_22_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_22_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_22_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_22_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_22_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_22_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_22_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_22_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_22_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_23_ap_clk,
    input wire                                           PEG_Yvec_23_ap_done,
    input wire                                           PEG_Yvec_23_ap_idle,
    input wire                                           PEG_Yvec_23_ap_ready,
    output wire                                          PEG_Yvec_23_ap_rst_n,
    output wire                                          PEG_Yvec_23_ap_start,
    input wire  [                                  64:0] PEG_Yvec_23_fifo_Y_out_din,
    output wire                                          PEG_Yvec_23_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_23_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_23_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_23_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_23_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_23_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_23_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_23_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_23_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_23_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_23_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_23_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_23_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_23_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_24_ap_clk,
    input wire                                           PEG_Yvec_24_ap_done,
    input wire                                           PEG_Yvec_24_ap_idle,
    input wire                                           PEG_Yvec_24_ap_ready,
    output wire                                          PEG_Yvec_24_ap_rst_n,
    output wire                                          PEG_Yvec_24_ap_start,
    input wire  [                                  64:0] PEG_Yvec_24_fifo_Y_out_din,
    output wire                                          PEG_Yvec_24_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_24_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_24_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_24_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_24_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_24_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_24_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_24_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_24_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_24_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_24_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_24_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_24_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_24_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_25_ap_clk,
    input wire                                           PEG_Yvec_25_ap_done,
    input wire                                           PEG_Yvec_25_ap_idle,
    input wire                                           PEG_Yvec_25_ap_ready,
    output wire                                          PEG_Yvec_25_ap_rst_n,
    output wire                                          PEG_Yvec_25_ap_start,
    input wire  [                                  64:0] PEG_Yvec_25_fifo_Y_out_din,
    output wire                                          PEG_Yvec_25_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_25_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_25_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_25_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_25_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_25_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_25_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_25_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_25_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_25_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_25_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_25_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_25_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_25_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_26_ap_clk,
    input wire                                           PEG_Yvec_26_ap_done,
    input wire                                           PEG_Yvec_26_ap_idle,
    input wire                                           PEG_Yvec_26_ap_ready,
    output wire                                          PEG_Yvec_26_ap_rst_n,
    output wire                                          PEG_Yvec_26_ap_start,
    input wire  [                                  64:0] PEG_Yvec_26_fifo_Y_out_din,
    output wire                                          PEG_Yvec_26_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_26_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_26_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_26_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_26_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_26_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_26_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_26_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_26_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_26_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_26_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_26_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_26_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_26_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_27_ap_clk,
    input wire                                           PEG_Yvec_27_ap_done,
    input wire                                           PEG_Yvec_27_ap_idle,
    input wire                                           PEG_Yvec_27_ap_ready,
    output wire                                          PEG_Yvec_27_ap_rst_n,
    output wire                                          PEG_Yvec_27_ap_start,
    input wire  [                                  64:0] PEG_Yvec_27_fifo_Y_out_din,
    output wire                                          PEG_Yvec_27_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_27_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_27_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_27_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_27_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_27_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_27_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_27_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_27_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_27_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_27_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_27_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_27_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_27_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_28_ap_clk,
    input wire                                           PEG_Yvec_28_ap_done,
    input wire                                           PEG_Yvec_28_ap_idle,
    input wire                                           PEG_Yvec_28_ap_ready,
    output wire                                          PEG_Yvec_28_ap_rst_n,
    output wire                                          PEG_Yvec_28_ap_start,
    input wire  [                                  64:0] PEG_Yvec_28_fifo_Y_out_din,
    output wire                                          PEG_Yvec_28_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_28_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_28_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_28_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_28_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_28_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_28_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_28_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_28_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_28_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_28_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_28_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_28_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_28_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_29_ap_clk,
    input wire                                           PEG_Yvec_29_ap_done,
    input wire                                           PEG_Yvec_29_ap_idle,
    input wire                                           PEG_Yvec_29_ap_ready,
    output wire                                          PEG_Yvec_29_ap_rst_n,
    output wire                                          PEG_Yvec_29_ap_start,
    input wire  [                                  64:0] PEG_Yvec_29_fifo_Y_out_din,
    output wire                                          PEG_Yvec_29_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_29_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_29_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_29_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_29_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_29_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_29_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_29_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_29_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_29_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_29_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_29_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_29_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_29_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_30_ap_clk,
    input wire                                           PEG_Yvec_30_ap_done,
    input wire                                           PEG_Yvec_30_ap_idle,
    input wire                                           PEG_Yvec_30_ap_ready,
    output wire                                          PEG_Yvec_30_ap_rst_n,
    output wire                                          PEG_Yvec_30_ap_start,
    input wire  [                                  64:0] PEG_Yvec_30_fifo_Y_out_din,
    output wire                                          PEG_Yvec_30_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_30_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_30_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_30_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_30_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_30_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_30_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_30_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_30_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_30_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_30_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_30_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_30_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_30_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_31_ap_clk,
    input wire                                           PEG_Yvec_31_ap_done,
    input wire                                           PEG_Yvec_31_ap_idle,
    input wire                                           PEG_Yvec_31_ap_ready,
    output wire                                          PEG_Yvec_31_ap_rst_n,
    output wire                                          PEG_Yvec_31_ap_start,
    input wire  [                                  64:0] PEG_Yvec_31_fifo_Y_out_din,
    output wire                                          PEG_Yvec_31_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_31_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_31_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_31_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_31_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_31_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_31_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_31_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_31_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_31_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_31_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_31_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_31_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_31_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_32_ap_clk,
    input wire                                           PEG_Yvec_32_ap_done,
    input wire                                           PEG_Yvec_32_ap_idle,
    input wire                                           PEG_Yvec_32_ap_ready,
    output wire                                          PEG_Yvec_32_ap_rst_n,
    output wire                                          PEG_Yvec_32_ap_start,
    input wire  [                                  64:0] PEG_Yvec_32_fifo_Y_out_din,
    output wire                                          PEG_Yvec_32_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_32_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_32_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_32_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_32_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_32_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_32_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_32_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_32_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_32_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_32_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_32_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_32_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_32_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_33_ap_clk,
    input wire                                           PEG_Yvec_33_ap_done,
    input wire                                           PEG_Yvec_33_ap_idle,
    input wire                                           PEG_Yvec_33_ap_ready,
    output wire                                          PEG_Yvec_33_ap_rst_n,
    output wire                                          PEG_Yvec_33_ap_start,
    input wire  [                                  64:0] PEG_Yvec_33_fifo_Y_out_din,
    output wire                                          PEG_Yvec_33_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_33_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_33_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_33_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_33_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_33_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_33_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_33_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_33_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_33_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_33_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_33_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_33_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_33_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_34_ap_clk,
    input wire                                           PEG_Yvec_34_ap_done,
    input wire                                           PEG_Yvec_34_ap_idle,
    input wire                                           PEG_Yvec_34_ap_ready,
    output wire                                          PEG_Yvec_34_ap_rst_n,
    output wire                                          PEG_Yvec_34_ap_start,
    input wire  [                                  64:0] PEG_Yvec_34_fifo_Y_out_din,
    output wire                                          PEG_Yvec_34_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_34_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_34_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_34_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_34_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_34_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_34_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_34_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_34_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_34_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_34_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_34_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_34_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_34_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_35_ap_clk,
    input wire                                           PEG_Yvec_35_ap_done,
    input wire                                           PEG_Yvec_35_ap_idle,
    input wire                                           PEG_Yvec_35_ap_ready,
    output wire                                          PEG_Yvec_35_ap_rst_n,
    output wire                                          PEG_Yvec_35_ap_start,
    input wire  [                                  64:0] PEG_Yvec_35_fifo_Y_out_din,
    output wire                                          PEG_Yvec_35_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_35_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_35_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_35_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_35_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_35_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_35_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_35_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_35_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_35_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_35_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_35_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_35_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_35_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_36_ap_clk,
    input wire                                           PEG_Yvec_36_ap_done,
    input wire                                           PEG_Yvec_36_ap_idle,
    input wire                                           PEG_Yvec_36_ap_ready,
    output wire                                          PEG_Yvec_36_ap_rst_n,
    output wire                                          PEG_Yvec_36_ap_start,
    input wire  [                                  64:0] PEG_Yvec_36_fifo_Y_out_din,
    output wire                                          PEG_Yvec_36_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_36_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_36_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_36_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_36_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_36_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_36_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_36_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_36_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_36_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_36_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_36_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_36_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_36_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_37_ap_clk,
    input wire                                           PEG_Yvec_37_ap_done,
    input wire                                           PEG_Yvec_37_ap_idle,
    input wire                                           PEG_Yvec_37_ap_ready,
    output wire                                          PEG_Yvec_37_ap_rst_n,
    output wire                                          PEG_Yvec_37_ap_start,
    input wire  [                                  64:0] PEG_Yvec_37_fifo_Y_out_din,
    output wire                                          PEG_Yvec_37_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_37_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_37_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_37_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_37_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_37_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_37_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_37_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_37_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_37_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_37_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_37_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_37_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_37_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_38_ap_clk,
    input wire                                           PEG_Yvec_38_ap_done,
    input wire                                           PEG_Yvec_38_ap_idle,
    input wire                                           PEG_Yvec_38_ap_ready,
    output wire                                          PEG_Yvec_38_ap_rst_n,
    output wire                                          PEG_Yvec_38_ap_start,
    input wire  [                                  64:0] PEG_Yvec_38_fifo_Y_out_din,
    output wire                                          PEG_Yvec_38_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_38_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_38_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_38_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_38_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_38_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_38_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_38_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_38_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_38_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_38_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_38_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_38_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_38_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_39_ap_clk,
    input wire                                           PEG_Yvec_39_ap_done,
    input wire                                           PEG_Yvec_39_ap_idle,
    input wire                                           PEG_Yvec_39_ap_ready,
    output wire                                          PEG_Yvec_39_ap_rst_n,
    output wire                                          PEG_Yvec_39_ap_start,
    input wire  [                                  64:0] PEG_Yvec_39_fifo_Y_out_din,
    output wire                                          PEG_Yvec_39_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_39_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_39_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_39_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_39_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_39_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_39_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_39_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_39_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_39_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_39_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_39_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_39_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_39_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_40_ap_clk,
    input wire                                           PEG_Yvec_40_ap_done,
    input wire                                           PEG_Yvec_40_ap_idle,
    input wire                                           PEG_Yvec_40_ap_ready,
    output wire                                          PEG_Yvec_40_ap_rst_n,
    output wire                                          PEG_Yvec_40_ap_start,
    input wire  [                                  64:0] PEG_Yvec_40_fifo_Y_out_din,
    output wire                                          PEG_Yvec_40_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_40_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_40_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_40_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_40_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_40_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_40_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_40_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_40_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_40_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_40_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_40_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_40_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_40_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_41_ap_clk,
    input wire                                           PEG_Yvec_41_ap_done,
    input wire                                           PEG_Yvec_41_ap_idle,
    input wire                                           PEG_Yvec_41_ap_ready,
    output wire                                          PEG_Yvec_41_ap_rst_n,
    output wire                                          PEG_Yvec_41_ap_start,
    input wire  [                                  64:0] PEG_Yvec_41_fifo_Y_out_din,
    output wire                                          PEG_Yvec_41_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_41_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_41_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_41_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_41_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_41_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_41_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_41_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_41_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_41_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_41_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_41_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_41_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_41_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_42_ap_clk,
    input wire                                           PEG_Yvec_42_ap_done,
    input wire                                           PEG_Yvec_42_ap_idle,
    input wire                                           PEG_Yvec_42_ap_ready,
    output wire                                          PEG_Yvec_42_ap_rst_n,
    output wire                                          PEG_Yvec_42_ap_start,
    input wire  [                                  64:0] PEG_Yvec_42_fifo_Y_out_din,
    output wire                                          PEG_Yvec_42_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_42_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_42_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_42_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_42_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_42_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_42_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_42_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_42_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_42_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_42_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_42_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_42_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_42_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_43_ap_clk,
    input wire                                           PEG_Yvec_43_ap_done,
    input wire                                           PEG_Yvec_43_ap_idle,
    input wire                                           PEG_Yvec_43_ap_ready,
    output wire                                          PEG_Yvec_43_ap_rst_n,
    output wire                                          PEG_Yvec_43_ap_start,
    input wire  [                                  64:0] PEG_Yvec_43_fifo_Y_out_din,
    output wire                                          PEG_Yvec_43_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_43_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_43_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_43_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_43_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_43_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_43_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_43_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_43_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_43_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_43_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_43_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_43_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_43_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_44_ap_clk,
    input wire                                           PEG_Yvec_44_ap_done,
    input wire                                           PEG_Yvec_44_ap_idle,
    input wire                                           PEG_Yvec_44_ap_ready,
    output wire                                          PEG_Yvec_44_ap_rst_n,
    output wire                                          PEG_Yvec_44_ap_start,
    input wire  [                                  64:0] PEG_Yvec_44_fifo_Y_out_din,
    output wire                                          PEG_Yvec_44_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_44_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_44_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_44_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_44_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_44_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_44_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_44_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_44_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_44_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_44_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_44_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_44_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_44_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_45_ap_clk,
    input wire                                           PEG_Yvec_45_ap_done,
    input wire                                           PEG_Yvec_45_ap_idle,
    input wire                                           PEG_Yvec_45_ap_ready,
    output wire                                          PEG_Yvec_45_ap_rst_n,
    output wire                                          PEG_Yvec_45_ap_start,
    input wire  [                                  64:0] PEG_Yvec_45_fifo_Y_out_din,
    output wire                                          PEG_Yvec_45_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_45_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_45_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_45_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_45_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_45_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_45_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_45_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_45_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_45_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_45_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_45_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_45_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_45_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_46_ap_clk,
    input wire                                           PEG_Yvec_46_ap_done,
    input wire                                           PEG_Yvec_46_ap_idle,
    input wire                                           PEG_Yvec_46_ap_ready,
    output wire                                          PEG_Yvec_46_ap_rst_n,
    output wire                                          PEG_Yvec_46_ap_start,
    input wire  [                                  64:0] PEG_Yvec_46_fifo_Y_out_din,
    output wire                                          PEG_Yvec_46_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_46_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_46_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_46_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_46_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_46_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_46_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_46_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_46_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_46_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_46_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_46_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_46_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_46_fifo_inst_in_s_read,
    output wire                                          PEG_Yvec_47_ap_clk,
    input wire                                           PEG_Yvec_47_ap_done,
    input wire                                           PEG_Yvec_47_ap_idle,
    input wire                                           PEG_Yvec_47_ap_ready,
    output wire                                          PEG_Yvec_47_ap_rst_n,
    output wire                                          PEG_Yvec_47_ap_start,
    input wire  [                                  64:0] PEG_Yvec_47_fifo_Y_out_din,
    output wire                                          PEG_Yvec_47_fifo_Y_out_full_n,
    input wire                                           PEG_Yvec_47_fifo_Y_out_write,
    output wire [                                 400:0] PEG_Yvec_47_fifo_aXvec_peek_dout,
    output wire                                          PEG_Yvec_47_fifo_aXvec_peek_empty_n,
    input wire                                           PEG_Yvec_47_fifo_aXvec_peek_read,
    output wire [                                 400:0] PEG_Yvec_47_fifo_aXvec_s_dout,
    output wire                                          PEG_Yvec_47_fifo_aXvec_s_empty_n,
    input wire                                           PEG_Yvec_47_fifo_aXvec_s_read,
    output wire [                                  32:0] PEG_Yvec_47_fifo_inst_in_peek_dout,
    output wire                                          PEG_Yvec_47_fifo_inst_in_peek_empty_n,
    input wire                                           PEG_Yvec_47_fifo_inst_in_peek_read,
    output wire [                                  32:0] PEG_Yvec_47_fifo_inst_in_s_dout,
    output wire                                          PEG_Yvec_47_fifo_inst_in_s_empty_n,
    input wire                                           PEG_Yvec_47_fifo_inst_in_s_read,
    output wire                                          black_hole_float_v16_0_ap_clk,
    input wire                                           black_hole_float_v16_0_ap_done,
    input wire                                           black_hole_float_v16_0_ap_idle,
    input wire                                           black_hole_float_v16_0_ap_ready,
    output wire                                          black_hole_float_v16_0_ap_rst_n,
    output wire                                          black_hole_float_v16_0_ap_start,
    output wire [                                 512:0] black_hole_float_v16_0_fifo_in_peek_dout,
    output wire                                          black_hole_float_v16_0_fifo_in_peek_empty_n,
    input wire                                           black_hole_float_v16_0_fifo_in_peek_read,
    output wire [                                 512:0] black_hole_float_v16_0_fifo_in_s_dout,
    output wire                                          black_hole_float_v16_0_fifo_in_s_empty_n,
    input wire                                           black_hole_float_v16_0_fifo_in_s_read,
    output wire                                          black_hole_int_0_ap_clk,
    input wire                                           black_hole_int_0_ap_done,
    input wire                                           black_hole_int_0_ap_idle,
    input wire                                           black_hole_int_0_ap_ready,
    output wire                                          black_hole_int_0_ap_rst_n,
    output wire                                          black_hole_int_0_ap_start,
    output wire [                                  32:0] black_hole_int_0_fifo_in_peek_dout,
    output wire                                          black_hole_int_0_fifo_in_peek_empty_n,
    input wire                                           black_hole_int_0_fifo_in_peek_read,
    output wire [                                  32:0] black_hole_int_0_fifo_in_s_dout,
    output wire                                          black_hole_int_0_fifo_in_s_empty_n,
    input wire                                           black_hole_int_0_fifo_in_s_read,
    output wire [                                  31:0] read_A_0_A_len,
    output wire [                                  63:0] read_A_0_A_read_addr_offset,
    input wire  [                                  63:0] read_A_0_A_read_addr_s_din,
    output wire                                          read_A_0_A_read_addr_s_full_n,
    input wire                                           read_A_0_A_read_addr_s_write,
    output wire [                                 256:0] read_A_0_A_read_data_peek_dout,
    output wire                                          read_A_0_A_read_data_peek_empty_n,
    input wire                                           read_A_0_A_read_data_peek_read,
    output wire [                                 256:0] read_A_0_A_read_data_s_dout,
    output wire                                          read_A_0_A_read_data_s_empty_n,
    input wire                                           read_A_0_A_read_data_s_read,
    output wire [                                  63:0] read_A_0_A_write_addr_offset,
    input wire  [                                  63:0] read_A_0_A_write_addr_s_din,
    output wire                                          read_A_0_A_write_addr_s_full_n,
    input wire                                           read_A_0_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_0_A_write_data_din,
    output wire                                          read_A_0_A_write_data_full_n,
    input wire                                           read_A_0_A_write_data_write,
    output wire [                                   8:0] read_A_0_A_write_resp_peek_dout,
    output wire                                          read_A_0_A_write_resp_peek_empty_n,
    input wire                                           read_A_0_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_0_A_write_resp_s_dout,
    output wire                                          read_A_0_A_write_resp_s_empty_n,
    input wire                                           read_A_0_A_write_resp_s_read,
    output wire [                                  31:0] read_A_0_P_N,
    output wire                                          read_A_0_ap_clk,
    input wire                                           read_A_0_ap_done,
    input wire                                           read_A_0_ap_idle,
    input wire                                           read_A_0_ap_ready,
    output wire                                          read_A_0_ap_rst_n,
    output wire                                          read_A_0_ap_start,
    input wire  [                                 512:0] read_A_0_fifo_A_din,
    output wire                                          read_A_0_fifo_A_full_n,
    input wire                                           read_A_0_fifo_A_write,
    output wire [                                  31:0] read_A_1_A_len,
    output wire [                                  63:0] read_A_1_A_read_addr_offset,
    input wire  [                                  63:0] read_A_1_A_read_addr_s_din,
    output wire                                          read_A_1_A_read_addr_s_full_n,
    input wire                                           read_A_1_A_read_addr_s_write,
    output wire [                                 256:0] read_A_1_A_read_data_peek_dout,
    output wire                                          read_A_1_A_read_data_peek_empty_n,
    input wire                                           read_A_1_A_read_data_peek_read,
    output wire [                                 256:0] read_A_1_A_read_data_s_dout,
    output wire                                          read_A_1_A_read_data_s_empty_n,
    input wire                                           read_A_1_A_read_data_s_read,
    output wire [                                  63:0] read_A_1_A_write_addr_offset,
    input wire  [                                  63:0] read_A_1_A_write_addr_s_din,
    output wire                                          read_A_1_A_write_addr_s_full_n,
    input wire                                           read_A_1_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_1_A_write_data_din,
    output wire                                          read_A_1_A_write_data_full_n,
    input wire                                           read_A_1_A_write_data_write,
    output wire [                                   8:0] read_A_1_A_write_resp_peek_dout,
    output wire                                          read_A_1_A_write_resp_peek_empty_n,
    input wire                                           read_A_1_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_1_A_write_resp_s_dout,
    output wire                                          read_A_1_A_write_resp_s_empty_n,
    input wire                                           read_A_1_A_write_resp_s_read,
    output wire [                                  31:0] read_A_1_P_N,
    output wire                                          read_A_1_ap_clk,
    input wire                                           read_A_1_ap_done,
    input wire                                           read_A_1_ap_idle,
    input wire                                           read_A_1_ap_ready,
    output wire                                          read_A_1_ap_rst_n,
    output wire                                          read_A_1_ap_start,
    input wire  [                                 512:0] read_A_1_fifo_A_din,
    output wire                                          read_A_1_fifo_A_full_n,
    input wire                                           read_A_1_fifo_A_write,
    output wire [                                  31:0] read_A_2_A_len,
    output wire [                                  63:0] read_A_2_A_read_addr_offset,
    input wire  [                                  63:0] read_A_2_A_read_addr_s_din,
    output wire                                          read_A_2_A_read_addr_s_full_n,
    input wire                                           read_A_2_A_read_addr_s_write,
    output wire [                                 256:0] read_A_2_A_read_data_peek_dout,
    output wire                                          read_A_2_A_read_data_peek_empty_n,
    input wire                                           read_A_2_A_read_data_peek_read,
    output wire [                                 256:0] read_A_2_A_read_data_s_dout,
    output wire                                          read_A_2_A_read_data_s_empty_n,
    input wire                                           read_A_2_A_read_data_s_read,
    output wire [                                  63:0] read_A_2_A_write_addr_offset,
    input wire  [                                  63:0] read_A_2_A_write_addr_s_din,
    output wire                                          read_A_2_A_write_addr_s_full_n,
    input wire                                           read_A_2_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_2_A_write_data_din,
    output wire                                          read_A_2_A_write_data_full_n,
    input wire                                           read_A_2_A_write_data_write,
    output wire [                                   8:0] read_A_2_A_write_resp_peek_dout,
    output wire                                          read_A_2_A_write_resp_peek_empty_n,
    input wire                                           read_A_2_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_2_A_write_resp_s_dout,
    output wire                                          read_A_2_A_write_resp_s_empty_n,
    input wire                                           read_A_2_A_write_resp_s_read,
    output wire [                                  31:0] read_A_2_P_N,
    output wire                                          read_A_2_ap_clk,
    input wire                                           read_A_2_ap_done,
    input wire                                           read_A_2_ap_idle,
    input wire                                           read_A_2_ap_ready,
    output wire                                          read_A_2_ap_rst_n,
    output wire                                          read_A_2_ap_start,
    input wire  [                                 512:0] read_A_2_fifo_A_din,
    output wire                                          read_A_2_fifo_A_full_n,
    input wire                                           read_A_2_fifo_A_write,
    output wire [                                  31:0] read_A_3_A_len,
    output wire [                                  63:0] read_A_3_A_read_addr_offset,
    input wire  [                                  63:0] read_A_3_A_read_addr_s_din,
    output wire                                          read_A_3_A_read_addr_s_full_n,
    input wire                                           read_A_3_A_read_addr_s_write,
    output wire [                                 256:0] read_A_3_A_read_data_peek_dout,
    output wire                                          read_A_3_A_read_data_peek_empty_n,
    input wire                                           read_A_3_A_read_data_peek_read,
    output wire [                                 256:0] read_A_3_A_read_data_s_dout,
    output wire                                          read_A_3_A_read_data_s_empty_n,
    input wire                                           read_A_3_A_read_data_s_read,
    output wire [                                  63:0] read_A_3_A_write_addr_offset,
    input wire  [                                  63:0] read_A_3_A_write_addr_s_din,
    output wire                                          read_A_3_A_write_addr_s_full_n,
    input wire                                           read_A_3_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_3_A_write_data_din,
    output wire                                          read_A_3_A_write_data_full_n,
    input wire                                           read_A_3_A_write_data_write,
    output wire [                                   8:0] read_A_3_A_write_resp_peek_dout,
    output wire                                          read_A_3_A_write_resp_peek_empty_n,
    input wire                                           read_A_3_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_3_A_write_resp_s_dout,
    output wire                                          read_A_3_A_write_resp_s_empty_n,
    input wire                                           read_A_3_A_write_resp_s_read,
    output wire [                                  31:0] read_A_3_P_N,
    output wire                                          read_A_3_ap_clk,
    input wire                                           read_A_3_ap_done,
    input wire                                           read_A_3_ap_idle,
    input wire                                           read_A_3_ap_ready,
    output wire                                          read_A_3_ap_rst_n,
    output wire                                          read_A_3_ap_start,
    input wire  [                                 512:0] read_A_3_fifo_A_din,
    output wire                                          read_A_3_fifo_A_full_n,
    input wire                                           read_A_3_fifo_A_write,
    output wire [                                  31:0] read_A_4_A_len,
    output wire [                                  63:0] read_A_4_A_read_addr_offset,
    input wire  [                                  63:0] read_A_4_A_read_addr_s_din,
    output wire                                          read_A_4_A_read_addr_s_full_n,
    input wire                                           read_A_4_A_read_addr_s_write,
    output wire [                                 256:0] read_A_4_A_read_data_peek_dout,
    output wire                                          read_A_4_A_read_data_peek_empty_n,
    input wire                                           read_A_4_A_read_data_peek_read,
    output wire [                                 256:0] read_A_4_A_read_data_s_dout,
    output wire                                          read_A_4_A_read_data_s_empty_n,
    input wire                                           read_A_4_A_read_data_s_read,
    output wire [                                  63:0] read_A_4_A_write_addr_offset,
    input wire  [                                  63:0] read_A_4_A_write_addr_s_din,
    output wire                                          read_A_4_A_write_addr_s_full_n,
    input wire                                           read_A_4_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_4_A_write_data_din,
    output wire                                          read_A_4_A_write_data_full_n,
    input wire                                           read_A_4_A_write_data_write,
    output wire [                                   8:0] read_A_4_A_write_resp_peek_dout,
    output wire                                          read_A_4_A_write_resp_peek_empty_n,
    input wire                                           read_A_4_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_4_A_write_resp_s_dout,
    output wire                                          read_A_4_A_write_resp_s_empty_n,
    input wire                                           read_A_4_A_write_resp_s_read,
    output wire [                                  31:0] read_A_4_P_N,
    output wire                                          read_A_4_ap_clk,
    input wire                                           read_A_4_ap_done,
    input wire                                           read_A_4_ap_idle,
    input wire                                           read_A_4_ap_ready,
    output wire                                          read_A_4_ap_rst_n,
    output wire                                          read_A_4_ap_start,
    input wire  [                                 512:0] read_A_4_fifo_A_din,
    output wire                                          read_A_4_fifo_A_full_n,
    input wire                                           read_A_4_fifo_A_write,
    output wire [                                  31:0] read_A_5_A_len,
    output wire [                                  63:0] read_A_5_A_read_addr_offset,
    input wire  [                                  63:0] read_A_5_A_read_addr_s_din,
    output wire                                          read_A_5_A_read_addr_s_full_n,
    input wire                                           read_A_5_A_read_addr_s_write,
    output wire [                                 256:0] read_A_5_A_read_data_peek_dout,
    output wire                                          read_A_5_A_read_data_peek_empty_n,
    input wire                                           read_A_5_A_read_data_peek_read,
    output wire [                                 256:0] read_A_5_A_read_data_s_dout,
    output wire                                          read_A_5_A_read_data_s_empty_n,
    input wire                                           read_A_5_A_read_data_s_read,
    output wire [                                  63:0] read_A_5_A_write_addr_offset,
    input wire  [                                  63:0] read_A_5_A_write_addr_s_din,
    output wire                                          read_A_5_A_write_addr_s_full_n,
    input wire                                           read_A_5_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_5_A_write_data_din,
    output wire                                          read_A_5_A_write_data_full_n,
    input wire                                           read_A_5_A_write_data_write,
    output wire [                                   8:0] read_A_5_A_write_resp_peek_dout,
    output wire                                          read_A_5_A_write_resp_peek_empty_n,
    input wire                                           read_A_5_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_5_A_write_resp_s_dout,
    output wire                                          read_A_5_A_write_resp_s_empty_n,
    input wire                                           read_A_5_A_write_resp_s_read,
    output wire [                                  31:0] read_A_5_P_N,
    output wire                                          read_A_5_ap_clk,
    input wire                                           read_A_5_ap_done,
    input wire                                           read_A_5_ap_idle,
    input wire                                           read_A_5_ap_ready,
    output wire                                          read_A_5_ap_rst_n,
    output wire                                          read_A_5_ap_start,
    input wire  [                                 512:0] read_A_5_fifo_A_din,
    output wire                                          read_A_5_fifo_A_full_n,
    input wire                                           read_A_5_fifo_A_write,
    output wire [                                  31:0] read_A_6_A_len,
    output wire [                                  63:0] read_A_6_A_read_addr_offset,
    input wire  [                                  63:0] read_A_6_A_read_addr_s_din,
    output wire                                          read_A_6_A_read_addr_s_full_n,
    input wire                                           read_A_6_A_read_addr_s_write,
    output wire [                                 256:0] read_A_6_A_read_data_peek_dout,
    output wire                                          read_A_6_A_read_data_peek_empty_n,
    input wire                                           read_A_6_A_read_data_peek_read,
    output wire [                                 256:0] read_A_6_A_read_data_s_dout,
    output wire                                          read_A_6_A_read_data_s_empty_n,
    input wire                                           read_A_6_A_read_data_s_read,
    output wire [                                  63:0] read_A_6_A_write_addr_offset,
    input wire  [                                  63:0] read_A_6_A_write_addr_s_din,
    output wire                                          read_A_6_A_write_addr_s_full_n,
    input wire                                           read_A_6_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_6_A_write_data_din,
    output wire                                          read_A_6_A_write_data_full_n,
    input wire                                           read_A_6_A_write_data_write,
    output wire [                                   8:0] read_A_6_A_write_resp_peek_dout,
    output wire                                          read_A_6_A_write_resp_peek_empty_n,
    input wire                                           read_A_6_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_6_A_write_resp_s_dout,
    output wire                                          read_A_6_A_write_resp_s_empty_n,
    input wire                                           read_A_6_A_write_resp_s_read,
    output wire [                                  31:0] read_A_6_P_N,
    output wire                                          read_A_6_ap_clk,
    input wire                                           read_A_6_ap_done,
    input wire                                           read_A_6_ap_idle,
    input wire                                           read_A_6_ap_ready,
    output wire                                          read_A_6_ap_rst_n,
    output wire                                          read_A_6_ap_start,
    input wire  [                                 512:0] read_A_6_fifo_A_din,
    output wire                                          read_A_6_fifo_A_full_n,
    input wire                                           read_A_6_fifo_A_write,
    output wire [                                  31:0] read_A_7_A_len,
    output wire [                                  63:0] read_A_7_A_read_addr_offset,
    input wire  [                                  63:0] read_A_7_A_read_addr_s_din,
    output wire                                          read_A_7_A_read_addr_s_full_n,
    input wire                                           read_A_7_A_read_addr_s_write,
    output wire [                                 256:0] read_A_7_A_read_data_peek_dout,
    output wire                                          read_A_7_A_read_data_peek_empty_n,
    input wire                                           read_A_7_A_read_data_peek_read,
    output wire [                                 256:0] read_A_7_A_read_data_s_dout,
    output wire                                          read_A_7_A_read_data_s_empty_n,
    input wire                                           read_A_7_A_read_data_s_read,
    output wire [                                  63:0] read_A_7_A_write_addr_offset,
    input wire  [                                  63:0] read_A_7_A_write_addr_s_din,
    output wire                                          read_A_7_A_write_addr_s_full_n,
    input wire                                           read_A_7_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_7_A_write_data_din,
    output wire                                          read_A_7_A_write_data_full_n,
    input wire                                           read_A_7_A_write_data_write,
    output wire [                                   8:0] read_A_7_A_write_resp_peek_dout,
    output wire                                          read_A_7_A_write_resp_peek_empty_n,
    input wire                                           read_A_7_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_7_A_write_resp_s_dout,
    output wire                                          read_A_7_A_write_resp_s_empty_n,
    input wire                                           read_A_7_A_write_resp_s_read,
    output wire [                                  31:0] read_A_7_P_N,
    output wire                                          read_A_7_ap_clk,
    input wire                                           read_A_7_ap_done,
    input wire                                           read_A_7_ap_idle,
    input wire                                           read_A_7_ap_ready,
    output wire                                          read_A_7_ap_rst_n,
    output wire                                          read_A_7_ap_start,
    input wire  [                                 512:0] read_A_7_fifo_A_din,
    output wire                                          read_A_7_fifo_A_full_n,
    input wire                                           read_A_7_fifo_A_write,
    output wire [                                  31:0] read_A_8_A_len,
    output wire [                                  63:0] read_A_8_A_read_addr_offset,
    input wire  [                                  63:0] read_A_8_A_read_addr_s_din,
    output wire                                          read_A_8_A_read_addr_s_full_n,
    input wire                                           read_A_8_A_read_addr_s_write,
    output wire [                                 256:0] read_A_8_A_read_data_peek_dout,
    output wire                                          read_A_8_A_read_data_peek_empty_n,
    input wire                                           read_A_8_A_read_data_peek_read,
    output wire [                                 256:0] read_A_8_A_read_data_s_dout,
    output wire                                          read_A_8_A_read_data_s_empty_n,
    input wire                                           read_A_8_A_read_data_s_read,
    output wire [                                  63:0] read_A_8_A_write_addr_offset,
    input wire  [                                  63:0] read_A_8_A_write_addr_s_din,
    output wire                                          read_A_8_A_write_addr_s_full_n,
    input wire                                           read_A_8_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_8_A_write_data_din,
    output wire                                          read_A_8_A_write_data_full_n,
    input wire                                           read_A_8_A_write_data_write,
    output wire [                                   8:0] read_A_8_A_write_resp_peek_dout,
    output wire                                          read_A_8_A_write_resp_peek_empty_n,
    input wire                                           read_A_8_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_8_A_write_resp_s_dout,
    output wire                                          read_A_8_A_write_resp_s_empty_n,
    input wire                                           read_A_8_A_write_resp_s_read,
    output wire [                                  31:0] read_A_8_P_N,
    output wire                                          read_A_8_ap_clk,
    input wire                                           read_A_8_ap_done,
    input wire                                           read_A_8_ap_idle,
    input wire                                           read_A_8_ap_ready,
    output wire                                          read_A_8_ap_rst_n,
    output wire                                          read_A_8_ap_start,
    input wire  [                                 512:0] read_A_8_fifo_A_din,
    output wire                                          read_A_8_fifo_A_full_n,
    input wire                                           read_A_8_fifo_A_write,
    output wire [                                  31:0] read_A_9_A_len,
    output wire [                                  63:0] read_A_9_A_read_addr_offset,
    input wire  [                                  63:0] read_A_9_A_read_addr_s_din,
    output wire                                          read_A_9_A_read_addr_s_full_n,
    input wire                                           read_A_9_A_read_addr_s_write,
    output wire [                                 256:0] read_A_9_A_read_data_peek_dout,
    output wire                                          read_A_9_A_read_data_peek_empty_n,
    input wire                                           read_A_9_A_read_data_peek_read,
    output wire [                                 256:0] read_A_9_A_read_data_s_dout,
    output wire                                          read_A_9_A_read_data_s_empty_n,
    input wire                                           read_A_9_A_read_data_s_read,
    output wire [                                  63:0] read_A_9_A_write_addr_offset,
    input wire  [                                  63:0] read_A_9_A_write_addr_s_din,
    output wire                                          read_A_9_A_write_addr_s_full_n,
    input wire                                           read_A_9_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_9_A_write_data_din,
    output wire                                          read_A_9_A_write_data_full_n,
    input wire                                           read_A_9_A_write_data_write,
    output wire [                                   8:0] read_A_9_A_write_resp_peek_dout,
    output wire                                          read_A_9_A_write_resp_peek_empty_n,
    input wire                                           read_A_9_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_9_A_write_resp_s_dout,
    output wire                                          read_A_9_A_write_resp_s_empty_n,
    input wire                                           read_A_9_A_write_resp_s_read,
    output wire [                                  31:0] read_A_9_P_N,
    output wire                                          read_A_9_ap_clk,
    input wire                                           read_A_9_ap_done,
    input wire                                           read_A_9_ap_idle,
    input wire                                           read_A_9_ap_ready,
    output wire                                          read_A_9_ap_rst_n,
    output wire                                          read_A_9_ap_start,
    input wire  [                                 512:0] read_A_9_fifo_A_din,
    output wire                                          read_A_9_fifo_A_full_n,
    input wire                                           read_A_9_fifo_A_write,
    output wire [                                  31:0] read_A_10_A_len,
    output wire [                                  63:0] read_A_10_A_read_addr_offset,
    input wire  [                                  63:0] read_A_10_A_read_addr_s_din,
    output wire                                          read_A_10_A_read_addr_s_full_n,
    input wire                                           read_A_10_A_read_addr_s_write,
    output wire [                                 256:0] read_A_10_A_read_data_peek_dout,
    output wire                                          read_A_10_A_read_data_peek_empty_n,
    input wire                                           read_A_10_A_read_data_peek_read,
    output wire [                                 256:0] read_A_10_A_read_data_s_dout,
    output wire                                          read_A_10_A_read_data_s_empty_n,
    input wire                                           read_A_10_A_read_data_s_read,
    output wire [                                  63:0] read_A_10_A_write_addr_offset,
    input wire  [                                  63:0] read_A_10_A_write_addr_s_din,
    output wire                                          read_A_10_A_write_addr_s_full_n,
    input wire                                           read_A_10_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_10_A_write_data_din,
    output wire                                          read_A_10_A_write_data_full_n,
    input wire                                           read_A_10_A_write_data_write,
    output wire [                                   8:0] read_A_10_A_write_resp_peek_dout,
    output wire                                          read_A_10_A_write_resp_peek_empty_n,
    input wire                                           read_A_10_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_10_A_write_resp_s_dout,
    output wire                                          read_A_10_A_write_resp_s_empty_n,
    input wire                                           read_A_10_A_write_resp_s_read,
    output wire [                                  31:0] read_A_10_P_N,
    output wire                                          read_A_10_ap_clk,
    input wire                                           read_A_10_ap_done,
    input wire                                           read_A_10_ap_idle,
    input wire                                           read_A_10_ap_ready,
    output wire                                          read_A_10_ap_rst_n,
    output wire                                          read_A_10_ap_start,
    input wire  [                                 512:0] read_A_10_fifo_A_din,
    output wire                                          read_A_10_fifo_A_full_n,
    input wire                                           read_A_10_fifo_A_write,
    output wire [                                  31:0] read_A_11_A_len,
    output wire [                                  63:0] read_A_11_A_read_addr_offset,
    input wire  [                                  63:0] read_A_11_A_read_addr_s_din,
    output wire                                          read_A_11_A_read_addr_s_full_n,
    input wire                                           read_A_11_A_read_addr_s_write,
    output wire [                                 256:0] read_A_11_A_read_data_peek_dout,
    output wire                                          read_A_11_A_read_data_peek_empty_n,
    input wire                                           read_A_11_A_read_data_peek_read,
    output wire [                                 256:0] read_A_11_A_read_data_s_dout,
    output wire                                          read_A_11_A_read_data_s_empty_n,
    input wire                                           read_A_11_A_read_data_s_read,
    output wire [                                  63:0] read_A_11_A_write_addr_offset,
    input wire  [                                  63:0] read_A_11_A_write_addr_s_din,
    output wire                                          read_A_11_A_write_addr_s_full_n,
    input wire                                           read_A_11_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_11_A_write_data_din,
    output wire                                          read_A_11_A_write_data_full_n,
    input wire                                           read_A_11_A_write_data_write,
    output wire [                                   8:0] read_A_11_A_write_resp_peek_dout,
    output wire                                          read_A_11_A_write_resp_peek_empty_n,
    input wire                                           read_A_11_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_11_A_write_resp_s_dout,
    output wire                                          read_A_11_A_write_resp_s_empty_n,
    input wire                                           read_A_11_A_write_resp_s_read,
    output wire [                                  31:0] read_A_11_P_N,
    output wire                                          read_A_11_ap_clk,
    input wire                                           read_A_11_ap_done,
    input wire                                           read_A_11_ap_idle,
    input wire                                           read_A_11_ap_ready,
    output wire                                          read_A_11_ap_rst_n,
    output wire                                          read_A_11_ap_start,
    input wire  [                                 512:0] read_A_11_fifo_A_din,
    output wire                                          read_A_11_fifo_A_full_n,
    input wire                                           read_A_11_fifo_A_write,
    output wire [                                  31:0] read_A_12_A_len,
    output wire [                                  63:0] read_A_12_A_read_addr_offset,
    input wire  [                                  63:0] read_A_12_A_read_addr_s_din,
    output wire                                          read_A_12_A_read_addr_s_full_n,
    input wire                                           read_A_12_A_read_addr_s_write,
    output wire [                                 256:0] read_A_12_A_read_data_peek_dout,
    output wire                                          read_A_12_A_read_data_peek_empty_n,
    input wire                                           read_A_12_A_read_data_peek_read,
    output wire [                                 256:0] read_A_12_A_read_data_s_dout,
    output wire                                          read_A_12_A_read_data_s_empty_n,
    input wire                                           read_A_12_A_read_data_s_read,
    output wire [                                  63:0] read_A_12_A_write_addr_offset,
    input wire  [                                  63:0] read_A_12_A_write_addr_s_din,
    output wire                                          read_A_12_A_write_addr_s_full_n,
    input wire                                           read_A_12_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_12_A_write_data_din,
    output wire                                          read_A_12_A_write_data_full_n,
    input wire                                           read_A_12_A_write_data_write,
    output wire [                                   8:0] read_A_12_A_write_resp_peek_dout,
    output wire                                          read_A_12_A_write_resp_peek_empty_n,
    input wire                                           read_A_12_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_12_A_write_resp_s_dout,
    output wire                                          read_A_12_A_write_resp_s_empty_n,
    input wire                                           read_A_12_A_write_resp_s_read,
    output wire [                                  31:0] read_A_12_P_N,
    output wire                                          read_A_12_ap_clk,
    input wire                                           read_A_12_ap_done,
    input wire                                           read_A_12_ap_idle,
    input wire                                           read_A_12_ap_ready,
    output wire                                          read_A_12_ap_rst_n,
    output wire                                          read_A_12_ap_start,
    input wire  [                                 512:0] read_A_12_fifo_A_din,
    output wire                                          read_A_12_fifo_A_full_n,
    input wire                                           read_A_12_fifo_A_write,
    output wire [                                  31:0] read_A_13_A_len,
    output wire [                                  63:0] read_A_13_A_read_addr_offset,
    input wire  [                                  63:0] read_A_13_A_read_addr_s_din,
    output wire                                          read_A_13_A_read_addr_s_full_n,
    input wire                                           read_A_13_A_read_addr_s_write,
    output wire [                                 256:0] read_A_13_A_read_data_peek_dout,
    output wire                                          read_A_13_A_read_data_peek_empty_n,
    input wire                                           read_A_13_A_read_data_peek_read,
    output wire [                                 256:0] read_A_13_A_read_data_s_dout,
    output wire                                          read_A_13_A_read_data_s_empty_n,
    input wire                                           read_A_13_A_read_data_s_read,
    output wire [                                  63:0] read_A_13_A_write_addr_offset,
    input wire  [                                  63:0] read_A_13_A_write_addr_s_din,
    output wire                                          read_A_13_A_write_addr_s_full_n,
    input wire                                           read_A_13_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_13_A_write_data_din,
    output wire                                          read_A_13_A_write_data_full_n,
    input wire                                           read_A_13_A_write_data_write,
    output wire [                                   8:0] read_A_13_A_write_resp_peek_dout,
    output wire                                          read_A_13_A_write_resp_peek_empty_n,
    input wire                                           read_A_13_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_13_A_write_resp_s_dout,
    output wire                                          read_A_13_A_write_resp_s_empty_n,
    input wire                                           read_A_13_A_write_resp_s_read,
    output wire [                                  31:0] read_A_13_P_N,
    output wire                                          read_A_13_ap_clk,
    input wire                                           read_A_13_ap_done,
    input wire                                           read_A_13_ap_idle,
    input wire                                           read_A_13_ap_ready,
    output wire                                          read_A_13_ap_rst_n,
    output wire                                          read_A_13_ap_start,
    input wire  [                                 512:0] read_A_13_fifo_A_din,
    output wire                                          read_A_13_fifo_A_full_n,
    input wire                                           read_A_13_fifo_A_write,
    output wire [                                  31:0] read_A_14_A_len,
    output wire [                                  63:0] read_A_14_A_read_addr_offset,
    input wire  [                                  63:0] read_A_14_A_read_addr_s_din,
    output wire                                          read_A_14_A_read_addr_s_full_n,
    input wire                                           read_A_14_A_read_addr_s_write,
    output wire [                                 256:0] read_A_14_A_read_data_peek_dout,
    output wire                                          read_A_14_A_read_data_peek_empty_n,
    input wire                                           read_A_14_A_read_data_peek_read,
    output wire [                                 256:0] read_A_14_A_read_data_s_dout,
    output wire                                          read_A_14_A_read_data_s_empty_n,
    input wire                                           read_A_14_A_read_data_s_read,
    output wire [                                  63:0] read_A_14_A_write_addr_offset,
    input wire  [                                  63:0] read_A_14_A_write_addr_s_din,
    output wire                                          read_A_14_A_write_addr_s_full_n,
    input wire                                           read_A_14_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_14_A_write_data_din,
    output wire                                          read_A_14_A_write_data_full_n,
    input wire                                           read_A_14_A_write_data_write,
    output wire [                                   8:0] read_A_14_A_write_resp_peek_dout,
    output wire                                          read_A_14_A_write_resp_peek_empty_n,
    input wire                                           read_A_14_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_14_A_write_resp_s_dout,
    output wire                                          read_A_14_A_write_resp_s_empty_n,
    input wire                                           read_A_14_A_write_resp_s_read,
    output wire [                                  31:0] read_A_14_P_N,
    output wire                                          read_A_14_ap_clk,
    input wire                                           read_A_14_ap_done,
    input wire                                           read_A_14_ap_idle,
    input wire                                           read_A_14_ap_ready,
    output wire                                          read_A_14_ap_rst_n,
    output wire                                          read_A_14_ap_start,
    input wire  [                                 512:0] read_A_14_fifo_A_din,
    output wire                                          read_A_14_fifo_A_full_n,
    input wire                                           read_A_14_fifo_A_write,
    output wire [                                  31:0] read_A_15_A_len,
    output wire [                                  63:0] read_A_15_A_read_addr_offset,
    input wire  [                                  63:0] read_A_15_A_read_addr_s_din,
    output wire                                          read_A_15_A_read_addr_s_full_n,
    input wire                                           read_A_15_A_read_addr_s_write,
    output wire [                                 256:0] read_A_15_A_read_data_peek_dout,
    output wire                                          read_A_15_A_read_data_peek_empty_n,
    input wire                                           read_A_15_A_read_data_peek_read,
    output wire [                                 256:0] read_A_15_A_read_data_s_dout,
    output wire                                          read_A_15_A_read_data_s_empty_n,
    input wire                                           read_A_15_A_read_data_s_read,
    output wire [                                  63:0] read_A_15_A_write_addr_offset,
    input wire  [                                  63:0] read_A_15_A_write_addr_s_din,
    output wire                                          read_A_15_A_write_addr_s_full_n,
    input wire                                           read_A_15_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_15_A_write_data_din,
    output wire                                          read_A_15_A_write_data_full_n,
    input wire                                           read_A_15_A_write_data_write,
    output wire [                                   8:0] read_A_15_A_write_resp_peek_dout,
    output wire                                          read_A_15_A_write_resp_peek_empty_n,
    input wire                                           read_A_15_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_15_A_write_resp_s_dout,
    output wire                                          read_A_15_A_write_resp_s_empty_n,
    input wire                                           read_A_15_A_write_resp_s_read,
    output wire [                                  31:0] read_A_15_P_N,
    output wire                                          read_A_15_ap_clk,
    input wire                                           read_A_15_ap_done,
    input wire                                           read_A_15_ap_idle,
    input wire                                           read_A_15_ap_ready,
    output wire                                          read_A_15_ap_rst_n,
    output wire                                          read_A_15_ap_start,
    input wire  [                                 512:0] read_A_15_fifo_A_din,
    output wire                                          read_A_15_fifo_A_full_n,
    input wire                                           read_A_15_fifo_A_write,
    output wire [                                  31:0] read_A_16_A_len,
    output wire [                                  63:0] read_A_16_A_read_addr_offset,
    input wire  [                                  63:0] read_A_16_A_read_addr_s_din,
    output wire                                          read_A_16_A_read_addr_s_full_n,
    input wire                                           read_A_16_A_read_addr_s_write,
    output wire [                                 256:0] read_A_16_A_read_data_peek_dout,
    output wire                                          read_A_16_A_read_data_peek_empty_n,
    input wire                                           read_A_16_A_read_data_peek_read,
    output wire [                                 256:0] read_A_16_A_read_data_s_dout,
    output wire                                          read_A_16_A_read_data_s_empty_n,
    input wire                                           read_A_16_A_read_data_s_read,
    output wire [                                  63:0] read_A_16_A_write_addr_offset,
    input wire  [                                  63:0] read_A_16_A_write_addr_s_din,
    output wire                                          read_A_16_A_write_addr_s_full_n,
    input wire                                           read_A_16_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_16_A_write_data_din,
    output wire                                          read_A_16_A_write_data_full_n,
    input wire                                           read_A_16_A_write_data_write,
    output wire [                                   8:0] read_A_16_A_write_resp_peek_dout,
    output wire                                          read_A_16_A_write_resp_peek_empty_n,
    input wire                                           read_A_16_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_16_A_write_resp_s_dout,
    output wire                                          read_A_16_A_write_resp_s_empty_n,
    input wire                                           read_A_16_A_write_resp_s_read,
    output wire [                                  31:0] read_A_16_P_N,
    output wire                                          read_A_16_ap_clk,
    input wire                                           read_A_16_ap_done,
    input wire                                           read_A_16_ap_idle,
    input wire                                           read_A_16_ap_ready,
    output wire                                          read_A_16_ap_rst_n,
    output wire                                          read_A_16_ap_start,
    input wire  [                                 512:0] read_A_16_fifo_A_din,
    output wire                                          read_A_16_fifo_A_full_n,
    input wire                                           read_A_16_fifo_A_write,
    output wire [                                  31:0] read_A_17_A_len,
    output wire [                                  63:0] read_A_17_A_read_addr_offset,
    input wire  [                                  63:0] read_A_17_A_read_addr_s_din,
    output wire                                          read_A_17_A_read_addr_s_full_n,
    input wire                                           read_A_17_A_read_addr_s_write,
    output wire [                                 256:0] read_A_17_A_read_data_peek_dout,
    output wire                                          read_A_17_A_read_data_peek_empty_n,
    input wire                                           read_A_17_A_read_data_peek_read,
    output wire [                                 256:0] read_A_17_A_read_data_s_dout,
    output wire                                          read_A_17_A_read_data_s_empty_n,
    input wire                                           read_A_17_A_read_data_s_read,
    output wire [                                  63:0] read_A_17_A_write_addr_offset,
    input wire  [                                  63:0] read_A_17_A_write_addr_s_din,
    output wire                                          read_A_17_A_write_addr_s_full_n,
    input wire                                           read_A_17_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_17_A_write_data_din,
    output wire                                          read_A_17_A_write_data_full_n,
    input wire                                           read_A_17_A_write_data_write,
    output wire [                                   8:0] read_A_17_A_write_resp_peek_dout,
    output wire                                          read_A_17_A_write_resp_peek_empty_n,
    input wire                                           read_A_17_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_17_A_write_resp_s_dout,
    output wire                                          read_A_17_A_write_resp_s_empty_n,
    input wire                                           read_A_17_A_write_resp_s_read,
    output wire [                                  31:0] read_A_17_P_N,
    output wire                                          read_A_17_ap_clk,
    input wire                                           read_A_17_ap_done,
    input wire                                           read_A_17_ap_idle,
    input wire                                           read_A_17_ap_ready,
    output wire                                          read_A_17_ap_rst_n,
    output wire                                          read_A_17_ap_start,
    input wire  [                                 512:0] read_A_17_fifo_A_din,
    output wire                                          read_A_17_fifo_A_full_n,
    input wire                                           read_A_17_fifo_A_write,
    output wire [                                  31:0] read_A_18_A_len,
    output wire [                                  63:0] read_A_18_A_read_addr_offset,
    input wire  [                                  63:0] read_A_18_A_read_addr_s_din,
    output wire                                          read_A_18_A_read_addr_s_full_n,
    input wire                                           read_A_18_A_read_addr_s_write,
    output wire [                                 256:0] read_A_18_A_read_data_peek_dout,
    output wire                                          read_A_18_A_read_data_peek_empty_n,
    input wire                                           read_A_18_A_read_data_peek_read,
    output wire [                                 256:0] read_A_18_A_read_data_s_dout,
    output wire                                          read_A_18_A_read_data_s_empty_n,
    input wire                                           read_A_18_A_read_data_s_read,
    output wire [                                  63:0] read_A_18_A_write_addr_offset,
    input wire  [                                  63:0] read_A_18_A_write_addr_s_din,
    output wire                                          read_A_18_A_write_addr_s_full_n,
    input wire                                           read_A_18_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_18_A_write_data_din,
    output wire                                          read_A_18_A_write_data_full_n,
    input wire                                           read_A_18_A_write_data_write,
    output wire [                                   8:0] read_A_18_A_write_resp_peek_dout,
    output wire                                          read_A_18_A_write_resp_peek_empty_n,
    input wire                                           read_A_18_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_18_A_write_resp_s_dout,
    output wire                                          read_A_18_A_write_resp_s_empty_n,
    input wire                                           read_A_18_A_write_resp_s_read,
    output wire [                                  31:0] read_A_18_P_N,
    output wire                                          read_A_18_ap_clk,
    input wire                                           read_A_18_ap_done,
    input wire                                           read_A_18_ap_idle,
    input wire                                           read_A_18_ap_ready,
    output wire                                          read_A_18_ap_rst_n,
    output wire                                          read_A_18_ap_start,
    input wire  [                                 512:0] read_A_18_fifo_A_din,
    output wire                                          read_A_18_fifo_A_full_n,
    input wire                                           read_A_18_fifo_A_write,
    output wire [                                  31:0] read_A_19_A_len,
    output wire [                                  63:0] read_A_19_A_read_addr_offset,
    input wire  [                                  63:0] read_A_19_A_read_addr_s_din,
    output wire                                          read_A_19_A_read_addr_s_full_n,
    input wire                                           read_A_19_A_read_addr_s_write,
    output wire [                                 256:0] read_A_19_A_read_data_peek_dout,
    output wire                                          read_A_19_A_read_data_peek_empty_n,
    input wire                                           read_A_19_A_read_data_peek_read,
    output wire [                                 256:0] read_A_19_A_read_data_s_dout,
    output wire                                          read_A_19_A_read_data_s_empty_n,
    input wire                                           read_A_19_A_read_data_s_read,
    output wire [                                  63:0] read_A_19_A_write_addr_offset,
    input wire  [                                  63:0] read_A_19_A_write_addr_s_din,
    output wire                                          read_A_19_A_write_addr_s_full_n,
    input wire                                           read_A_19_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_19_A_write_data_din,
    output wire                                          read_A_19_A_write_data_full_n,
    input wire                                           read_A_19_A_write_data_write,
    output wire [                                   8:0] read_A_19_A_write_resp_peek_dout,
    output wire                                          read_A_19_A_write_resp_peek_empty_n,
    input wire                                           read_A_19_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_19_A_write_resp_s_dout,
    output wire                                          read_A_19_A_write_resp_s_empty_n,
    input wire                                           read_A_19_A_write_resp_s_read,
    output wire [                                  31:0] read_A_19_P_N,
    output wire                                          read_A_19_ap_clk,
    input wire                                           read_A_19_ap_done,
    input wire                                           read_A_19_ap_idle,
    input wire                                           read_A_19_ap_ready,
    output wire                                          read_A_19_ap_rst_n,
    output wire                                          read_A_19_ap_start,
    input wire  [                                 512:0] read_A_19_fifo_A_din,
    output wire                                          read_A_19_fifo_A_full_n,
    input wire                                           read_A_19_fifo_A_write,
    output wire [                                  31:0] read_A_20_A_len,
    output wire [                                  63:0] read_A_20_A_read_addr_offset,
    input wire  [                                  63:0] read_A_20_A_read_addr_s_din,
    output wire                                          read_A_20_A_read_addr_s_full_n,
    input wire                                           read_A_20_A_read_addr_s_write,
    output wire [                                 256:0] read_A_20_A_read_data_peek_dout,
    output wire                                          read_A_20_A_read_data_peek_empty_n,
    input wire                                           read_A_20_A_read_data_peek_read,
    output wire [                                 256:0] read_A_20_A_read_data_s_dout,
    output wire                                          read_A_20_A_read_data_s_empty_n,
    input wire                                           read_A_20_A_read_data_s_read,
    output wire [                                  63:0] read_A_20_A_write_addr_offset,
    input wire  [                                  63:0] read_A_20_A_write_addr_s_din,
    output wire                                          read_A_20_A_write_addr_s_full_n,
    input wire                                           read_A_20_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_20_A_write_data_din,
    output wire                                          read_A_20_A_write_data_full_n,
    input wire                                           read_A_20_A_write_data_write,
    output wire [                                   8:0] read_A_20_A_write_resp_peek_dout,
    output wire                                          read_A_20_A_write_resp_peek_empty_n,
    input wire                                           read_A_20_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_20_A_write_resp_s_dout,
    output wire                                          read_A_20_A_write_resp_s_empty_n,
    input wire                                           read_A_20_A_write_resp_s_read,
    output wire [                                  31:0] read_A_20_P_N,
    output wire                                          read_A_20_ap_clk,
    input wire                                           read_A_20_ap_done,
    input wire                                           read_A_20_ap_idle,
    input wire                                           read_A_20_ap_ready,
    output wire                                          read_A_20_ap_rst_n,
    output wire                                          read_A_20_ap_start,
    input wire  [                                 512:0] read_A_20_fifo_A_din,
    output wire                                          read_A_20_fifo_A_full_n,
    input wire                                           read_A_20_fifo_A_write,
    output wire [                                  31:0] read_A_21_A_len,
    output wire [                                  63:0] read_A_21_A_read_addr_offset,
    input wire  [                                  63:0] read_A_21_A_read_addr_s_din,
    output wire                                          read_A_21_A_read_addr_s_full_n,
    input wire                                           read_A_21_A_read_addr_s_write,
    output wire [                                 256:0] read_A_21_A_read_data_peek_dout,
    output wire                                          read_A_21_A_read_data_peek_empty_n,
    input wire                                           read_A_21_A_read_data_peek_read,
    output wire [                                 256:0] read_A_21_A_read_data_s_dout,
    output wire                                          read_A_21_A_read_data_s_empty_n,
    input wire                                           read_A_21_A_read_data_s_read,
    output wire [                                  63:0] read_A_21_A_write_addr_offset,
    input wire  [                                  63:0] read_A_21_A_write_addr_s_din,
    output wire                                          read_A_21_A_write_addr_s_full_n,
    input wire                                           read_A_21_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_21_A_write_data_din,
    output wire                                          read_A_21_A_write_data_full_n,
    input wire                                           read_A_21_A_write_data_write,
    output wire [                                   8:0] read_A_21_A_write_resp_peek_dout,
    output wire                                          read_A_21_A_write_resp_peek_empty_n,
    input wire                                           read_A_21_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_21_A_write_resp_s_dout,
    output wire                                          read_A_21_A_write_resp_s_empty_n,
    input wire                                           read_A_21_A_write_resp_s_read,
    output wire [                                  31:0] read_A_21_P_N,
    output wire                                          read_A_21_ap_clk,
    input wire                                           read_A_21_ap_done,
    input wire                                           read_A_21_ap_idle,
    input wire                                           read_A_21_ap_ready,
    output wire                                          read_A_21_ap_rst_n,
    output wire                                          read_A_21_ap_start,
    input wire  [                                 512:0] read_A_21_fifo_A_din,
    output wire                                          read_A_21_fifo_A_full_n,
    input wire                                           read_A_21_fifo_A_write,
    output wire [                                  31:0] read_A_22_A_len,
    output wire [                                  63:0] read_A_22_A_read_addr_offset,
    input wire  [                                  63:0] read_A_22_A_read_addr_s_din,
    output wire                                          read_A_22_A_read_addr_s_full_n,
    input wire                                           read_A_22_A_read_addr_s_write,
    output wire [                                 256:0] read_A_22_A_read_data_peek_dout,
    output wire                                          read_A_22_A_read_data_peek_empty_n,
    input wire                                           read_A_22_A_read_data_peek_read,
    output wire [                                 256:0] read_A_22_A_read_data_s_dout,
    output wire                                          read_A_22_A_read_data_s_empty_n,
    input wire                                           read_A_22_A_read_data_s_read,
    output wire [                                  63:0] read_A_22_A_write_addr_offset,
    input wire  [                                  63:0] read_A_22_A_write_addr_s_din,
    output wire                                          read_A_22_A_write_addr_s_full_n,
    input wire                                           read_A_22_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_22_A_write_data_din,
    output wire                                          read_A_22_A_write_data_full_n,
    input wire                                           read_A_22_A_write_data_write,
    output wire [                                   8:0] read_A_22_A_write_resp_peek_dout,
    output wire                                          read_A_22_A_write_resp_peek_empty_n,
    input wire                                           read_A_22_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_22_A_write_resp_s_dout,
    output wire                                          read_A_22_A_write_resp_s_empty_n,
    input wire                                           read_A_22_A_write_resp_s_read,
    output wire [                                  31:0] read_A_22_P_N,
    output wire                                          read_A_22_ap_clk,
    input wire                                           read_A_22_ap_done,
    input wire                                           read_A_22_ap_idle,
    input wire                                           read_A_22_ap_ready,
    output wire                                          read_A_22_ap_rst_n,
    output wire                                          read_A_22_ap_start,
    input wire  [                                 512:0] read_A_22_fifo_A_din,
    output wire                                          read_A_22_fifo_A_full_n,
    input wire                                           read_A_22_fifo_A_write,
    output wire [                                  31:0] read_A_23_A_len,
    output wire [                                  63:0] read_A_23_A_read_addr_offset,
    input wire  [                                  63:0] read_A_23_A_read_addr_s_din,
    output wire                                          read_A_23_A_read_addr_s_full_n,
    input wire                                           read_A_23_A_read_addr_s_write,
    output wire [                                 256:0] read_A_23_A_read_data_peek_dout,
    output wire                                          read_A_23_A_read_data_peek_empty_n,
    input wire                                           read_A_23_A_read_data_peek_read,
    output wire [                                 256:0] read_A_23_A_read_data_s_dout,
    output wire                                          read_A_23_A_read_data_s_empty_n,
    input wire                                           read_A_23_A_read_data_s_read,
    output wire [                                  63:0] read_A_23_A_write_addr_offset,
    input wire  [                                  63:0] read_A_23_A_write_addr_s_din,
    output wire                                          read_A_23_A_write_addr_s_full_n,
    input wire                                           read_A_23_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_23_A_write_data_din,
    output wire                                          read_A_23_A_write_data_full_n,
    input wire                                           read_A_23_A_write_data_write,
    output wire [                                   8:0] read_A_23_A_write_resp_peek_dout,
    output wire                                          read_A_23_A_write_resp_peek_empty_n,
    input wire                                           read_A_23_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_23_A_write_resp_s_dout,
    output wire                                          read_A_23_A_write_resp_s_empty_n,
    input wire                                           read_A_23_A_write_resp_s_read,
    output wire [                                  31:0] read_A_23_P_N,
    output wire                                          read_A_23_ap_clk,
    input wire                                           read_A_23_ap_done,
    input wire                                           read_A_23_ap_idle,
    input wire                                           read_A_23_ap_ready,
    output wire                                          read_A_23_ap_rst_n,
    output wire                                          read_A_23_ap_start,
    input wire  [                                 512:0] read_A_23_fifo_A_din,
    output wire                                          read_A_23_fifo_A_full_n,
    input wire                                           read_A_23_fifo_A_write,
    output wire [                                  31:0] read_A_24_A_len,
    output wire [                                  63:0] read_A_24_A_read_addr_offset,
    input wire  [                                  63:0] read_A_24_A_read_addr_s_din,
    output wire                                          read_A_24_A_read_addr_s_full_n,
    input wire                                           read_A_24_A_read_addr_s_write,
    output wire [                                 256:0] read_A_24_A_read_data_peek_dout,
    output wire                                          read_A_24_A_read_data_peek_empty_n,
    input wire                                           read_A_24_A_read_data_peek_read,
    output wire [                                 256:0] read_A_24_A_read_data_s_dout,
    output wire                                          read_A_24_A_read_data_s_empty_n,
    input wire                                           read_A_24_A_read_data_s_read,
    output wire [                                  63:0] read_A_24_A_write_addr_offset,
    input wire  [                                  63:0] read_A_24_A_write_addr_s_din,
    output wire                                          read_A_24_A_write_addr_s_full_n,
    input wire                                           read_A_24_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_24_A_write_data_din,
    output wire                                          read_A_24_A_write_data_full_n,
    input wire                                           read_A_24_A_write_data_write,
    output wire [                                   8:0] read_A_24_A_write_resp_peek_dout,
    output wire                                          read_A_24_A_write_resp_peek_empty_n,
    input wire                                           read_A_24_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_24_A_write_resp_s_dout,
    output wire                                          read_A_24_A_write_resp_s_empty_n,
    input wire                                           read_A_24_A_write_resp_s_read,
    output wire [                                  31:0] read_A_24_P_N,
    output wire                                          read_A_24_ap_clk,
    input wire                                           read_A_24_ap_done,
    input wire                                           read_A_24_ap_idle,
    input wire                                           read_A_24_ap_ready,
    output wire                                          read_A_24_ap_rst_n,
    output wire                                          read_A_24_ap_start,
    input wire  [                                 512:0] read_A_24_fifo_A_din,
    output wire                                          read_A_24_fifo_A_full_n,
    input wire                                           read_A_24_fifo_A_write,
    output wire [                                  31:0] read_A_25_A_len,
    output wire [                                  63:0] read_A_25_A_read_addr_offset,
    input wire  [                                  63:0] read_A_25_A_read_addr_s_din,
    output wire                                          read_A_25_A_read_addr_s_full_n,
    input wire                                           read_A_25_A_read_addr_s_write,
    output wire [                                 256:0] read_A_25_A_read_data_peek_dout,
    output wire                                          read_A_25_A_read_data_peek_empty_n,
    input wire                                           read_A_25_A_read_data_peek_read,
    output wire [                                 256:0] read_A_25_A_read_data_s_dout,
    output wire                                          read_A_25_A_read_data_s_empty_n,
    input wire                                           read_A_25_A_read_data_s_read,
    output wire [                                  63:0] read_A_25_A_write_addr_offset,
    input wire  [                                  63:0] read_A_25_A_write_addr_s_din,
    output wire                                          read_A_25_A_write_addr_s_full_n,
    input wire                                           read_A_25_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_25_A_write_data_din,
    output wire                                          read_A_25_A_write_data_full_n,
    input wire                                           read_A_25_A_write_data_write,
    output wire [                                   8:0] read_A_25_A_write_resp_peek_dout,
    output wire                                          read_A_25_A_write_resp_peek_empty_n,
    input wire                                           read_A_25_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_25_A_write_resp_s_dout,
    output wire                                          read_A_25_A_write_resp_s_empty_n,
    input wire                                           read_A_25_A_write_resp_s_read,
    output wire [                                  31:0] read_A_25_P_N,
    output wire                                          read_A_25_ap_clk,
    input wire                                           read_A_25_ap_done,
    input wire                                           read_A_25_ap_idle,
    input wire                                           read_A_25_ap_ready,
    output wire                                          read_A_25_ap_rst_n,
    output wire                                          read_A_25_ap_start,
    input wire  [                                 512:0] read_A_25_fifo_A_din,
    output wire                                          read_A_25_fifo_A_full_n,
    input wire                                           read_A_25_fifo_A_write,
    output wire [                                  31:0] read_A_26_A_len,
    output wire [                                  63:0] read_A_26_A_read_addr_offset,
    input wire  [                                  63:0] read_A_26_A_read_addr_s_din,
    output wire                                          read_A_26_A_read_addr_s_full_n,
    input wire                                           read_A_26_A_read_addr_s_write,
    output wire [                                 256:0] read_A_26_A_read_data_peek_dout,
    output wire                                          read_A_26_A_read_data_peek_empty_n,
    input wire                                           read_A_26_A_read_data_peek_read,
    output wire [                                 256:0] read_A_26_A_read_data_s_dout,
    output wire                                          read_A_26_A_read_data_s_empty_n,
    input wire                                           read_A_26_A_read_data_s_read,
    output wire [                                  63:0] read_A_26_A_write_addr_offset,
    input wire  [                                  63:0] read_A_26_A_write_addr_s_din,
    output wire                                          read_A_26_A_write_addr_s_full_n,
    input wire                                           read_A_26_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_26_A_write_data_din,
    output wire                                          read_A_26_A_write_data_full_n,
    input wire                                           read_A_26_A_write_data_write,
    output wire [                                   8:0] read_A_26_A_write_resp_peek_dout,
    output wire                                          read_A_26_A_write_resp_peek_empty_n,
    input wire                                           read_A_26_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_26_A_write_resp_s_dout,
    output wire                                          read_A_26_A_write_resp_s_empty_n,
    input wire                                           read_A_26_A_write_resp_s_read,
    output wire [                                  31:0] read_A_26_P_N,
    output wire                                          read_A_26_ap_clk,
    input wire                                           read_A_26_ap_done,
    input wire                                           read_A_26_ap_idle,
    input wire                                           read_A_26_ap_ready,
    output wire                                          read_A_26_ap_rst_n,
    output wire                                          read_A_26_ap_start,
    input wire  [                                 512:0] read_A_26_fifo_A_din,
    output wire                                          read_A_26_fifo_A_full_n,
    input wire                                           read_A_26_fifo_A_write,
    output wire [                                  31:0] read_A_27_A_len,
    output wire [                                  63:0] read_A_27_A_read_addr_offset,
    input wire  [                                  63:0] read_A_27_A_read_addr_s_din,
    output wire                                          read_A_27_A_read_addr_s_full_n,
    input wire                                           read_A_27_A_read_addr_s_write,
    output wire [                                 256:0] read_A_27_A_read_data_peek_dout,
    output wire                                          read_A_27_A_read_data_peek_empty_n,
    input wire                                           read_A_27_A_read_data_peek_read,
    output wire [                                 256:0] read_A_27_A_read_data_s_dout,
    output wire                                          read_A_27_A_read_data_s_empty_n,
    input wire                                           read_A_27_A_read_data_s_read,
    output wire [                                  63:0] read_A_27_A_write_addr_offset,
    input wire  [                                  63:0] read_A_27_A_write_addr_s_din,
    output wire                                          read_A_27_A_write_addr_s_full_n,
    input wire                                           read_A_27_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_27_A_write_data_din,
    output wire                                          read_A_27_A_write_data_full_n,
    input wire                                           read_A_27_A_write_data_write,
    output wire [                                   8:0] read_A_27_A_write_resp_peek_dout,
    output wire                                          read_A_27_A_write_resp_peek_empty_n,
    input wire                                           read_A_27_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_27_A_write_resp_s_dout,
    output wire                                          read_A_27_A_write_resp_s_empty_n,
    input wire                                           read_A_27_A_write_resp_s_read,
    output wire [                                  31:0] read_A_27_P_N,
    output wire                                          read_A_27_ap_clk,
    input wire                                           read_A_27_ap_done,
    input wire                                           read_A_27_ap_idle,
    input wire                                           read_A_27_ap_ready,
    output wire                                          read_A_27_ap_rst_n,
    output wire                                          read_A_27_ap_start,
    input wire  [                                 512:0] read_A_27_fifo_A_din,
    output wire                                          read_A_27_fifo_A_full_n,
    input wire                                           read_A_27_fifo_A_write,
    output wire [                                  31:0] read_A_28_A_len,
    output wire [                                  63:0] read_A_28_A_read_addr_offset,
    input wire  [                                  63:0] read_A_28_A_read_addr_s_din,
    output wire                                          read_A_28_A_read_addr_s_full_n,
    input wire                                           read_A_28_A_read_addr_s_write,
    output wire [                                 256:0] read_A_28_A_read_data_peek_dout,
    output wire                                          read_A_28_A_read_data_peek_empty_n,
    input wire                                           read_A_28_A_read_data_peek_read,
    output wire [                                 256:0] read_A_28_A_read_data_s_dout,
    output wire                                          read_A_28_A_read_data_s_empty_n,
    input wire                                           read_A_28_A_read_data_s_read,
    output wire [                                  63:0] read_A_28_A_write_addr_offset,
    input wire  [                                  63:0] read_A_28_A_write_addr_s_din,
    output wire                                          read_A_28_A_write_addr_s_full_n,
    input wire                                           read_A_28_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_28_A_write_data_din,
    output wire                                          read_A_28_A_write_data_full_n,
    input wire                                           read_A_28_A_write_data_write,
    output wire [                                   8:0] read_A_28_A_write_resp_peek_dout,
    output wire                                          read_A_28_A_write_resp_peek_empty_n,
    input wire                                           read_A_28_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_28_A_write_resp_s_dout,
    output wire                                          read_A_28_A_write_resp_s_empty_n,
    input wire                                           read_A_28_A_write_resp_s_read,
    output wire [                                  31:0] read_A_28_P_N,
    output wire                                          read_A_28_ap_clk,
    input wire                                           read_A_28_ap_done,
    input wire                                           read_A_28_ap_idle,
    input wire                                           read_A_28_ap_ready,
    output wire                                          read_A_28_ap_rst_n,
    output wire                                          read_A_28_ap_start,
    input wire  [                                 512:0] read_A_28_fifo_A_din,
    output wire                                          read_A_28_fifo_A_full_n,
    input wire                                           read_A_28_fifo_A_write,
    output wire [                                  31:0] read_A_29_A_len,
    output wire [                                  63:0] read_A_29_A_read_addr_offset,
    input wire  [                                  63:0] read_A_29_A_read_addr_s_din,
    output wire                                          read_A_29_A_read_addr_s_full_n,
    input wire                                           read_A_29_A_read_addr_s_write,
    output wire [                                 256:0] read_A_29_A_read_data_peek_dout,
    output wire                                          read_A_29_A_read_data_peek_empty_n,
    input wire                                           read_A_29_A_read_data_peek_read,
    output wire [                                 256:0] read_A_29_A_read_data_s_dout,
    output wire                                          read_A_29_A_read_data_s_empty_n,
    input wire                                           read_A_29_A_read_data_s_read,
    output wire [                                  63:0] read_A_29_A_write_addr_offset,
    input wire  [                                  63:0] read_A_29_A_write_addr_s_din,
    output wire                                          read_A_29_A_write_addr_s_full_n,
    input wire                                           read_A_29_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_29_A_write_data_din,
    output wire                                          read_A_29_A_write_data_full_n,
    input wire                                           read_A_29_A_write_data_write,
    output wire [                                   8:0] read_A_29_A_write_resp_peek_dout,
    output wire                                          read_A_29_A_write_resp_peek_empty_n,
    input wire                                           read_A_29_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_29_A_write_resp_s_dout,
    output wire                                          read_A_29_A_write_resp_s_empty_n,
    input wire                                           read_A_29_A_write_resp_s_read,
    output wire [                                  31:0] read_A_29_P_N,
    output wire                                          read_A_29_ap_clk,
    input wire                                           read_A_29_ap_done,
    input wire                                           read_A_29_ap_idle,
    input wire                                           read_A_29_ap_ready,
    output wire                                          read_A_29_ap_rst_n,
    output wire                                          read_A_29_ap_start,
    input wire  [                                 512:0] read_A_29_fifo_A_din,
    output wire                                          read_A_29_fifo_A_full_n,
    input wire                                           read_A_29_fifo_A_write,
    output wire [                                  31:0] read_A_30_A_len,
    output wire [                                  63:0] read_A_30_A_read_addr_offset,
    input wire  [                                  63:0] read_A_30_A_read_addr_s_din,
    output wire                                          read_A_30_A_read_addr_s_full_n,
    input wire                                           read_A_30_A_read_addr_s_write,
    output wire [                                 256:0] read_A_30_A_read_data_peek_dout,
    output wire                                          read_A_30_A_read_data_peek_empty_n,
    input wire                                           read_A_30_A_read_data_peek_read,
    output wire [                                 256:0] read_A_30_A_read_data_s_dout,
    output wire                                          read_A_30_A_read_data_s_empty_n,
    input wire                                           read_A_30_A_read_data_s_read,
    output wire [                                  63:0] read_A_30_A_write_addr_offset,
    input wire  [                                  63:0] read_A_30_A_write_addr_s_din,
    output wire                                          read_A_30_A_write_addr_s_full_n,
    input wire                                           read_A_30_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_30_A_write_data_din,
    output wire                                          read_A_30_A_write_data_full_n,
    input wire                                           read_A_30_A_write_data_write,
    output wire [                                   8:0] read_A_30_A_write_resp_peek_dout,
    output wire                                          read_A_30_A_write_resp_peek_empty_n,
    input wire                                           read_A_30_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_30_A_write_resp_s_dout,
    output wire                                          read_A_30_A_write_resp_s_empty_n,
    input wire                                           read_A_30_A_write_resp_s_read,
    output wire [                                  31:0] read_A_30_P_N,
    output wire                                          read_A_30_ap_clk,
    input wire                                           read_A_30_ap_done,
    input wire                                           read_A_30_ap_idle,
    input wire                                           read_A_30_ap_ready,
    output wire                                          read_A_30_ap_rst_n,
    output wire                                          read_A_30_ap_start,
    input wire  [                                 512:0] read_A_30_fifo_A_din,
    output wire                                          read_A_30_fifo_A_full_n,
    input wire                                           read_A_30_fifo_A_write,
    output wire [                                  31:0] read_A_31_A_len,
    output wire [                                  63:0] read_A_31_A_read_addr_offset,
    input wire  [                                  63:0] read_A_31_A_read_addr_s_din,
    output wire                                          read_A_31_A_read_addr_s_full_n,
    input wire                                           read_A_31_A_read_addr_s_write,
    output wire [                                 256:0] read_A_31_A_read_data_peek_dout,
    output wire                                          read_A_31_A_read_data_peek_empty_n,
    input wire                                           read_A_31_A_read_data_peek_read,
    output wire [                                 256:0] read_A_31_A_read_data_s_dout,
    output wire                                          read_A_31_A_read_data_s_empty_n,
    input wire                                           read_A_31_A_read_data_s_read,
    output wire [                                  63:0] read_A_31_A_write_addr_offset,
    input wire  [                                  63:0] read_A_31_A_write_addr_s_din,
    output wire                                          read_A_31_A_write_addr_s_full_n,
    input wire                                           read_A_31_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_31_A_write_data_din,
    output wire                                          read_A_31_A_write_data_full_n,
    input wire                                           read_A_31_A_write_data_write,
    output wire [                                   8:0] read_A_31_A_write_resp_peek_dout,
    output wire                                          read_A_31_A_write_resp_peek_empty_n,
    input wire                                           read_A_31_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_31_A_write_resp_s_dout,
    output wire                                          read_A_31_A_write_resp_s_empty_n,
    input wire                                           read_A_31_A_write_resp_s_read,
    output wire [                                  31:0] read_A_31_P_N,
    output wire                                          read_A_31_ap_clk,
    input wire                                           read_A_31_ap_done,
    input wire                                           read_A_31_ap_idle,
    input wire                                           read_A_31_ap_ready,
    output wire                                          read_A_31_ap_rst_n,
    output wire                                          read_A_31_ap_start,
    input wire  [                                 512:0] read_A_31_fifo_A_din,
    output wire                                          read_A_31_fifo_A_full_n,
    input wire                                           read_A_31_fifo_A_write,
    output wire [                                  31:0] read_A_32_A_len,
    output wire [                                  63:0] read_A_32_A_read_addr_offset,
    input wire  [                                  63:0] read_A_32_A_read_addr_s_din,
    output wire                                          read_A_32_A_read_addr_s_full_n,
    input wire                                           read_A_32_A_read_addr_s_write,
    output wire [                                 256:0] read_A_32_A_read_data_peek_dout,
    output wire                                          read_A_32_A_read_data_peek_empty_n,
    input wire                                           read_A_32_A_read_data_peek_read,
    output wire [                                 256:0] read_A_32_A_read_data_s_dout,
    output wire                                          read_A_32_A_read_data_s_empty_n,
    input wire                                           read_A_32_A_read_data_s_read,
    output wire [                                  63:0] read_A_32_A_write_addr_offset,
    input wire  [                                  63:0] read_A_32_A_write_addr_s_din,
    output wire                                          read_A_32_A_write_addr_s_full_n,
    input wire                                           read_A_32_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_32_A_write_data_din,
    output wire                                          read_A_32_A_write_data_full_n,
    input wire                                           read_A_32_A_write_data_write,
    output wire [                                   8:0] read_A_32_A_write_resp_peek_dout,
    output wire                                          read_A_32_A_write_resp_peek_empty_n,
    input wire                                           read_A_32_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_32_A_write_resp_s_dout,
    output wire                                          read_A_32_A_write_resp_s_empty_n,
    input wire                                           read_A_32_A_write_resp_s_read,
    output wire [                                  31:0] read_A_32_P_N,
    output wire                                          read_A_32_ap_clk,
    input wire                                           read_A_32_ap_done,
    input wire                                           read_A_32_ap_idle,
    input wire                                           read_A_32_ap_ready,
    output wire                                          read_A_32_ap_rst_n,
    output wire                                          read_A_32_ap_start,
    input wire  [                                 512:0] read_A_32_fifo_A_din,
    output wire                                          read_A_32_fifo_A_full_n,
    input wire                                           read_A_32_fifo_A_write,
    output wire [                                  31:0] read_A_33_A_len,
    output wire [                                  63:0] read_A_33_A_read_addr_offset,
    input wire  [                                  63:0] read_A_33_A_read_addr_s_din,
    output wire                                          read_A_33_A_read_addr_s_full_n,
    input wire                                           read_A_33_A_read_addr_s_write,
    output wire [                                 256:0] read_A_33_A_read_data_peek_dout,
    output wire                                          read_A_33_A_read_data_peek_empty_n,
    input wire                                           read_A_33_A_read_data_peek_read,
    output wire [                                 256:0] read_A_33_A_read_data_s_dout,
    output wire                                          read_A_33_A_read_data_s_empty_n,
    input wire                                           read_A_33_A_read_data_s_read,
    output wire [                                  63:0] read_A_33_A_write_addr_offset,
    input wire  [                                  63:0] read_A_33_A_write_addr_s_din,
    output wire                                          read_A_33_A_write_addr_s_full_n,
    input wire                                           read_A_33_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_33_A_write_data_din,
    output wire                                          read_A_33_A_write_data_full_n,
    input wire                                           read_A_33_A_write_data_write,
    output wire [                                   8:0] read_A_33_A_write_resp_peek_dout,
    output wire                                          read_A_33_A_write_resp_peek_empty_n,
    input wire                                           read_A_33_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_33_A_write_resp_s_dout,
    output wire                                          read_A_33_A_write_resp_s_empty_n,
    input wire                                           read_A_33_A_write_resp_s_read,
    output wire [                                  31:0] read_A_33_P_N,
    output wire                                          read_A_33_ap_clk,
    input wire                                           read_A_33_ap_done,
    input wire                                           read_A_33_ap_idle,
    input wire                                           read_A_33_ap_ready,
    output wire                                          read_A_33_ap_rst_n,
    output wire                                          read_A_33_ap_start,
    input wire  [                                 512:0] read_A_33_fifo_A_din,
    output wire                                          read_A_33_fifo_A_full_n,
    input wire                                           read_A_33_fifo_A_write,
    output wire [                                  31:0] read_A_34_A_len,
    output wire [                                  63:0] read_A_34_A_read_addr_offset,
    input wire  [                                  63:0] read_A_34_A_read_addr_s_din,
    output wire                                          read_A_34_A_read_addr_s_full_n,
    input wire                                           read_A_34_A_read_addr_s_write,
    output wire [                                 256:0] read_A_34_A_read_data_peek_dout,
    output wire                                          read_A_34_A_read_data_peek_empty_n,
    input wire                                           read_A_34_A_read_data_peek_read,
    output wire [                                 256:0] read_A_34_A_read_data_s_dout,
    output wire                                          read_A_34_A_read_data_s_empty_n,
    input wire                                           read_A_34_A_read_data_s_read,
    output wire [                                  63:0] read_A_34_A_write_addr_offset,
    input wire  [                                  63:0] read_A_34_A_write_addr_s_din,
    output wire                                          read_A_34_A_write_addr_s_full_n,
    input wire                                           read_A_34_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_34_A_write_data_din,
    output wire                                          read_A_34_A_write_data_full_n,
    input wire                                           read_A_34_A_write_data_write,
    output wire [                                   8:0] read_A_34_A_write_resp_peek_dout,
    output wire                                          read_A_34_A_write_resp_peek_empty_n,
    input wire                                           read_A_34_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_34_A_write_resp_s_dout,
    output wire                                          read_A_34_A_write_resp_s_empty_n,
    input wire                                           read_A_34_A_write_resp_s_read,
    output wire [                                  31:0] read_A_34_P_N,
    output wire                                          read_A_34_ap_clk,
    input wire                                           read_A_34_ap_done,
    input wire                                           read_A_34_ap_idle,
    input wire                                           read_A_34_ap_ready,
    output wire                                          read_A_34_ap_rst_n,
    output wire                                          read_A_34_ap_start,
    input wire  [                                 512:0] read_A_34_fifo_A_din,
    output wire                                          read_A_34_fifo_A_full_n,
    input wire                                           read_A_34_fifo_A_write,
    output wire [                                  31:0] read_A_35_A_len,
    output wire [                                  63:0] read_A_35_A_read_addr_offset,
    input wire  [                                  63:0] read_A_35_A_read_addr_s_din,
    output wire                                          read_A_35_A_read_addr_s_full_n,
    input wire                                           read_A_35_A_read_addr_s_write,
    output wire [                                 256:0] read_A_35_A_read_data_peek_dout,
    output wire                                          read_A_35_A_read_data_peek_empty_n,
    input wire                                           read_A_35_A_read_data_peek_read,
    output wire [                                 256:0] read_A_35_A_read_data_s_dout,
    output wire                                          read_A_35_A_read_data_s_empty_n,
    input wire                                           read_A_35_A_read_data_s_read,
    output wire [                                  63:0] read_A_35_A_write_addr_offset,
    input wire  [                                  63:0] read_A_35_A_write_addr_s_din,
    output wire                                          read_A_35_A_write_addr_s_full_n,
    input wire                                           read_A_35_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_35_A_write_data_din,
    output wire                                          read_A_35_A_write_data_full_n,
    input wire                                           read_A_35_A_write_data_write,
    output wire [                                   8:0] read_A_35_A_write_resp_peek_dout,
    output wire                                          read_A_35_A_write_resp_peek_empty_n,
    input wire                                           read_A_35_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_35_A_write_resp_s_dout,
    output wire                                          read_A_35_A_write_resp_s_empty_n,
    input wire                                           read_A_35_A_write_resp_s_read,
    output wire [                                  31:0] read_A_35_P_N,
    output wire                                          read_A_35_ap_clk,
    input wire                                           read_A_35_ap_done,
    input wire                                           read_A_35_ap_idle,
    input wire                                           read_A_35_ap_ready,
    output wire                                          read_A_35_ap_rst_n,
    output wire                                          read_A_35_ap_start,
    input wire  [                                 512:0] read_A_35_fifo_A_din,
    output wire                                          read_A_35_fifo_A_full_n,
    input wire                                           read_A_35_fifo_A_write,
    output wire [                                  31:0] read_A_36_A_len,
    output wire [                                  63:0] read_A_36_A_read_addr_offset,
    input wire  [                                  63:0] read_A_36_A_read_addr_s_din,
    output wire                                          read_A_36_A_read_addr_s_full_n,
    input wire                                           read_A_36_A_read_addr_s_write,
    output wire [                                 256:0] read_A_36_A_read_data_peek_dout,
    output wire                                          read_A_36_A_read_data_peek_empty_n,
    input wire                                           read_A_36_A_read_data_peek_read,
    output wire [                                 256:0] read_A_36_A_read_data_s_dout,
    output wire                                          read_A_36_A_read_data_s_empty_n,
    input wire                                           read_A_36_A_read_data_s_read,
    output wire [                                  63:0] read_A_36_A_write_addr_offset,
    input wire  [                                  63:0] read_A_36_A_write_addr_s_din,
    output wire                                          read_A_36_A_write_addr_s_full_n,
    input wire                                           read_A_36_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_36_A_write_data_din,
    output wire                                          read_A_36_A_write_data_full_n,
    input wire                                           read_A_36_A_write_data_write,
    output wire [                                   8:0] read_A_36_A_write_resp_peek_dout,
    output wire                                          read_A_36_A_write_resp_peek_empty_n,
    input wire                                           read_A_36_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_36_A_write_resp_s_dout,
    output wire                                          read_A_36_A_write_resp_s_empty_n,
    input wire                                           read_A_36_A_write_resp_s_read,
    output wire [                                  31:0] read_A_36_P_N,
    output wire                                          read_A_36_ap_clk,
    input wire                                           read_A_36_ap_done,
    input wire                                           read_A_36_ap_idle,
    input wire                                           read_A_36_ap_ready,
    output wire                                          read_A_36_ap_rst_n,
    output wire                                          read_A_36_ap_start,
    input wire  [                                 512:0] read_A_36_fifo_A_din,
    output wire                                          read_A_36_fifo_A_full_n,
    input wire                                           read_A_36_fifo_A_write,
    output wire [                                  31:0] read_A_37_A_len,
    output wire [                                  63:0] read_A_37_A_read_addr_offset,
    input wire  [                                  63:0] read_A_37_A_read_addr_s_din,
    output wire                                          read_A_37_A_read_addr_s_full_n,
    input wire                                           read_A_37_A_read_addr_s_write,
    output wire [                                 256:0] read_A_37_A_read_data_peek_dout,
    output wire                                          read_A_37_A_read_data_peek_empty_n,
    input wire                                           read_A_37_A_read_data_peek_read,
    output wire [                                 256:0] read_A_37_A_read_data_s_dout,
    output wire                                          read_A_37_A_read_data_s_empty_n,
    input wire                                           read_A_37_A_read_data_s_read,
    output wire [                                  63:0] read_A_37_A_write_addr_offset,
    input wire  [                                  63:0] read_A_37_A_write_addr_s_din,
    output wire                                          read_A_37_A_write_addr_s_full_n,
    input wire                                           read_A_37_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_37_A_write_data_din,
    output wire                                          read_A_37_A_write_data_full_n,
    input wire                                           read_A_37_A_write_data_write,
    output wire [                                   8:0] read_A_37_A_write_resp_peek_dout,
    output wire                                          read_A_37_A_write_resp_peek_empty_n,
    input wire                                           read_A_37_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_37_A_write_resp_s_dout,
    output wire                                          read_A_37_A_write_resp_s_empty_n,
    input wire                                           read_A_37_A_write_resp_s_read,
    output wire [                                  31:0] read_A_37_P_N,
    output wire                                          read_A_37_ap_clk,
    input wire                                           read_A_37_ap_done,
    input wire                                           read_A_37_ap_idle,
    input wire                                           read_A_37_ap_ready,
    output wire                                          read_A_37_ap_rst_n,
    output wire                                          read_A_37_ap_start,
    input wire  [                                 512:0] read_A_37_fifo_A_din,
    output wire                                          read_A_37_fifo_A_full_n,
    input wire                                           read_A_37_fifo_A_write,
    output wire [                                  31:0] read_A_38_A_len,
    output wire [                                  63:0] read_A_38_A_read_addr_offset,
    input wire  [                                  63:0] read_A_38_A_read_addr_s_din,
    output wire                                          read_A_38_A_read_addr_s_full_n,
    input wire                                           read_A_38_A_read_addr_s_write,
    output wire [                                 256:0] read_A_38_A_read_data_peek_dout,
    output wire                                          read_A_38_A_read_data_peek_empty_n,
    input wire                                           read_A_38_A_read_data_peek_read,
    output wire [                                 256:0] read_A_38_A_read_data_s_dout,
    output wire                                          read_A_38_A_read_data_s_empty_n,
    input wire                                           read_A_38_A_read_data_s_read,
    output wire [                                  63:0] read_A_38_A_write_addr_offset,
    input wire  [                                  63:0] read_A_38_A_write_addr_s_din,
    output wire                                          read_A_38_A_write_addr_s_full_n,
    input wire                                           read_A_38_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_38_A_write_data_din,
    output wire                                          read_A_38_A_write_data_full_n,
    input wire                                           read_A_38_A_write_data_write,
    output wire [                                   8:0] read_A_38_A_write_resp_peek_dout,
    output wire                                          read_A_38_A_write_resp_peek_empty_n,
    input wire                                           read_A_38_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_38_A_write_resp_s_dout,
    output wire                                          read_A_38_A_write_resp_s_empty_n,
    input wire                                           read_A_38_A_write_resp_s_read,
    output wire [                                  31:0] read_A_38_P_N,
    output wire                                          read_A_38_ap_clk,
    input wire                                           read_A_38_ap_done,
    input wire                                           read_A_38_ap_idle,
    input wire                                           read_A_38_ap_ready,
    output wire                                          read_A_38_ap_rst_n,
    output wire                                          read_A_38_ap_start,
    input wire  [                                 512:0] read_A_38_fifo_A_din,
    output wire                                          read_A_38_fifo_A_full_n,
    input wire                                           read_A_38_fifo_A_write,
    output wire [                                  31:0] read_A_39_A_len,
    output wire [                                  63:0] read_A_39_A_read_addr_offset,
    input wire  [                                  63:0] read_A_39_A_read_addr_s_din,
    output wire                                          read_A_39_A_read_addr_s_full_n,
    input wire                                           read_A_39_A_read_addr_s_write,
    output wire [                                 256:0] read_A_39_A_read_data_peek_dout,
    output wire                                          read_A_39_A_read_data_peek_empty_n,
    input wire                                           read_A_39_A_read_data_peek_read,
    output wire [                                 256:0] read_A_39_A_read_data_s_dout,
    output wire                                          read_A_39_A_read_data_s_empty_n,
    input wire                                           read_A_39_A_read_data_s_read,
    output wire [                                  63:0] read_A_39_A_write_addr_offset,
    input wire  [                                  63:0] read_A_39_A_write_addr_s_din,
    output wire                                          read_A_39_A_write_addr_s_full_n,
    input wire                                           read_A_39_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_39_A_write_data_din,
    output wire                                          read_A_39_A_write_data_full_n,
    input wire                                           read_A_39_A_write_data_write,
    output wire [                                   8:0] read_A_39_A_write_resp_peek_dout,
    output wire                                          read_A_39_A_write_resp_peek_empty_n,
    input wire                                           read_A_39_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_39_A_write_resp_s_dout,
    output wire                                          read_A_39_A_write_resp_s_empty_n,
    input wire                                           read_A_39_A_write_resp_s_read,
    output wire [                                  31:0] read_A_39_P_N,
    output wire                                          read_A_39_ap_clk,
    input wire                                           read_A_39_ap_done,
    input wire                                           read_A_39_ap_idle,
    input wire                                           read_A_39_ap_ready,
    output wire                                          read_A_39_ap_rst_n,
    output wire                                          read_A_39_ap_start,
    input wire  [                                 512:0] read_A_39_fifo_A_din,
    output wire                                          read_A_39_fifo_A_full_n,
    input wire                                           read_A_39_fifo_A_write,
    output wire [                                  31:0] read_A_40_A_len,
    output wire [                                  63:0] read_A_40_A_read_addr_offset,
    input wire  [                                  63:0] read_A_40_A_read_addr_s_din,
    output wire                                          read_A_40_A_read_addr_s_full_n,
    input wire                                           read_A_40_A_read_addr_s_write,
    output wire [                                 256:0] read_A_40_A_read_data_peek_dout,
    output wire                                          read_A_40_A_read_data_peek_empty_n,
    input wire                                           read_A_40_A_read_data_peek_read,
    output wire [                                 256:0] read_A_40_A_read_data_s_dout,
    output wire                                          read_A_40_A_read_data_s_empty_n,
    input wire                                           read_A_40_A_read_data_s_read,
    output wire [                                  63:0] read_A_40_A_write_addr_offset,
    input wire  [                                  63:0] read_A_40_A_write_addr_s_din,
    output wire                                          read_A_40_A_write_addr_s_full_n,
    input wire                                           read_A_40_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_40_A_write_data_din,
    output wire                                          read_A_40_A_write_data_full_n,
    input wire                                           read_A_40_A_write_data_write,
    output wire [                                   8:0] read_A_40_A_write_resp_peek_dout,
    output wire                                          read_A_40_A_write_resp_peek_empty_n,
    input wire                                           read_A_40_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_40_A_write_resp_s_dout,
    output wire                                          read_A_40_A_write_resp_s_empty_n,
    input wire                                           read_A_40_A_write_resp_s_read,
    output wire [                                  31:0] read_A_40_P_N,
    output wire                                          read_A_40_ap_clk,
    input wire                                           read_A_40_ap_done,
    input wire                                           read_A_40_ap_idle,
    input wire                                           read_A_40_ap_ready,
    output wire                                          read_A_40_ap_rst_n,
    output wire                                          read_A_40_ap_start,
    input wire  [                                 512:0] read_A_40_fifo_A_din,
    output wire                                          read_A_40_fifo_A_full_n,
    input wire                                           read_A_40_fifo_A_write,
    output wire [                                  31:0] read_A_41_A_len,
    output wire [                                  63:0] read_A_41_A_read_addr_offset,
    input wire  [                                  63:0] read_A_41_A_read_addr_s_din,
    output wire                                          read_A_41_A_read_addr_s_full_n,
    input wire                                           read_A_41_A_read_addr_s_write,
    output wire [                                 256:0] read_A_41_A_read_data_peek_dout,
    output wire                                          read_A_41_A_read_data_peek_empty_n,
    input wire                                           read_A_41_A_read_data_peek_read,
    output wire [                                 256:0] read_A_41_A_read_data_s_dout,
    output wire                                          read_A_41_A_read_data_s_empty_n,
    input wire                                           read_A_41_A_read_data_s_read,
    output wire [                                  63:0] read_A_41_A_write_addr_offset,
    input wire  [                                  63:0] read_A_41_A_write_addr_s_din,
    output wire                                          read_A_41_A_write_addr_s_full_n,
    input wire                                           read_A_41_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_41_A_write_data_din,
    output wire                                          read_A_41_A_write_data_full_n,
    input wire                                           read_A_41_A_write_data_write,
    output wire [                                   8:0] read_A_41_A_write_resp_peek_dout,
    output wire                                          read_A_41_A_write_resp_peek_empty_n,
    input wire                                           read_A_41_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_41_A_write_resp_s_dout,
    output wire                                          read_A_41_A_write_resp_s_empty_n,
    input wire                                           read_A_41_A_write_resp_s_read,
    output wire [                                  31:0] read_A_41_P_N,
    output wire                                          read_A_41_ap_clk,
    input wire                                           read_A_41_ap_done,
    input wire                                           read_A_41_ap_idle,
    input wire                                           read_A_41_ap_ready,
    output wire                                          read_A_41_ap_rst_n,
    output wire                                          read_A_41_ap_start,
    input wire  [                                 512:0] read_A_41_fifo_A_din,
    output wire                                          read_A_41_fifo_A_full_n,
    input wire                                           read_A_41_fifo_A_write,
    output wire [                                  31:0] read_A_42_A_len,
    output wire [                                  63:0] read_A_42_A_read_addr_offset,
    input wire  [                                  63:0] read_A_42_A_read_addr_s_din,
    output wire                                          read_A_42_A_read_addr_s_full_n,
    input wire                                           read_A_42_A_read_addr_s_write,
    output wire [                                 256:0] read_A_42_A_read_data_peek_dout,
    output wire                                          read_A_42_A_read_data_peek_empty_n,
    input wire                                           read_A_42_A_read_data_peek_read,
    output wire [                                 256:0] read_A_42_A_read_data_s_dout,
    output wire                                          read_A_42_A_read_data_s_empty_n,
    input wire                                           read_A_42_A_read_data_s_read,
    output wire [                                  63:0] read_A_42_A_write_addr_offset,
    input wire  [                                  63:0] read_A_42_A_write_addr_s_din,
    output wire                                          read_A_42_A_write_addr_s_full_n,
    input wire                                           read_A_42_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_42_A_write_data_din,
    output wire                                          read_A_42_A_write_data_full_n,
    input wire                                           read_A_42_A_write_data_write,
    output wire [                                   8:0] read_A_42_A_write_resp_peek_dout,
    output wire                                          read_A_42_A_write_resp_peek_empty_n,
    input wire                                           read_A_42_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_42_A_write_resp_s_dout,
    output wire                                          read_A_42_A_write_resp_s_empty_n,
    input wire                                           read_A_42_A_write_resp_s_read,
    output wire [                                  31:0] read_A_42_P_N,
    output wire                                          read_A_42_ap_clk,
    input wire                                           read_A_42_ap_done,
    input wire                                           read_A_42_ap_idle,
    input wire                                           read_A_42_ap_ready,
    output wire                                          read_A_42_ap_rst_n,
    output wire                                          read_A_42_ap_start,
    input wire  [                                 512:0] read_A_42_fifo_A_din,
    output wire                                          read_A_42_fifo_A_full_n,
    input wire                                           read_A_42_fifo_A_write,
    output wire [                                  31:0] read_A_43_A_len,
    output wire [                                  63:0] read_A_43_A_read_addr_offset,
    input wire  [                                  63:0] read_A_43_A_read_addr_s_din,
    output wire                                          read_A_43_A_read_addr_s_full_n,
    input wire                                           read_A_43_A_read_addr_s_write,
    output wire [                                 256:0] read_A_43_A_read_data_peek_dout,
    output wire                                          read_A_43_A_read_data_peek_empty_n,
    input wire                                           read_A_43_A_read_data_peek_read,
    output wire [                                 256:0] read_A_43_A_read_data_s_dout,
    output wire                                          read_A_43_A_read_data_s_empty_n,
    input wire                                           read_A_43_A_read_data_s_read,
    output wire [                                  63:0] read_A_43_A_write_addr_offset,
    input wire  [                                  63:0] read_A_43_A_write_addr_s_din,
    output wire                                          read_A_43_A_write_addr_s_full_n,
    input wire                                           read_A_43_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_43_A_write_data_din,
    output wire                                          read_A_43_A_write_data_full_n,
    input wire                                           read_A_43_A_write_data_write,
    output wire [                                   8:0] read_A_43_A_write_resp_peek_dout,
    output wire                                          read_A_43_A_write_resp_peek_empty_n,
    input wire                                           read_A_43_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_43_A_write_resp_s_dout,
    output wire                                          read_A_43_A_write_resp_s_empty_n,
    input wire                                           read_A_43_A_write_resp_s_read,
    output wire [                                  31:0] read_A_43_P_N,
    output wire                                          read_A_43_ap_clk,
    input wire                                           read_A_43_ap_done,
    input wire                                           read_A_43_ap_idle,
    input wire                                           read_A_43_ap_ready,
    output wire                                          read_A_43_ap_rst_n,
    output wire                                          read_A_43_ap_start,
    input wire  [                                 512:0] read_A_43_fifo_A_din,
    output wire                                          read_A_43_fifo_A_full_n,
    input wire                                           read_A_43_fifo_A_write,
    output wire [                                  31:0] read_A_44_A_len,
    output wire [                                  63:0] read_A_44_A_read_addr_offset,
    input wire  [                                  63:0] read_A_44_A_read_addr_s_din,
    output wire                                          read_A_44_A_read_addr_s_full_n,
    input wire                                           read_A_44_A_read_addr_s_write,
    output wire [                                 256:0] read_A_44_A_read_data_peek_dout,
    output wire                                          read_A_44_A_read_data_peek_empty_n,
    input wire                                           read_A_44_A_read_data_peek_read,
    output wire [                                 256:0] read_A_44_A_read_data_s_dout,
    output wire                                          read_A_44_A_read_data_s_empty_n,
    input wire                                           read_A_44_A_read_data_s_read,
    output wire [                                  63:0] read_A_44_A_write_addr_offset,
    input wire  [                                  63:0] read_A_44_A_write_addr_s_din,
    output wire                                          read_A_44_A_write_addr_s_full_n,
    input wire                                           read_A_44_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_44_A_write_data_din,
    output wire                                          read_A_44_A_write_data_full_n,
    input wire                                           read_A_44_A_write_data_write,
    output wire [                                   8:0] read_A_44_A_write_resp_peek_dout,
    output wire                                          read_A_44_A_write_resp_peek_empty_n,
    input wire                                           read_A_44_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_44_A_write_resp_s_dout,
    output wire                                          read_A_44_A_write_resp_s_empty_n,
    input wire                                           read_A_44_A_write_resp_s_read,
    output wire [                                  31:0] read_A_44_P_N,
    output wire                                          read_A_44_ap_clk,
    input wire                                           read_A_44_ap_done,
    input wire                                           read_A_44_ap_idle,
    input wire                                           read_A_44_ap_ready,
    output wire                                          read_A_44_ap_rst_n,
    output wire                                          read_A_44_ap_start,
    input wire  [                                 512:0] read_A_44_fifo_A_din,
    output wire                                          read_A_44_fifo_A_full_n,
    input wire                                           read_A_44_fifo_A_write,
    output wire [                                  31:0] read_A_45_A_len,
    output wire [                                  63:0] read_A_45_A_read_addr_offset,
    input wire  [                                  63:0] read_A_45_A_read_addr_s_din,
    output wire                                          read_A_45_A_read_addr_s_full_n,
    input wire                                           read_A_45_A_read_addr_s_write,
    output wire [                                 256:0] read_A_45_A_read_data_peek_dout,
    output wire                                          read_A_45_A_read_data_peek_empty_n,
    input wire                                           read_A_45_A_read_data_peek_read,
    output wire [                                 256:0] read_A_45_A_read_data_s_dout,
    output wire                                          read_A_45_A_read_data_s_empty_n,
    input wire                                           read_A_45_A_read_data_s_read,
    output wire [                                  63:0] read_A_45_A_write_addr_offset,
    input wire  [                                  63:0] read_A_45_A_write_addr_s_din,
    output wire                                          read_A_45_A_write_addr_s_full_n,
    input wire                                           read_A_45_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_45_A_write_data_din,
    output wire                                          read_A_45_A_write_data_full_n,
    input wire                                           read_A_45_A_write_data_write,
    output wire [                                   8:0] read_A_45_A_write_resp_peek_dout,
    output wire                                          read_A_45_A_write_resp_peek_empty_n,
    input wire                                           read_A_45_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_45_A_write_resp_s_dout,
    output wire                                          read_A_45_A_write_resp_s_empty_n,
    input wire                                           read_A_45_A_write_resp_s_read,
    output wire [                                  31:0] read_A_45_P_N,
    output wire                                          read_A_45_ap_clk,
    input wire                                           read_A_45_ap_done,
    input wire                                           read_A_45_ap_idle,
    input wire                                           read_A_45_ap_ready,
    output wire                                          read_A_45_ap_rst_n,
    output wire                                          read_A_45_ap_start,
    input wire  [                                 512:0] read_A_45_fifo_A_din,
    output wire                                          read_A_45_fifo_A_full_n,
    input wire                                           read_A_45_fifo_A_write,
    output wire [                                  31:0] read_A_46_A_len,
    output wire [                                  63:0] read_A_46_A_read_addr_offset,
    input wire  [                                  63:0] read_A_46_A_read_addr_s_din,
    output wire                                          read_A_46_A_read_addr_s_full_n,
    input wire                                           read_A_46_A_read_addr_s_write,
    output wire [                                 256:0] read_A_46_A_read_data_peek_dout,
    output wire                                          read_A_46_A_read_data_peek_empty_n,
    input wire                                           read_A_46_A_read_data_peek_read,
    output wire [                                 256:0] read_A_46_A_read_data_s_dout,
    output wire                                          read_A_46_A_read_data_s_empty_n,
    input wire                                           read_A_46_A_read_data_s_read,
    output wire [                                  63:0] read_A_46_A_write_addr_offset,
    input wire  [                                  63:0] read_A_46_A_write_addr_s_din,
    output wire                                          read_A_46_A_write_addr_s_full_n,
    input wire                                           read_A_46_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_46_A_write_data_din,
    output wire                                          read_A_46_A_write_data_full_n,
    input wire                                           read_A_46_A_write_data_write,
    output wire [                                   8:0] read_A_46_A_write_resp_peek_dout,
    output wire                                          read_A_46_A_write_resp_peek_empty_n,
    input wire                                           read_A_46_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_46_A_write_resp_s_dout,
    output wire                                          read_A_46_A_write_resp_s_empty_n,
    input wire                                           read_A_46_A_write_resp_s_read,
    output wire [                                  31:0] read_A_46_P_N,
    output wire                                          read_A_46_ap_clk,
    input wire                                           read_A_46_ap_done,
    input wire                                           read_A_46_ap_idle,
    input wire                                           read_A_46_ap_ready,
    output wire                                          read_A_46_ap_rst_n,
    output wire                                          read_A_46_ap_start,
    input wire  [                                 512:0] read_A_46_fifo_A_din,
    output wire                                          read_A_46_fifo_A_full_n,
    input wire                                           read_A_46_fifo_A_write,
    output wire [                                  31:0] read_A_47_A_len,
    output wire [                                  63:0] read_A_47_A_read_addr_offset,
    input wire  [                                  63:0] read_A_47_A_read_addr_s_din,
    output wire                                          read_A_47_A_read_addr_s_full_n,
    input wire                                           read_A_47_A_read_addr_s_write,
    output wire [                                 256:0] read_A_47_A_read_data_peek_dout,
    output wire                                          read_A_47_A_read_data_peek_empty_n,
    input wire                                           read_A_47_A_read_data_peek_read,
    output wire [                                 256:0] read_A_47_A_read_data_s_dout,
    output wire                                          read_A_47_A_read_data_s_empty_n,
    input wire                                           read_A_47_A_read_data_s_read,
    output wire [                                  63:0] read_A_47_A_write_addr_offset,
    input wire  [                                  63:0] read_A_47_A_write_addr_s_din,
    output wire                                          read_A_47_A_write_addr_s_full_n,
    input wire                                           read_A_47_A_write_addr_s_write,
    input wire  [                                 256:0] read_A_47_A_write_data_din,
    output wire                                          read_A_47_A_write_data_full_n,
    input wire                                           read_A_47_A_write_data_write,
    output wire [                                   8:0] read_A_47_A_write_resp_peek_dout,
    output wire                                          read_A_47_A_write_resp_peek_empty_n,
    input wire                                           read_A_47_A_write_resp_peek_read,
    output wire [                                   8:0] read_A_47_A_write_resp_s_dout,
    output wire                                          read_A_47_A_write_resp_s_empty_n,
    input wire                                           read_A_47_A_write_resp_s_read,
    output wire [                                  31:0] read_A_47_P_N,
    output wire                                          read_A_47_ap_clk,
    input wire                                           read_A_47_ap_done,
    input wire                                           read_A_47_ap_idle,
    input wire                                           read_A_47_ap_ready,
    output wire                                          read_A_47_ap_rst_n,
    output wire                                          read_A_47_ap_start,
    input wire  [                                 512:0] read_A_47_fifo_A_din,
    output wire                                          read_A_47_fifo_A_full_n,
    input wire                                           read_A_47_fifo_A_write,
    output wire [                                  31:0] read_X_0_K,
    output wire [                                  31:0] read_X_0_P_N,
    output wire                                          read_X_0_ap_clk,
    input wire                                           read_X_0_ap_done,
    input wire                                           read_X_0_ap_idle,
    input wire                                           read_X_0_ap_ready,
    output wire                                          read_X_0_ap_rst_n,
    output wire                                          read_X_0_ap_start,
    input wire  [                                 512:0] read_X_0_fifo_X_din,
    output wire                                          read_X_0_fifo_X_full_n,
    input wire                                           read_X_0_fifo_X_write,
    output wire [                                  63:0] read_X_0_vec_X_read_addr_offset,
    input wire  [                                  63:0] read_X_0_vec_X_read_addr_s_din,
    output wire                                          read_X_0_vec_X_read_addr_s_full_n,
    input wire                                           read_X_0_vec_X_read_addr_s_write,
    output wire [                                 256:0] read_X_0_vec_X_read_data_peek_dout,
    output wire                                          read_X_0_vec_X_read_data_peek_empty_n,
    input wire                                           read_X_0_vec_X_read_data_peek_read,
    output wire [                                 256:0] read_X_0_vec_X_read_data_s_dout,
    output wire                                          read_X_0_vec_X_read_data_s_empty_n,
    input wire                                           read_X_0_vec_X_read_data_s_read,
    output wire [                                  63:0] read_X_0_vec_X_write_addr_offset,
    input wire  [                                  63:0] read_X_0_vec_X_write_addr_s_din,
    output wire                                          read_X_0_vec_X_write_addr_s_full_n,
    input wire                                           read_X_0_vec_X_write_addr_s_write,
    input wire  [                                 256:0] read_X_0_vec_X_write_data_din,
    output wire                                          read_X_0_vec_X_write_data_full_n,
    input wire                                           read_X_0_vec_X_write_data_write,
    output wire [                                   8:0] read_X_0_vec_X_write_resp_peek_dout,
    output wire                                          read_X_0_vec_X_write_resp_peek_empty_n,
    input wire                                           read_X_0_vec_X_write_resp_peek_read,
    output wire [                                   8:0] read_X_0_vec_X_write_resp_s_dout,
    output wire                                          read_X_0_vec_X_write_resp_s_empty_n,
    input wire                                           read_X_0_vec_X_write_resp_s_read,
    output wire [                                  31:0] read_Y_0_M,
    output wire [                                  31:0] read_Y_0_P_N,
    output wire [                                  63:0] read_Y_0_Y_read_addr_offset,
    input wire  [                                  63:0] read_Y_0_Y_read_addr_s_din,
    output wire                                          read_Y_0_Y_read_addr_s_full_n,
    input wire                                           read_Y_0_Y_read_addr_s_write,
    output wire [                                 256:0] read_Y_0_Y_read_data_peek_dout,
    output wire                                          read_Y_0_Y_read_data_peek_empty_n,
    input wire                                           read_Y_0_Y_read_data_peek_read,
    output wire [                                 256:0] read_Y_0_Y_read_data_s_dout,
    output wire                                          read_Y_0_Y_read_data_s_empty_n,
    input wire                                           read_Y_0_Y_read_data_s_read,
    output wire [                                  63:0] read_Y_0_Y_write_addr_offset,
    input wire  [                                  63:0] read_Y_0_Y_write_addr_s_din,
    output wire                                          read_Y_0_Y_write_addr_s_full_n,
    input wire                                           read_Y_0_Y_write_addr_s_write,
    input wire  [                                 256:0] read_Y_0_Y_write_data_din,
    output wire                                          read_Y_0_Y_write_data_full_n,
    input wire                                           read_Y_0_Y_write_data_write,
    output wire [                                   8:0] read_Y_0_Y_write_resp_peek_dout,
    output wire                                          read_Y_0_Y_write_resp_peek_empty_n,
    input wire                                           read_Y_0_Y_write_resp_peek_read,
    output wire [                                   8:0] read_Y_0_Y_write_resp_s_dout,
    output wire                                          read_Y_0_Y_write_resp_s_empty_n,
    input wire                                           read_Y_0_Y_write_resp_s_read,
    output wire                                          read_Y_0_ap_clk,
    input wire                                           read_Y_0_ap_done,
    input wire                                           read_Y_0_ap_idle,
    input wire                                           read_Y_0_ap_ready,
    output wire                                          read_Y_0_ap_rst_n,
    output wire                                          read_Y_0_ap_start,
    input wire  [                                 512:0] read_Y_0_fifo_Y_din,
    output wire                                          read_Y_0_fifo_Y_full_n,
    input wire                                           read_Y_0_fifo_Y_write,
    output wire [                                  31:0] read_edge_list_ptr_0_K,
    output wire [                                  31:0] read_edge_list_ptr_0_M,
    input wire  [                                  32:0] read_edge_list_ptr_0_PE_inst_din,
    output wire                                          read_edge_list_ptr_0_PE_inst_full_n,
    input wire                                           read_edge_list_ptr_0_PE_inst_write,
    output wire [                                  31:0] read_edge_list_ptr_0_P_N,
    output wire                                          read_edge_list_ptr_0_ap_clk,
    input wire                                           read_edge_list_ptr_0_ap_done,
    input wire                                           read_edge_list_ptr_0_ap_idle,
    input wire                                           read_edge_list_ptr_0_ap_ready,
    output wire                                          read_edge_list_ptr_0_ap_rst_n,
    output wire                                          read_edge_list_ptr_0_ap_start,
    output wire [                                  63:0] read_edge_list_ptr_0_edge_list_ptr_read_addr_offset,
    input wire  [                                  63:0] read_edge_list_ptr_0_edge_list_ptr_read_addr_s_din,
    output wire                                          read_edge_list_ptr_0_edge_list_ptr_read_addr_s_full_n,
    input wire                                           read_edge_list_ptr_0_edge_list_ptr_read_addr_s_write,
    output wire [                                  32:0] read_edge_list_ptr_0_edge_list_ptr_read_data_peek_dout,
    output wire                                          read_edge_list_ptr_0_edge_list_ptr_read_data_peek_empty_n,
    input wire                                           read_edge_list_ptr_0_edge_list_ptr_read_data_peek_read,
    output wire [                                  32:0] read_edge_list_ptr_0_edge_list_ptr_read_data_s_dout,
    output wire                                          read_edge_list_ptr_0_edge_list_ptr_read_data_s_empty_n,
    input wire                                           read_edge_list_ptr_0_edge_list_ptr_read_data_s_read,
    output wire [                                  63:0] read_edge_list_ptr_0_edge_list_ptr_write_addr_offset,
    input wire  [                                  63:0] read_edge_list_ptr_0_edge_list_ptr_write_addr_s_din,
    output wire                                          read_edge_list_ptr_0_edge_list_ptr_write_addr_s_full_n,
    input wire                                           read_edge_list_ptr_0_edge_list_ptr_write_addr_s_write,
    input wire  [                                  32:0] read_edge_list_ptr_0_edge_list_ptr_write_data_din,
    output wire                                          read_edge_list_ptr_0_edge_list_ptr_write_data_full_n,
    input wire                                           read_edge_list_ptr_0_edge_list_ptr_write_data_write,
    output wire [                                   8:0] read_edge_list_ptr_0_edge_list_ptr_write_resp_peek_dout,
    output wire                                          read_edge_list_ptr_0_edge_list_ptr_write_resp_peek_empty_n,
    input wire                                           read_edge_list_ptr_0_edge_list_ptr_write_resp_peek_read,
    output wire [                                   8:0] read_edge_list_ptr_0_edge_list_ptr_write_resp_s_dout,
    output wire                                          read_edge_list_ptr_0_edge_list_ptr_write_resp_s_empty_n,
    input wire                                           read_edge_list_ptr_0_edge_list_ptr_write_resp_s_read,
    output wire [                                  31:0] read_edge_list_ptr_0_num_ite,
    output wire [                                  31:0] write_Y_0_M,
    output wire [                                  31:0] write_Y_0_P_N,
    output wire [                                  63:0] write_Y_0_Y_out_read_addr_offset,
    input wire  [                                  63:0] write_Y_0_Y_out_read_addr_s_din,
    output wire                                          write_Y_0_Y_out_read_addr_s_full_n,
    input wire                                           write_Y_0_Y_out_read_addr_s_write,
    output wire [                                 256:0] write_Y_0_Y_out_read_data_peek_dout,
    output wire                                          write_Y_0_Y_out_read_data_peek_empty_n,
    input wire                                           write_Y_0_Y_out_read_data_peek_read,
    output wire [                                 256:0] write_Y_0_Y_out_read_data_s_dout,
    output wire                                          write_Y_0_Y_out_read_data_s_empty_n,
    input wire                                           write_Y_0_Y_out_read_data_s_read,
    output wire [                                  63:0] write_Y_0_Y_out_write_addr_offset,
    input wire  [                                  63:0] write_Y_0_Y_out_write_addr_s_din,
    output wire                                          write_Y_0_Y_out_write_addr_s_full_n,
    input wire                                           write_Y_0_Y_out_write_addr_s_write,
    input wire  [                                 256:0] write_Y_0_Y_out_write_data_din,
    output wire                                          write_Y_0_Y_out_write_data_full_n,
    input wire                                           write_Y_0_Y_out_write_data_write,
    output wire [                                   8:0] write_Y_0_Y_out_write_resp_peek_dout,
    output wire                                          write_Y_0_Y_out_write_resp_peek_empty_n,
    input wire                                           write_Y_0_Y_out_write_resp_peek_read,
    output wire [                                   8:0] write_Y_0_Y_out_write_resp_s_dout,
    output wire                                          write_Y_0_Y_out_write_resp_s_empty_n,
    input wire                                           write_Y_0_Y_out_write_resp_s_read,
    output wire                                          write_Y_0_ap_clk,
    input wire                                           write_Y_0_ap_done,
    input wire                                           write_Y_0_ap_idle,
    input wire                                           write_Y_0_ap_ready,
    output wire                                          write_Y_0_ap_rst_n,
    output wire                                          write_Y_0_ap_start,
    output wire [                                 512:0] write_Y_0_fifo_Y_peek_dout,
    output wire                                          write_Y_0_fifo_Y_peek_empty_n,
    input wire                                           write_Y_0_fifo_Y_peek_read,
    output wire [                                 512:0] write_Y_0_fifo_Y_s_dout,
    output wire                                          write_Y_0_fifo_Y_s_empty_n,
    input wire                                           write_Y_0_fifo_Y_s_read,
    output wire                                          edge_list_ch_0__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_0__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_0__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_0__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_0__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_0__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_0__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_0__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_0__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_0__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_0__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_0__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_0__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_0__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_0__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_0__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_0__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_0__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_0__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_0__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_0__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_0__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_0__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_0__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_0__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_0__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_0__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_0__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_0__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_0__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_0__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_0__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_0__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_0__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_0__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_0__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_0__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_0__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_0__m_axi_read_addr_din,
    input wire                                           edge_list_ch_0__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_0__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_0__m_axi_read_data_dout,
    input wire                                           edge_list_ch_0__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_0__m_axi_read_data_read,
    output wire                                          edge_list_ch_0__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_0__m_axi_write_addr_din,
    input wire                                           edge_list_ch_0__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_0__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_0__m_axi_write_data_din,
    input wire                                           edge_list_ch_0__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_0__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_0__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_0__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_0__m_axi_write_resp_read,
    output wire                                          edge_list_ch_1__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_1__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_1__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_1__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_1__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_1__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_1__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_1__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_1__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_1__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_1__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_1__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_1__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_1__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_1__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_1__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_1__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_1__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_1__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_1__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_1__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_1__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_1__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_1__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_1__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_1__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_1__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_1__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_1__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_1__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_1__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_1__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_1__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_1__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_1__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_1__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_1__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_1__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_1__m_axi_read_addr_din,
    input wire                                           edge_list_ch_1__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_1__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_1__m_axi_read_data_dout,
    input wire                                           edge_list_ch_1__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_1__m_axi_read_data_read,
    output wire                                          edge_list_ch_1__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_1__m_axi_write_addr_din,
    input wire                                           edge_list_ch_1__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_1__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_1__m_axi_write_data_din,
    input wire                                           edge_list_ch_1__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_1__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_1__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_1__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_1__m_axi_write_resp_read,
    output wire                                          edge_list_ch_2__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_2__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_2__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_2__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_2__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_2__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_2__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_2__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_2__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_2__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_2__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_2__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_2__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_2__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_2__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_2__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_2__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_2__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_2__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_2__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_2__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_2__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_2__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_2__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_2__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_2__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_2__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_2__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_2__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_2__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_2__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_2__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_2__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_2__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_2__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_2__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_2__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_2__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_2__m_axi_read_addr_din,
    input wire                                           edge_list_ch_2__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_2__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_2__m_axi_read_data_dout,
    input wire                                           edge_list_ch_2__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_2__m_axi_read_data_read,
    output wire                                          edge_list_ch_2__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_2__m_axi_write_addr_din,
    input wire                                           edge_list_ch_2__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_2__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_2__m_axi_write_data_din,
    input wire                                           edge_list_ch_2__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_2__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_2__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_2__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_2__m_axi_write_resp_read,
    output wire                                          edge_list_ch_3__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_3__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_3__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_3__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_3__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_3__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_3__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_3__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_3__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_3__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_3__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_3__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_3__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_3__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_3__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_3__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_3__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_3__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_3__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_3__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_3__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_3__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_3__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_3__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_3__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_3__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_3__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_3__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_3__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_3__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_3__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_3__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_3__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_3__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_3__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_3__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_3__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_3__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_3__m_axi_read_addr_din,
    input wire                                           edge_list_ch_3__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_3__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_3__m_axi_read_data_dout,
    input wire                                           edge_list_ch_3__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_3__m_axi_read_data_read,
    output wire                                          edge_list_ch_3__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_3__m_axi_write_addr_din,
    input wire                                           edge_list_ch_3__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_3__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_3__m_axi_write_data_din,
    input wire                                           edge_list_ch_3__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_3__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_3__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_3__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_3__m_axi_write_resp_read,
    output wire                                          edge_list_ch_4__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_4__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_4__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_4__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_4__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_4__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_4__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_4__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_4__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_4__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_4__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_4__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_4__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_4__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_4__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_4__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_4__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_4__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_4__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_4__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_4__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_4__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_4__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_4__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_4__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_4__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_4__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_4__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_4__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_4__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_4__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_4__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_4__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_4__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_4__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_4__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_4__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_4__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_4__m_axi_read_addr_din,
    input wire                                           edge_list_ch_4__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_4__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_4__m_axi_read_data_dout,
    input wire                                           edge_list_ch_4__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_4__m_axi_read_data_read,
    output wire                                          edge_list_ch_4__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_4__m_axi_write_addr_din,
    input wire                                           edge_list_ch_4__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_4__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_4__m_axi_write_data_din,
    input wire                                           edge_list_ch_4__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_4__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_4__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_4__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_4__m_axi_write_resp_read,
    output wire                                          edge_list_ch_5__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_5__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_5__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_5__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_5__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_5__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_5__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_5__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_5__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_5__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_5__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_5__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_5__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_5__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_5__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_5__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_5__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_5__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_5__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_5__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_5__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_5__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_5__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_5__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_5__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_5__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_5__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_5__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_5__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_5__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_5__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_5__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_5__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_5__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_5__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_5__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_5__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_5__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_5__m_axi_read_addr_din,
    input wire                                           edge_list_ch_5__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_5__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_5__m_axi_read_data_dout,
    input wire                                           edge_list_ch_5__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_5__m_axi_read_data_read,
    output wire                                          edge_list_ch_5__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_5__m_axi_write_addr_din,
    input wire                                           edge_list_ch_5__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_5__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_5__m_axi_write_data_din,
    input wire                                           edge_list_ch_5__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_5__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_5__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_5__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_5__m_axi_write_resp_read,
    output wire                                          edge_list_ch_6__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_6__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_6__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_6__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_6__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_6__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_6__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_6__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_6__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_6__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_6__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_6__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_6__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_6__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_6__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_6__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_6__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_6__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_6__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_6__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_6__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_6__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_6__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_6__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_6__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_6__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_6__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_6__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_6__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_6__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_6__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_6__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_6__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_6__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_6__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_6__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_6__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_6__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_6__m_axi_read_addr_din,
    input wire                                           edge_list_ch_6__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_6__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_6__m_axi_read_data_dout,
    input wire                                           edge_list_ch_6__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_6__m_axi_read_data_read,
    output wire                                          edge_list_ch_6__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_6__m_axi_write_addr_din,
    input wire                                           edge_list_ch_6__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_6__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_6__m_axi_write_data_din,
    input wire                                           edge_list_ch_6__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_6__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_6__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_6__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_6__m_axi_write_resp_read,
    output wire                                          edge_list_ch_7__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_7__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_7__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_7__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_7__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_7__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_7__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_7__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_7__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_7__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_7__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_7__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_7__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_7__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_7__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_7__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_7__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_7__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_7__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_7__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_7__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_7__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_7__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_7__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_7__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_7__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_7__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_7__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_7__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_7__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_7__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_7__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_7__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_7__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_7__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_7__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_7__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_7__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_7__m_axi_read_addr_din,
    input wire                                           edge_list_ch_7__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_7__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_7__m_axi_read_data_dout,
    input wire                                           edge_list_ch_7__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_7__m_axi_read_data_read,
    output wire                                          edge_list_ch_7__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_7__m_axi_write_addr_din,
    input wire                                           edge_list_ch_7__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_7__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_7__m_axi_write_data_din,
    input wire                                           edge_list_ch_7__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_7__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_7__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_7__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_7__m_axi_write_resp_read,
    output wire                                          edge_list_ch_8__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_8__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_8__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_8__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_8__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_8__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_8__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_8__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_8__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_8__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_8__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_8__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_8__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_8__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_8__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_8__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_8__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_8__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_8__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_8__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_8__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_8__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_8__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_8__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_8__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_8__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_8__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_8__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_8__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_8__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_8__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_8__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_8__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_8__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_8__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_8__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_8__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_8__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_8__m_axi_read_addr_din,
    input wire                                           edge_list_ch_8__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_8__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_8__m_axi_read_data_dout,
    input wire                                           edge_list_ch_8__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_8__m_axi_read_data_read,
    output wire                                          edge_list_ch_8__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_8__m_axi_write_addr_din,
    input wire                                           edge_list_ch_8__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_8__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_8__m_axi_write_data_din,
    input wire                                           edge_list_ch_8__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_8__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_8__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_8__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_8__m_axi_write_resp_read,
    output wire                                          edge_list_ch_9__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_9__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_9__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_9__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_9__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_9__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_9__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_9__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_9__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_9__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_9__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_9__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_9__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_9__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_9__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_9__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_9__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_9__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_9__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_9__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_9__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_9__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_9__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_9__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_9__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_9__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_9__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_9__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_9__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_9__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_9__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_9__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_9__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_9__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_9__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_9__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_9__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_9__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_9__m_axi_read_addr_din,
    input wire                                           edge_list_ch_9__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_9__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_9__m_axi_read_data_dout,
    input wire                                           edge_list_ch_9__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_9__m_axi_read_data_read,
    output wire                                          edge_list_ch_9__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_9__m_axi_write_addr_din,
    input wire                                           edge_list_ch_9__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_9__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_9__m_axi_write_data_din,
    input wire                                           edge_list_ch_9__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_9__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_9__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_9__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_9__m_axi_write_resp_read,
    output wire                                          edge_list_ch_10__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_10__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_10__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_10__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_10__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_10__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_10__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_10__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_10__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_10__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_10__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_10__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_10__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_10__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_10__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_10__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_10__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_10__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_10__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_10__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_10__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_10__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_10__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_10__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_10__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_10__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_10__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_10__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_10__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_10__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_10__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_10__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_10__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_10__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_10__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_10__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_10__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_10__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_10__m_axi_read_addr_din,
    input wire                                           edge_list_ch_10__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_10__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_10__m_axi_read_data_dout,
    input wire                                           edge_list_ch_10__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_10__m_axi_read_data_read,
    output wire                                          edge_list_ch_10__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_10__m_axi_write_addr_din,
    input wire                                           edge_list_ch_10__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_10__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_10__m_axi_write_data_din,
    input wire                                           edge_list_ch_10__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_10__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_10__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_10__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_10__m_axi_write_resp_read,
    output wire                                          edge_list_ch_11__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_11__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_11__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_11__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_11__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_11__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_11__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_11__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_11__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_11__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_11__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_11__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_11__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_11__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_11__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_11__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_11__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_11__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_11__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_11__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_11__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_11__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_11__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_11__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_11__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_11__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_11__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_11__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_11__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_11__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_11__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_11__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_11__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_11__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_11__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_11__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_11__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_11__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_11__m_axi_read_addr_din,
    input wire                                           edge_list_ch_11__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_11__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_11__m_axi_read_data_dout,
    input wire                                           edge_list_ch_11__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_11__m_axi_read_data_read,
    output wire                                          edge_list_ch_11__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_11__m_axi_write_addr_din,
    input wire                                           edge_list_ch_11__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_11__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_11__m_axi_write_data_din,
    input wire                                           edge_list_ch_11__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_11__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_11__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_11__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_11__m_axi_write_resp_read,
    output wire                                          edge_list_ch_12__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_12__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_12__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_12__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_12__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_12__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_12__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_12__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_12__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_12__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_12__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_12__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_12__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_12__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_12__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_12__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_12__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_12__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_12__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_12__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_12__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_12__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_12__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_12__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_12__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_12__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_12__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_12__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_12__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_12__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_12__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_12__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_12__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_12__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_12__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_12__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_12__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_12__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_12__m_axi_read_addr_din,
    input wire                                           edge_list_ch_12__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_12__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_12__m_axi_read_data_dout,
    input wire                                           edge_list_ch_12__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_12__m_axi_read_data_read,
    output wire                                          edge_list_ch_12__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_12__m_axi_write_addr_din,
    input wire                                           edge_list_ch_12__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_12__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_12__m_axi_write_data_din,
    input wire                                           edge_list_ch_12__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_12__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_12__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_12__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_12__m_axi_write_resp_read,
    output wire                                          edge_list_ch_13__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_13__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_13__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_13__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_13__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_13__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_13__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_13__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_13__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_13__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_13__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_13__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_13__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_13__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_13__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_13__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_13__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_13__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_13__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_13__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_13__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_13__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_13__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_13__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_13__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_13__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_13__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_13__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_13__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_13__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_13__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_13__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_13__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_13__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_13__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_13__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_13__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_13__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_13__m_axi_read_addr_din,
    input wire                                           edge_list_ch_13__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_13__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_13__m_axi_read_data_dout,
    input wire                                           edge_list_ch_13__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_13__m_axi_read_data_read,
    output wire                                          edge_list_ch_13__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_13__m_axi_write_addr_din,
    input wire                                           edge_list_ch_13__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_13__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_13__m_axi_write_data_din,
    input wire                                           edge_list_ch_13__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_13__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_13__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_13__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_13__m_axi_write_resp_read,
    output wire                                          edge_list_ch_14__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_14__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_14__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_14__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_14__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_14__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_14__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_14__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_14__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_14__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_14__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_14__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_14__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_14__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_14__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_14__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_14__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_14__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_14__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_14__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_14__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_14__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_14__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_14__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_14__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_14__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_14__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_14__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_14__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_14__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_14__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_14__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_14__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_14__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_14__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_14__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_14__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_14__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_14__m_axi_read_addr_din,
    input wire                                           edge_list_ch_14__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_14__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_14__m_axi_read_data_dout,
    input wire                                           edge_list_ch_14__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_14__m_axi_read_data_read,
    output wire                                          edge_list_ch_14__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_14__m_axi_write_addr_din,
    input wire                                           edge_list_ch_14__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_14__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_14__m_axi_write_data_din,
    input wire                                           edge_list_ch_14__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_14__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_14__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_14__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_14__m_axi_write_resp_read,
    output wire                                          edge_list_ch_15__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_15__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_15__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_15__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_15__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_15__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_15__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_15__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_15__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_15__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_15__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_15__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_15__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_15__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_15__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_15__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_15__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_15__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_15__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_15__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_15__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_15__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_15__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_15__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_15__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_15__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_15__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_15__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_15__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_15__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_15__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_15__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_15__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_15__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_15__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_15__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_15__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_15__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_15__m_axi_read_addr_din,
    input wire                                           edge_list_ch_15__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_15__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_15__m_axi_read_data_dout,
    input wire                                           edge_list_ch_15__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_15__m_axi_read_data_read,
    output wire                                          edge_list_ch_15__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_15__m_axi_write_addr_din,
    input wire                                           edge_list_ch_15__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_15__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_15__m_axi_write_data_din,
    input wire                                           edge_list_ch_15__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_15__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_15__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_15__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_15__m_axi_write_resp_read,
    output wire                                          edge_list_ch_16__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_16__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_16__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_16__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_16__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_16__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_16__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_16__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_16__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_16__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_16__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_16__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_16__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_16__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_16__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_16__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_16__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_16__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_16__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_16__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_16__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_16__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_16__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_16__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_16__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_16__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_16__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_16__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_16__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_16__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_16__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_16__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_16__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_16__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_16__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_16__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_16__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_16__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_16__m_axi_read_addr_din,
    input wire                                           edge_list_ch_16__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_16__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_16__m_axi_read_data_dout,
    input wire                                           edge_list_ch_16__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_16__m_axi_read_data_read,
    output wire                                          edge_list_ch_16__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_16__m_axi_write_addr_din,
    input wire                                           edge_list_ch_16__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_16__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_16__m_axi_write_data_din,
    input wire                                           edge_list_ch_16__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_16__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_16__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_16__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_16__m_axi_write_resp_read,
    output wire                                          edge_list_ch_17__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_17__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_17__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_17__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_17__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_17__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_17__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_17__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_17__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_17__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_17__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_17__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_17__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_17__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_17__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_17__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_17__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_17__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_17__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_17__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_17__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_17__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_17__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_17__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_17__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_17__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_17__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_17__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_17__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_17__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_17__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_17__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_17__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_17__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_17__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_17__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_17__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_17__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_17__m_axi_read_addr_din,
    input wire                                           edge_list_ch_17__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_17__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_17__m_axi_read_data_dout,
    input wire                                           edge_list_ch_17__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_17__m_axi_read_data_read,
    output wire                                          edge_list_ch_17__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_17__m_axi_write_addr_din,
    input wire                                           edge_list_ch_17__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_17__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_17__m_axi_write_data_din,
    input wire                                           edge_list_ch_17__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_17__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_17__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_17__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_17__m_axi_write_resp_read,
    output wire                                          edge_list_ch_18__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_18__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_18__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_18__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_18__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_18__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_18__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_18__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_18__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_18__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_18__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_18__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_18__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_18__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_18__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_18__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_18__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_18__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_18__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_18__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_18__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_18__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_18__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_18__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_18__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_18__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_18__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_18__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_18__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_18__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_18__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_18__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_18__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_18__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_18__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_18__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_18__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_18__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_18__m_axi_read_addr_din,
    input wire                                           edge_list_ch_18__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_18__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_18__m_axi_read_data_dout,
    input wire                                           edge_list_ch_18__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_18__m_axi_read_data_read,
    output wire                                          edge_list_ch_18__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_18__m_axi_write_addr_din,
    input wire                                           edge_list_ch_18__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_18__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_18__m_axi_write_data_din,
    input wire                                           edge_list_ch_18__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_18__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_18__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_18__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_18__m_axi_write_resp_read,
    output wire                                          edge_list_ch_19__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_19__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_19__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_19__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_19__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_19__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_19__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_19__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_19__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_19__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_19__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_19__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_19__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_19__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_19__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_19__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_19__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_19__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_19__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_19__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_19__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_19__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_19__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_19__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_19__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_19__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_19__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_19__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_19__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_19__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_19__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_19__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_19__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_19__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_19__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_19__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_19__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_19__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_19__m_axi_read_addr_din,
    input wire                                           edge_list_ch_19__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_19__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_19__m_axi_read_data_dout,
    input wire                                           edge_list_ch_19__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_19__m_axi_read_data_read,
    output wire                                          edge_list_ch_19__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_19__m_axi_write_addr_din,
    input wire                                           edge_list_ch_19__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_19__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_19__m_axi_write_data_din,
    input wire                                           edge_list_ch_19__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_19__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_19__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_19__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_19__m_axi_write_resp_read,
    output wire                                          edge_list_ch_20__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_20__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_20__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_20__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_20__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_20__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_20__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_20__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_20__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_20__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_20__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_20__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_20__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_20__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_20__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_20__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_20__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_20__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_20__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_20__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_20__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_20__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_20__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_20__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_20__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_20__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_20__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_20__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_20__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_20__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_20__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_20__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_20__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_20__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_20__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_20__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_20__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_20__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_20__m_axi_read_addr_din,
    input wire                                           edge_list_ch_20__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_20__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_20__m_axi_read_data_dout,
    input wire                                           edge_list_ch_20__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_20__m_axi_read_data_read,
    output wire                                          edge_list_ch_20__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_20__m_axi_write_addr_din,
    input wire                                           edge_list_ch_20__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_20__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_20__m_axi_write_data_din,
    input wire                                           edge_list_ch_20__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_20__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_20__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_20__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_20__m_axi_write_resp_read,
    output wire                                          edge_list_ch_21__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_21__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_21__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_21__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_21__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_21__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_21__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_21__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_21__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_21__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_21__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_21__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_21__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_21__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_21__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_21__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_21__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_21__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_21__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_21__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_21__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_21__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_21__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_21__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_21__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_21__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_21__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_21__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_21__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_21__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_21__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_21__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_21__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_21__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_21__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_21__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_21__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_21__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_21__m_axi_read_addr_din,
    input wire                                           edge_list_ch_21__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_21__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_21__m_axi_read_data_dout,
    input wire                                           edge_list_ch_21__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_21__m_axi_read_data_read,
    output wire                                          edge_list_ch_21__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_21__m_axi_write_addr_din,
    input wire                                           edge_list_ch_21__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_21__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_21__m_axi_write_data_din,
    input wire                                           edge_list_ch_21__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_21__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_21__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_21__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_21__m_axi_write_resp_read,
    output wire                                          edge_list_ch_22__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_22__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_22__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_22__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_22__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_22__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_22__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_22__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_22__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_22__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_22__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_22__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_22__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_22__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_22__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_22__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_22__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_22__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_22__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_22__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_22__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_22__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_22__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_22__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_22__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_22__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_22__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_22__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_22__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_22__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_22__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_22__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_22__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_22__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_22__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_22__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_22__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_22__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_22__m_axi_read_addr_din,
    input wire                                           edge_list_ch_22__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_22__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_22__m_axi_read_data_dout,
    input wire                                           edge_list_ch_22__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_22__m_axi_read_data_read,
    output wire                                          edge_list_ch_22__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_22__m_axi_write_addr_din,
    input wire                                           edge_list_ch_22__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_22__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_22__m_axi_write_data_din,
    input wire                                           edge_list_ch_22__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_22__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_22__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_22__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_22__m_axi_write_resp_read,
    output wire                                          edge_list_ch_23__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_23__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_23__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_23__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_23__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_23__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_23__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_23__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_23__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_23__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_23__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_23__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_23__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_23__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_23__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_23__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_23__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_23__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_23__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_23__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_23__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_23__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_23__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_23__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_23__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_23__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_23__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_23__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_23__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_23__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_23__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_23__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_23__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_23__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_23__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_23__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_23__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_23__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_23__m_axi_read_addr_din,
    input wire                                           edge_list_ch_23__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_23__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_23__m_axi_read_data_dout,
    input wire                                           edge_list_ch_23__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_23__m_axi_read_data_read,
    output wire                                          edge_list_ch_23__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_23__m_axi_write_addr_din,
    input wire                                           edge_list_ch_23__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_23__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_23__m_axi_write_data_din,
    input wire                                           edge_list_ch_23__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_23__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_23__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_23__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_23__m_axi_write_resp_read,
    output wire                                          edge_list_ch_24__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_24__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_24__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_24__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_24__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_24__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_24__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_24__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_24__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_24__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_24__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_24__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_24__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_24__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_24__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_24__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_24__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_24__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_24__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_24__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_24__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_24__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_24__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_24__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_24__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_24__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_24__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_24__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_24__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_24__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_24__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_24__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_24__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_24__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_24__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_24__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_24__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_24__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_24__m_axi_read_addr_din,
    input wire                                           edge_list_ch_24__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_24__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_24__m_axi_read_data_dout,
    input wire                                           edge_list_ch_24__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_24__m_axi_read_data_read,
    output wire                                          edge_list_ch_24__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_24__m_axi_write_addr_din,
    input wire                                           edge_list_ch_24__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_24__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_24__m_axi_write_data_din,
    input wire                                           edge_list_ch_24__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_24__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_24__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_24__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_24__m_axi_write_resp_read,
    output wire                                          edge_list_ch_25__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_25__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_25__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_25__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_25__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_25__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_25__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_25__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_25__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_25__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_25__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_25__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_25__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_25__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_25__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_25__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_25__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_25__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_25__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_25__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_25__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_25__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_25__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_25__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_25__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_25__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_25__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_25__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_25__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_25__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_25__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_25__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_25__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_25__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_25__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_25__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_25__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_25__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_25__m_axi_read_addr_din,
    input wire                                           edge_list_ch_25__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_25__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_25__m_axi_read_data_dout,
    input wire                                           edge_list_ch_25__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_25__m_axi_read_data_read,
    output wire                                          edge_list_ch_25__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_25__m_axi_write_addr_din,
    input wire                                           edge_list_ch_25__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_25__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_25__m_axi_write_data_din,
    input wire                                           edge_list_ch_25__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_25__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_25__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_25__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_25__m_axi_write_resp_read,
    output wire                                          edge_list_ch_26__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_26__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_26__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_26__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_26__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_26__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_26__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_26__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_26__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_26__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_26__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_26__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_26__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_26__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_26__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_26__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_26__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_26__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_26__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_26__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_26__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_26__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_26__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_26__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_26__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_26__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_26__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_26__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_26__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_26__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_26__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_26__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_26__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_26__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_26__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_26__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_26__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_26__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_26__m_axi_read_addr_din,
    input wire                                           edge_list_ch_26__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_26__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_26__m_axi_read_data_dout,
    input wire                                           edge_list_ch_26__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_26__m_axi_read_data_read,
    output wire                                          edge_list_ch_26__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_26__m_axi_write_addr_din,
    input wire                                           edge_list_ch_26__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_26__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_26__m_axi_write_data_din,
    input wire                                           edge_list_ch_26__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_26__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_26__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_26__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_26__m_axi_write_resp_read,
    output wire                                          edge_list_ch_27__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_27__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_27__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_27__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_27__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_27__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_27__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_27__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_27__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_27__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_27__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_27__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_27__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_27__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_27__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_27__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_27__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_27__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_27__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_27__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_27__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_27__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_27__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_27__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_27__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_27__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_27__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_27__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_27__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_27__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_27__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_27__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_27__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_27__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_27__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_27__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_27__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_27__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_27__m_axi_read_addr_din,
    input wire                                           edge_list_ch_27__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_27__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_27__m_axi_read_data_dout,
    input wire                                           edge_list_ch_27__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_27__m_axi_read_data_read,
    output wire                                          edge_list_ch_27__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_27__m_axi_write_addr_din,
    input wire                                           edge_list_ch_27__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_27__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_27__m_axi_write_data_din,
    input wire                                           edge_list_ch_27__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_27__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_27__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_27__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_27__m_axi_write_resp_read,
    output wire                                          edge_list_ch_28__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_28__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_28__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_28__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_28__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_28__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_28__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_28__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_28__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_28__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_28__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_28__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_28__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_28__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_28__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_28__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_28__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_28__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_28__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_28__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_28__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_28__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_28__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_28__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_28__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_28__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_28__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_28__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_28__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_28__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_28__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_28__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_28__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_28__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_28__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_28__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_28__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_28__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_28__m_axi_read_addr_din,
    input wire                                           edge_list_ch_28__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_28__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_28__m_axi_read_data_dout,
    input wire                                           edge_list_ch_28__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_28__m_axi_read_data_read,
    output wire                                          edge_list_ch_28__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_28__m_axi_write_addr_din,
    input wire                                           edge_list_ch_28__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_28__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_28__m_axi_write_data_din,
    input wire                                           edge_list_ch_28__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_28__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_28__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_28__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_28__m_axi_write_resp_read,
    output wire                                          edge_list_ch_29__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_29__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_29__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_29__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_29__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_29__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_29__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_29__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_29__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_29__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_29__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_29__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_29__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_29__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_29__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_29__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_29__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_29__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_29__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_29__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_29__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_29__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_29__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_29__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_29__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_29__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_29__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_29__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_29__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_29__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_29__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_29__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_29__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_29__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_29__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_29__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_29__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_29__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_29__m_axi_read_addr_din,
    input wire                                           edge_list_ch_29__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_29__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_29__m_axi_read_data_dout,
    input wire                                           edge_list_ch_29__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_29__m_axi_read_data_read,
    output wire                                          edge_list_ch_29__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_29__m_axi_write_addr_din,
    input wire                                           edge_list_ch_29__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_29__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_29__m_axi_write_data_din,
    input wire                                           edge_list_ch_29__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_29__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_29__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_29__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_29__m_axi_write_resp_read,
    output wire                                          edge_list_ch_30__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_30__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_30__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_30__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_30__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_30__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_30__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_30__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_30__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_30__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_30__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_30__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_30__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_30__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_30__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_30__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_30__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_30__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_30__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_30__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_30__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_30__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_30__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_30__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_30__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_30__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_30__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_30__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_30__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_30__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_30__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_30__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_30__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_30__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_30__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_30__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_30__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_30__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_30__m_axi_read_addr_din,
    input wire                                           edge_list_ch_30__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_30__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_30__m_axi_read_data_dout,
    input wire                                           edge_list_ch_30__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_30__m_axi_read_data_read,
    output wire                                          edge_list_ch_30__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_30__m_axi_write_addr_din,
    input wire                                           edge_list_ch_30__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_30__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_30__m_axi_write_data_din,
    input wire                                           edge_list_ch_30__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_30__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_30__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_30__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_30__m_axi_write_resp_read,
    output wire                                          edge_list_ch_31__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_31__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_31__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_31__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_31__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_31__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_31__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_31__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_31__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_31__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_31__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_31__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_31__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_31__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_31__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_31__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_31__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_31__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_31__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_31__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_31__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_31__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_31__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_31__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_31__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_31__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_31__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_31__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_31__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_31__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_31__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_31__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_31__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_31__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_31__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_31__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_31__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_31__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_31__m_axi_read_addr_din,
    input wire                                           edge_list_ch_31__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_31__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_31__m_axi_read_data_dout,
    input wire                                           edge_list_ch_31__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_31__m_axi_read_data_read,
    output wire                                          edge_list_ch_31__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_31__m_axi_write_addr_din,
    input wire                                           edge_list_ch_31__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_31__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_31__m_axi_write_data_din,
    input wire                                           edge_list_ch_31__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_31__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_31__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_31__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_31__m_axi_write_resp_read,
    output wire                                          edge_list_ch_32__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_32__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_32__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_32__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_32__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_32__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_32__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_32__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_32__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_32__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_32__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_32__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_32__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_32__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_32__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_32__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_32__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_32__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_32__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_32__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_32__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_32__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_32__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_32__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_32__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_32__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_32__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_32__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_32__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_32__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_32__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_32__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_32__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_32__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_32__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_32__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_32__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_32__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_32__m_axi_read_addr_din,
    input wire                                           edge_list_ch_32__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_32__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_32__m_axi_read_data_dout,
    input wire                                           edge_list_ch_32__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_32__m_axi_read_data_read,
    output wire                                          edge_list_ch_32__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_32__m_axi_write_addr_din,
    input wire                                           edge_list_ch_32__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_32__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_32__m_axi_write_data_din,
    input wire                                           edge_list_ch_32__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_32__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_32__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_32__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_32__m_axi_write_resp_read,
    output wire                                          edge_list_ch_33__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_33__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_33__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_33__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_33__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_33__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_33__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_33__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_33__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_33__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_33__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_33__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_33__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_33__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_33__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_33__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_33__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_33__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_33__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_33__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_33__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_33__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_33__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_33__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_33__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_33__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_33__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_33__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_33__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_33__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_33__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_33__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_33__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_33__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_33__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_33__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_33__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_33__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_33__m_axi_read_addr_din,
    input wire                                           edge_list_ch_33__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_33__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_33__m_axi_read_data_dout,
    input wire                                           edge_list_ch_33__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_33__m_axi_read_data_read,
    output wire                                          edge_list_ch_33__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_33__m_axi_write_addr_din,
    input wire                                           edge_list_ch_33__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_33__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_33__m_axi_write_data_din,
    input wire                                           edge_list_ch_33__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_33__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_33__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_33__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_33__m_axi_write_resp_read,
    output wire                                          edge_list_ch_34__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_34__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_34__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_34__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_34__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_34__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_34__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_34__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_34__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_34__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_34__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_34__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_34__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_34__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_34__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_34__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_34__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_34__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_34__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_34__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_34__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_34__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_34__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_34__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_34__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_34__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_34__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_34__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_34__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_34__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_34__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_34__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_34__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_34__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_34__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_34__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_34__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_34__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_34__m_axi_read_addr_din,
    input wire                                           edge_list_ch_34__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_34__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_34__m_axi_read_data_dout,
    input wire                                           edge_list_ch_34__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_34__m_axi_read_data_read,
    output wire                                          edge_list_ch_34__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_34__m_axi_write_addr_din,
    input wire                                           edge_list_ch_34__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_34__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_34__m_axi_write_data_din,
    input wire                                           edge_list_ch_34__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_34__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_34__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_34__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_34__m_axi_write_resp_read,
    output wire                                          edge_list_ch_35__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_35__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_35__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_35__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_35__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_35__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_35__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_35__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_35__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_35__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_35__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_35__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_35__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_35__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_35__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_35__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_35__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_35__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_35__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_35__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_35__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_35__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_35__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_35__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_35__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_35__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_35__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_35__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_35__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_35__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_35__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_35__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_35__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_35__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_35__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_35__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_35__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_35__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_35__m_axi_read_addr_din,
    input wire                                           edge_list_ch_35__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_35__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_35__m_axi_read_data_dout,
    input wire                                           edge_list_ch_35__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_35__m_axi_read_data_read,
    output wire                                          edge_list_ch_35__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_35__m_axi_write_addr_din,
    input wire                                           edge_list_ch_35__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_35__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_35__m_axi_write_data_din,
    input wire                                           edge_list_ch_35__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_35__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_35__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_35__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_35__m_axi_write_resp_read,
    output wire                                          edge_list_ch_36__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_36__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_36__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_36__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_36__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_36__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_36__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_36__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_36__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_36__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_36__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_36__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_36__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_36__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_36__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_36__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_36__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_36__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_36__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_36__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_36__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_36__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_36__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_36__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_36__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_36__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_36__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_36__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_36__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_36__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_36__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_36__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_36__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_36__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_36__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_36__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_36__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_36__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_36__m_axi_read_addr_din,
    input wire                                           edge_list_ch_36__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_36__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_36__m_axi_read_data_dout,
    input wire                                           edge_list_ch_36__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_36__m_axi_read_data_read,
    output wire                                          edge_list_ch_36__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_36__m_axi_write_addr_din,
    input wire                                           edge_list_ch_36__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_36__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_36__m_axi_write_data_din,
    input wire                                           edge_list_ch_36__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_36__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_36__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_36__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_36__m_axi_write_resp_read,
    output wire                                          edge_list_ch_37__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_37__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_37__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_37__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_37__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_37__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_37__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_37__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_37__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_37__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_37__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_37__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_37__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_37__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_37__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_37__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_37__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_37__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_37__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_37__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_37__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_37__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_37__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_37__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_37__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_37__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_37__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_37__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_37__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_37__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_37__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_37__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_37__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_37__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_37__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_37__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_37__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_37__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_37__m_axi_read_addr_din,
    input wire                                           edge_list_ch_37__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_37__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_37__m_axi_read_data_dout,
    input wire                                           edge_list_ch_37__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_37__m_axi_read_data_read,
    output wire                                          edge_list_ch_37__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_37__m_axi_write_addr_din,
    input wire                                           edge_list_ch_37__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_37__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_37__m_axi_write_data_din,
    input wire                                           edge_list_ch_37__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_37__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_37__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_37__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_37__m_axi_write_resp_read,
    output wire                                          edge_list_ch_38__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_38__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_38__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_38__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_38__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_38__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_38__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_38__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_38__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_38__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_38__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_38__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_38__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_38__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_38__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_38__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_38__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_38__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_38__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_38__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_38__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_38__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_38__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_38__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_38__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_38__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_38__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_38__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_38__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_38__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_38__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_38__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_38__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_38__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_38__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_38__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_38__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_38__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_38__m_axi_read_addr_din,
    input wire                                           edge_list_ch_38__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_38__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_38__m_axi_read_data_dout,
    input wire                                           edge_list_ch_38__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_38__m_axi_read_data_read,
    output wire                                          edge_list_ch_38__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_38__m_axi_write_addr_din,
    input wire                                           edge_list_ch_38__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_38__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_38__m_axi_write_data_din,
    input wire                                           edge_list_ch_38__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_38__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_38__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_38__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_38__m_axi_write_resp_read,
    output wire                                          edge_list_ch_39__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_39__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_39__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_39__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_39__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_39__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_39__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_39__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_39__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_39__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_39__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_39__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_39__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_39__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_39__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_39__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_39__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_39__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_39__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_39__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_39__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_39__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_39__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_39__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_39__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_39__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_39__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_39__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_39__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_39__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_39__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_39__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_39__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_39__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_39__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_39__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_39__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_39__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_39__m_axi_read_addr_din,
    input wire                                           edge_list_ch_39__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_39__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_39__m_axi_read_data_dout,
    input wire                                           edge_list_ch_39__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_39__m_axi_read_data_read,
    output wire                                          edge_list_ch_39__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_39__m_axi_write_addr_din,
    input wire                                           edge_list_ch_39__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_39__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_39__m_axi_write_data_din,
    input wire                                           edge_list_ch_39__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_39__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_39__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_39__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_39__m_axi_write_resp_read,
    output wire                                          edge_list_ch_40__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_40__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_40__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_40__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_40__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_40__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_40__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_40__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_40__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_40__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_40__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_40__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_40__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_40__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_40__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_40__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_40__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_40__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_40__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_40__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_40__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_40__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_40__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_40__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_40__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_40__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_40__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_40__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_40__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_40__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_40__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_40__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_40__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_40__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_40__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_40__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_40__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_40__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_40__m_axi_read_addr_din,
    input wire                                           edge_list_ch_40__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_40__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_40__m_axi_read_data_dout,
    input wire                                           edge_list_ch_40__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_40__m_axi_read_data_read,
    output wire                                          edge_list_ch_40__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_40__m_axi_write_addr_din,
    input wire                                           edge_list_ch_40__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_40__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_40__m_axi_write_data_din,
    input wire                                           edge_list_ch_40__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_40__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_40__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_40__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_40__m_axi_write_resp_read,
    output wire                                          edge_list_ch_41__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_41__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_41__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_41__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_41__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_41__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_41__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_41__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_41__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_41__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_41__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_41__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_41__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_41__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_41__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_41__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_41__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_41__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_41__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_41__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_41__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_41__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_41__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_41__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_41__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_41__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_41__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_41__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_41__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_41__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_41__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_41__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_41__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_41__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_41__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_41__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_41__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_41__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_41__m_axi_read_addr_din,
    input wire                                           edge_list_ch_41__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_41__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_41__m_axi_read_data_dout,
    input wire                                           edge_list_ch_41__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_41__m_axi_read_data_read,
    output wire                                          edge_list_ch_41__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_41__m_axi_write_addr_din,
    input wire                                           edge_list_ch_41__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_41__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_41__m_axi_write_data_din,
    input wire                                           edge_list_ch_41__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_41__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_41__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_41__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_41__m_axi_write_resp_read,
    output wire                                          edge_list_ch_42__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_42__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_42__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_42__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_42__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_42__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_42__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_42__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_42__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_42__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_42__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_42__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_42__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_42__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_42__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_42__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_42__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_42__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_42__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_42__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_42__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_42__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_42__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_42__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_42__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_42__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_42__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_42__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_42__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_42__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_42__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_42__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_42__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_42__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_42__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_42__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_42__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_42__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_42__m_axi_read_addr_din,
    input wire                                           edge_list_ch_42__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_42__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_42__m_axi_read_data_dout,
    input wire                                           edge_list_ch_42__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_42__m_axi_read_data_read,
    output wire                                          edge_list_ch_42__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_42__m_axi_write_addr_din,
    input wire                                           edge_list_ch_42__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_42__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_42__m_axi_write_data_din,
    input wire                                           edge_list_ch_42__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_42__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_42__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_42__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_42__m_axi_write_resp_read,
    output wire                                          edge_list_ch_43__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_43__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_43__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_43__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_43__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_43__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_43__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_43__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_43__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_43__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_43__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_43__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_43__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_43__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_43__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_43__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_43__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_43__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_43__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_43__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_43__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_43__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_43__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_43__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_43__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_43__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_43__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_43__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_43__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_43__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_43__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_43__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_43__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_43__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_43__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_43__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_43__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_43__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_43__m_axi_read_addr_din,
    input wire                                           edge_list_ch_43__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_43__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_43__m_axi_read_data_dout,
    input wire                                           edge_list_ch_43__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_43__m_axi_read_data_read,
    output wire                                          edge_list_ch_43__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_43__m_axi_write_addr_din,
    input wire                                           edge_list_ch_43__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_43__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_43__m_axi_write_data_din,
    input wire                                           edge_list_ch_43__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_43__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_43__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_43__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_43__m_axi_write_resp_read,
    output wire                                          edge_list_ch_44__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_44__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_44__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_44__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_44__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_44__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_44__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_44__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_44__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_44__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_44__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_44__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_44__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_44__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_44__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_44__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_44__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_44__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_44__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_44__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_44__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_44__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_44__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_44__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_44__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_44__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_44__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_44__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_44__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_44__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_44__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_44__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_44__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_44__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_44__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_44__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_44__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_44__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_44__m_axi_read_addr_din,
    input wire                                           edge_list_ch_44__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_44__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_44__m_axi_read_data_dout,
    input wire                                           edge_list_ch_44__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_44__m_axi_read_data_read,
    output wire                                          edge_list_ch_44__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_44__m_axi_write_addr_din,
    input wire                                           edge_list_ch_44__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_44__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_44__m_axi_write_data_din,
    input wire                                           edge_list_ch_44__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_44__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_44__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_44__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_44__m_axi_write_resp_read,
    output wire                                          edge_list_ch_45__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_45__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_45__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_45__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_45__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_45__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_45__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_45__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_45__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_45__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_45__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_45__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_45__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_45__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_45__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_45__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_45__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_45__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_45__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_45__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_45__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_45__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_45__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_45__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_45__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_45__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_45__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_45__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_45__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_45__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_45__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_45__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_45__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_45__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_45__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_45__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_45__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_45__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_45__m_axi_read_addr_din,
    input wire                                           edge_list_ch_45__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_45__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_45__m_axi_read_data_dout,
    input wire                                           edge_list_ch_45__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_45__m_axi_read_data_read,
    output wire                                          edge_list_ch_45__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_45__m_axi_write_addr_din,
    input wire                                           edge_list_ch_45__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_45__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_45__m_axi_write_data_din,
    input wire                                           edge_list_ch_45__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_45__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_45__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_45__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_45__m_axi_write_resp_read,
    output wire                                          edge_list_ch_46__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_46__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_46__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_46__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_46__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_46__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_46__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_46__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_46__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_46__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_46__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_46__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_46__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_46__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_46__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_46__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_46__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_46__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_46__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_46__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_46__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_46__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_46__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_46__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_46__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_46__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_46__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_46__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_46__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_46__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_46__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_46__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_46__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_46__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_46__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_46__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_46__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_46__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_46__m_axi_read_addr_din,
    input wire                                           edge_list_ch_46__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_46__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_46__m_axi_read_data_dout,
    input wire                                           edge_list_ch_46__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_46__m_axi_read_data_read,
    output wire                                          edge_list_ch_46__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_46__m_axi_write_addr_din,
    input wire                                           edge_list_ch_46__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_46__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_46__m_axi_write_data_din,
    input wire                                           edge_list_ch_46__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_46__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_46__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_46__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_46__m_axi_write_resp_read,
    output wire                                          edge_list_ch_47__m_axi_clk,
    input wire  [                                  63:0] edge_list_ch_47__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ch_47__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ch_47__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ch_47__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ch_47__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ch_47__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ch_47__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ch_47__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ch_47__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ch_47__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ch_47__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ch_47__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ch_47__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ch_47__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ch_47__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ch_47__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ch_47__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ch_47__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ch_47__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ch_47__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ch_47__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ch_47__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ch_47__m_axi_m_axi_BID,
    input wire                                           edge_list_ch_47__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ch_47__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ch_47__m_axi_m_axi_BVALID,
    output wire [                                 255:0] edge_list_ch_47__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ch_47__m_axi_m_axi_RID,
    output wire                                          edge_list_ch_47__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ch_47__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ch_47__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ch_47__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] edge_list_ch_47__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ch_47__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ch_47__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] edge_list_ch_47__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ch_47__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ch_47__m_axi_read_addr_din,
    input wire                                           edge_list_ch_47__m_axi_read_addr_full_n,
    output wire                                          edge_list_ch_47__m_axi_read_addr_write,
    input wire  [                                 255:0] edge_list_ch_47__m_axi_read_data_dout,
    input wire                                           edge_list_ch_47__m_axi_read_data_empty_n,
    output wire                                          edge_list_ch_47__m_axi_read_data_read,
    output wire                                          edge_list_ch_47__m_axi_rst,
    output wire [                                  63:0] edge_list_ch_47__m_axi_write_addr_din,
    input wire                                           edge_list_ch_47__m_axi_write_addr_full_n,
    output wire                                          edge_list_ch_47__m_axi_write_addr_write,
    output wire [                                 255:0] edge_list_ch_47__m_axi_write_data_din,
    input wire                                           edge_list_ch_47__m_axi_write_data_full_n,
    output wire                                          edge_list_ch_47__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ch_47__m_axi_write_resp_dout,
    input wire                                           edge_list_ch_47__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ch_47__m_axi_write_resp_read,
    output wire                                          vec_X__m_axi_clk,
    input wire  [                                  63:0] vec_X__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] vec_X__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] vec_X__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] vec_X__m_axi_m_axi_ARID,
    input wire  [                                   7:0] vec_X__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] vec_X__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] vec_X__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] vec_X__m_axi_m_axi_ARQOS,
    output wire                                          vec_X__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] vec_X__m_axi_m_axi_ARSIZE,
    input wire                                           vec_X__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] vec_X__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] vec_X__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] vec_X__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] vec_X__m_axi_m_axi_AWID,
    input wire  [                                   7:0] vec_X__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] vec_X__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] vec_X__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] vec_X__m_axi_m_axi_AWQOS,
    output wire                                          vec_X__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] vec_X__m_axi_m_axi_AWSIZE,
    input wire                                           vec_X__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] vec_X__m_axi_m_axi_BID,
    input wire                                           vec_X__m_axi_m_axi_BREADY,
    output wire [                                   1:0] vec_X__m_axi_m_axi_BRESP,
    output wire                                          vec_X__m_axi_m_axi_BVALID,
    output wire [                                 255:0] vec_X__m_axi_m_axi_RDATA,
    output wire [                                   0:0] vec_X__m_axi_m_axi_RID,
    output wire                                          vec_X__m_axi_m_axi_RLAST,
    input wire                                           vec_X__m_axi_m_axi_RREADY,
    output wire [                                   1:0] vec_X__m_axi_m_axi_RRESP,
    output wire                                          vec_X__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] vec_X__m_axi_m_axi_WDATA,
    input wire                                           vec_X__m_axi_m_axi_WLAST,
    output wire                                          vec_X__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] vec_X__m_axi_m_axi_WSTRB,
    input wire                                           vec_X__m_axi_m_axi_WVALID,
    output wire [                                  63:0] vec_X__m_axi_read_addr_din,
    input wire                                           vec_X__m_axi_read_addr_full_n,
    output wire                                          vec_X__m_axi_read_addr_write,
    input wire  [                                 255:0] vec_X__m_axi_read_data_dout,
    input wire                                           vec_X__m_axi_read_data_empty_n,
    output wire                                          vec_X__m_axi_read_data_read,
    output wire                                          vec_X__m_axi_rst,
    output wire [                                  63:0] vec_X__m_axi_write_addr_din,
    input wire                                           vec_X__m_axi_write_addr_full_n,
    output wire                                          vec_X__m_axi_write_addr_write,
    output wire [                                 255:0] vec_X__m_axi_write_data_din,
    input wire                                           vec_X__m_axi_write_data_full_n,
    output wire                                          vec_X__m_axi_write_data_write,
    input wire  [                                   7:0] vec_X__m_axi_write_resp_dout,
    input wire                                           vec_X__m_axi_write_resp_empty_n,
    output wire                                          vec_X__m_axi_write_resp_read,
    output wire                                          vec_Y__m_axi_clk,
    input wire  [                                  63:0] vec_Y__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] vec_Y__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] vec_Y__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] vec_Y__m_axi_m_axi_ARID,
    input wire  [                                   7:0] vec_Y__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] vec_Y__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] vec_Y__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] vec_Y__m_axi_m_axi_ARQOS,
    output wire                                          vec_Y__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] vec_Y__m_axi_m_axi_ARSIZE,
    input wire                                           vec_Y__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] vec_Y__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] vec_Y__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] vec_Y__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] vec_Y__m_axi_m_axi_AWID,
    input wire  [                                   7:0] vec_Y__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] vec_Y__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] vec_Y__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] vec_Y__m_axi_m_axi_AWQOS,
    output wire                                          vec_Y__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] vec_Y__m_axi_m_axi_AWSIZE,
    input wire                                           vec_Y__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] vec_Y__m_axi_m_axi_BID,
    input wire                                           vec_Y__m_axi_m_axi_BREADY,
    output wire [                                   1:0] vec_Y__m_axi_m_axi_BRESP,
    output wire                                          vec_Y__m_axi_m_axi_BVALID,
    output wire [                                 255:0] vec_Y__m_axi_m_axi_RDATA,
    output wire [                                   0:0] vec_Y__m_axi_m_axi_RID,
    output wire                                          vec_Y__m_axi_m_axi_RLAST,
    input wire                                           vec_Y__m_axi_m_axi_RREADY,
    output wire [                                   1:0] vec_Y__m_axi_m_axi_RRESP,
    output wire                                          vec_Y__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] vec_Y__m_axi_m_axi_WDATA,
    input wire                                           vec_Y__m_axi_m_axi_WLAST,
    output wire                                          vec_Y__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] vec_Y__m_axi_m_axi_WSTRB,
    input wire                                           vec_Y__m_axi_m_axi_WVALID,
    output wire [                                  63:0] vec_Y__m_axi_read_addr_din,
    input wire                                           vec_Y__m_axi_read_addr_full_n,
    output wire                                          vec_Y__m_axi_read_addr_write,
    input wire  [                                 255:0] vec_Y__m_axi_read_data_dout,
    input wire                                           vec_Y__m_axi_read_data_empty_n,
    output wire                                          vec_Y__m_axi_read_data_read,
    output wire                                          vec_Y__m_axi_rst,
    output wire [                                  63:0] vec_Y__m_axi_write_addr_din,
    input wire                                           vec_Y__m_axi_write_addr_full_n,
    output wire                                          vec_Y__m_axi_write_addr_write,
    output wire [                                 255:0] vec_Y__m_axi_write_data_din,
    input wire                                           vec_Y__m_axi_write_data_full_n,
    output wire                                          vec_Y__m_axi_write_data_write,
    input wire  [                                   7:0] vec_Y__m_axi_write_resp_dout,
    input wire                                           vec_Y__m_axi_write_resp_empty_n,
    output wire                                          vec_Y__m_axi_write_resp_read,
    output wire                                          edge_list_ptr__m_axi_clk,
    input wire  [                                  63:0] edge_list_ptr__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] edge_list_ptr__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] edge_list_ptr__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] edge_list_ptr__m_axi_m_axi_ARID,
    input wire  [                                   7:0] edge_list_ptr__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] edge_list_ptr__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] edge_list_ptr__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] edge_list_ptr__m_axi_m_axi_ARQOS,
    output wire                                          edge_list_ptr__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] edge_list_ptr__m_axi_m_axi_ARSIZE,
    input wire                                           edge_list_ptr__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] edge_list_ptr__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] edge_list_ptr__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] edge_list_ptr__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] edge_list_ptr__m_axi_m_axi_AWID,
    input wire  [                                   7:0] edge_list_ptr__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] edge_list_ptr__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] edge_list_ptr__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] edge_list_ptr__m_axi_m_axi_AWQOS,
    output wire                                          edge_list_ptr__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] edge_list_ptr__m_axi_m_axi_AWSIZE,
    input wire                                           edge_list_ptr__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] edge_list_ptr__m_axi_m_axi_BID,
    input wire                                           edge_list_ptr__m_axi_m_axi_BREADY,
    output wire [                                   1:0] edge_list_ptr__m_axi_m_axi_BRESP,
    output wire                                          edge_list_ptr__m_axi_m_axi_BVALID,
    output wire [                                  31:0] edge_list_ptr__m_axi_m_axi_RDATA,
    output wire [                                   0:0] edge_list_ptr__m_axi_m_axi_RID,
    output wire                                          edge_list_ptr__m_axi_m_axi_RLAST,
    input wire                                           edge_list_ptr__m_axi_m_axi_RREADY,
    output wire [                                   1:0] edge_list_ptr__m_axi_m_axi_RRESP,
    output wire                                          edge_list_ptr__m_axi_m_axi_RVALID,
    input wire  [                                  31:0] edge_list_ptr__m_axi_m_axi_WDATA,
    input wire                                           edge_list_ptr__m_axi_m_axi_WLAST,
    output wire                                          edge_list_ptr__m_axi_m_axi_WREADY,
    input wire  [                                   3:0] edge_list_ptr__m_axi_m_axi_WSTRB,
    input wire                                           edge_list_ptr__m_axi_m_axi_WVALID,
    output wire [                                  63:0] edge_list_ptr__m_axi_read_addr_din,
    input wire                                           edge_list_ptr__m_axi_read_addr_full_n,
    output wire                                          edge_list_ptr__m_axi_read_addr_write,
    input wire  [                                  31:0] edge_list_ptr__m_axi_read_data_dout,
    input wire                                           edge_list_ptr__m_axi_read_data_empty_n,
    output wire                                          edge_list_ptr__m_axi_read_data_read,
    output wire                                          edge_list_ptr__m_axi_rst,
    output wire [                                  63:0] edge_list_ptr__m_axi_write_addr_din,
    input wire                                           edge_list_ptr__m_axi_write_addr_full_n,
    output wire                                          edge_list_ptr__m_axi_write_addr_write,
    output wire [                                  31:0] edge_list_ptr__m_axi_write_data_din,
    input wire                                           edge_list_ptr__m_axi_write_data_full_n,
    output wire                                          edge_list_ptr__m_axi_write_data_write,
    input wire  [                                   7:0] edge_list_ptr__m_axi_write_resp_dout,
    input wire                                           edge_list_ptr__m_axi_write_resp_empty_n,
    output wire                                          edge_list_ptr__m_axi_write_resp_read,
    output wire                                          vec_Y_out__m_axi_clk,
    input wire  [                                  63:0] vec_Y_out__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] vec_Y_out__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] vec_Y_out__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] vec_Y_out__m_axi_m_axi_ARID,
    input wire  [                                   7:0] vec_Y_out__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] vec_Y_out__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] vec_Y_out__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] vec_Y_out__m_axi_m_axi_ARQOS,
    output wire                                          vec_Y_out__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] vec_Y_out__m_axi_m_axi_ARSIZE,
    input wire                                           vec_Y_out__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] vec_Y_out__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] vec_Y_out__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] vec_Y_out__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] vec_Y_out__m_axi_m_axi_AWID,
    input wire  [                                   7:0] vec_Y_out__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] vec_Y_out__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] vec_Y_out__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] vec_Y_out__m_axi_m_axi_AWQOS,
    output wire                                          vec_Y_out__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] vec_Y_out__m_axi_m_axi_AWSIZE,
    input wire                                           vec_Y_out__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] vec_Y_out__m_axi_m_axi_BID,
    input wire                                           vec_Y_out__m_axi_m_axi_BREADY,
    output wire [                                   1:0] vec_Y_out__m_axi_m_axi_BRESP,
    output wire                                          vec_Y_out__m_axi_m_axi_BVALID,
    output wire [                                 255:0] vec_Y_out__m_axi_m_axi_RDATA,
    output wire [                                   0:0] vec_Y_out__m_axi_m_axi_RID,
    output wire                                          vec_Y_out__m_axi_m_axi_RLAST,
    input wire                                           vec_Y_out__m_axi_m_axi_RREADY,
    output wire [                                   1:0] vec_Y_out__m_axi_m_axi_RRESP,
    output wire                                          vec_Y_out__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] vec_Y_out__m_axi_m_axi_WDATA,
    input wire                                           vec_Y_out__m_axi_m_axi_WLAST,
    output wire                                          vec_Y_out__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] vec_Y_out__m_axi_m_axi_WSTRB,
    input wire                                           vec_Y_out__m_axi_m_axi_WVALID,
    output wire [                                  63:0] vec_Y_out__m_axi_read_addr_din,
    input wire                                           vec_Y_out__m_axi_read_addr_full_n,
    output wire                                          vec_Y_out__m_axi_read_addr_write,
    input wire  [                                 255:0] vec_Y_out__m_axi_read_data_dout,
    input wire                                           vec_Y_out__m_axi_read_data_empty_n,
    output wire                                          vec_Y_out__m_axi_read_data_read,
    output wire                                          vec_Y_out__m_axi_rst,
    output wire [                                  63:0] vec_Y_out__m_axi_write_addr_din,
    input wire                                           vec_Y_out__m_axi_write_addr_full_n,
    output wire                                          vec_Y_out__m_axi_write_addr_write,
    output wire [                                 255:0] vec_Y_out__m_axi_write_data_din,
    input wire                                           vec_Y_out__m_axi_write_data_full_n,
    output wire                                          vec_Y_out__m_axi_write_data_write,
    input wire  [                                   7:0] vec_Y_out__m_axi_write_resp_dout,
    input wire                                           vec_Y_out__m_axi_write_resp_empty_n,
    output wire                                          vec_Y_out__m_axi_write_resp_read,
    input wire  [                                  31:0] __tapa_fsm_unit_Arbiter_Y_0___M__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_Arbiter_Y_0___P_N__q0,
    output wire                                          __tapa_fsm_unit_Arbiter_Y_0__ap_done,
    output wire                                          __tapa_fsm_unit_Arbiter_Y_0__ap_idle,
    output wire                                          __tapa_fsm_unit_Arbiter_Y_0__ap_ready,
    input wire                                           __tapa_fsm_unit_Arbiter_Y_0__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_Arbiter_Y_1___M__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_Arbiter_Y_1___P_N__q0,
    output wire                                          __tapa_fsm_unit_Arbiter_Y_1__ap_done,
    output wire                                          __tapa_fsm_unit_Arbiter_Y_1__ap_idle,
    output wire                                          __tapa_fsm_unit_Arbiter_Y_1__ap_ready,
    input wire                                           __tapa_fsm_unit_Arbiter_Y_1__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_Arbiter_Y_2___M__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_Arbiter_Y_2___P_N__q0,
    output wire                                          __tapa_fsm_unit_Arbiter_Y_2__ap_done,
    output wire                                          __tapa_fsm_unit_Arbiter_Y_2__ap_idle,
    output wire                                          __tapa_fsm_unit_Arbiter_Y_2__ap_ready,
    input wire                                           __tapa_fsm_unit_Arbiter_Y_2__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_Arbiter_Y_3___M__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_Arbiter_Y_3___P_N__q0,
    output wire                                          __tapa_fsm_unit_Arbiter_Y_3__ap_done,
    output wire                                          __tapa_fsm_unit_Arbiter_Y_3__ap_idle,
    output wire                                          __tapa_fsm_unit_Arbiter_Y_3__ap_ready,
    input wire                                           __tapa_fsm_unit_Arbiter_Y_3__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_Arbiter_Y_4___M__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_Arbiter_Y_4___P_N__q0,
    output wire                                          __tapa_fsm_unit_Arbiter_Y_4__ap_done,
    output wire                                          __tapa_fsm_unit_Arbiter_Y_4__ap_idle,
    output wire                                          __tapa_fsm_unit_Arbiter_Y_4__ap_ready,
    input wire                                           __tapa_fsm_unit_Arbiter_Y_4__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_Arbiter_Y_5___M__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_Arbiter_Y_5___P_N__q0,
    output wire                                          __tapa_fsm_unit_Arbiter_Y_5__ap_done,
    output wire                                          __tapa_fsm_unit_Arbiter_Y_5__ap_idle,
    output wire                                          __tapa_fsm_unit_Arbiter_Y_5__ap_ready,
    input wire                                           __tapa_fsm_unit_Arbiter_Y_5__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_Arbiter_Y_6___M__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_Arbiter_Y_6___P_N__q0,
    output wire                                          __tapa_fsm_unit_Arbiter_Y_6__ap_done,
    output wire                                          __tapa_fsm_unit_Arbiter_Y_6__ap_idle,
    output wire                                          __tapa_fsm_unit_Arbiter_Y_6__ap_ready,
    input wire                                           __tapa_fsm_unit_Arbiter_Y_6__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_Arbiter_Y_7___M__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_Arbiter_Y_7___P_N__q0,
    output wire                                          __tapa_fsm_unit_Arbiter_Y_7__ap_done,
    output wire                                          __tapa_fsm_unit_Arbiter_Y_7__ap_idle,
    output wire                                          __tapa_fsm_unit_Arbiter_Y_7__ap_ready,
    input wire                                           __tapa_fsm_unit_Arbiter_Y_7__ap_start,
    input wire                                           __tapa_fsm_unit_FloatvAddFloatv_0__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_FloatvMultConst_0___M__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_FloatvMultConst_0___P_N__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_FloatvMultConst_0___alpha_u__q0,
    output wire                                          __tapa_fsm_unit_FloatvMultConst_0__ap_done,
    output wire                                          __tapa_fsm_unit_FloatvMultConst_0__ap_idle,
    output wire                                          __tapa_fsm_unit_FloatvMultConst_0__ap_ready,
    input wire                                           __tapa_fsm_unit_FloatvMultConst_0__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_FloatvMultConst_1___M__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_FloatvMultConst_1___P_N__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_FloatvMultConst_1___beta_u__q0,
    output wire                                          __tapa_fsm_unit_FloatvMultConst_1__ap_done,
    output wire                                          __tapa_fsm_unit_FloatvMultConst_1__ap_idle,
    output wire                                          __tapa_fsm_unit_FloatvMultConst_1__ap_ready,
    input wire                                           __tapa_fsm_unit_FloatvMultConst_1__ap_start,
    output wire [                                  31:0] __tapa_fsm_unit_K,
    output wire [                                  31:0] __tapa_fsm_unit_M,
    input wire                                           __tapa_fsm_unit_Merger_Y_0__ap_start,
    output wire [                                  31:0] __tapa_fsm_unit_NUM_A_LEN,
    output wire [                                  31:0] __tapa_fsm_unit_NUM_ITE,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_0__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_0__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_0__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_0__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_10__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_10__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_10__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_10__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_11__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_11__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_11__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_11__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_12__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_12__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_12__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_12__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_13__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_13__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_13__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_13__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_14__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_14__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_14__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_14__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_15__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_15__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_15__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_15__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_16__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_16__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_16__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_16__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_17__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_17__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_17__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_17__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_18__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_18__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_18__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_18__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_19__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_19__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_19__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_19__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_1__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_1__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_1__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_1__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_20__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_20__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_20__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_20__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_21__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_21__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_21__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_21__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_22__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_22__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_22__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_22__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_23__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_23__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_23__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_23__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_24__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_24__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_24__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_24__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_25__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_25__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_25__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_25__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_26__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_26__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_26__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_26__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_27__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_27__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_27__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_27__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_28__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_28__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_28__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_28__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_29__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_29__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_29__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_29__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_2__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_2__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_2__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_2__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_30__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_30__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_30__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_30__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_31__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_31__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_31__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_31__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_32__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_32__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_32__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_32__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_33__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_33__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_33__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_33__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_34__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_34__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_34__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_34__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_35__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_35__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_35__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_35__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_36__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_36__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_36__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_36__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_37__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_37__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_37__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_37__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_38__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_38__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_38__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_38__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_39__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_39__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_39__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_39__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_3__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_3__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_3__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_3__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_40__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_40__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_40__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_40__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_41__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_41__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_41__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_41__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_42__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_42__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_42__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_42__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_43__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_43__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_43__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_43__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_44__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_44__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_44__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_44__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_45__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_45__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_45__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_45__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_46__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_46__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_46__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_46__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_47__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_47__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_47__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_47__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_4__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_4__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_4__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_4__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_5__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_5__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_5__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_5__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_6__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_6__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_6__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_6__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_7__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_7__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_7__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_7__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_8__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_8__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_8__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_8__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_9__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_9__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Xvec_9__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Xvec_9__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_0__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_0__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_0__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_0__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_10__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_10__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_10__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_10__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_11__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_11__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_11__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_11__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_12__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_12__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_12__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_12__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_13__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_13__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_13__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_13__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_14__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_14__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_14__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_14__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_15__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_15__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_15__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_15__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_16__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_16__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_16__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_16__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_17__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_17__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_17__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_17__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_18__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_18__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_18__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_18__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_19__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_19__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_19__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_19__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_1__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_1__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_1__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_1__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_20__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_20__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_20__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_20__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_21__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_21__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_21__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_21__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_22__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_22__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_22__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_22__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_23__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_23__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_23__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_23__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_24__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_24__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_24__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_24__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_25__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_25__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_25__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_25__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_26__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_26__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_26__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_26__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_27__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_27__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_27__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_27__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_28__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_28__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_28__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_28__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_29__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_29__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_29__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_29__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_2__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_2__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_2__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_2__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_30__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_30__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_30__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_30__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_31__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_31__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_31__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_31__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_32__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_32__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_32__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_32__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_33__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_33__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_33__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_33__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_34__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_34__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_34__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_34__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_35__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_35__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_35__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_35__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_36__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_36__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_36__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_36__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_37__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_37__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_37__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_37__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_38__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_38__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_38__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_38__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_39__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_39__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_39__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_39__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_3__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_3__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_3__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_3__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_40__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_40__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_40__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_40__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_41__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_41__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_41__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_41__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_42__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_42__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_42__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_42__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_43__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_43__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_43__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_43__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_44__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_44__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_44__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_44__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_45__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_45__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_45__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_45__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_46__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_46__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_46__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_46__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_47__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_47__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_47__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_47__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_4__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_4__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_4__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_4__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_5__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_5__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_5__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_5__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_6__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_6__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_6__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_6__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_7__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_7__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_7__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_7__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_8__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_8__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_8__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_8__ap_start,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_9__ap_done,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_9__ap_idle,
    output wire                                          __tapa_fsm_unit_PEG_Yvec_9__ap_ready,
    input wire                                           __tapa_fsm_unit_PEG_Yvec_9__ap_start,
    output wire [                                  31:0] __tapa_fsm_unit_P_N,
    output wire [                                  31:0] __tapa_fsm_unit_alpha_u,
    output wire                                          __tapa_fsm_unit_ap_clk,
    input wire                                           __tapa_fsm_unit_ap_done,
    input wire                                           __tapa_fsm_unit_ap_idle,
    input wire                                           __tapa_fsm_unit_ap_ready,
    output wire                                          __tapa_fsm_unit_ap_rst_n,
    output wire                                          __tapa_fsm_unit_ap_start,
    output wire [                                  31:0] __tapa_fsm_unit_beta_u,
    input wire                                           __tapa_fsm_unit_black_hole_float_v16_0__ap_start,
    input wire                                           __tapa_fsm_unit_black_hole_int_0__ap_start,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_0,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_1,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_10,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_11,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_12,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_13,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_14,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_15,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_16,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_17,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_18,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_19,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_2,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_20,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_21,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_22,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_23,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_24,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_25,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_26,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_27,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_28,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_29,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_3,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_30,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_31,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_32,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_33,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_34,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_35,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_36,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_37,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_38,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_39,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_4,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_40,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_41,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_42,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_43,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_44,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_45,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_46,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_47,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_5,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_6,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_7,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_8,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ch_9,
    output wire [                                  63:0] __tapa_fsm_unit_edge_list_ptr,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_0___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_0___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_0___edge_list_ch_0__q0,
    output wire                                          __tapa_fsm_unit_read_A_0__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_0__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_0__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_0__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_10___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_10___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_10___edge_list_ch_10__q0,
    output wire                                          __tapa_fsm_unit_read_A_10__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_10__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_10__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_10__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_11___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_11___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_11___edge_list_ch_11__q0,
    output wire                                          __tapa_fsm_unit_read_A_11__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_11__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_11__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_11__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_12___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_12___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_12___edge_list_ch_12__q0,
    output wire                                          __tapa_fsm_unit_read_A_12__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_12__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_12__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_12__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_13___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_13___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_13___edge_list_ch_13__q0,
    output wire                                          __tapa_fsm_unit_read_A_13__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_13__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_13__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_13__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_14___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_14___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_14___edge_list_ch_14__q0,
    output wire                                          __tapa_fsm_unit_read_A_14__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_14__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_14__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_14__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_15___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_15___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_15___edge_list_ch_15__q0,
    output wire                                          __tapa_fsm_unit_read_A_15__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_15__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_15__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_15__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_16___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_16___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_16___edge_list_ch_16__q0,
    output wire                                          __tapa_fsm_unit_read_A_16__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_16__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_16__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_16__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_17___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_17___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_17___edge_list_ch_17__q0,
    output wire                                          __tapa_fsm_unit_read_A_17__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_17__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_17__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_17__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_18___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_18___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_18___edge_list_ch_18__q0,
    output wire                                          __tapa_fsm_unit_read_A_18__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_18__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_18__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_18__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_19___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_19___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_19___edge_list_ch_19__q0,
    output wire                                          __tapa_fsm_unit_read_A_19__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_19__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_19__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_19__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_1___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_1___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_1___edge_list_ch_1__q0,
    output wire                                          __tapa_fsm_unit_read_A_1__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_1__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_1__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_1__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_20___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_20___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_20___edge_list_ch_20__q0,
    output wire                                          __tapa_fsm_unit_read_A_20__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_20__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_20__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_20__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_21___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_21___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_21___edge_list_ch_21__q0,
    output wire                                          __tapa_fsm_unit_read_A_21__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_21__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_21__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_21__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_22___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_22___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_22___edge_list_ch_22__q0,
    output wire                                          __tapa_fsm_unit_read_A_22__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_22__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_22__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_22__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_23___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_23___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_23___edge_list_ch_23__q0,
    output wire                                          __tapa_fsm_unit_read_A_23__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_23__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_23__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_23__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_24___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_24___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_24___edge_list_ch_24__q0,
    output wire                                          __tapa_fsm_unit_read_A_24__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_24__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_24__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_24__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_25___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_25___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_25___edge_list_ch_25__q0,
    output wire                                          __tapa_fsm_unit_read_A_25__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_25__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_25__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_25__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_26___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_26___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_26___edge_list_ch_26__q0,
    output wire                                          __tapa_fsm_unit_read_A_26__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_26__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_26__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_26__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_27___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_27___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_27___edge_list_ch_27__q0,
    output wire                                          __tapa_fsm_unit_read_A_27__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_27__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_27__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_27__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_28___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_28___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_28___edge_list_ch_28__q0,
    output wire                                          __tapa_fsm_unit_read_A_28__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_28__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_28__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_28__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_29___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_29___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_29___edge_list_ch_29__q0,
    output wire                                          __tapa_fsm_unit_read_A_29__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_29__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_29__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_29__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_2___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_2___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_2___edge_list_ch_2__q0,
    output wire                                          __tapa_fsm_unit_read_A_2__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_2__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_2__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_2__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_30___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_30___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_30___edge_list_ch_30__q0,
    output wire                                          __tapa_fsm_unit_read_A_30__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_30__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_30__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_30__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_31___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_31___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_31___edge_list_ch_31__q0,
    output wire                                          __tapa_fsm_unit_read_A_31__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_31__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_31__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_31__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_32___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_32___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_32___edge_list_ch_32__q0,
    output wire                                          __tapa_fsm_unit_read_A_32__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_32__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_32__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_32__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_33___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_33___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_33___edge_list_ch_33__q0,
    output wire                                          __tapa_fsm_unit_read_A_33__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_33__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_33__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_33__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_34___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_34___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_34___edge_list_ch_34__q0,
    output wire                                          __tapa_fsm_unit_read_A_34__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_34__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_34__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_34__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_35___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_35___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_35___edge_list_ch_35__q0,
    output wire                                          __tapa_fsm_unit_read_A_35__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_35__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_35__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_35__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_36___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_36___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_36___edge_list_ch_36__q0,
    output wire                                          __tapa_fsm_unit_read_A_36__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_36__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_36__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_36__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_37___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_37___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_37___edge_list_ch_37__q0,
    output wire                                          __tapa_fsm_unit_read_A_37__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_37__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_37__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_37__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_38___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_38___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_38___edge_list_ch_38__q0,
    output wire                                          __tapa_fsm_unit_read_A_38__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_38__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_38__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_38__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_39___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_39___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_39___edge_list_ch_39__q0,
    output wire                                          __tapa_fsm_unit_read_A_39__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_39__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_39__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_39__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_3___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_3___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_3___edge_list_ch_3__q0,
    output wire                                          __tapa_fsm_unit_read_A_3__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_3__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_3__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_3__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_40___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_40___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_40___edge_list_ch_40__q0,
    output wire                                          __tapa_fsm_unit_read_A_40__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_40__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_40__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_40__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_41___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_41___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_41___edge_list_ch_41__q0,
    output wire                                          __tapa_fsm_unit_read_A_41__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_41__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_41__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_41__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_42___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_42___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_42___edge_list_ch_42__q0,
    output wire                                          __tapa_fsm_unit_read_A_42__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_42__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_42__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_42__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_43___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_43___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_43___edge_list_ch_43__q0,
    output wire                                          __tapa_fsm_unit_read_A_43__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_43__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_43__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_43__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_44___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_44___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_44___edge_list_ch_44__q0,
    output wire                                          __tapa_fsm_unit_read_A_44__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_44__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_44__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_44__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_45___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_45___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_45___edge_list_ch_45__q0,
    output wire                                          __tapa_fsm_unit_read_A_45__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_45__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_45__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_45__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_46___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_46___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_46___edge_list_ch_46__q0,
    output wire                                          __tapa_fsm_unit_read_A_46__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_46__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_46__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_46__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_47___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_47___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_47___edge_list_ch_47__q0,
    output wire                                          __tapa_fsm_unit_read_A_47__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_47__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_47__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_47__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_4___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_4___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_4___edge_list_ch_4__q0,
    output wire                                          __tapa_fsm_unit_read_A_4__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_4__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_4__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_4__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_5___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_5___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_5___edge_list_ch_5__q0,
    output wire                                          __tapa_fsm_unit_read_A_5__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_5__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_5__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_5__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_6___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_6___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_6___edge_list_ch_6__q0,
    output wire                                          __tapa_fsm_unit_read_A_6__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_6__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_6__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_6__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_7___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_7___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_7___edge_list_ch_7__q0,
    output wire                                          __tapa_fsm_unit_read_A_7__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_7__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_7__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_7__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_8___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_8___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_8___edge_list_ch_8__q0,
    output wire                                          __tapa_fsm_unit_read_A_8__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_8__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_8__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_8__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_9___NUM_A_LEN__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_A_9___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_A_9___edge_list_ch_9__q0,
    output wire                                          __tapa_fsm_unit_read_A_9__ap_done,
    output wire                                          __tapa_fsm_unit_read_A_9__ap_idle,
    output wire                                          __tapa_fsm_unit_read_A_9__ap_ready,
    input wire                                           __tapa_fsm_unit_read_A_9__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_X_0___K__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_X_0___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_X_0___vec_X__q0,
    output wire                                          __tapa_fsm_unit_read_X_0__ap_done,
    output wire                                          __tapa_fsm_unit_read_X_0__ap_idle,
    output wire                                          __tapa_fsm_unit_read_X_0__ap_ready,
    input wire                                           __tapa_fsm_unit_read_X_0__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_Y_0___M__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_Y_0___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_Y_0___vec_Y__q0,
    output wire                                          __tapa_fsm_unit_read_Y_0__ap_done,
    output wire                                          __tapa_fsm_unit_read_Y_0__ap_idle,
    output wire                                          __tapa_fsm_unit_read_Y_0__ap_ready,
    input wire                                           __tapa_fsm_unit_read_Y_0__ap_start,
    input wire  [                                  31:0] __tapa_fsm_unit_read_edge_list_ptr_0___K__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_edge_list_ptr_0___M__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_edge_list_ptr_0___NUM_ITE__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_read_edge_list_ptr_0___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_read_edge_list_ptr_0___edge_list_ptr__q0,
    output wire                                          __tapa_fsm_unit_read_edge_list_ptr_0__ap_done,
    output wire                                          __tapa_fsm_unit_read_edge_list_ptr_0__ap_idle,
    output wire                                          __tapa_fsm_unit_read_edge_list_ptr_0__ap_ready,
    input wire                                           __tapa_fsm_unit_read_edge_list_ptr_0__ap_start,
    output wire [                                  63:0] __tapa_fsm_unit_vec_X,
    output wire [                                  63:0] __tapa_fsm_unit_vec_Y,
    output wire [                                  63:0] __tapa_fsm_unit_vec_Y_out,
    input wire  [                                  31:0] __tapa_fsm_unit_write_Y_0___M__q0,
    input wire  [                                  31:0] __tapa_fsm_unit_write_Y_0___P_N__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_write_Y_0___vec_Y_out__q0,
    output wire                                          __tapa_fsm_unit_write_Y_0__ap_done,
    output wire                                          __tapa_fsm_unit_write_Y_0__ap_idle,
    output wire                                          __tapa_fsm_unit_write_Y_0__ap_ready,
    input wire                                           __tapa_fsm_unit_write_Y_0__ap_start
);
  wire ap_start;
  wire [63:0] edge_list_ptr;
  wire [63:0] edge_list_ch_0;
  wire [63:0] edge_list_ch_1;
  wire [63:0] edge_list_ch_2;
  wire [63:0] edge_list_ch_3;
  wire [63:0] edge_list_ch_4;
  wire [63:0] edge_list_ch_5;
  wire [63:0] edge_list_ch_6;
  wire [63:0] edge_list_ch_7;
  wire [63:0] edge_list_ch_8;
  wire [63:0] edge_list_ch_9;
  wire [63:0] edge_list_ch_10;
  wire [63:0] edge_list_ch_11;
  wire [63:0] edge_list_ch_12;
  wire [63:0] edge_list_ch_13;
  wire [63:0] edge_list_ch_14;
  wire [63:0] edge_list_ch_15;
  wire [63:0] edge_list_ch_16;
  wire [63:0] edge_list_ch_17;
  wire [63:0] edge_list_ch_18;
  wire [63:0] edge_list_ch_19;
  wire [63:0] edge_list_ch_20;
  wire [63:0] edge_list_ch_21;
  wire [63:0] edge_list_ch_22;
  wire [63:0] edge_list_ch_23;
  wire [63:0] edge_list_ch_24;
  wire [63:0] edge_list_ch_25;
  wire [63:0] edge_list_ch_26;
  wire [63:0] edge_list_ch_27;
  wire [63:0] edge_list_ch_28;
  wire [63:0] edge_list_ch_29;
  wire [63:0] edge_list_ch_30;
  wire [63:0] edge_list_ch_31;
  wire [63:0] edge_list_ch_32;
  wire [63:0] edge_list_ch_33;
  wire [63:0] edge_list_ch_34;
  wire [63:0] edge_list_ch_35;
  wire [63:0] edge_list_ch_36;
  wire [63:0] edge_list_ch_37;
  wire [63:0] edge_list_ch_38;
  wire [63:0] edge_list_ch_39;
  wire [63:0] edge_list_ch_40;
  wire [63:0] edge_list_ch_41;
  wire [63:0] edge_list_ch_42;
  wire [63:0] edge_list_ch_43;
  wire [63:0] edge_list_ch_44;
  wire [63:0] edge_list_ch_45;
  wire [63:0] edge_list_ch_46;
  wire [63:0] edge_list_ch_47;
  wire [63:0] vec_X;
  wire [63:0] vec_Y;
  wire [63:0] vec_Y_out;
  wire [31:0] NUM_ITE;
  wire [31:0] NUM_A_LEN;
  wire [31:0] M;
  wire [31:0] K;
  wire [31:0] P_N;
  wire [31:0] alpha_u;
  wire [31:0] beta_u;
  wire [32:0] PE_inst_0__dout;
  wire PE_inst_0__empty_n;
  wire PE_inst_0__read;
  wire [32:0] PE_inst_0__din;
  wire PE_inst_0__full_n;
  wire PE_inst_0__write;
  wire [32:0] PE_inst_10__dout;
  wire PE_inst_10__empty_n;
  wire PE_inst_10__read;
  wire [32:0] PE_inst_10__din;
  wire PE_inst_10__full_n;
  wire PE_inst_10__write;
  wire [32:0] PE_inst_11__dout;
  wire PE_inst_11__empty_n;
  wire PE_inst_11__read;
  wire [32:0] PE_inst_11__din;
  wire PE_inst_11__full_n;
  wire PE_inst_11__write;
  wire [32:0] PE_inst_12__dout;
  wire PE_inst_12__empty_n;
  wire PE_inst_12__read;
  wire [32:0] PE_inst_12__din;
  wire PE_inst_12__full_n;
  wire PE_inst_12__write;
  wire [32:0] PE_inst_13__dout;
  wire PE_inst_13__empty_n;
  wire PE_inst_13__read;
  wire [32:0] PE_inst_13__din;
  wire PE_inst_13__full_n;
  wire PE_inst_13__write;
  wire [32:0] PE_inst_14__dout;
  wire PE_inst_14__empty_n;
  wire PE_inst_14__read;
  wire [32:0] PE_inst_14__din;
  wire PE_inst_14__full_n;
  wire PE_inst_14__write;
  wire [32:0] PE_inst_15__dout;
  wire PE_inst_15__empty_n;
  wire PE_inst_15__read;
  wire [32:0] PE_inst_15__din;
  wire PE_inst_15__full_n;
  wire PE_inst_15__write;
  wire [32:0] PE_inst_16__dout;
  wire PE_inst_16__empty_n;
  wire PE_inst_16__read;
  wire [32:0] PE_inst_16__din;
  wire PE_inst_16__full_n;
  wire PE_inst_16__write;
  wire [32:0] PE_inst_17__dout;
  wire PE_inst_17__empty_n;
  wire PE_inst_17__read;
  wire [32:0] PE_inst_17__din;
  wire PE_inst_17__full_n;
  wire PE_inst_17__write;
  wire [32:0] PE_inst_18__dout;
  wire PE_inst_18__empty_n;
  wire PE_inst_18__read;
  wire [32:0] PE_inst_18__din;
  wire PE_inst_18__full_n;
  wire PE_inst_18__write;
  wire [32:0] PE_inst_19__dout;
  wire PE_inst_19__empty_n;
  wire PE_inst_19__read;
  wire [32:0] PE_inst_19__din;
  wire PE_inst_19__full_n;
  wire PE_inst_19__write;
  wire [32:0] PE_inst_1__dout;
  wire PE_inst_1__empty_n;
  wire PE_inst_1__read;
  wire [32:0] PE_inst_1__din;
  wire PE_inst_1__full_n;
  wire PE_inst_1__write;
  wire [32:0] PE_inst_20__dout;
  wire PE_inst_20__empty_n;
  wire PE_inst_20__read;
  wire [32:0] PE_inst_20__din;
  wire PE_inst_20__full_n;
  wire PE_inst_20__write;
  wire [32:0] PE_inst_21__dout;
  wire PE_inst_21__empty_n;
  wire PE_inst_21__read;
  wire [32:0] PE_inst_21__din;
  wire PE_inst_21__full_n;
  wire PE_inst_21__write;
  wire [32:0] PE_inst_22__dout;
  wire PE_inst_22__empty_n;
  wire PE_inst_22__read;
  wire [32:0] PE_inst_22__din;
  wire PE_inst_22__full_n;
  wire PE_inst_22__write;
  wire [32:0] PE_inst_23__dout;
  wire PE_inst_23__empty_n;
  wire PE_inst_23__read;
  wire [32:0] PE_inst_23__din;
  wire PE_inst_23__full_n;
  wire PE_inst_23__write;
  wire [32:0] PE_inst_24__dout;
  wire PE_inst_24__empty_n;
  wire PE_inst_24__read;
  wire [32:0] PE_inst_24__din;
  wire PE_inst_24__full_n;
  wire PE_inst_24__write;
  wire [32:0] PE_inst_25__dout;
  wire PE_inst_25__empty_n;
  wire PE_inst_25__read;
  wire [32:0] PE_inst_25__din;
  wire PE_inst_25__full_n;
  wire PE_inst_25__write;
  wire [32:0] PE_inst_26__dout;
  wire PE_inst_26__empty_n;
  wire PE_inst_26__read;
  wire [32:0] PE_inst_26__din;
  wire PE_inst_26__full_n;
  wire PE_inst_26__write;
  wire [32:0] PE_inst_27__dout;
  wire PE_inst_27__empty_n;
  wire PE_inst_27__read;
  wire [32:0] PE_inst_27__din;
  wire PE_inst_27__full_n;
  wire PE_inst_27__write;
  wire [32:0] PE_inst_28__dout;
  wire PE_inst_28__empty_n;
  wire PE_inst_28__read;
  wire [32:0] PE_inst_28__din;
  wire PE_inst_28__full_n;
  wire PE_inst_28__write;
  wire [32:0] PE_inst_29__dout;
  wire PE_inst_29__empty_n;
  wire PE_inst_29__read;
  wire [32:0] PE_inst_29__din;
  wire PE_inst_29__full_n;
  wire PE_inst_29__write;
  wire [32:0] PE_inst_2__dout;
  wire PE_inst_2__empty_n;
  wire PE_inst_2__read;
  wire [32:0] PE_inst_2__din;
  wire PE_inst_2__full_n;
  wire PE_inst_2__write;
  wire [32:0] PE_inst_30__dout;
  wire PE_inst_30__empty_n;
  wire PE_inst_30__read;
  wire [32:0] PE_inst_30__din;
  wire PE_inst_30__full_n;
  wire PE_inst_30__write;
  wire [32:0] PE_inst_31__dout;
  wire PE_inst_31__empty_n;
  wire PE_inst_31__read;
  wire [32:0] PE_inst_31__din;
  wire PE_inst_31__full_n;
  wire PE_inst_31__write;
  wire [32:0] PE_inst_32__dout;
  wire PE_inst_32__empty_n;
  wire PE_inst_32__read;
  wire [32:0] PE_inst_32__din;
  wire PE_inst_32__full_n;
  wire PE_inst_32__write;
  wire [32:0] PE_inst_33__dout;
  wire PE_inst_33__empty_n;
  wire PE_inst_33__read;
  wire [32:0] PE_inst_33__din;
  wire PE_inst_33__full_n;
  wire PE_inst_33__write;
  wire [32:0] PE_inst_34__dout;
  wire PE_inst_34__empty_n;
  wire PE_inst_34__read;
  wire [32:0] PE_inst_34__din;
  wire PE_inst_34__full_n;
  wire PE_inst_34__write;
  wire [32:0] PE_inst_35__dout;
  wire PE_inst_35__empty_n;
  wire PE_inst_35__read;
  wire [32:0] PE_inst_35__din;
  wire PE_inst_35__full_n;
  wire PE_inst_35__write;
  wire [32:0] PE_inst_36__dout;
  wire PE_inst_36__empty_n;
  wire PE_inst_36__read;
  wire [32:0] PE_inst_36__din;
  wire PE_inst_36__full_n;
  wire PE_inst_36__write;
  wire [32:0] PE_inst_37__dout;
  wire PE_inst_37__empty_n;
  wire PE_inst_37__read;
  wire [32:0] PE_inst_37__din;
  wire PE_inst_37__full_n;
  wire PE_inst_37__write;
  wire [32:0] PE_inst_38__dout;
  wire PE_inst_38__empty_n;
  wire PE_inst_38__read;
  wire [32:0] PE_inst_38__din;
  wire PE_inst_38__full_n;
  wire PE_inst_38__write;
  wire [32:0] PE_inst_39__dout;
  wire PE_inst_39__empty_n;
  wire PE_inst_39__read;
  wire [32:0] PE_inst_39__din;
  wire PE_inst_39__full_n;
  wire PE_inst_39__write;
  wire [32:0] PE_inst_3__dout;
  wire PE_inst_3__empty_n;
  wire PE_inst_3__read;
  wire [32:0] PE_inst_3__din;
  wire PE_inst_3__full_n;
  wire PE_inst_3__write;
  wire [32:0] PE_inst_40__dout;
  wire PE_inst_40__empty_n;
  wire PE_inst_40__read;
  wire [32:0] PE_inst_40__din;
  wire PE_inst_40__full_n;
  wire PE_inst_40__write;
  wire [32:0] PE_inst_41__dout;
  wire PE_inst_41__empty_n;
  wire PE_inst_41__read;
  wire [32:0] PE_inst_41__din;
  wire PE_inst_41__full_n;
  wire PE_inst_41__write;
  wire [32:0] PE_inst_42__dout;
  wire PE_inst_42__empty_n;
  wire PE_inst_42__read;
  wire [32:0] PE_inst_42__din;
  wire PE_inst_42__full_n;
  wire PE_inst_42__write;
  wire [32:0] PE_inst_43__dout;
  wire PE_inst_43__empty_n;
  wire PE_inst_43__read;
  wire [32:0] PE_inst_43__din;
  wire PE_inst_43__full_n;
  wire PE_inst_43__write;
  wire [32:0] PE_inst_44__dout;
  wire PE_inst_44__empty_n;
  wire PE_inst_44__read;
  wire [32:0] PE_inst_44__din;
  wire PE_inst_44__full_n;
  wire PE_inst_44__write;
  wire [32:0] PE_inst_45__dout;
  wire PE_inst_45__empty_n;
  wire PE_inst_45__read;
  wire [32:0] PE_inst_45__din;
  wire PE_inst_45__full_n;
  wire PE_inst_45__write;
  wire [32:0] PE_inst_46__dout;
  wire PE_inst_46__empty_n;
  wire PE_inst_46__read;
  wire [32:0] PE_inst_46__din;
  wire PE_inst_46__full_n;
  wire PE_inst_46__write;
  wire [32:0] PE_inst_47__dout;
  wire PE_inst_47__empty_n;
  wire PE_inst_47__read;
  wire [32:0] PE_inst_47__din;
  wire PE_inst_47__full_n;
  wire PE_inst_47__write;
  wire [32:0] PE_inst_48__dout;
  wire PE_inst_48__empty_n;
  wire PE_inst_48__read;
  wire [32:0] PE_inst_48__din;
  wire PE_inst_48__full_n;
  wire PE_inst_48__write;
  wire [32:0] PE_inst_4__dout;
  wire PE_inst_4__empty_n;
  wire PE_inst_4__read;
  wire [32:0] PE_inst_4__din;
  wire PE_inst_4__full_n;
  wire PE_inst_4__write;
  wire [32:0] PE_inst_5__dout;
  wire PE_inst_5__empty_n;
  wire PE_inst_5__read;
  wire [32:0] PE_inst_5__din;
  wire PE_inst_5__full_n;
  wire PE_inst_5__write;
  wire [32:0] PE_inst_6__dout;
  wire PE_inst_6__empty_n;
  wire PE_inst_6__read;
  wire [32:0] PE_inst_6__din;
  wire PE_inst_6__full_n;
  wire PE_inst_6__write;
  wire [32:0] PE_inst_7__dout;
  wire PE_inst_7__empty_n;
  wire PE_inst_7__read;
  wire [32:0] PE_inst_7__din;
  wire PE_inst_7__full_n;
  wire PE_inst_7__write;
  wire [32:0] PE_inst_8__dout;
  wire PE_inst_8__empty_n;
  wire PE_inst_8__read;
  wire [32:0] PE_inst_8__din;
  wire PE_inst_8__full_n;
  wire PE_inst_8__write;
  wire [32:0] PE_inst_9__dout;
  wire PE_inst_9__empty_n;
  wire PE_inst_9__read;
  wire [32:0] PE_inst_9__din;
  wire PE_inst_9__full_n;
  wire PE_inst_9__write;
  wire [32:0] Yvec_inst_0__dout;
  wire Yvec_inst_0__empty_n;
  wire Yvec_inst_0__read;
  wire [32:0] Yvec_inst_0__din;
  wire Yvec_inst_0__full_n;
  wire Yvec_inst_0__write;
  wire [32:0] Yvec_inst_10__dout;
  wire Yvec_inst_10__empty_n;
  wire Yvec_inst_10__read;
  wire [32:0] Yvec_inst_10__din;
  wire Yvec_inst_10__full_n;
  wire Yvec_inst_10__write;
  wire [32:0] Yvec_inst_11__dout;
  wire Yvec_inst_11__empty_n;
  wire Yvec_inst_11__read;
  wire [32:0] Yvec_inst_11__din;
  wire Yvec_inst_11__full_n;
  wire Yvec_inst_11__write;
  wire [32:0] Yvec_inst_12__dout;
  wire Yvec_inst_12__empty_n;
  wire Yvec_inst_12__read;
  wire [32:0] Yvec_inst_12__din;
  wire Yvec_inst_12__full_n;
  wire Yvec_inst_12__write;
  wire [32:0] Yvec_inst_13__dout;
  wire Yvec_inst_13__empty_n;
  wire Yvec_inst_13__read;
  wire [32:0] Yvec_inst_13__din;
  wire Yvec_inst_13__full_n;
  wire Yvec_inst_13__write;
  wire [32:0] Yvec_inst_14__dout;
  wire Yvec_inst_14__empty_n;
  wire Yvec_inst_14__read;
  wire [32:0] Yvec_inst_14__din;
  wire Yvec_inst_14__full_n;
  wire Yvec_inst_14__write;
  wire [32:0] Yvec_inst_15__dout;
  wire Yvec_inst_15__empty_n;
  wire Yvec_inst_15__read;
  wire [32:0] Yvec_inst_15__din;
  wire Yvec_inst_15__full_n;
  wire Yvec_inst_15__write;
  wire [32:0] Yvec_inst_16__dout;
  wire Yvec_inst_16__empty_n;
  wire Yvec_inst_16__read;
  wire [32:0] Yvec_inst_16__din;
  wire Yvec_inst_16__full_n;
  wire Yvec_inst_16__write;
  wire [32:0] Yvec_inst_17__dout;
  wire Yvec_inst_17__empty_n;
  wire Yvec_inst_17__read;
  wire [32:0] Yvec_inst_17__din;
  wire Yvec_inst_17__full_n;
  wire Yvec_inst_17__write;
  wire [32:0] Yvec_inst_18__dout;
  wire Yvec_inst_18__empty_n;
  wire Yvec_inst_18__read;
  wire [32:0] Yvec_inst_18__din;
  wire Yvec_inst_18__full_n;
  wire Yvec_inst_18__write;
  wire [32:0] Yvec_inst_19__dout;
  wire Yvec_inst_19__empty_n;
  wire Yvec_inst_19__read;
  wire [32:0] Yvec_inst_19__din;
  wire Yvec_inst_19__full_n;
  wire Yvec_inst_19__write;
  wire [32:0] Yvec_inst_1__dout;
  wire Yvec_inst_1__empty_n;
  wire Yvec_inst_1__read;
  wire [32:0] Yvec_inst_1__din;
  wire Yvec_inst_1__full_n;
  wire Yvec_inst_1__write;
  wire [32:0] Yvec_inst_20__dout;
  wire Yvec_inst_20__empty_n;
  wire Yvec_inst_20__read;
  wire [32:0] Yvec_inst_20__din;
  wire Yvec_inst_20__full_n;
  wire Yvec_inst_20__write;
  wire [32:0] Yvec_inst_21__dout;
  wire Yvec_inst_21__empty_n;
  wire Yvec_inst_21__read;
  wire [32:0] Yvec_inst_21__din;
  wire Yvec_inst_21__full_n;
  wire Yvec_inst_21__write;
  wire [32:0] Yvec_inst_22__dout;
  wire Yvec_inst_22__empty_n;
  wire Yvec_inst_22__read;
  wire [32:0] Yvec_inst_22__din;
  wire Yvec_inst_22__full_n;
  wire Yvec_inst_22__write;
  wire [32:0] Yvec_inst_23__dout;
  wire Yvec_inst_23__empty_n;
  wire Yvec_inst_23__read;
  wire [32:0] Yvec_inst_23__din;
  wire Yvec_inst_23__full_n;
  wire Yvec_inst_23__write;
  wire [32:0] Yvec_inst_24__dout;
  wire Yvec_inst_24__empty_n;
  wire Yvec_inst_24__read;
  wire [32:0] Yvec_inst_24__din;
  wire Yvec_inst_24__full_n;
  wire Yvec_inst_24__write;
  wire [32:0] Yvec_inst_25__dout;
  wire Yvec_inst_25__empty_n;
  wire Yvec_inst_25__read;
  wire [32:0] Yvec_inst_25__din;
  wire Yvec_inst_25__full_n;
  wire Yvec_inst_25__write;
  wire [32:0] Yvec_inst_26__dout;
  wire Yvec_inst_26__empty_n;
  wire Yvec_inst_26__read;
  wire [32:0] Yvec_inst_26__din;
  wire Yvec_inst_26__full_n;
  wire Yvec_inst_26__write;
  wire [32:0] Yvec_inst_27__dout;
  wire Yvec_inst_27__empty_n;
  wire Yvec_inst_27__read;
  wire [32:0] Yvec_inst_27__din;
  wire Yvec_inst_27__full_n;
  wire Yvec_inst_27__write;
  wire [32:0] Yvec_inst_28__dout;
  wire Yvec_inst_28__empty_n;
  wire Yvec_inst_28__read;
  wire [32:0] Yvec_inst_28__din;
  wire Yvec_inst_28__full_n;
  wire Yvec_inst_28__write;
  wire [32:0] Yvec_inst_29__dout;
  wire Yvec_inst_29__empty_n;
  wire Yvec_inst_29__read;
  wire [32:0] Yvec_inst_29__din;
  wire Yvec_inst_29__full_n;
  wire Yvec_inst_29__write;
  wire [32:0] Yvec_inst_2__dout;
  wire Yvec_inst_2__empty_n;
  wire Yvec_inst_2__read;
  wire [32:0] Yvec_inst_2__din;
  wire Yvec_inst_2__full_n;
  wire Yvec_inst_2__write;
  wire [32:0] Yvec_inst_30__dout;
  wire Yvec_inst_30__empty_n;
  wire Yvec_inst_30__read;
  wire [32:0] Yvec_inst_30__din;
  wire Yvec_inst_30__full_n;
  wire Yvec_inst_30__write;
  wire [32:0] Yvec_inst_31__dout;
  wire Yvec_inst_31__empty_n;
  wire Yvec_inst_31__read;
  wire [32:0] Yvec_inst_31__din;
  wire Yvec_inst_31__full_n;
  wire Yvec_inst_31__write;
  wire [32:0] Yvec_inst_32__dout;
  wire Yvec_inst_32__empty_n;
  wire Yvec_inst_32__read;
  wire [32:0] Yvec_inst_32__din;
  wire Yvec_inst_32__full_n;
  wire Yvec_inst_32__write;
  wire [32:0] Yvec_inst_33__dout;
  wire Yvec_inst_33__empty_n;
  wire Yvec_inst_33__read;
  wire [32:0] Yvec_inst_33__din;
  wire Yvec_inst_33__full_n;
  wire Yvec_inst_33__write;
  wire [32:0] Yvec_inst_34__dout;
  wire Yvec_inst_34__empty_n;
  wire Yvec_inst_34__read;
  wire [32:0] Yvec_inst_34__din;
  wire Yvec_inst_34__full_n;
  wire Yvec_inst_34__write;
  wire [32:0] Yvec_inst_35__dout;
  wire Yvec_inst_35__empty_n;
  wire Yvec_inst_35__read;
  wire [32:0] Yvec_inst_35__din;
  wire Yvec_inst_35__full_n;
  wire Yvec_inst_35__write;
  wire [32:0] Yvec_inst_36__dout;
  wire Yvec_inst_36__empty_n;
  wire Yvec_inst_36__read;
  wire [32:0] Yvec_inst_36__din;
  wire Yvec_inst_36__full_n;
  wire Yvec_inst_36__write;
  wire [32:0] Yvec_inst_37__dout;
  wire Yvec_inst_37__empty_n;
  wire Yvec_inst_37__read;
  wire [32:0] Yvec_inst_37__din;
  wire Yvec_inst_37__full_n;
  wire Yvec_inst_37__write;
  wire [32:0] Yvec_inst_38__dout;
  wire Yvec_inst_38__empty_n;
  wire Yvec_inst_38__read;
  wire [32:0] Yvec_inst_38__din;
  wire Yvec_inst_38__full_n;
  wire Yvec_inst_38__write;
  wire [32:0] Yvec_inst_39__dout;
  wire Yvec_inst_39__empty_n;
  wire Yvec_inst_39__read;
  wire [32:0] Yvec_inst_39__din;
  wire Yvec_inst_39__full_n;
  wire Yvec_inst_39__write;
  wire [32:0] Yvec_inst_3__dout;
  wire Yvec_inst_3__empty_n;
  wire Yvec_inst_3__read;
  wire [32:0] Yvec_inst_3__din;
  wire Yvec_inst_3__full_n;
  wire Yvec_inst_3__write;
  wire [32:0] Yvec_inst_40__dout;
  wire Yvec_inst_40__empty_n;
  wire Yvec_inst_40__read;
  wire [32:0] Yvec_inst_40__din;
  wire Yvec_inst_40__full_n;
  wire Yvec_inst_40__write;
  wire [32:0] Yvec_inst_41__dout;
  wire Yvec_inst_41__empty_n;
  wire Yvec_inst_41__read;
  wire [32:0] Yvec_inst_41__din;
  wire Yvec_inst_41__full_n;
  wire Yvec_inst_41__write;
  wire [32:0] Yvec_inst_42__dout;
  wire Yvec_inst_42__empty_n;
  wire Yvec_inst_42__read;
  wire [32:0] Yvec_inst_42__din;
  wire Yvec_inst_42__full_n;
  wire Yvec_inst_42__write;
  wire [32:0] Yvec_inst_43__dout;
  wire Yvec_inst_43__empty_n;
  wire Yvec_inst_43__read;
  wire [32:0] Yvec_inst_43__din;
  wire Yvec_inst_43__full_n;
  wire Yvec_inst_43__write;
  wire [32:0] Yvec_inst_44__dout;
  wire Yvec_inst_44__empty_n;
  wire Yvec_inst_44__read;
  wire [32:0] Yvec_inst_44__din;
  wire Yvec_inst_44__full_n;
  wire Yvec_inst_44__write;
  wire [32:0] Yvec_inst_45__dout;
  wire Yvec_inst_45__empty_n;
  wire Yvec_inst_45__read;
  wire [32:0] Yvec_inst_45__din;
  wire Yvec_inst_45__full_n;
  wire Yvec_inst_45__write;
  wire [32:0] Yvec_inst_46__dout;
  wire Yvec_inst_46__empty_n;
  wire Yvec_inst_46__read;
  wire [32:0] Yvec_inst_46__din;
  wire Yvec_inst_46__full_n;
  wire Yvec_inst_46__write;
  wire [32:0] Yvec_inst_47__dout;
  wire Yvec_inst_47__empty_n;
  wire Yvec_inst_47__read;
  wire [32:0] Yvec_inst_47__din;
  wire Yvec_inst_47__full_n;
  wire Yvec_inst_47__write;
  wire [32:0] Yvec_inst_4__dout;
  wire Yvec_inst_4__empty_n;
  wire Yvec_inst_4__read;
  wire [32:0] Yvec_inst_4__din;
  wire Yvec_inst_4__full_n;
  wire Yvec_inst_4__write;
  wire [32:0] Yvec_inst_5__dout;
  wire Yvec_inst_5__empty_n;
  wire Yvec_inst_5__read;
  wire [32:0] Yvec_inst_5__din;
  wire Yvec_inst_5__full_n;
  wire Yvec_inst_5__write;
  wire [32:0] Yvec_inst_6__dout;
  wire Yvec_inst_6__empty_n;
  wire Yvec_inst_6__read;
  wire [32:0] Yvec_inst_6__din;
  wire Yvec_inst_6__full_n;
  wire Yvec_inst_6__write;
  wire [32:0] Yvec_inst_7__dout;
  wire Yvec_inst_7__empty_n;
  wire Yvec_inst_7__read;
  wire [32:0] Yvec_inst_7__din;
  wire Yvec_inst_7__full_n;
  wire Yvec_inst_7__write;
  wire [32:0] Yvec_inst_8__dout;
  wire Yvec_inst_8__empty_n;
  wire Yvec_inst_8__read;
  wire [32:0] Yvec_inst_8__din;
  wire Yvec_inst_8__full_n;
  wire Yvec_inst_8__write;
  wire [32:0] Yvec_inst_9__dout;
  wire Yvec_inst_9__empty_n;
  wire Yvec_inst_9__read;
  wire [32:0] Yvec_inst_9__din;
  wire Yvec_inst_9__full_n;
  wire Yvec_inst_9__write;
  wire [512:0] fifo_A_0__dout;
  wire fifo_A_0__empty_n;
  wire fifo_A_0__read;
  wire [512:0] fifo_A_0__din;
  wire fifo_A_0__full_n;
  wire fifo_A_0__write;
  wire [512:0] fifo_A_10__dout;
  wire fifo_A_10__empty_n;
  wire fifo_A_10__read;
  wire [512:0] fifo_A_10__din;
  wire fifo_A_10__full_n;
  wire fifo_A_10__write;
  wire [512:0] fifo_A_11__dout;
  wire fifo_A_11__empty_n;
  wire fifo_A_11__read;
  wire [512:0] fifo_A_11__din;
  wire fifo_A_11__full_n;
  wire fifo_A_11__write;
  wire [512:0] fifo_A_12__dout;
  wire fifo_A_12__empty_n;
  wire fifo_A_12__read;
  wire [512:0] fifo_A_12__din;
  wire fifo_A_12__full_n;
  wire fifo_A_12__write;
  wire [512:0] fifo_A_13__dout;
  wire fifo_A_13__empty_n;
  wire fifo_A_13__read;
  wire [512:0] fifo_A_13__din;
  wire fifo_A_13__full_n;
  wire fifo_A_13__write;
  wire [512:0] fifo_A_14__dout;
  wire fifo_A_14__empty_n;
  wire fifo_A_14__read;
  wire [512:0] fifo_A_14__din;
  wire fifo_A_14__full_n;
  wire fifo_A_14__write;
  wire [512:0] fifo_A_15__dout;
  wire fifo_A_15__empty_n;
  wire fifo_A_15__read;
  wire [512:0] fifo_A_15__din;
  wire fifo_A_15__full_n;
  wire fifo_A_15__write;
  wire [512:0] fifo_A_16__dout;
  wire fifo_A_16__empty_n;
  wire fifo_A_16__read;
  wire [512:0] fifo_A_16__din;
  wire fifo_A_16__full_n;
  wire fifo_A_16__write;
  wire [512:0] fifo_A_17__dout;
  wire fifo_A_17__empty_n;
  wire fifo_A_17__read;
  wire [512:0] fifo_A_17__din;
  wire fifo_A_17__full_n;
  wire fifo_A_17__write;
  wire [512:0] fifo_A_18__dout;
  wire fifo_A_18__empty_n;
  wire fifo_A_18__read;
  wire [512:0] fifo_A_18__din;
  wire fifo_A_18__full_n;
  wire fifo_A_18__write;
  wire [512:0] fifo_A_19__dout;
  wire fifo_A_19__empty_n;
  wire fifo_A_19__read;
  wire [512:0] fifo_A_19__din;
  wire fifo_A_19__full_n;
  wire fifo_A_19__write;
  wire [512:0] fifo_A_1__dout;
  wire fifo_A_1__empty_n;
  wire fifo_A_1__read;
  wire [512:0] fifo_A_1__din;
  wire fifo_A_1__full_n;
  wire fifo_A_1__write;
  wire [512:0] fifo_A_20__dout;
  wire fifo_A_20__empty_n;
  wire fifo_A_20__read;
  wire [512:0] fifo_A_20__din;
  wire fifo_A_20__full_n;
  wire fifo_A_20__write;
  wire [512:0] fifo_A_21__dout;
  wire fifo_A_21__empty_n;
  wire fifo_A_21__read;
  wire [512:0] fifo_A_21__din;
  wire fifo_A_21__full_n;
  wire fifo_A_21__write;
  wire [512:0] fifo_A_22__dout;
  wire fifo_A_22__empty_n;
  wire fifo_A_22__read;
  wire [512:0] fifo_A_22__din;
  wire fifo_A_22__full_n;
  wire fifo_A_22__write;
  wire [512:0] fifo_A_23__dout;
  wire fifo_A_23__empty_n;
  wire fifo_A_23__read;
  wire [512:0] fifo_A_23__din;
  wire fifo_A_23__full_n;
  wire fifo_A_23__write;
  wire [512:0] fifo_A_24__dout;
  wire fifo_A_24__empty_n;
  wire fifo_A_24__read;
  wire [512:0] fifo_A_24__din;
  wire fifo_A_24__full_n;
  wire fifo_A_24__write;
  wire [512:0] fifo_A_25__dout;
  wire fifo_A_25__empty_n;
  wire fifo_A_25__read;
  wire [512:0] fifo_A_25__din;
  wire fifo_A_25__full_n;
  wire fifo_A_25__write;
  wire [512:0] fifo_A_26__dout;
  wire fifo_A_26__empty_n;
  wire fifo_A_26__read;
  wire [512:0] fifo_A_26__din;
  wire fifo_A_26__full_n;
  wire fifo_A_26__write;
  wire [512:0] fifo_A_27__dout;
  wire fifo_A_27__empty_n;
  wire fifo_A_27__read;
  wire [512:0] fifo_A_27__din;
  wire fifo_A_27__full_n;
  wire fifo_A_27__write;
  wire [512:0] fifo_A_28__dout;
  wire fifo_A_28__empty_n;
  wire fifo_A_28__read;
  wire [512:0] fifo_A_28__din;
  wire fifo_A_28__full_n;
  wire fifo_A_28__write;
  wire [512:0] fifo_A_29__dout;
  wire fifo_A_29__empty_n;
  wire fifo_A_29__read;
  wire [512:0] fifo_A_29__din;
  wire fifo_A_29__full_n;
  wire fifo_A_29__write;
  wire [512:0] fifo_A_2__dout;
  wire fifo_A_2__empty_n;
  wire fifo_A_2__read;
  wire [512:0] fifo_A_2__din;
  wire fifo_A_2__full_n;
  wire fifo_A_2__write;
  wire [512:0] fifo_A_30__dout;
  wire fifo_A_30__empty_n;
  wire fifo_A_30__read;
  wire [512:0] fifo_A_30__din;
  wire fifo_A_30__full_n;
  wire fifo_A_30__write;
  wire [512:0] fifo_A_31__dout;
  wire fifo_A_31__empty_n;
  wire fifo_A_31__read;
  wire [512:0] fifo_A_31__din;
  wire fifo_A_31__full_n;
  wire fifo_A_31__write;
  wire [512:0] fifo_A_32__dout;
  wire fifo_A_32__empty_n;
  wire fifo_A_32__read;
  wire [512:0] fifo_A_32__din;
  wire fifo_A_32__full_n;
  wire fifo_A_32__write;
  wire [512:0] fifo_A_33__dout;
  wire fifo_A_33__empty_n;
  wire fifo_A_33__read;
  wire [512:0] fifo_A_33__din;
  wire fifo_A_33__full_n;
  wire fifo_A_33__write;
  wire [512:0] fifo_A_34__dout;
  wire fifo_A_34__empty_n;
  wire fifo_A_34__read;
  wire [512:0] fifo_A_34__din;
  wire fifo_A_34__full_n;
  wire fifo_A_34__write;
  wire [512:0] fifo_A_35__dout;
  wire fifo_A_35__empty_n;
  wire fifo_A_35__read;
  wire [512:0] fifo_A_35__din;
  wire fifo_A_35__full_n;
  wire fifo_A_35__write;
  wire [512:0] fifo_A_36__dout;
  wire fifo_A_36__empty_n;
  wire fifo_A_36__read;
  wire [512:0] fifo_A_36__din;
  wire fifo_A_36__full_n;
  wire fifo_A_36__write;
  wire [512:0] fifo_A_37__dout;
  wire fifo_A_37__empty_n;
  wire fifo_A_37__read;
  wire [512:0] fifo_A_37__din;
  wire fifo_A_37__full_n;
  wire fifo_A_37__write;
  wire [512:0] fifo_A_38__dout;
  wire fifo_A_38__empty_n;
  wire fifo_A_38__read;
  wire [512:0] fifo_A_38__din;
  wire fifo_A_38__full_n;
  wire fifo_A_38__write;
  wire [512:0] fifo_A_39__dout;
  wire fifo_A_39__empty_n;
  wire fifo_A_39__read;
  wire [512:0] fifo_A_39__din;
  wire fifo_A_39__full_n;
  wire fifo_A_39__write;
  wire [512:0] fifo_A_3__dout;
  wire fifo_A_3__empty_n;
  wire fifo_A_3__read;
  wire [512:0] fifo_A_3__din;
  wire fifo_A_3__full_n;
  wire fifo_A_3__write;
  wire [512:0] fifo_A_40__dout;
  wire fifo_A_40__empty_n;
  wire fifo_A_40__read;
  wire [512:0] fifo_A_40__din;
  wire fifo_A_40__full_n;
  wire fifo_A_40__write;
  wire [512:0] fifo_A_41__dout;
  wire fifo_A_41__empty_n;
  wire fifo_A_41__read;
  wire [512:0] fifo_A_41__din;
  wire fifo_A_41__full_n;
  wire fifo_A_41__write;
  wire [512:0] fifo_A_42__dout;
  wire fifo_A_42__empty_n;
  wire fifo_A_42__read;
  wire [512:0] fifo_A_42__din;
  wire fifo_A_42__full_n;
  wire fifo_A_42__write;
  wire [512:0] fifo_A_43__dout;
  wire fifo_A_43__empty_n;
  wire fifo_A_43__read;
  wire [512:0] fifo_A_43__din;
  wire fifo_A_43__full_n;
  wire fifo_A_43__write;
  wire [512:0] fifo_A_44__dout;
  wire fifo_A_44__empty_n;
  wire fifo_A_44__read;
  wire [512:0] fifo_A_44__din;
  wire fifo_A_44__full_n;
  wire fifo_A_44__write;
  wire [512:0] fifo_A_45__dout;
  wire fifo_A_45__empty_n;
  wire fifo_A_45__read;
  wire [512:0] fifo_A_45__din;
  wire fifo_A_45__full_n;
  wire fifo_A_45__write;
  wire [512:0] fifo_A_46__dout;
  wire fifo_A_46__empty_n;
  wire fifo_A_46__read;
  wire [512:0] fifo_A_46__din;
  wire fifo_A_46__full_n;
  wire fifo_A_46__write;
  wire [512:0] fifo_A_47__dout;
  wire fifo_A_47__empty_n;
  wire fifo_A_47__read;
  wire [512:0] fifo_A_47__din;
  wire fifo_A_47__full_n;
  wire fifo_A_47__write;
  wire [512:0] fifo_A_4__dout;
  wire fifo_A_4__empty_n;
  wire fifo_A_4__read;
  wire [512:0] fifo_A_4__din;
  wire fifo_A_4__full_n;
  wire fifo_A_4__write;
  wire [512:0] fifo_A_5__dout;
  wire fifo_A_5__empty_n;
  wire fifo_A_5__read;
  wire [512:0] fifo_A_5__din;
  wire fifo_A_5__full_n;
  wire fifo_A_5__write;
  wire [512:0] fifo_A_6__dout;
  wire fifo_A_6__empty_n;
  wire fifo_A_6__read;
  wire [512:0] fifo_A_6__din;
  wire fifo_A_6__full_n;
  wire fifo_A_6__write;
  wire [512:0] fifo_A_7__dout;
  wire fifo_A_7__empty_n;
  wire fifo_A_7__read;
  wire [512:0] fifo_A_7__din;
  wire fifo_A_7__full_n;
  wire fifo_A_7__write;
  wire [512:0] fifo_A_8__dout;
  wire fifo_A_8__empty_n;
  wire fifo_A_8__read;
  wire [512:0] fifo_A_8__din;
  wire fifo_A_8__full_n;
  wire fifo_A_8__write;
  wire [512:0] fifo_A_9__dout;
  wire fifo_A_9__empty_n;
  wire fifo_A_9__read;
  wire [512:0] fifo_A_9__din;
  wire fifo_A_9__full_n;
  wire fifo_A_9__write;
  wire [512:0] fifo_X_pe_0__dout;
  wire fifo_X_pe_0__empty_n;
  wire fifo_X_pe_0__read;
  wire [512:0] fifo_X_pe_0__din;
  wire fifo_X_pe_0__full_n;
  wire fifo_X_pe_0__write;
  wire [512:0] fifo_X_pe_10__dout;
  wire fifo_X_pe_10__empty_n;
  wire fifo_X_pe_10__read;
  wire [512:0] fifo_X_pe_10__din;
  wire fifo_X_pe_10__full_n;
  wire fifo_X_pe_10__write;
  wire [512:0] fifo_X_pe_11__dout;
  wire fifo_X_pe_11__empty_n;
  wire fifo_X_pe_11__read;
  wire [512:0] fifo_X_pe_11__din;
  wire fifo_X_pe_11__full_n;
  wire fifo_X_pe_11__write;
  wire [512:0] fifo_X_pe_12__dout;
  wire fifo_X_pe_12__empty_n;
  wire fifo_X_pe_12__read;
  wire [512:0] fifo_X_pe_12__din;
  wire fifo_X_pe_12__full_n;
  wire fifo_X_pe_12__write;
  wire [512:0] fifo_X_pe_13__dout;
  wire fifo_X_pe_13__empty_n;
  wire fifo_X_pe_13__read;
  wire [512:0] fifo_X_pe_13__din;
  wire fifo_X_pe_13__full_n;
  wire fifo_X_pe_13__write;
  wire [512:0] fifo_X_pe_14__dout;
  wire fifo_X_pe_14__empty_n;
  wire fifo_X_pe_14__read;
  wire [512:0] fifo_X_pe_14__din;
  wire fifo_X_pe_14__full_n;
  wire fifo_X_pe_14__write;
  wire [512:0] fifo_X_pe_15__dout;
  wire fifo_X_pe_15__empty_n;
  wire fifo_X_pe_15__read;
  wire [512:0] fifo_X_pe_15__din;
  wire fifo_X_pe_15__full_n;
  wire fifo_X_pe_15__write;
  wire [512:0] fifo_X_pe_16__dout;
  wire fifo_X_pe_16__empty_n;
  wire fifo_X_pe_16__read;
  wire [512:0] fifo_X_pe_16__din;
  wire fifo_X_pe_16__full_n;
  wire fifo_X_pe_16__write;
  wire [512:0] fifo_X_pe_17__dout;
  wire fifo_X_pe_17__empty_n;
  wire fifo_X_pe_17__read;
  wire [512:0] fifo_X_pe_17__din;
  wire fifo_X_pe_17__full_n;
  wire fifo_X_pe_17__write;
  wire [512:0] fifo_X_pe_18__dout;
  wire fifo_X_pe_18__empty_n;
  wire fifo_X_pe_18__read;
  wire [512:0] fifo_X_pe_18__din;
  wire fifo_X_pe_18__full_n;
  wire fifo_X_pe_18__write;
  wire [512:0] fifo_X_pe_19__dout;
  wire fifo_X_pe_19__empty_n;
  wire fifo_X_pe_19__read;
  wire [512:0] fifo_X_pe_19__din;
  wire fifo_X_pe_19__full_n;
  wire fifo_X_pe_19__write;
  wire [512:0] fifo_X_pe_1__dout;
  wire fifo_X_pe_1__empty_n;
  wire fifo_X_pe_1__read;
  wire [512:0] fifo_X_pe_1__din;
  wire fifo_X_pe_1__full_n;
  wire fifo_X_pe_1__write;
  wire [512:0] fifo_X_pe_20__dout;
  wire fifo_X_pe_20__empty_n;
  wire fifo_X_pe_20__read;
  wire [512:0] fifo_X_pe_20__din;
  wire fifo_X_pe_20__full_n;
  wire fifo_X_pe_20__write;
  wire [512:0] fifo_X_pe_21__dout;
  wire fifo_X_pe_21__empty_n;
  wire fifo_X_pe_21__read;
  wire [512:0] fifo_X_pe_21__din;
  wire fifo_X_pe_21__full_n;
  wire fifo_X_pe_21__write;
  wire [512:0] fifo_X_pe_22__dout;
  wire fifo_X_pe_22__empty_n;
  wire fifo_X_pe_22__read;
  wire [512:0] fifo_X_pe_22__din;
  wire fifo_X_pe_22__full_n;
  wire fifo_X_pe_22__write;
  wire [512:0] fifo_X_pe_23__dout;
  wire fifo_X_pe_23__empty_n;
  wire fifo_X_pe_23__read;
  wire [512:0] fifo_X_pe_23__din;
  wire fifo_X_pe_23__full_n;
  wire fifo_X_pe_23__write;
  wire [512:0] fifo_X_pe_24__dout;
  wire fifo_X_pe_24__empty_n;
  wire fifo_X_pe_24__read;
  wire [512:0] fifo_X_pe_24__din;
  wire fifo_X_pe_24__full_n;
  wire fifo_X_pe_24__write;
  wire [512:0] fifo_X_pe_25__dout;
  wire fifo_X_pe_25__empty_n;
  wire fifo_X_pe_25__read;
  wire [512:0] fifo_X_pe_25__din;
  wire fifo_X_pe_25__full_n;
  wire fifo_X_pe_25__write;
  wire [512:0] fifo_X_pe_26__dout;
  wire fifo_X_pe_26__empty_n;
  wire fifo_X_pe_26__read;
  wire [512:0] fifo_X_pe_26__din;
  wire fifo_X_pe_26__full_n;
  wire fifo_X_pe_26__write;
  wire [512:0] fifo_X_pe_27__dout;
  wire fifo_X_pe_27__empty_n;
  wire fifo_X_pe_27__read;
  wire [512:0] fifo_X_pe_27__din;
  wire fifo_X_pe_27__full_n;
  wire fifo_X_pe_27__write;
  wire [512:0] fifo_X_pe_28__dout;
  wire fifo_X_pe_28__empty_n;
  wire fifo_X_pe_28__read;
  wire [512:0] fifo_X_pe_28__din;
  wire fifo_X_pe_28__full_n;
  wire fifo_X_pe_28__write;
  wire [512:0] fifo_X_pe_29__dout;
  wire fifo_X_pe_29__empty_n;
  wire fifo_X_pe_29__read;
  wire [512:0] fifo_X_pe_29__din;
  wire fifo_X_pe_29__full_n;
  wire fifo_X_pe_29__write;
  wire [512:0] fifo_X_pe_2__dout;
  wire fifo_X_pe_2__empty_n;
  wire fifo_X_pe_2__read;
  wire [512:0] fifo_X_pe_2__din;
  wire fifo_X_pe_2__full_n;
  wire fifo_X_pe_2__write;
  wire [512:0] fifo_X_pe_30__dout;
  wire fifo_X_pe_30__empty_n;
  wire fifo_X_pe_30__read;
  wire [512:0] fifo_X_pe_30__din;
  wire fifo_X_pe_30__full_n;
  wire fifo_X_pe_30__write;
  wire [512:0] fifo_X_pe_31__dout;
  wire fifo_X_pe_31__empty_n;
  wire fifo_X_pe_31__read;
  wire [512:0] fifo_X_pe_31__din;
  wire fifo_X_pe_31__full_n;
  wire fifo_X_pe_31__write;
  wire [512:0] fifo_X_pe_32__dout;
  wire fifo_X_pe_32__empty_n;
  wire fifo_X_pe_32__read;
  wire [512:0] fifo_X_pe_32__din;
  wire fifo_X_pe_32__full_n;
  wire fifo_X_pe_32__write;
  wire [512:0] fifo_X_pe_33__dout;
  wire fifo_X_pe_33__empty_n;
  wire fifo_X_pe_33__read;
  wire [512:0] fifo_X_pe_33__din;
  wire fifo_X_pe_33__full_n;
  wire fifo_X_pe_33__write;
  wire [512:0] fifo_X_pe_34__dout;
  wire fifo_X_pe_34__empty_n;
  wire fifo_X_pe_34__read;
  wire [512:0] fifo_X_pe_34__din;
  wire fifo_X_pe_34__full_n;
  wire fifo_X_pe_34__write;
  wire [512:0] fifo_X_pe_35__dout;
  wire fifo_X_pe_35__empty_n;
  wire fifo_X_pe_35__read;
  wire [512:0] fifo_X_pe_35__din;
  wire fifo_X_pe_35__full_n;
  wire fifo_X_pe_35__write;
  wire [512:0] fifo_X_pe_36__dout;
  wire fifo_X_pe_36__empty_n;
  wire fifo_X_pe_36__read;
  wire [512:0] fifo_X_pe_36__din;
  wire fifo_X_pe_36__full_n;
  wire fifo_X_pe_36__write;
  wire [512:0] fifo_X_pe_37__dout;
  wire fifo_X_pe_37__empty_n;
  wire fifo_X_pe_37__read;
  wire [512:0] fifo_X_pe_37__din;
  wire fifo_X_pe_37__full_n;
  wire fifo_X_pe_37__write;
  wire [512:0] fifo_X_pe_38__dout;
  wire fifo_X_pe_38__empty_n;
  wire fifo_X_pe_38__read;
  wire [512:0] fifo_X_pe_38__din;
  wire fifo_X_pe_38__full_n;
  wire fifo_X_pe_38__write;
  wire [512:0] fifo_X_pe_39__dout;
  wire fifo_X_pe_39__empty_n;
  wire fifo_X_pe_39__read;
  wire [512:0] fifo_X_pe_39__din;
  wire fifo_X_pe_39__full_n;
  wire fifo_X_pe_39__write;
  wire [512:0] fifo_X_pe_3__dout;
  wire fifo_X_pe_3__empty_n;
  wire fifo_X_pe_3__read;
  wire [512:0] fifo_X_pe_3__din;
  wire fifo_X_pe_3__full_n;
  wire fifo_X_pe_3__write;
  wire [512:0] fifo_X_pe_40__dout;
  wire fifo_X_pe_40__empty_n;
  wire fifo_X_pe_40__read;
  wire [512:0] fifo_X_pe_40__din;
  wire fifo_X_pe_40__full_n;
  wire fifo_X_pe_40__write;
  wire [512:0] fifo_X_pe_41__dout;
  wire fifo_X_pe_41__empty_n;
  wire fifo_X_pe_41__read;
  wire [512:0] fifo_X_pe_41__din;
  wire fifo_X_pe_41__full_n;
  wire fifo_X_pe_41__write;
  wire [512:0] fifo_X_pe_42__dout;
  wire fifo_X_pe_42__empty_n;
  wire fifo_X_pe_42__read;
  wire [512:0] fifo_X_pe_42__din;
  wire fifo_X_pe_42__full_n;
  wire fifo_X_pe_42__write;
  wire [512:0] fifo_X_pe_43__dout;
  wire fifo_X_pe_43__empty_n;
  wire fifo_X_pe_43__read;
  wire [512:0] fifo_X_pe_43__din;
  wire fifo_X_pe_43__full_n;
  wire fifo_X_pe_43__write;
  wire [512:0] fifo_X_pe_44__dout;
  wire fifo_X_pe_44__empty_n;
  wire fifo_X_pe_44__read;
  wire [512:0] fifo_X_pe_44__din;
  wire fifo_X_pe_44__full_n;
  wire fifo_X_pe_44__write;
  wire [512:0] fifo_X_pe_45__dout;
  wire fifo_X_pe_45__empty_n;
  wire fifo_X_pe_45__read;
  wire [512:0] fifo_X_pe_45__din;
  wire fifo_X_pe_45__full_n;
  wire fifo_X_pe_45__write;
  wire [512:0] fifo_X_pe_46__dout;
  wire fifo_X_pe_46__empty_n;
  wire fifo_X_pe_46__read;
  wire [512:0] fifo_X_pe_46__din;
  wire fifo_X_pe_46__full_n;
  wire fifo_X_pe_46__write;
  wire [512:0] fifo_X_pe_47__dout;
  wire fifo_X_pe_47__empty_n;
  wire fifo_X_pe_47__read;
  wire [512:0] fifo_X_pe_47__din;
  wire fifo_X_pe_47__full_n;
  wire fifo_X_pe_47__write;
  wire [512:0] fifo_X_pe_48__dout;
  wire fifo_X_pe_48__empty_n;
  wire fifo_X_pe_48__read;
  wire [512:0] fifo_X_pe_48__din;
  wire fifo_X_pe_48__full_n;
  wire fifo_X_pe_48__write;
  wire [512:0] fifo_X_pe_4__dout;
  wire fifo_X_pe_4__empty_n;
  wire fifo_X_pe_4__read;
  wire [512:0] fifo_X_pe_4__din;
  wire fifo_X_pe_4__full_n;
  wire fifo_X_pe_4__write;
  wire [512:0] fifo_X_pe_5__dout;
  wire fifo_X_pe_5__empty_n;
  wire fifo_X_pe_5__read;
  wire [512:0] fifo_X_pe_5__din;
  wire fifo_X_pe_5__full_n;
  wire fifo_X_pe_5__write;
  wire [512:0] fifo_X_pe_6__dout;
  wire fifo_X_pe_6__empty_n;
  wire fifo_X_pe_6__read;
  wire [512:0] fifo_X_pe_6__din;
  wire fifo_X_pe_6__full_n;
  wire fifo_X_pe_6__write;
  wire [512:0] fifo_X_pe_7__dout;
  wire fifo_X_pe_7__empty_n;
  wire fifo_X_pe_7__read;
  wire [512:0] fifo_X_pe_7__din;
  wire fifo_X_pe_7__full_n;
  wire fifo_X_pe_7__write;
  wire [512:0] fifo_X_pe_8__dout;
  wire fifo_X_pe_8__empty_n;
  wire fifo_X_pe_8__read;
  wire [512:0] fifo_X_pe_8__din;
  wire fifo_X_pe_8__full_n;
  wire fifo_X_pe_8__write;
  wire [512:0] fifo_X_pe_9__dout;
  wire fifo_X_pe_9__empty_n;
  wire fifo_X_pe_9__read;
  wire [512:0] fifo_X_pe_9__din;
  wire fifo_X_pe_9__full_n;
  wire fifo_X_pe_9__write;
  wire [512:0] fifo_Y_AX__dout;
  wire fifo_Y_AX__empty_n;
  wire fifo_Y_AX__read;
  wire [512:0] fifo_Y_AX__din;
  wire fifo_Y_AX__full_n;
  wire fifo_Y_AX__write;
  wire [512:0] fifo_Y_alpha_AX__dout;
  wire fifo_Y_alpha_AX__empty_n;
  wire fifo_Y_alpha_AX__read;
  wire [512:0] fifo_Y_alpha_AX__din;
  wire fifo_Y_alpha_AX__full_n;
  wire fifo_Y_alpha_AX__write;
  wire [512:0] fifo_Y_in__dout;
  wire fifo_Y_in__empty_n;
  wire fifo_Y_in__read;
  wire [512:0] fifo_Y_in__din;
  wire fifo_Y_in__full_n;
  wire fifo_Y_in__write;
  wire [512:0] fifo_Y_in_beta__dout;
  wire fifo_Y_in_beta__empty_n;
  wire fifo_Y_in_beta__read;
  wire [512:0] fifo_Y_in_beta__din;
  wire fifo_Y_in_beta__full_n;
  wire fifo_Y_in_beta__write;
  wire [512:0] fifo_Y_out__dout;
  wire fifo_Y_out__empty_n;
  wire fifo_Y_out__read;
  wire [512:0] fifo_Y_out__din;
  wire fifo_Y_out__full_n;
  wire fifo_Y_out__write;
  wire [64:0] fifo_Y_pe_0__dout;
  wire fifo_Y_pe_0__empty_n;
  wire fifo_Y_pe_0__read;
  wire [64:0] fifo_Y_pe_0__din;
  wire fifo_Y_pe_0__full_n;
  wire fifo_Y_pe_0__write;
  wire [64:0] fifo_Y_pe_10__dout;
  wire fifo_Y_pe_10__empty_n;
  wire fifo_Y_pe_10__read;
  wire [64:0] fifo_Y_pe_10__din;
  wire fifo_Y_pe_10__full_n;
  wire fifo_Y_pe_10__write;
  wire [64:0] fifo_Y_pe_11__dout;
  wire fifo_Y_pe_11__empty_n;
  wire fifo_Y_pe_11__read;
  wire [64:0] fifo_Y_pe_11__din;
  wire fifo_Y_pe_11__full_n;
  wire fifo_Y_pe_11__write;
  wire [64:0] fifo_Y_pe_12__dout;
  wire fifo_Y_pe_12__empty_n;
  wire fifo_Y_pe_12__read;
  wire [64:0] fifo_Y_pe_12__din;
  wire fifo_Y_pe_12__full_n;
  wire fifo_Y_pe_12__write;
  wire [64:0] fifo_Y_pe_13__dout;
  wire fifo_Y_pe_13__empty_n;
  wire fifo_Y_pe_13__read;
  wire [64:0] fifo_Y_pe_13__din;
  wire fifo_Y_pe_13__full_n;
  wire fifo_Y_pe_13__write;
  wire [64:0] fifo_Y_pe_14__dout;
  wire fifo_Y_pe_14__empty_n;
  wire fifo_Y_pe_14__read;
  wire [64:0] fifo_Y_pe_14__din;
  wire fifo_Y_pe_14__full_n;
  wire fifo_Y_pe_14__write;
  wire [64:0] fifo_Y_pe_15__dout;
  wire fifo_Y_pe_15__empty_n;
  wire fifo_Y_pe_15__read;
  wire [64:0] fifo_Y_pe_15__din;
  wire fifo_Y_pe_15__full_n;
  wire fifo_Y_pe_15__write;
  wire [64:0] fifo_Y_pe_16__dout;
  wire fifo_Y_pe_16__empty_n;
  wire fifo_Y_pe_16__read;
  wire [64:0] fifo_Y_pe_16__din;
  wire fifo_Y_pe_16__full_n;
  wire fifo_Y_pe_16__write;
  wire [64:0] fifo_Y_pe_17__dout;
  wire fifo_Y_pe_17__empty_n;
  wire fifo_Y_pe_17__read;
  wire [64:0] fifo_Y_pe_17__din;
  wire fifo_Y_pe_17__full_n;
  wire fifo_Y_pe_17__write;
  wire [64:0] fifo_Y_pe_18__dout;
  wire fifo_Y_pe_18__empty_n;
  wire fifo_Y_pe_18__read;
  wire [64:0] fifo_Y_pe_18__din;
  wire fifo_Y_pe_18__full_n;
  wire fifo_Y_pe_18__write;
  wire [64:0] fifo_Y_pe_19__dout;
  wire fifo_Y_pe_19__empty_n;
  wire fifo_Y_pe_19__read;
  wire [64:0] fifo_Y_pe_19__din;
  wire fifo_Y_pe_19__full_n;
  wire fifo_Y_pe_19__write;
  wire [64:0] fifo_Y_pe_1__dout;
  wire fifo_Y_pe_1__empty_n;
  wire fifo_Y_pe_1__read;
  wire [64:0] fifo_Y_pe_1__din;
  wire fifo_Y_pe_1__full_n;
  wire fifo_Y_pe_1__write;
  wire [64:0] fifo_Y_pe_20__dout;
  wire fifo_Y_pe_20__empty_n;
  wire fifo_Y_pe_20__read;
  wire [64:0] fifo_Y_pe_20__din;
  wire fifo_Y_pe_20__full_n;
  wire fifo_Y_pe_20__write;
  wire [64:0] fifo_Y_pe_21__dout;
  wire fifo_Y_pe_21__empty_n;
  wire fifo_Y_pe_21__read;
  wire [64:0] fifo_Y_pe_21__din;
  wire fifo_Y_pe_21__full_n;
  wire fifo_Y_pe_21__write;
  wire [64:0] fifo_Y_pe_22__dout;
  wire fifo_Y_pe_22__empty_n;
  wire fifo_Y_pe_22__read;
  wire [64:0] fifo_Y_pe_22__din;
  wire fifo_Y_pe_22__full_n;
  wire fifo_Y_pe_22__write;
  wire [64:0] fifo_Y_pe_23__dout;
  wire fifo_Y_pe_23__empty_n;
  wire fifo_Y_pe_23__read;
  wire [64:0] fifo_Y_pe_23__din;
  wire fifo_Y_pe_23__full_n;
  wire fifo_Y_pe_23__write;
  wire [64:0] fifo_Y_pe_24__dout;
  wire fifo_Y_pe_24__empty_n;
  wire fifo_Y_pe_24__read;
  wire [64:0] fifo_Y_pe_24__din;
  wire fifo_Y_pe_24__full_n;
  wire fifo_Y_pe_24__write;
  wire [64:0] fifo_Y_pe_25__dout;
  wire fifo_Y_pe_25__empty_n;
  wire fifo_Y_pe_25__read;
  wire [64:0] fifo_Y_pe_25__din;
  wire fifo_Y_pe_25__full_n;
  wire fifo_Y_pe_25__write;
  wire [64:0] fifo_Y_pe_26__dout;
  wire fifo_Y_pe_26__empty_n;
  wire fifo_Y_pe_26__read;
  wire [64:0] fifo_Y_pe_26__din;
  wire fifo_Y_pe_26__full_n;
  wire fifo_Y_pe_26__write;
  wire [64:0] fifo_Y_pe_27__dout;
  wire fifo_Y_pe_27__empty_n;
  wire fifo_Y_pe_27__read;
  wire [64:0] fifo_Y_pe_27__din;
  wire fifo_Y_pe_27__full_n;
  wire fifo_Y_pe_27__write;
  wire [64:0] fifo_Y_pe_28__dout;
  wire fifo_Y_pe_28__empty_n;
  wire fifo_Y_pe_28__read;
  wire [64:0] fifo_Y_pe_28__din;
  wire fifo_Y_pe_28__full_n;
  wire fifo_Y_pe_28__write;
  wire [64:0] fifo_Y_pe_29__dout;
  wire fifo_Y_pe_29__empty_n;
  wire fifo_Y_pe_29__read;
  wire [64:0] fifo_Y_pe_29__din;
  wire fifo_Y_pe_29__full_n;
  wire fifo_Y_pe_29__write;
  wire [64:0] fifo_Y_pe_2__dout;
  wire fifo_Y_pe_2__empty_n;
  wire fifo_Y_pe_2__read;
  wire [64:0] fifo_Y_pe_2__din;
  wire fifo_Y_pe_2__full_n;
  wire fifo_Y_pe_2__write;
  wire [64:0] fifo_Y_pe_30__dout;
  wire fifo_Y_pe_30__empty_n;
  wire fifo_Y_pe_30__read;
  wire [64:0] fifo_Y_pe_30__din;
  wire fifo_Y_pe_30__full_n;
  wire fifo_Y_pe_30__write;
  wire [64:0] fifo_Y_pe_31__dout;
  wire fifo_Y_pe_31__empty_n;
  wire fifo_Y_pe_31__read;
  wire [64:0] fifo_Y_pe_31__din;
  wire fifo_Y_pe_31__full_n;
  wire fifo_Y_pe_31__write;
  wire [64:0] fifo_Y_pe_32__dout;
  wire fifo_Y_pe_32__empty_n;
  wire fifo_Y_pe_32__read;
  wire [64:0] fifo_Y_pe_32__din;
  wire fifo_Y_pe_32__full_n;
  wire fifo_Y_pe_32__write;
  wire [64:0] fifo_Y_pe_33__dout;
  wire fifo_Y_pe_33__empty_n;
  wire fifo_Y_pe_33__read;
  wire [64:0] fifo_Y_pe_33__din;
  wire fifo_Y_pe_33__full_n;
  wire fifo_Y_pe_33__write;
  wire [64:0] fifo_Y_pe_34__dout;
  wire fifo_Y_pe_34__empty_n;
  wire fifo_Y_pe_34__read;
  wire [64:0] fifo_Y_pe_34__din;
  wire fifo_Y_pe_34__full_n;
  wire fifo_Y_pe_34__write;
  wire [64:0] fifo_Y_pe_35__dout;
  wire fifo_Y_pe_35__empty_n;
  wire fifo_Y_pe_35__read;
  wire [64:0] fifo_Y_pe_35__din;
  wire fifo_Y_pe_35__full_n;
  wire fifo_Y_pe_35__write;
  wire [64:0] fifo_Y_pe_36__dout;
  wire fifo_Y_pe_36__empty_n;
  wire fifo_Y_pe_36__read;
  wire [64:0] fifo_Y_pe_36__din;
  wire fifo_Y_pe_36__full_n;
  wire fifo_Y_pe_36__write;
  wire [64:0] fifo_Y_pe_37__dout;
  wire fifo_Y_pe_37__empty_n;
  wire fifo_Y_pe_37__read;
  wire [64:0] fifo_Y_pe_37__din;
  wire fifo_Y_pe_37__full_n;
  wire fifo_Y_pe_37__write;
  wire [64:0] fifo_Y_pe_38__dout;
  wire fifo_Y_pe_38__empty_n;
  wire fifo_Y_pe_38__read;
  wire [64:0] fifo_Y_pe_38__din;
  wire fifo_Y_pe_38__full_n;
  wire fifo_Y_pe_38__write;
  wire [64:0] fifo_Y_pe_39__dout;
  wire fifo_Y_pe_39__empty_n;
  wire fifo_Y_pe_39__read;
  wire [64:0] fifo_Y_pe_39__din;
  wire fifo_Y_pe_39__full_n;
  wire fifo_Y_pe_39__write;
  wire [64:0] fifo_Y_pe_3__dout;
  wire fifo_Y_pe_3__empty_n;
  wire fifo_Y_pe_3__read;
  wire [64:0] fifo_Y_pe_3__din;
  wire fifo_Y_pe_3__full_n;
  wire fifo_Y_pe_3__write;
  wire [64:0] fifo_Y_pe_40__dout;
  wire fifo_Y_pe_40__empty_n;
  wire fifo_Y_pe_40__read;
  wire [64:0] fifo_Y_pe_40__din;
  wire fifo_Y_pe_40__full_n;
  wire fifo_Y_pe_40__write;
  wire [64:0] fifo_Y_pe_41__dout;
  wire fifo_Y_pe_41__empty_n;
  wire fifo_Y_pe_41__read;
  wire [64:0] fifo_Y_pe_41__din;
  wire fifo_Y_pe_41__full_n;
  wire fifo_Y_pe_41__write;
  wire [64:0] fifo_Y_pe_42__dout;
  wire fifo_Y_pe_42__empty_n;
  wire fifo_Y_pe_42__read;
  wire [64:0] fifo_Y_pe_42__din;
  wire fifo_Y_pe_42__full_n;
  wire fifo_Y_pe_42__write;
  wire [64:0] fifo_Y_pe_43__dout;
  wire fifo_Y_pe_43__empty_n;
  wire fifo_Y_pe_43__read;
  wire [64:0] fifo_Y_pe_43__din;
  wire fifo_Y_pe_43__full_n;
  wire fifo_Y_pe_43__write;
  wire [64:0] fifo_Y_pe_44__dout;
  wire fifo_Y_pe_44__empty_n;
  wire fifo_Y_pe_44__read;
  wire [64:0] fifo_Y_pe_44__din;
  wire fifo_Y_pe_44__full_n;
  wire fifo_Y_pe_44__write;
  wire [64:0] fifo_Y_pe_45__dout;
  wire fifo_Y_pe_45__empty_n;
  wire fifo_Y_pe_45__read;
  wire [64:0] fifo_Y_pe_45__din;
  wire fifo_Y_pe_45__full_n;
  wire fifo_Y_pe_45__write;
  wire [64:0] fifo_Y_pe_46__dout;
  wire fifo_Y_pe_46__empty_n;
  wire fifo_Y_pe_46__read;
  wire [64:0] fifo_Y_pe_46__din;
  wire fifo_Y_pe_46__full_n;
  wire fifo_Y_pe_46__write;
  wire [64:0] fifo_Y_pe_47__dout;
  wire fifo_Y_pe_47__empty_n;
  wire fifo_Y_pe_47__read;
  wire [64:0] fifo_Y_pe_47__din;
  wire fifo_Y_pe_47__full_n;
  wire fifo_Y_pe_47__write;
  wire [64:0] fifo_Y_pe_4__dout;
  wire fifo_Y_pe_4__empty_n;
  wire fifo_Y_pe_4__read;
  wire [64:0] fifo_Y_pe_4__din;
  wire fifo_Y_pe_4__full_n;
  wire fifo_Y_pe_4__write;
  wire [64:0] fifo_Y_pe_5__dout;
  wire fifo_Y_pe_5__empty_n;
  wire fifo_Y_pe_5__read;
  wire [64:0] fifo_Y_pe_5__din;
  wire fifo_Y_pe_5__full_n;
  wire fifo_Y_pe_5__write;
  wire [64:0] fifo_Y_pe_6__dout;
  wire fifo_Y_pe_6__empty_n;
  wire fifo_Y_pe_6__read;
  wire [64:0] fifo_Y_pe_6__din;
  wire fifo_Y_pe_6__full_n;
  wire fifo_Y_pe_6__write;
  wire [64:0] fifo_Y_pe_7__dout;
  wire fifo_Y_pe_7__empty_n;
  wire fifo_Y_pe_7__read;
  wire [64:0] fifo_Y_pe_7__din;
  wire fifo_Y_pe_7__full_n;
  wire fifo_Y_pe_7__write;
  wire [64:0] fifo_Y_pe_8__dout;
  wire fifo_Y_pe_8__empty_n;
  wire fifo_Y_pe_8__read;
  wire [64:0] fifo_Y_pe_8__din;
  wire fifo_Y_pe_8__full_n;
  wire fifo_Y_pe_8__write;
  wire [64:0] fifo_Y_pe_9__dout;
  wire fifo_Y_pe_9__empty_n;
  wire fifo_Y_pe_9__read;
  wire [64:0] fifo_Y_pe_9__din;
  wire fifo_Y_pe_9__full_n;
  wire fifo_Y_pe_9__write;
  wire [64:0] fifo_Y_pe_abd_0__dout;
  wire fifo_Y_pe_abd_0__empty_n;
  wire fifo_Y_pe_abd_0__read;
  wire [64:0] fifo_Y_pe_abd_0__din;
  wire fifo_Y_pe_abd_0__full_n;
  wire fifo_Y_pe_abd_0__write;
  wire [64:0] fifo_Y_pe_abd_1__dout;
  wire fifo_Y_pe_abd_1__empty_n;
  wire fifo_Y_pe_abd_1__read;
  wire [64:0] fifo_Y_pe_abd_1__din;
  wire fifo_Y_pe_abd_1__full_n;
  wire fifo_Y_pe_abd_1__write;
  wire [64:0] fifo_Y_pe_abd_2__dout;
  wire fifo_Y_pe_abd_2__empty_n;
  wire fifo_Y_pe_abd_2__read;
  wire [64:0] fifo_Y_pe_abd_2__din;
  wire fifo_Y_pe_abd_2__full_n;
  wire fifo_Y_pe_abd_2__write;
  wire [64:0] fifo_Y_pe_abd_3__dout;
  wire fifo_Y_pe_abd_3__empty_n;
  wire fifo_Y_pe_abd_3__read;
  wire [64:0] fifo_Y_pe_abd_3__din;
  wire fifo_Y_pe_abd_3__full_n;
  wire fifo_Y_pe_abd_3__write;
  wire [64:0] fifo_Y_pe_abd_4__dout;
  wire fifo_Y_pe_abd_4__empty_n;
  wire fifo_Y_pe_abd_4__read;
  wire [64:0] fifo_Y_pe_abd_4__din;
  wire fifo_Y_pe_abd_4__full_n;
  wire fifo_Y_pe_abd_4__write;
  wire [64:0] fifo_Y_pe_abd_5__dout;
  wire fifo_Y_pe_abd_5__empty_n;
  wire fifo_Y_pe_abd_5__read;
  wire [64:0] fifo_Y_pe_abd_5__din;
  wire fifo_Y_pe_abd_5__full_n;
  wire fifo_Y_pe_abd_5__write;
  wire [64:0] fifo_Y_pe_abd_6__dout;
  wire fifo_Y_pe_abd_6__empty_n;
  wire fifo_Y_pe_abd_6__read;
  wire [64:0] fifo_Y_pe_abd_6__din;
  wire fifo_Y_pe_abd_6__full_n;
  wire fifo_Y_pe_abd_6__write;
  wire [64:0] fifo_Y_pe_abd_7__dout;
  wire fifo_Y_pe_abd_7__empty_n;
  wire fifo_Y_pe_abd_7__read;
  wire [64:0] fifo_Y_pe_abd_7__din;
  wire fifo_Y_pe_abd_7__full_n;
  wire fifo_Y_pe_abd_7__write;
  wire [400:0] fifo_aXvec_0__dout;
  wire fifo_aXvec_0__empty_n;
  wire fifo_aXvec_0__read;
  wire [400:0] fifo_aXvec_0__din;
  wire fifo_aXvec_0__full_n;
  wire fifo_aXvec_0__write;
  wire [400:0] fifo_aXvec_10__dout;
  wire fifo_aXvec_10__empty_n;
  wire fifo_aXvec_10__read;
  wire [400:0] fifo_aXvec_10__din;
  wire fifo_aXvec_10__full_n;
  wire fifo_aXvec_10__write;
  wire [400:0] fifo_aXvec_11__dout;
  wire fifo_aXvec_11__empty_n;
  wire fifo_aXvec_11__read;
  wire [400:0] fifo_aXvec_11__din;
  wire fifo_aXvec_11__full_n;
  wire fifo_aXvec_11__write;
  wire [400:0] fifo_aXvec_12__dout;
  wire fifo_aXvec_12__empty_n;
  wire fifo_aXvec_12__read;
  wire [400:0] fifo_aXvec_12__din;
  wire fifo_aXvec_12__full_n;
  wire fifo_aXvec_12__write;
  wire [400:0] fifo_aXvec_13__dout;
  wire fifo_aXvec_13__empty_n;
  wire fifo_aXvec_13__read;
  wire [400:0] fifo_aXvec_13__din;
  wire fifo_aXvec_13__full_n;
  wire fifo_aXvec_13__write;
  wire [400:0] fifo_aXvec_14__dout;
  wire fifo_aXvec_14__empty_n;
  wire fifo_aXvec_14__read;
  wire [400:0] fifo_aXvec_14__din;
  wire fifo_aXvec_14__full_n;
  wire fifo_aXvec_14__write;
  wire [400:0] fifo_aXvec_15__dout;
  wire fifo_aXvec_15__empty_n;
  wire fifo_aXvec_15__read;
  wire [400:0] fifo_aXvec_15__din;
  wire fifo_aXvec_15__full_n;
  wire fifo_aXvec_15__write;
  wire [400:0] fifo_aXvec_16__dout;
  wire fifo_aXvec_16__empty_n;
  wire fifo_aXvec_16__read;
  wire [400:0] fifo_aXvec_16__din;
  wire fifo_aXvec_16__full_n;
  wire fifo_aXvec_16__write;
  wire [400:0] fifo_aXvec_17__dout;
  wire fifo_aXvec_17__empty_n;
  wire fifo_aXvec_17__read;
  wire [400:0] fifo_aXvec_17__din;
  wire fifo_aXvec_17__full_n;
  wire fifo_aXvec_17__write;
  wire [400:0] fifo_aXvec_18__dout;
  wire fifo_aXvec_18__empty_n;
  wire fifo_aXvec_18__read;
  wire [400:0] fifo_aXvec_18__din;
  wire fifo_aXvec_18__full_n;
  wire fifo_aXvec_18__write;
  wire [400:0] fifo_aXvec_19__dout;
  wire fifo_aXvec_19__empty_n;
  wire fifo_aXvec_19__read;
  wire [400:0] fifo_aXvec_19__din;
  wire fifo_aXvec_19__full_n;
  wire fifo_aXvec_19__write;
  wire [400:0] fifo_aXvec_1__dout;
  wire fifo_aXvec_1__empty_n;
  wire fifo_aXvec_1__read;
  wire [400:0] fifo_aXvec_1__din;
  wire fifo_aXvec_1__full_n;
  wire fifo_aXvec_1__write;
  wire [400:0] fifo_aXvec_20__dout;
  wire fifo_aXvec_20__empty_n;
  wire fifo_aXvec_20__read;
  wire [400:0] fifo_aXvec_20__din;
  wire fifo_aXvec_20__full_n;
  wire fifo_aXvec_20__write;
  wire [400:0] fifo_aXvec_21__dout;
  wire fifo_aXvec_21__empty_n;
  wire fifo_aXvec_21__read;
  wire [400:0] fifo_aXvec_21__din;
  wire fifo_aXvec_21__full_n;
  wire fifo_aXvec_21__write;
  wire [400:0] fifo_aXvec_22__dout;
  wire fifo_aXvec_22__empty_n;
  wire fifo_aXvec_22__read;
  wire [400:0] fifo_aXvec_22__din;
  wire fifo_aXvec_22__full_n;
  wire fifo_aXvec_22__write;
  wire [400:0] fifo_aXvec_23__dout;
  wire fifo_aXvec_23__empty_n;
  wire fifo_aXvec_23__read;
  wire [400:0] fifo_aXvec_23__din;
  wire fifo_aXvec_23__full_n;
  wire fifo_aXvec_23__write;
  wire [400:0] fifo_aXvec_24__dout;
  wire fifo_aXvec_24__empty_n;
  wire fifo_aXvec_24__read;
  wire [400:0] fifo_aXvec_24__din;
  wire fifo_aXvec_24__full_n;
  wire fifo_aXvec_24__write;
  wire [400:0] fifo_aXvec_25__dout;
  wire fifo_aXvec_25__empty_n;
  wire fifo_aXvec_25__read;
  wire [400:0] fifo_aXvec_25__din;
  wire fifo_aXvec_25__full_n;
  wire fifo_aXvec_25__write;
  wire [400:0] fifo_aXvec_26__dout;
  wire fifo_aXvec_26__empty_n;
  wire fifo_aXvec_26__read;
  wire [400:0] fifo_aXvec_26__din;
  wire fifo_aXvec_26__full_n;
  wire fifo_aXvec_26__write;
  wire [400:0] fifo_aXvec_27__dout;
  wire fifo_aXvec_27__empty_n;
  wire fifo_aXvec_27__read;
  wire [400:0] fifo_aXvec_27__din;
  wire fifo_aXvec_27__full_n;
  wire fifo_aXvec_27__write;
  wire [400:0] fifo_aXvec_28__dout;
  wire fifo_aXvec_28__empty_n;
  wire fifo_aXvec_28__read;
  wire [400:0] fifo_aXvec_28__din;
  wire fifo_aXvec_28__full_n;
  wire fifo_aXvec_28__write;
  wire [400:0] fifo_aXvec_29__dout;
  wire fifo_aXvec_29__empty_n;
  wire fifo_aXvec_29__read;
  wire [400:0] fifo_aXvec_29__din;
  wire fifo_aXvec_29__full_n;
  wire fifo_aXvec_29__write;
  wire [400:0] fifo_aXvec_2__dout;
  wire fifo_aXvec_2__empty_n;
  wire fifo_aXvec_2__read;
  wire [400:0] fifo_aXvec_2__din;
  wire fifo_aXvec_2__full_n;
  wire fifo_aXvec_2__write;
  wire [400:0] fifo_aXvec_30__dout;
  wire fifo_aXvec_30__empty_n;
  wire fifo_aXvec_30__read;
  wire [400:0] fifo_aXvec_30__din;
  wire fifo_aXvec_30__full_n;
  wire fifo_aXvec_30__write;
  wire [400:0] fifo_aXvec_31__dout;
  wire fifo_aXvec_31__empty_n;
  wire fifo_aXvec_31__read;
  wire [400:0] fifo_aXvec_31__din;
  wire fifo_aXvec_31__full_n;
  wire fifo_aXvec_31__write;
  wire [400:0] fifo_aXvec_32__dout;
  wire fifo_aXvec_32__empty_n;
  wire fifo_aXvec_32__read;
  wire [400:0] fifo_aXvec_32__din;
  wire fifo_aXvec_32__full_n;
  wire fifo_aXvec_32__write;
  wire [400:0] fifo_aXvec_33__dout;
  wire fifo_aXvec_33__empty_n;
  wire fifo_aXvec_33__read;
  wire [400:0] fifo_aXvec_33__din;
  wire fifo_aXvec_33__full_n;
  wire fifo_aXvec_33__write;
  wire [400:0] fifo_aXvec_34__dout;
  wire fifo_aXvec_34__empty_n;
  wire fifo_aXvec_34__read;
  wire [400:0] fifo_aXvec_34__din;
  wire fifo_aXvec_34__full_n;
  wire fifo_aXvec_34__write;
  wire [400:0] fifo_aXvec_35__dout;
  wire fifo_aXvec_35__empty_n;
  wire fifo_aXvec_35__read;
  wire [400:0] fifo_aXvec_35__din;
  wire fifo_aXvec_35__full_n;
  wire fifo_aXvec_35__write;
  wire [400:0] fifo_aXvec_36__dout;
  wire fifo_aXvec_36__empty_n;
  wire fifo_aXvec_36__read;
  wire [400:0] fifo_aXvec_36__din;
  wire fifo_aXvec_36__full_n;
  wire fifo_aXvec_36__write;
  wire [400:0] fifo_aXvec_37__dout;
  wire fifo_aXvec_37__empty_n;
  wire fifo_aXvec_37__read;
  wire [400:0] fifo_aXvec_37__din;
  wire fifo_aXvec_37__full_n;
  wire fifo_aXvec_37__write;
  wire [400:0] fifo_aXvec_38__dout;
  wire fifo_aXvec_38__empty_n;
  wire fifo_aXvec_38__read;
  wire [400:0] fifo_aXvec_38__din;
  wire fifo_aXvec_38__full_n;
  wire fifo_aXvec_38__write;
  wire [400:0] fifo_aXvec_39__dout;
  wire fifo_aXvec_39__empty_n;
  wire fifo_aXvec_39__read;
  wire [400:0] fifo_aXvec_39__din;
  wire fifo_aXvec_39__full_n;
  wire fifo_aXvec_39__write;
  wire [400:0] fifo_aXvec_3__dout;
  wire fifo_aXvec_3__empty_n;
  wire fifo_aXvec_3__read;
  wire [400:0] fifo_aXvec_3__din;
  wire fifo_aXvec_3__full_n;
  wire fifo_aXvec_3__write;
  wire [400:0] fifo_aXvec_40__dout;
  wire fifo_aXvec_40__empty_n;
  wire fifo_aXvec_40__read;
  wire [400:0] fifo_aXvec_40__din;
  wire fifo_aXvec_40__full_n;
  wire fifo_aXvec_40__write;
  wire [400:0] fifo_aXvec_41__dout;
  wire fifo_aXvec_41__empty_n;
  wire fifo_aXvec_41__read;
  wire [400:0] fifo_aXvec_41__din;
  wire fifo_aXvec_41__full_n;
  wire fifo_aXvec_41__write;
  wire [400:0] fifo_aXvec_42__dout;
  wire fifo_aXvec_42__empty_n;
  wire fifo_aXvec_42__read;
  wire [400:0] fifo_aXvec_42__din;
  wire fifo_aXvec_42__full_n;
  wire fifo_aXvec_42__write;
  wire [400:0] fifo_aXvec_43__dout;
  wire fifo_aXvec_43__empty_n;
  wire fifo_aXvec_43__read;
  wire [400:0] fifo_aXvec_43__din;
  wire fifo_aXvec_43__full_n;
  wire fifo_aXvec_43__write;
  wire [400:0] fifo_aXvec_44__dout;
  wire fifo_aXvec_44__empty_n;
  wire fifo_aXvec_44__read;
  wire [400:0] fifo_aXvec_44__din;
  wire fifo_aXvec_44__full_n;
  wire fifo_aXvec_44__write;
  wire [400:0] fifo_aXvec_45__dout;
  wire fifo_aXvec_45__empty_n;
  wire fifo_aXvec_45__read;
  wire [400:0] fifo_aXvec_45__din;
  wire fifo_aXvec_45__full_n;
  wire fifo_aXvec_45__write;
  wire [400:0] fifo_aXvec_46__dout;
  wire fifo_aXvec_46__empty_n;
  wire fifo_aXvec_46__read;
  wire [400:0] fifo_aXvec_46__din;
  wire fifo_aXvec_46__full_n;
  wire fifo_aXvec_46__write;
  wire [400:0] fifo_aXvec_47__dout;
  wire fifo_aXvec_47__empty_n;
  wire fifo_aXvec_47__read;
  wire [400:0] fifo_aXvec_47__din;
  wire fifo_aXvec_47__full_n;
  wire fifo_aXvec_47__write;
  wire [400:0] fifo_aXvec_4__dout;
  wire fifo_aXvec_4__empty_n;
  wire fifo_aXvec_4__read;
  wire [400:0] fifo_aXvec_4__din;
  wire fifo_aXvec_4__full_n;
  wire fifo_aXvec_4__write;
  wire [400:0] fifo_aXvec_5__dout;
  wire fifo_aXvec_5__empty_n;
  wire fifo_aXvec_5__read;
  wire [400:0] fifo_aXvec_5__din;
  wire fifo_aXvec_5__full_n;
  wire fifo_aXvec_5__write;
  wire [400:0] fifo_aXvec_6__dout;
  wire fifo_aXvec_6__empty_n;
  wire fifo_aXvec_6__read;
  wire [400:0] fifo_aXvec_6__din;
  wire fifo_aXvec_6__full_n;
  wire fifo_aXvec_6__write;
  wire [400:0] fifo_aXvec_7__dout;
  wire fifo_aXvec_7__empty_n;
  wire fifo_aXvec_7__read;
  wire [400:0] fifo_aXvec_7__din;
  wire fifo_aXvec_7__full_n;
  wire fifo_aXvec_7__write;
  wire [400:0] fifo_aXvec_8__dout;
  wire fifo_aXvec_8__empty_n;
  wire fifo_aXvec_8__read;
  wire [400:0] fifo_aXvec_8__din;
  wire fifo_aXvec_8__full_n;
  wire fifo_aXvec_8__write;
  wire [400:0] fifo_aXvec_9__dout;
  wire fifo_aXvec_9__empty_n;
  wire fifo_aXvec_9__read;
  wire [400:0] fifo_aXvec_9__din;
  wire fifo_aXvec_9__full_n;
  wire fifo_aXvec_9__write;
  wire [31:0] Arbiter_Y_0___M__q0;
  wire [31:0] Arbiter_Y_0___P_N__q0;
  wire Arbiter_Y_0__ap_start;
  wire Arbiter_Y_0__ap_ready;
  wire Arbiter_Y_0__ap_done;
  wire Arbiter_Y_0__ap_idle;
  wire [31:0] Arbiter_Y_1___M__q0;
  wire [31:0] Arbiter_Y_1___P_N__q0;
  wire Arbiter_Y_1__ap_start;
  wire Arbiter_Y_1__ap_ready;
  wire Arbiter_Y_1__ap_done;
  wire Arbiter_Y_1__ap_idle;
  wire [31:0] Arbiter_Y_2___M__q0;
  wire [31:0] Arbiter_Y_2___P_N__q0;
  wire Arbiter_Y_2__ap_start;
  wire Arbiter_Y_2__ap_ready;
  wire Arbiter_Y_2__ap_done;
  wire Arbiter_Y_2__ap_idle;
  wire [31:0] Arbiter_Y_3___M__q0;
  wire [31:0] Arbiter_Y_3___P_N__q0;
  wire Arbiter_Y_3__ap_start;
  wire Arbiter_Y_3__ap_ready;
  wire Arbiter_Y_3__ap_done;
  wire Arbiter_Y_3__ap_idle;
  wire [31:0] Arbiter_Y_4___M__q0;
  wire [31:0] Arbiter_Y_4___P_N__q0;
  wire Arbiter_Y_4__ap_start;
  wire Arbiter_Y_4__ap_ready;
  wire Arbiter_Y_4__ap_done;
  wire Arbiter_Y_4__ap_idle;
  wire [31:0] Arbiter_Y_5___M__q0;
  wire [31:0] Arbiter_Y_5___P_N__q0;
  wire Arbiter_Y_5__ap_start;
  wire Arbiter_Y_5__ap_ready;
  wire Arbiter_Y_5__ap_done;
  wire Arbiter_Y_5__ap_idle;
  wire [31:0] Arbiter_Y_6___M__q0;
  wire [31:0] Arbiter_Y_6___P_N__q0;
  wire Arbiter_Y_6__ap_start;
  wire Arbiter_Y_6__ap_ready;
  wire Arbiter_Y_6__ap_done;
  wire Arbiter_Y_6__ap_idle;
  wire [31:0] Arbiter_Y_7___M__q0;
  wire [31:0] Arbiter_Y_7___P_N__q0;
  wire Arbiter_Y_7__ap_start;
  wire Arbiter_Y_7__ap_ready;
  wire Arbiter_Y_7__ap_done;
  wire Arbiter_Y_7__ap_idle;
  wire FloatvAddFloatv_0__ap_start;
  wire [31:0] FloatvMultConst_0___M__q0;
  wire [31:0] FloatvMultConst_0___P_N__q0;
  wire [31:0] FloatvMultConst_0___alpha_u__q0;
  wire FloatvMultConst_0__ap_start;
  wire FloatvMultConst_0__ap_ready;
  wire FloatvMultConst_0__ap_done;
  wire FloatvMultConst_0__ap_idle;
  wire [31:0] FloatvMultConst_1___M__q0;
  wire [31:0] FloatvMultConst_1___P_N__q0;
  wire [31:0] FloatvMultConst_1___beta_u__q0;
  wire FloatvMultConst_1__ap_start;
  wire FloatvMultConst_1__ap_ready;
  wire FloatvMultConst_1__ap_done;
  wire FloatvMultConst_1__ap_idle;
  wire Merger_Y_0__ap_start;
  wire PEG_Xvec_0__ap_start;
  wire PEG_Xvec_0__ap_ready;
  wire PEG_Xvec_0__ap_done;
  wire PEG_Xvec_0__ap_idle;
  wire PEG_Xvec_1__ap_start;
  wire PEG_Xvec_1__ap_ready;
  wire PEG_Xvec_1__ap_done;
  wire PEG_Xvec_1__ap_idle;
  wire PEG_Xvec_2__ap_start;
  wire PEG_Xvec_2__ap_ready;
  wire PEG_Xvec_2__ap_done;
  wire PEG_Xvec_2__ap_idle;
  wire PEG_Xvec_3__ap_start;
  wire PEG_Xvec_3__ap_ready;
  wire PEG_Xvec_3__ap_done;
  wire PEG_Xvec_3__ap_idle;
  wire PEG_Xvec_4__ap_start;
  wire PEG_Xvec_4__ap_ready;
  wire PEG_Xvec_4__ap_done;
  wire PEG_Xvec_4__ap_idle;
  wire PEG_Xvec_5__ap_start;
  wire PEG_Xvec_5__ap_ready;
  wire PEG_Xvec_5__ap_done;
  wire PEG_Xvec_5__ap_idle;
  wire PEG_Xvec_6__ap_start;
  wire PEG_Xvec_6__ap_ready;
  wire PEG_Xvec_6__ap_done;
  wire PEG_Xvec_6__ap_idle;
  wire PEG_Xvec_7__ap_start;
  wire PEG_Xvec_7__ap_ready;
  wire PEG_Xvec_7__ap_done;
  wire PEG_Xvec_7__ap_idle;
  wire PEG_Xvec_8__ap_start;
  wire PEG_Xvec_8__ap_ready;
  wire PEG_Xvec_8__ap_done;
  wire PEG_Xvec_8__ap_idle;
  wire PEG_Xvec_9__ap_start;
  wire PEG_Xvec_9__ap_ready;
  wire PEG_Xvec_9__ap_done;
  wire PEG_Xvec_9__ap_idle;
  wire PEG_Xvec_10__ap_start;
  wire PEG_Xvec_10__ap_ready;
  wire PEG_Xvec_10__ap_done;
  wire PEG_Xvec_10__ap_idle;
  wire PEG_Xvec_11__ap_start;
  wire PEG_Xvec_11__ap_ready;
  wire PEG_Xvec_11__ap_done;
  wire PEG_Xvec_11__ap_idle;
  wire PEG_Xvec_12__ap_start;
  wire PEG_Xvec_12__ap_ready;
  wire PEG_Xvec_12__ap_done;
  wire PEG_Xvec_12__ap_idle;
  wire PEG_Xvec_13__ap_start;
  wire PEG_Xvec_13__ap_ready;
  wire PEG_Xvec_13__ap_done;
  wire PEG_Xvec_13__ap_idle;
  wire PEG_Xvec_14__ap_start;
  wire PEG_Xvec_14__ap_ready;
  wire PEG_Xvec_14__ap_done;
  wire PEG_Xvec_14__ap_idle;
  wire PEG_Xvec_15__ap_start;
  wire PEG_Xvec_15__ap_ready;
  wire PEG_Xvec_15__ap_done;
  wire PEG_Xvec_15__ap_idle;
  wire PEG_Xvec_16__ap_start;
  wire PEG_Xvec_16__ap_ready;
  wire PEG_Xvec_16__ap_done;
  wire PEG_Xvec_16__ap_idle;
  wire PEG_Xvec_17__ap_start;
  wire PEG_Xvec_17__ap_ready;
  wire PEG_Xvec_17__ap_done;
  wire PEG_Xvec_17__ap_idle;
  wire PEG_Xvec_18__ap_start;
  wire PEG_Xvec_18__ap_ready;
  wire PEG_Xvec_18__ap_done;
  wire PEG_Xvec_18__ap_idle;
  wire PEG_Xvec_19__ap_start;
  wire PEG_Xvec_19__ap_ready;
  wire PEG_Xvec_19__ap_done;
  wire PEG_Xvec_19__ap_idle;
  wire PEG_Xvec_20__ap_start;
  wire PEG_Xvec_20__ap_ready;
  wire PEG_Xvec_20__ap_done;
  wire PEG_Xvec_20__ap_idle;
  wire PEG_Xvec_21__ap_start;
  wire PEG_Xvec_21__ap_ready;
  wire PEG_Xvec_21__ap_done;
  wire PEG_Xvec_21__ap_idle;
  wire PEG_Xvec_22__ap_start;
  wire PEG_Xvec_22__ap_ready;
  wire PEG_Xvec_22__ap_done;
  wire PEG_Xvec_22__ap_idle;
  wire PEG_Xvec_23__ap_start;
  wire PEG_Xvec_23__ap_ready;
  wire PEG_Xvec_23__ap_done;
  wire PEG_Xvec_23__ap_idle;
  wire PEG_Xvec_24__ap_start;
  wire PEG_Xvec_24__ap_ready;
  wire PEG_Xvec_24__ap_done;
  wire PEG_Xvec_24__ap_idle;
  wire PEG_Xvec_25__ap_start;
  wire PEG_Xvec_25__ap_ready;
  wire PEG_Xvec_25__ap_done;
  wire PEG_Xvec_25__ap_idle;
  wire PEG_Xvec_26__ap_start;
  wire PEG_Xvec_26__ap_ready;
  wire PEG_Xvec_26__ap_done;
  wire PEG_Xvec_26__ap_idle;
  wire PEG_Xvec_27__ap_start;
  wire PEG_Xvec_27__ap_ready;
  wire PEG_Xvec_27__ap_done;
  wire PEG_Xvec_27__ap_idle;
  wire PEG_Xvec_28__ap_start;
  wire PEG_Xvec_28__ap_ready;
  wire PEG_Xvec_28__ap_done;
  wire PEG_Xvec_28__ap_idle;
  wire PEG_Xvec_29__ap_start;
  wire PEG_Xvec_29__ap_ready;
  wire PEG_Xvec_29__ap_done;
  wire PEG_Xvec_29__ap_idle;
  wire PEG_Xvec_30__ap_start;
  wire PEG_Xvec_30__ap_ready;
  wire PEG_Xvec_30__ap_done;
  wire PEG_Xvec_30__ap_idle;
  wire PEG_Xvec_31__ap_start;
  wire PEG_Xvec_31__ap_ready;
  wire PEG_Xvec_31__ap_done;
  wire PEG_Xvec_31__ap_idle;
  wire PEG_Xvec_32__ap_start;
  wire PEG_Xvec_32__ap_ready;
  wire PEG_Xvec_32__ap_done;
  wire PEG_Xvec_32__ap_idle;
  wire PEG_Xvec_33__ap_start;
  wire PEG_Xvec_33__ap_ready;
  wire PEG_Xvec_33__ap_done;
  wire PEG_Xvec_33__ap_idle;
  wire PEG_Xvec_34__ap_start;
  wire PEG_Xvec_34__ap_ready;
  wire PEG_Xvec_34__ap_done;
  wire PEG_Xvec_34__ap_idle;
  wire PEG_Xvec_35__ap_start;
  wire PEG_Xvec_35__ap_ready;
  wire PEG_Xvec_35__ap_done;
  wire PEG_Xvec_35__ap_idle;
  wire PEG_Xvec_36__ap_start;
  wire PEG_Xvec_36__ap_ready;
  wire PEG_Xvec_36__ap_done;
  wire PEG_Xvec_36__ap_idle;
  wire PEG_Xvec_37__ap_start;
  wire PEG_Xvec_37__ap_ready;
  wire PEG_Xvec_37__ap_done;
  wire PEG_Xvec_37__ap_idle;
  wire PEG_Xvec_38__ap_start;
  wire PEG_Xvec_38__ap_ready;
  wire PEG_Xvec_38__ap_done;
  wire PEG_Xvec_38__ap_idle;
  wire PEG_Xvec_39__ap_start;
  wire PEG_Xvec_39__ap_ready;
  wire PEG_Xvec_39__ap_done;
  wire PEG_Xvec_39__ap_idle;
  wire PEG_Xvec_40__ap_start;
  wire PEG_Xvec_40__ap_ready;
  wire PEG_Xvec_40__ap_done;
  wire PEG_Xvec_40__ap_idle;
  wire PEG_Xvec_41__ap_start;
  wire PEG_Xvec_41__ap_ready;
  wire PEG_Xvec_41__ap_done;
  wire PEG_Xvec_41__ap_idle;
  wire PEG_Xvec_42__ap_start;
  wire PEG_Xvec_42__ap_ready;
  wire PEG_Xvec_42__ap_done;
  wire PEG_Xvec_42__ap_idle;
  wire PEG_Xvec_43__ap_start;
  wire PEG_Xvec_43__ap_ready;
  wire PEG_Xvec_43__ap_done;
  wire PEG_Xvec_43__ap_idle;
  wire PEG_Xvec_44__ap_start;
  wire PEG_Xvec_44__ap_ready;
  wire PEG_Xvec_44__ap_done;
  wire PEG_Xvec_44__ap_idle;
  wire PEG_Xvec_45__ap_start;
  wire PEG_Xvec_45__ap_ready;
  wire PEG_Xvec_45__ap_done;
  wire PEG_Xvec_45__ap_idle;
  wire PEG_Xvec_46__ap_start;
  wire PEG_Xvec_46__ap_ready;
  wire PEG_Xvec_46__ap_done;
  wire PEG_Xvec_46__ap_idle;
  wire PEG_Xvec_47__ap_start;
  wire PEG_Xvec_47__ap_ready;
  wire PEG_Xvec_47__ap_done;
  wire PEG_Xvec_47__ap_idle;
  wire PEG_Yvec_0__ap_start;
  wire PEG_Yvec_0__ap_ready;
  wire PEG_Yvec_0__ap_done;
  wire PEG_Yvec_0__ap_idle;
  wire PEG_Yvec_1__ap_start;
  wire PEG_Yvec_1__ap_ready;
  wire PEG_Yvec_1__ap_done;
  wire PEG_Yvec_1__ap_idle;
  wire PEG_Yvec_2__ap_start;
  wire PEG_Yvec_2__ap_ready;
  wire PEG_Yvec_2__ap_done;
  wire PEG_Yvec_2__ap_idle;
  wire PEG_Yvec_3__ap_start;
  wire PEG_Yvec_3__ap_ready;
  wire PEG_Yvec_3__ap_done;
  wire PEG_Yvec_3__ap_idle;
  wire PEG_Yvec_4__ap_start;
  wire PEG_Yvec_4__ap_ready;
  wire PEG_Yvec_4__ap_done;
  wire PEG_Yvec_4__ap_idle;
  wire PEG_Yvec_5__ap_start;
  wire PEG_Yvec_5__ap_ready;
  wire PEG_Yvec_5__ap_done;
  wire PEG_Yvec_5__ap_idle;
  wire PEG_Yvec_6__ap_start;
  wire PEG_Yvec_6__ap_ready;
  wire PEG_Yvec_6__ap_done;
  wire PEG_Yvec_6__ap_idle;
  wire PEG_Yvec_7__ap_start;
  wire PEG_Yvec_7__ap_ready;
  wire PEG_Yvec_7__ap_done;
  wire PEG_Yvec_7__ap_idle;
  wire PEG_Yvec_8__ap_start;
  wire PEG_Yvec_8__ap_ready;
  wire PEG_Yvec_8__ap_done;
  wire PEG_Yvec_8__ap_idle;
  wire PEG_Yvec_9__ap_start;
  wire PEG_Yvec_9__ap_ready;
  wire PEG_Yvec_9__ap_done;
  wire PEG_Yvec_9__ap_idle;
  wire PEG_Yvec_10__ap_start;
  wire PEG_Yvec_10__ap_ready;
  wire PEG_Yvec_10__ap_done;
  wire PEG_Yvec_10__ap_idle;
  wire PEG_Yvec_11__ap_start;
  wire PEG_Yvec_11__ap_ready;
  wire PEG_Yvec_11__ap_done;
  wire PEG_Yvec_11__ap_idle;
  wire PEG_Yvec_12__ap_start;
  wire PEG_Yvec_12__ap_ready;
  wire PEG_Yvec_12__ap_done;
  wire PEG_Yvec_12__ap_idle;
  wire PEG_Yvec_13__ap_start;
  wire PEG_Yvec_13__ap_ready;
  wire PEG_Yvec_13__ap_done;
  wire PEG_Yvec_13__ap_idle;
  wire PEG_Yvec_14__ap_start;
  wire PEG_Yvec_14__ap_ready;
  wire PEG_Yvec_14__ap_done;
  wire PEG_Yvec_14__ap_idle;
  wire PEG_Yvec_15__ap_start;
  wire PEG_Yvec_15__ap_ready;
  wire PEG_Yvec_15__ap_done;
  wire PEG_Yvec_15__ap_idle;
  wire PEG_Yvec_16__ap_start;
  wire PEG_Yvec_16__ap_ready;
  wire PEG_Yvec_16__ap_done;
  wire PEG_Yvec_16__ap_idle;
  wire PEG_Yvec_17__ap_start;
  wire PEG_Yvec_17__ap_ready;
  wire PEG_Yvec_17__ap_done;
  wire PEG_Yvec_17__ap_idle;
  wire PEG_Yvec_18__ap_start;
  wire PEG_Yvec_18__ap_ready;
  wire PEG_Yvec_18__ap_done;
  wire PEG_Yvec_18__ap_idle;
  wire PEG_Yvec_19__ap_start;
  wire PEG_Yvec_19__ap_ready;
  wire PEG_Yvec_19__ap_done;
  wire PEG_Yvec_19__ap_idle;
  wire PEG_Yvec_20__ap_start;
  wire PEG_Yvec_20__ap_ready;
  wire PEG_Yvec_20__ap_done;
  wire PEG_Yvec_20__ap_idle;
  wire PEG_Yvec_21__ap_start;
  wire PEG_Yvec_21__ap_ready;
  wire PEG_Yvec_21__ap_done;
  wire PEG_Yvec_21__ap_idle;
  wire PEG_Yvec_22__ap_start;
  wire PEG_Yvec_22__ap_ready;
  wire PEG_Yvec_22__ap_done;
  wire PEG_Yvec_22__ap_idle;
  wire PEG_Yvec_23__ap_start;
  wire PEG_Yvec_23__ap_ready;
  wire PEG_Yvec_23__ap_done;
  wire PEG_Yvec_23__ap_idle;
  wire PEG_Yvec_24__ap_start;
  wire PEG_Yvec_24__ap_ready;
  wire PEG_Yvec_24__ap_done;
  wire PEG_Yvec_24__ap_idle;
  wire PEG_Yvec_25__ap_start;
  wire PEG_Yvec_25__ap_ready;
  wire PEG_Yvec_25__ap_done;
  wire PEG_Yvec_25__ap_idle;
  wire PEG_Yvec_26__ap_start;
  wire PEG_Yvec_26__ap_ready;
  wire PEG_Yvec_26__ap_done;
  wire PEG_Yvec_26__ap_idle;
  wire PEG_Yvec_27__ap_start;
  wire PEG_Yvec_27__ap_ready;
  wire PEG_Yvec_27__ap_done;
  wire PEG_Yvec_27__ap_idle;
  wire PEG_Yvec_28__ap_start;
  wire PEG_Yvec_28__ap_ready;
  wire PEG_Yvec_28__ap_done;
  wire PEG_Yvec_28__ap_idle;
  wire PEG_Yvec_29__ap_start;
  wire PEG_Yvec_29__ap_ready;
  wire PEG_Yvec_29__ap_done;
  wire PEG_Yvec_29__ap_idle;
  wire PEG_Yvec_30__ap_start;
  wire PEG_Yvec_30__ap_ready;
  wire PEG_Yvec_30__ap_done;
  wire PEG_Yvec_30__ap_idle;
  wire PEG_Yvec_31__ap_start;
  wire PEG_Yvec_31__ap_ready;
  wire PEG_Yvec_31__ap_done;
  wire PEG_Yvec_31__ap_idle;
  wire PEG_Yvec_32__ap_start;
  wire PEG_Yvec_32__ap_ready;
  wire PEG_Yvec_32__ap_done;
  wire PEG_Yvec_32__ap_idle;
  wire PEG_Yvec_33__ap_start;
  wire PEG_Yvec_33__ap_ready;
  wire PEG_Yvec_33__ap_done;
  wire PEG_Yvec_33__ap_idle;
  wire PEG_Yvec_34__ap_start;
  wire PEG_Yvec_34__ap_ready;
  wire PEG_Yvec_34__ap_done;
  wire PEG_Yvec_34__ap_idle;
  wire PEG_Yvec_35__ap_start;
  wire PEG_Yvec_35__ap_ready;
  wire PEG_Yvec_35__ap_done;
  wire PEG_Yvec_35__ap_idle;
  wire PEG_Yvec_36__ap_start;
  wire PEG_Yvec_36__ap_ready;
  wire PEG_Yvec_36__ap_done;
  wire PEG_Yvec_36__ap_idle;
  wire PEG_Yvec_37__ap_start;
  wire PEG_Yvec_37__ap_ready;
  wire PEG_Yvec_37__ap_done;
  wire PEG_Yvec_37__ap_idle;
  wire PEG_Yvec_38__ap_start;
  wire PEG_Yvec_38__ap_ready;
  wire PEG_Yvec_38__ap_done;
  wire PEG_Yvec_38__ap_idle;
  wire PEG_Yvec_39__ap_start;
  wire PEG_Yvec_39__ap_ready;
  wire PEG_Yvec_39__ap_done;
  wire PEG_Yvec_39__ap_idle;
  wire PEG_Yvec_40__ap_start;
  wire PEG_Yvec_40__ap_ready;
  wire PEG_Yvec_40__ap_done;
  wire PEG_Yvec_40__ap_idle;
  wire PEG_Yvec_41__ap_start;
  wire PEG_Yvec_41__ap_ready;
  wire PEG_Yvec_41__ap_done;
  wire PEG_Yvec_41__ap_idle;
  wire PEG_Yvec_42__ap_start;
  wire PEG_Yvec_42__ap_ready;
  wire PEG_Yvec_42__ap_done;
  wire PEG_Yvec_42__ap_idle;
  wire PEG_Yvec_43__ap_start;
  wire PEG_Yvec_43__ap_ready;
  wire PEG_Yvec_43__ap_done;
  wire PEG_Yvec_43__ap_idle;
  wire PEG_Yvec_44__ap_start;
  wire PEG_Yvec_44__ap_ready;
  wire PEG_Yvec_44__ap_done;
  wire PEG_Yvec_44__ap_idle;
  wire PEG_Yvec_45__ap_start;
  wire PEG_Yvec_45__ap_ready;
  wire PEG_Yvec_45__ap_done;
  wire PEG_Yvec_45__ap_idle;
  wire PEG_Yvec_46__ap_start;
  wire PEG_Yvec_46__ap_ready;
  wire PEG_Yvec_46__ap_done;
  wire PEG_Yvec_46__ap_idle;
  wire PEG_Yvec_47__ap_start;
  wire PEG_Yvec_47__ap_ready;
  wire PEG_Yvec_47__ap_done;
  wire PEG_Yvec_47__ap_idle;
  wire black_hole_float_v16_0__ap_start;
  wire black_hole_int_0__ap_start;
  wire [31:0] read_A_0___NUM_A_LEN__q0;
  wire [31:0] read_A_0___P_N__q0;
  wire [63:0] read_A_0___edge_list_ch_0__q0;
  wire [63:0] edge_list_ch_0_read_addr__din;
  wire edge_list_ch_0_read_addr__full_n;
  wire edge_list_ch_0_read_addr__write;
  wire [255:0] edge_list_ch_0_read_data__dout;
  wire edge_list_ch_0_read_data__empty_n;
  wire edge_list_ch_0_read_data__read;
  wire [63:0] edge_list_ch_0_write_addr__din;
  wire edge_list_ch_0_write_addr__full_n;
  wire edge_list_ch_0_write_addr__write;
  wire [255:0] edge_list_ch_0_write_data__din;
  wire edge_list_ch_0_write_data__full_n;
  wire edge_list_ch_0_write_data__write;
  wire [7:0] edge_list_ch_0_write_resp__dout;
  wire edge_list_ch_0_write_resp__empty_n;
  wire edge_list_ch_0_write_resp__read;
  wire read_A_0__ap_start;
  wire read_A_0__ap_ready;
  wire read_A_0__ap_done;
  wire read_A_0__ap_idle;
  wire [31:0] read_A_1___NUM_A_LEN__q0;
  wire [31:0] read_A_1___P_N__q0;
  wire [63:0] read_A_1___edge_list_ch_1__q0;
  wire [63:0] edge_list_ch_1_read_addr__din;
  wire edge_list_ch_1_read_addr__full_n;
  wire edge_list_ch_1_read_addr__write;
  wire [255:0] edge_list_ch_1_read_data__dout;
  wire edge_list_ch_1_read_data__empty_n;
  wire edge_list_ch_1_read_data__read;
  wire [63:0] edge_list_ch_1_write_addr__din;
  wire edge_list_ch_1_write_addr__full_n;
  wire edge_list_ch_1_write_addr__write;
  wire [255:0] edge_list_ch_1_write_data__din;
  wire edge_list_ch_1_write_data__full_n;
  wire edge_list_ch_1_write_data__write;
  wire [7:0] edge_list_ch_1_write_resp__dout;
  wire edge_list_ch_1_write_resp__empty_n;
  wire edge_list_ch_1_write_resp__read;
  wire read_A_1__ap_start;
  wire read_A_1__ap_ready;
  wire read_A_1__ap_done;
  wire read_A_1__ap_idle;
  wire [31:0] read_A_2___NUM_A_LEN__q0;
  wire [31:0] read_A_2___P_N__q0;
  wire [63:0] read_A_2___edge_list_ch_2__q0;
  wire [63:0] edge_list_ch_2_read_addr__din;
  wire edge_list_ch_2_read_addr__full_n;
  wire edge_list_ch_2_read_addr__write;
  wire [255:0] edge_list_ch_2_read_data__dout;
  wire edge_list_ch_2_read_data__empty_n;
  wire edge_list_ch_2_read_data__read;
  wire [63:0] edge_list_ch_2_write_addr__din;
  wire edge_list_ch_2_write_addr__full_n;
  wire edge_list_ch_2_write_addr__write;
  wire [255:0] edge_list_ch_2_write_data__din;
  wire edge_list_ch_2_write_data__full_n;
  wire edge_list_ch_2_write_data__write;
  wire [7:0] edge_list_ch_2_write_resp__dout;
  wire edge_list_ch_2_write_resp__empty_n;
  wire edge_list_ch_2_write_resp__read;
  wire read_A_2__ap_start;
  wire read_A_2__ap_ready;
  wire read_A_2__ap_done;
  wire read_A_2__ap_idle;
  wire [31:0] read_A_3___NUM_A_LEN__q0;
  wire [31:0] read_A_3___P_N__q0;
  wire [63:0] read_A_3___edge_list_ch_3__q0;
  wire [63:0] edge_list_ch_3_read_addr__din;
  wire edge_list_ch_3_read_addr__full_n;
  wire edge_list_ch_3_read_addr__write;
  wire [255:0] edge_list_ch_3_read_data__dout;
  wire edge_list_ch_3_read_data__empty_n;
  wire edge_list_ch_3_read_data__read;
  wire [63:0] edge_list_ch_3_write_addr__din;
  wire edge_list_ch_3_write_addr__full_n;
  wire edge_list_ch_3_write_addr__write;
  wire [255:0] edge_list_ch_3_write_data__din;
  wire edge_list_ch_3_write_data__full_n;
  wire edge_list_ch_3_write_data__write;
  wire [7:0] edge_list_ch_3_write_resp__dout;
  wire edge_list_ch_3_write_resp__empty_n;
  wire edge_list_ch_3_write_resp__read;
  wire read_A_3__ap_start;
  wire read_A_3__ap_ready;
  wire read_A_3__ap_done;
  wire read_A_3__ap_idle;
  wire [31:0] read_A_4___NUM_A_LEN__q0;
  wire [31:0] read_A_4___P_N__q0;
  wire [63:0] read_A_4___edge_list_ch_4__q0;
  wire [63:0] edge_list_ch_4_read_addr__din;
  wire edge_list_ch_4_read_addr__full_n;
  wire edge_list_ch_4_read_addr__write;
  wire [255:0] edge_list_ch_4_read_data__dout;
  wire edge_list_ch_4_read_data__empty_n;
  wire edge_list_ch_4_read_data__read;
  wire [63:0] edge_list_ch_4_write_addr__din;
  wire edge_list_ch_4_write_addr__full_n;
  wire edge_list_ch_4_write_addr__write;
  wire [255:0] edge_list_ch_4_write_data__din;
  wire edge_list_ch_4_write_data__full_n;
  wire edge_list_ch_4_write_data__write;
  wire [7:0] edge_list_ch_4_write_resp__dout;
  wire edge_list_ch_4_write_resp__empty_n;
  wire edge_list_ch_4_write_resp__read;
  wire read_A_4__ap_start;
  wire read_A_4__ap_ready;
  wire read_A_4__ap_done;
  wire read_A_4__ap_idle;
  wire [31:0] read_A_5___NUM_A_LEN__q0;
  wire [31:0] read_A_5___P_N__q0;
  wire [63:0] read_A_5___edge_list_ch_5__q0;
  wire [63:0] edge_list_ch_5_read_addr__din;
  wire edge_list_ch_5_read_addr__full_n;
  wire edge_list_ch_5_read_addr__write;
  wire [255:0] edge_list_ch_5_read_data__dout;
  wire edge_list_ch_5_read_data__empty_n;
  wire edge_list_ch_5_read_data__read;
  wire [63:0] edge_list_ch_5_write_addr__din;
  wire edge_list_ch_5_write_addr__full_n;
  wire edge_list_ch_5_write_addr__write;
  wire [255:0] edge_list_ch_5_write_data__din;
  wire edge_list_ch_5_write_data__full_n;
  wire edge_list_ch_5_write_data__write;
  wire [7:0] edge_list_ch_5_write_resp__dout;
  wire edge_list_ch_5_write_resp__empty_n;
  wire edge_list_ch_5_write_resp__read;
  wire read_A_5__ap_start;
  wire read_A_5__ap_ready;
  wire read_A_5__ap_done;
  wire read_A_5__ap_idle;
  wire [31:0] read_A_6___NUM_A_LEN__q0;
  wire [31:0] read_A_6___P_N__q0;
  wire [63:0] read_A_6___edge_list_ch_6__q0;
  wire [63:0] edge_list_ch_6_read_addr__din;
  wire edge_list_ch_6_read_addr__full_n;
  wire edge_list_ch_6_read_addr__write;
  wire [255:0] edge_list_ch_6_read_data__dout;
  wire edge_list_ch_6_read_data__empty_n;
  wire edge_list_ch_6_read_data__read;
  wire [63:0] edge_list_ch_6_write_addr__din;
  wire edge_list_ch_6_write_addr__full_n;
  wire edge_list_ch_6_write_addr__write;
  wire [255:0] edge_list_ch_6_write_data__din;
  wire edge_list_ch_6_write_data__full_n;
  wire edge_list_ch_6_write_data__write;
  wire [7:0] edge_list_ch_6_write_resp__dout;
  wire edge_list_ch_6_write_resp__empty_n;
  wire edge_list_ch_6_write_resp__read;
  wire read_A_6__ap_start;
  wire read_A_6__ap_ready;
  wire read_A_6__ap_done;
  wire read_A_6__ap_idle;
  wire [31:0] read_A_7___NUM_A_LEN__q0;
  wire [31:0] read_A_7___P_N__q0;
  wire [63:0] read_A_7___edge_list_ch_7__q0;
  wire [63:0] edge_list_ch_7_read_addr__din;
  wire edge_list_ch_7_read_addr__full_n;
  wire edge_list_ch_7_read_addr__write;
  wire [255:0] edge_list_ch_7_read_data__dout;
  wire edge_list_ch_7_read_data__empty_n;
  wire edge_list_ch_7_read_data__read;
  wire [63:0] edge_list_ch_7_write_addr__din;
  wire edge_list_ch_7_write_addr__full_n;
  wire edge_list_ch_7_write_addr__write;
  wire [255:0] edge_list_ch_7_write_data__din;
  wire edge_list_ch_7_write_data__full_n;
  wire edge_list_ch_7_write_data__write;
  wire [7:0] edge_list_ch_7_write_resp__dout;
  wire edge_list_ch_7_write_resp__empty_n;
  wire edge_list_ch_7_write_resp__read;
  wire read_A_7__ap_start;
  wire read_A_7__ap_ready;
  wire read_A_7__ap_done;
  wire read_A_7__ap_idle;
  wire [31:0] read_A_8___NUM_A_LEN__q0;
  wire [31:0] read_A_8___P_N__q0;
  wire [63:0] read_A_8___edge_list_ch_8__q0;
  wire [63:0] edge_list_ch_8_read_addr__din;
  wire edge_list_ch_8_read_addr__full_n;
  wire edge_list_ch_8_read_addr__write;
  wire [255:0] edge_list_ch_8_read_data__dout;
  wire edge_list_ch_8_read_data__empty_n;
  wire edge_list_ch_8_read_data__read;
  wire [63:0] edge_list_ch_8_write_addr__din;
  wire edge_list_ch_8_write_addr__full_n;
  wire edge_list_ch_8_write_addr__write;
  wire [255:0] edge_list_ch_8_write_data__din;
  wire edge_list_ch_8_write_data__full_n;
  wire edge_list_ch_8_write_data__write;
  wire [7:0] edge_list_ch_8_write_resp__dout;
  wire edge_list_ch_8_write_resp__empty_n;
  wire edge_list_ch_8_write_resp__read;
  wire read_A_8__ap_start;
  wire read_A_8__ap_ready;
  wire read_A_8__ap_done;
  wire read_A_8__ap_idle;
  wire [31:0] read_A_9___NUM_A_LEN__q0;
  wire [31:0] read_A_9___P_N__q0;
  wire [63:0] read_A_9___edge_list_ch_9__q0;
  wire [63:0] edge_list_ch_9_read_addr__din;
  wire edge_list_ch_9_read_addr__full_n;
  wire edge_list_ch_9_read_addr__write;
  wire [255:0] edge_list_ch_9_read_data__dout;
  wire edge_list_ch_9_read_data__empty_n;
  wire edge_list_ch_9_read_data__read;
  wire [63:0] edge_list_ch_9_write_addr__din;
  wire edge_list_ch_9_write_addr__full_n;
  wire edge_list_ch_9_write_addr__write;
  wire [255:0] edge_list_ch_9_write_data__din;
  wire edge_list_ch_9_write_data__full_n;
  wire edge_list_ch_9_write_data__write;
  wire [7:0] edge_list_ch_9_write_resp__dout;
  wire edge_list_ch_9_write_resp__empty_n;
  wire edge_list_ch_9_write_resp__read;
  wire read_A_9__ap_start;
  wire read_A_9__ap_ready;
  wire read_A_9__ap_done;
  wire read_A_9__ap_idle;
  wire [31:0] read_A_10___NUM_A_LEN__q0;
  wire [31:0] read_A_10___P_N__q0;
  wire [63:0] read_A_10___edge_list_ch_10__q0;
  wire [63:0] edge_list_ch_10_read_addr__din;
  wire edge_list_ch_10_read_addr__full_n;
  wire edge_list_ch_10_read_addr__write;
  wire [255:0] edge_list_ch_10_read_data__dout;
  wire edge_list_ch_10_read_data__empty_n;
  wire edge_list_ch_10_read_data__read;
  wire [63:0] edge_list_ch_10_write_addr__din;
  wire edge_list_ch_10_write_addr__full_n;
  wire edge_list_ch_10_write_addr__write;
  wire [255:0] edge_list_ch_10_write_data__din;
  wire edge_list_ch_10_write_data__full_n;
  wire edge_list_ch_10_write_data__write;
  wire [7:0] edge_list_ch_10_write_resp__dout;
  wire edge_list_ch_10_write_resp__empty_n;
  wire edge_list_ch_10_write_resp__read;
  wire read_A_10__ap_start;
  wire read_A_10__ap_ready;
  wire read_A_10__ap_done;
  wire read_A_10__ap_idle;
  wire [31:0] read_A_11___NUM_A_LEN__q0;
  wire [31:0] read_A_11___P_N__q0;
  wire [63:0] read_A_11___edge_list_ch_11__q0;
  wire [63:0] edge_list_ch_11_read_addr__din;
  wire edge_list_ch_11_read_addr__full_n;
  wire edge_list_ch_11_read_addr__write;
  wire [255:0] edge_list_ch_11_read_data__dout;
  wire edge_list_ch_11_read_data__empty_n;
  wire edge_list_ch_11_read_data__read;
  wire [63:0] edge_list_ch_11_write_addr__din;
  wire edge_list_ch_11_write_addr__full_n;
  wire edge_list_ch_11_write_addr__write;
  wire [255:0] edge_list_ch_11_write_data__din;
  wire edge_list_ch_11_write_data__full_n;
  wire edge_list_ch_11_write_data__write;
  wire [7:0] edge_list_ch_11_write_resp__dout;
  wire edge_list_ch_11_write_resp__empty_n;
  wire edge_list_ch_11_write_resp__read;
  wire read_A_11__ap_start;
  wire read_A_11__ap_ready;
  wire read_A_11__ap_done;
  wire read_A_11__ap_idle;
  wire [31:0] read_A_12___NUM_A_LEN__q0;
  wire [31:0] read_A_12___P_N__q0;
  wire [63:0] read_A_12___edge_list_ch_12__q0;
  wire [63:0] edge_list_ch_12_read_addr__din;
  wire edge_list_ch_12_read_addr__full_n;
  wire edge_list_ch_12_read_addr__write;
  wire [255:0] edge_list_ch_12_read_data__dout;
  wire edge_list_ch_12_read_data__empty_n;
  wire edge_list_ch_12_read_data__read;
  wire [63:0] edge_list_ch_12_write_addr__din;
  wire edge_list_ch_12_write_addr__full_n;
  wire edge_list_ch_12_write_addr__write;
  wire [255:0] edge_list_ch_12_write_data__din;
  wire edge_list_ch_12_write_data__full_n;
  wire edge_list_ch_12_write_data__write;
  wire [7:0] edge_list_ch_12_write_resp__dout;
  wire edge_list_ch_12_write_resp__empty_n;
  wire edge_list_ch_12_write_resp__read;
  wire read_A_12__ap_start;
  wire read_A_12__ap_ready;
  wire read_A_12__ap_done;
  wire read_A_12__ap_idle;
  wire [31:0] read_A_13___NUM_A_LEN__q0;
  wire [31:0] read_A_13___P_N__q0;
  wire [63:0] read_A_13___edge_list_ch_13__q0;
  wire [63:0] edge_list_ch_13_read_addr__din;
  wire edge_list_ch_13_read_addr__full_n;
  wire edge_list_ch_13_read_addr__write;
  wire [255:0] edge_list_ch_13_read_data__dout;
  wire edge_list_ch_13_read_data__empty_n;
  wire edge_list_ch_13_read_data__read;
  wire [63:0] edge_list_ch_13_write_addr__din;
  wire edge_list_ch_13_write_addr__full_n;
  wire edge_list_ch_13_write_addr__write;
  wire [255:0] edge_list_ch_13_write_data__din;
  wire edge_list_ch_13_write_data__full_n;
  wire edge_list_ch_13_write_data__write;
  wire [7:0] edge_list_ch_13_write_resp__dout;
  wire edge_list_ch_13_write_resp__empty_n;
  wire edge_list_ch_13_write_resp__read;
  wire read_A_13__ap_start;
  wire read_A_13__ap_ready;
  wire read_A_13__ap_done;
  wire read_A_13__ap_idle;
  wire [31:0] read_A_14___NUM_A_LEN__q0;
  wire [31:0] read_A_14___P_N__q0;
  wire [63:0] read_A_14___edge_list_ch_14__q0;
  wire [63:0] edge_list_ch_14_read_addr__din;
  wire edge_list_ch_14_read_addr__full_n;
  wire edge_list_ch_14_read_addr__write;
  wire [255:0] edge_list_ch_14_read_data__dout;
  wire edge_list_ch_14_read_data__empty_n;
  wire edge_list_ch_14_read_data__read;
  wire [63:0] edge_list_ch_14_write_addr__din;
  wire edge_list_ch_14_write_addr__full_n;
  wire edge_list_ch_14_write_addr__write;
  wire [255:0] edge_list_ch_14_write_data__din;
  wire edge_list_ch_14_write_data__full_n;
  wire edge_list_ch_14_write_data__write;
  wire [7:0] edge_list_ch_14_write_resp__dout;
  wire edge_list_ch_14_write_resp__empty_n;
  wire edge_list_ch_14_write_resp__read;
  wire read_A_14__ap_start;
  wire read_A_14__ap_ready;
  wire read_A_14__ap_done;
  wire read_A_14__ap_idle;
  wire [31:0] read_A_15___NUM_A_LEN__q0;
  wire [31:0] read_A_15___P_N__q0;
  wire [63:0] read_A_15___edge_list_ch_15__q0;
  wire [63:0] edge_list_ch_15_read_addr__din;
  wire edge_list_ch_15_read_addr__full_n;
  wire edge_list_ch_15_read_addr__write;
  wire [255:0] edge_list_ch_15_read_data__dout;
  wire edge_list_ch_15_read_data__empty_n;
  wire edge_list_ch_15_read_data__read;
  wire [63:0] edge_list_ch_15_write_addr__din;
  wire edge_list_ch_15_write_addr__full_n;
  wire edge_list_ch_15_write_addr__write;
  wire [255:0] edge_list_ch_15_write_data__din;
  wire edge_list_ch_15_write_data__full_n;
  wire edge_list_ch_15_write_data__write;
  wire [7:0] edge_list_ch_15_write_resp__dout;
  wire edge_list_ch_15_write_resp__empty_n;
  wire edge_list_ch_15_write_resp__read;
  wire read_A_15__ap_start;
  wire read_A_15__ap_ready;
  wire read_A_15__ap_done;
  wire read_A_15__ap_idle;
  wire [31:0] read_A_16___NUM_A_LEN__q0;
  wire [31:0] read_A_16___P_N__q0;
  wire [63:0] read_A_16___edge_list_ch_16__q0;
  wire [63:0] edge_list_ch_16_read_addr__din;
  wire edge_list_ch_16_read_addr__full_n;
  wire edge_list_ch_16_read_addr__write;
  wire [255:0] edge_list_ch_16_read_data__dout;
  wire edge_list_ch_16_read_data__empty_n;
  wire edge_list_ch_16_read_data__read;
  wire [63:0] edge_list_ch_16_write_addr__din;
  wire edge_list_ch_16_write_addr__full_n;
  wire edge_list_ch_16_write_addr__write;
  wire [255:0] edge_list_ch_16_write_data__din;
  wire edge_list_ch_16_write_data__full_n;
  wire edge_list_ch_16_write_data__write;
  wire [7:0] edge_list_ch_16_write_resp__dout;
  wire edge_list_ch_16_write_resp__empty_n;
  wire edge_list_ch_16_write_resp__read;
  wire read_A_16__ap_start;
  wire read_A_16__ap_ready;
  wire read_A_16__ap_done;
  wire read_A_16__ap_idle;
  wire [31:0] read_A_17___NUM_A_LEN__q0;
  wire [31:0] read_A_17___P_N__q0;
  wire [63:0] read_A_17___edge_list_ch_17__q0;
  wire [63:0] edge_list_ch_17_read_addr__din;
  wire edge_list_ch_17_read_addr__full_n;
  wire edge_list_ch_17_read_addr__write;
  wire [255:0] edge_list_ch_17_read_data__dout;
  wire edge_list_ch_17_read_data__empty_n;
  wire edge_list_ch_17_read_data__read;
  wire [63:0] edge_list_ch_17_write_addr__din;
  wire edge_list_ch_17_write_addr__full_n;
  wire edge_list_ch_17_write_addr__write;
  wire [255:0] edge_list_ch_17_write_data__din;
  wire edge_list_ch_17_write_data__full_n;
  wire edge_list_ch_17_write_data__write;
  wire [7:0] edge_list_ch_17_write_resp__dout;
  wire edge_list_ch_17_write_resp__empty_n;
  wire edge_list_ch_17_write_resp__read;
  wire read_A_17__ap_start;
  wire read_A_17__ap_ready;
  wire read_A_17__ap_done;
  wire read_A_17__ap_idle;
  wire [31:0] read_A_18___NUM_A_LEN__q0;
  wire [31:0] read_A_18___P_N__q0;
  wire [63:0] read_A_18___edge_list_ch_18__q0;
  wire [63:0] edge_list_ch_18_read_addr__din;
  wire edge_list_ch_18_read_addr__full_n;
  wire edge_list_ch_18_read_addr__write;
  wire [255:0] edge_list_ch_18_read_data__dout;
  wire edge_list_ch_18_read_data__empty_n;
  wire edge_list_ch_18_read_data__read;
  wire [63:0] edge_list_ch_18_write_addr__din;
  wire edge_list_ch_18_write_addr__full_n;
  wire edge_list_ch_18_write_addr__write;
  wire [255:0] edge_list_ch_18_write_data__din;
  wire edge_list_ch_18_write_data__full_n;
  wire edge_list_ch_18_write_data__write;
  wire [7:0] edge_list_ch_18_write_resp__dout;
  wire edge_list_ch_18_write_resp__empty_n;
  wire edge_list_ch_18_write_resp__read;
  wire read_A_18__ap_start;
  wire read_A_18__ap_ready;
  wire read_A_18__ap_done;
  wire read_A_18__ap_idle;
  wire [31:0] read_A_19___NUM_A_LEN__q0;
  wire [31:0] read_A_19___P_N__q0;
  wire [63:0] read_A_19___edge_list_ch_19__q0;
  wire [63:0] edge_list_ch_19_read_addr__din;
  wire edge_list_ch_19_read_addr__full_n;
  wire edge_list_ch_19_read_addr__write;
  wire [255:0] edge_list_ch_19_read_data__dout;
  wire edge_list_ch_19_read_data__empty_n;
  wire edge_list_ch_19_read_data__read;
  wire [63:0] edge_list_ch_19_write_addr__din;
  wire edge_list_ch_19_write_addr__full_n;
  wire edge_list_ch_19_write_addr__write;
  wire [255:0] edge_list_ch_19_write_data__din;
  wire edge_list_ch_19_write_data__full_n;
  wire edge_list_ch_19_write_data__write;
  wire [7:0] edge_list_ch_19_write_resp__dout;
  wire edge_list_ch_19_write_resp__empty_n;
  wire edge_list_ch_19_write_resp__read;
  wire read_A_19__ap_start;
  wire read_A_19__ap_ready;
  wire read_A_19__ap_done;
  wire read_A_19__ap_idle;
  wire [31:0] read_A_20___NUM_A_LEN__q0;
  wire [31:0] read_A_20___P_N__q0;
  wire [63:0] read_A_20___edge_list_ch_20__q0;
  wire [63:0] edge_list_ch_20_read_addr__din;
  wire edge_list_ch_20_read_addr__full_n;
  wire edge_list_ch_20_read_addr__write;
  wire [255:0] edge_list_ch_20_read_data__dout;
  wire edge_list_ch_20_read_data__empty_n;
  wire edge_list_ch_20_read_data__read;
  wire [63:0] edge_list_ch_20_write_addr__din;
  wire edge_list_ch_20_write_addr__full_n;
  wire edge_list_ch_20_write_addr__write;
  wire [255:0] edge_list_ch_20_write_data__din;
  wire edge_list_ch_20_write_data__full_n;
  wire edge_list_ch_20_write_data__write;
  wire [7:0] edge_list_ch_20_write_resp__dout;
  wire edge_list_ch_20_write_resp__empty_n;
  wire edge_list_ch_20_write_resp__read;
  wire read_A_20__ap_start;
  wire read_A_20__ap_ready;
  wire read_A_20__ap_done;
  wire read_A_20__ap_idle;
  wire [31:0] read_A_21___NUM_A_LEN__q0;
  wire [31:0] read_A_21___P_N__q0;
  wire [63:0] read_A_21___edge_list_ch_21__q0;
  wire [63:0] edge_list_ch_21_read_addr__din;
  wire edge_list_ch_21_read_addr__full_n;
  wire edge_list_ch_21_read_addr__write;
  wire [255:0] edge_list_ch_21_read_data__dout;
  wire edge_list_ch_21_read_data__empty_n;
  wire edge_list_ch_21_read_data__read;
  wire [63:0] edge_list_ch_21_write_addr__din;
  wire edge_list_ch_21_write_addr__full_n;
  wire edge_list_ch_21_write_addr__write;
  wire [255:0] edge_list_ch_21_write_data__din;
  wire edge_list_ch_21_write_data__full_n;
  wire edge_list_ch_21_write_data__write;
  wire [7:0] edge_list_ch_21_write_resp__dout;
  wire edge_list_ch_21_write_resp__empty_n;
  wire edge_list_ch_21_write_resp__read;
  wire read_A_21__ap_start;
  wire read_A_21__ap_ready;
  wire read_A_21__ap_done;
  wire read_A_21__ap_idle;
  wire [31:0] read_A_22___NUM_A_LEN__q0;
  wire [31:0] read_A_22___P_N__q0;
  wire [63:0] read_A_22___edge_list_ch_22__q0;
  wire [63:0] edge_list_ch_22_read_addr__din;
  wire edge_list_ch_22_read_addr__full_n;
  wire edge_list_ch_22_read_addr__write;
  wire [255:0] edge_list_ch_22_read_data__dout;
  wire edge_list_ch_22_read_data__empty_n;
  wire edge_list_ch_22_read_data__read;
  wire [63:0] edge_list_ch_22_write_addr__din;
  wire edge_list_ch_22_write_addr__full_n;
  wire edge_list_ch_22_write_addr__write;
  wire [255:0] edge_list_ch_22_write_data__din;
  wire edge_list_ch_22_write_data__full_n;
  wire edge_list_ch_22_write_data__write;
  wire [7:0] edge_list_ch_22_write_resp__dout;
  wire edge_list_ch_22_write_resp__empty_n;
  wire edge_list_ch_22_write_resp__read;
  wire read_A_22__ap_start;
  wire read_A_22__ap_ready;
  wire read_A_22__ap_done;
  wire read_A_22__ap_idle;
  wire [31:0] read_A_23___NUM_A_LEN__q0;
  wire [31:0] read_A_23___P_N__q0;
  wire [63:0] read_A_23___edge_list_ch_23__q0;
  wire [63:0] edge_list_ch_23_read_addr__din;
  wire edge_list_ch_23_read_addr__full_n;
  wire edge_list_ch_23_read_addr__write;
  wire [255:0] edge_list_ch_23_read_data__dout;
  wire edge_list_ch_23_read_data__empty_n;
  wire edge_list_ch_23_read_data__read;
  wire [63:0] edge_list_ch_23_write_addr__din;
  wire edge_list_ch_23_write_addr__full_n;
  wire edge_list_ch_23_write_addr__write;
  wire [255:0] edge_list_ch_23_write_data__din;
  wire edge_list_ch_23_write_data__full_n;
  wire edge_list_ch_23_write_data__write;
  wire [7:0] edge_list_ch_23_write_resp__dout;
  wire edge_list_ch_23_write_resp__empty_n;
  wire edge_list_ch_23_write_resp__read;
  wire read_A_23__ap_start;
  wire read_A_23__ap_ready;
  wire read_A_23__ap_done;
  wire read_A_23__ap_idle;
  wire [31:0] read_A_24___NUM_A_LEN__q0;
  wire [31:0] read_A_24___P_N__q0;
  wire [63:0] read_A_24___edge_list_ch_24__q0;
  wire [63:0] edge_list_ch_24_read_addr__din;
  wire edge_list_ch_24_read_addr__full_n;
  wire edge_list_ch_24_read_addr__write;
  wire [255:0] edge_list_ch_24_read_data__dout;
  wire edge_list_ch_24_read_data__empty_n;
  wire edge_list_ch_24_read_data__read;
  wire [63:0] edge_list_ch_24_write_addr__din;
  wire edge_list_ch_24_write_addr__full_n;
  wire edge_list_ch_24_write_addr__write;
  wire [255:0] edge_list_ch_24_write_data__din;
  wire edge_list_ch_24_write_data__full_n;
  wire edge_list_ch_24_write_data__write;
  wire [7:0] edge_list_ch_24_write_resp__dout;
  wire edge_list_ch_24_write_resp__empty_n;
  wire edge_list_ch_24_write_resp__read;
  wire read_A_24__ap_start;
  wire read_A_24__ap_ready;
  wire read_A_24__ap_done;
  wire read_A_24__ap_idle;
  wire [31:0] read_A_25___NUM_A_LEN__q0;
  wire [31:0] read_A_25___P_N__q0;
  wire [63:0] read_A_25___edge_list_ch_25__q0;
  wire [63:0] edge_list_ch_25_read_addr__din;
  wire edge_list_ch_25_read_addr__full_n;
  wire edge_list_ch_25_read_addr__write;
  wire [255:0] edge_list_ch_25_read_data__dout;
  wire edge_list_ch_25_read_data__empty_n;
  wire edge_list_ch_25_read_data__read;
  wire [63:0] edge_list_ch_25_write_addr__din;
  wire edge_list_ch_25_write_addr__full_n;
  wire edge_list_ch_25_write_addr__write;
  wire [255:0] edge_list_ch_25_write_data__din;
  wire edge_list_ch_25_write_data__full_n;
  wire edge_list_ch_25_write_data__write;
  wire [7:0] edge_list_ch_25_write_resp__dout;
  wire edge_list_ch_25_write_resp__empty_n;
  wire edge_list_ch_25_write_resp__read;
  wire read_A_25__ap_start;
  wire read_A_25__ap_ready;
  wire read_A_25__ap_done;
  wire read_A_25__ap_idle;
  wire [31:0] read_A_26___NUM_A_LEN__q0;
  wire [31:0] read_A_26___P_N__q0;
  wire [63:0] read_A_26___edge_list_ch_26__q0;
  wire [63:0] edge_list_ch_26_read_addr__din;
  wire edge_list_ch_26_read_addr__full_n;
  wire edge_list_ch_26_read_addr__write;
  wire [255:0] edge_list_ch_26_read_data__dout;
  wire edge_list_ch_26_read_data__empty_n;
  wire edge_list_ch_26_read_data__read;
  wire [63:0] edge_list_ch_26_write_addr__din;
  wire edge_list_ch_26_write_addr__full_n;
  wire edge_list_ch_26_write_addr__write;
  wire [255:0] edge_list_ch_26_write_data__din;
  wire edge_list_ch_26_write_data__full_n;
  wire edge_list_ch_26_write_data__write;
  wire [7:0] edge_list_ch_26_write_resp__dout;
  wire edge_list_ch_26_write_resp__empty_n;
  wire edge_list_ch_26_write_resp__read;
  wire read_A_26__ap_start;
  wire read_A_26__ap_ready;
  wire read_A_26__ap_done;
  wire read_A_26__ap_idle;
  wire [31:0] read_A_27___NUM_A_LEN__q0;
  wire [31:0] read_A_27___P_N__q0;
  wire [63:0] read_A_27___edge_list_ch_27__q0;
  wire [63:0] edge_list_ch_27_read_addr__din;
  wire edge_list_ch_27_read_addr__full_n;
  wire edge_list_ch_27_read_addr__write;
  wire [255:0] edge_list_ch_27_read_data__dout;
  wire edge_list_ch_27_read_data__empty_n;
  wire edge_list_ch_27_read_data__read;
  wire [63:0] edge_list_ch_27_write_addr__din;
  wire edge_list_ch_27_write_addr__full_n;
  wire edge_list_ch_27_write_addr__write;
  wire [255:0] edge_list_ch_27_write_data__din;
  wire edge_list_ch_27_write_data__full_n;
  wire edge_list_ch_27_write_data__write;
  wire [7:0] edge_list_ch_27_write_resp__dout;
  wire edge_list_ch_27_write_resp__empty_n;
  wire edge_list_ch_27_write_resp__read;
  wire read_A_27__ap_start;
  wire read_A_27__ap_ready;
  wire read_A_27__ap_done;
  wire read_A_27__ap_idle;
  wire [31:0] read_A_28___NUM_A_LEN__q0;
  wire [31:0] read_A_28___P_N__q0;
  wire [63:0] read_A_28___edge_list_ch_28__q0;
  wire [63:0] edge_list_ch_28_read_addr__din;
  wire edge_list_ch_28_read_addr__full_n;
  wire edge_list_ch_28_read_addr__write;
  wire [255:0] edge_list_ch_28_read_data__dout;
  wire edge_list_ch_28_read_data__empty_n;
  wire edge_list_ch_28_read_data__read;
  wire [63:0] edge_list_ch_28_write_addr__din;
  wire edge_list_ch_28_write_addr__full_n;
  wire edge_list_ch_28_write_addr__write;
  wire [255:0] edge_list_ch_28_write_data__din;
  wire edge_list_ch_28_write_data__full_n;
  wire edge_list_ch_28_write_data__write;
  wire [7:0] edge_list_ch_28_write_resp__dout;
  wire edge_list_ch_28_write_resp__empty_n;
  wire edge_list_ch_28_write_resp__read;
  wire read_A_28__ap_start;
  wire read_A_28__ap_ready;
  wire read_A_28__ap_done;
  wire read_A_28__ap_idle;
  wire [31:0] read_A_29___NUM_A_LEN__q0;
  wire [31:0] read_A_29___P_N__q0;
  wire [63:0] read_A_29___edge_list_ch_29__q0;
  wire [63:0] edge_list_ch_29_read_addr__din;
  wire edge_list_ch_29_read_addr__full_n;
  wire edge_list_ch_29_read_addr__write;
  wire [255:0] edge_list_ch_29_read_data__dout;
  wire edge_list_ch_29_read_data__empty_n;
  wire edge_list_ch_29_read_data__read;
  wire [63:0] edge_list_ch_29_write_addr__din;
  wire edge_list_ch_29_write_addr__full_n;
  wire edge_list_ch_29_write_addr__write;
  wire [255:0] edge_list_ch_29_write_data__din;
  wire edge_list_ch_29_write_data__full_n;
  wire edge_list_ch_29_write_data__write;
  wire [7:0] edge_list_ch_29_write_resp__dout;
  wire edge_list_ch_29_write_resp__empty_n;
  wire edge_list_ch_29_write_resp__read;
  wire read_A_29__ap_start;
  wire read_A_29__ap_ready;
  wire read_A_29__ap_done;
  wire read_A_29__ap_idle;
  wire [31:0] read_A_30___NUM_A_LEN__q0;
  wire [31:0] read_A_30___P_N__q0;
  wire [63:0] read_A_30___edge_list_ch_30__q0;
  wire [63:0] edge_list_ch_30_read_addr__din;
  wire edge_list_ch_30_read_addr__full_n;
  wire edge_list_ch_30_read_addr__write;
  wire [255:0] edge_list_ch_30_read_data__dout;
  wire edge_list_ch_30_read_data__empty_n;
  wire edge_list_ch_30_read_data__read;
  wire [63:0] edge_list_ch_30_write_addr__din;
  wire edge_list_ch_30_write_addr__full_n;
  wire edge_list_ch_30_write_addr__write;
  wire [255:0] edge_list_ch_30_write_data__din;
  wire edge_list_ch_30_write_data__full_n;
  wire edge_list_ch_30_write_data__write;
  wire [7:0] edge_list_ch_30_write_resp__dout;
  wire edge_list_ch_30_write_resp__empty_n;
  wire edge_list_ch_30_write_resp__read;
  wire read_A_30__ap_start;
  wire read_A_30__ap_ready;
  wire read_A_30__ap_done;
  wire read_A_30__ap_idle;
  wire [31:0] read_A_31___NUM_A_LEN__q0;
  wire [31:0] read_A_31___P_N__q0;
  wire [63:0] read_A_31___edge_list_ch_31__q0;
  wire [63:0] edge_list_ch_31_read_addr__din;
  wire edge_list_ch_31_read_addr__full_n;
  wire edge_list_ch_31_read_addr__write;
  wire [255:0] edge_list_ch_31_read_data__dout;
  wire edge_list_ch_31_read_data__empty_n;
  wire edge_list_ch_31_read_data__read;
  wire [63:0] edge_list_ch_31_write_addr__din;
  wire edge_list_ch_31_write_addr__full_n;
  wire edge_list_ch_31_write_addr__write;
  wire [255:0] edge_list_ch_31_write_data__din;
  wire edge_list_ch_31_write_data__full_n;
  wire edge_list_ch_31_write_data__write;
  wire [7:0] edge_list_ch_31_write_resp__dout;
  wire edge_list_ch_31_write_resp__empty_n;
  wire edge_list_ch_31_write_resp__read;
  wire read_A_31__ap_start;
  wire read_A_31__ap_ready;
  wire read_A_31__ap_done;
  wire read_A_31__ap_idle;
  wire [31:0] read_A_32___NUM_A_LEN__q0;
  wire [31:0] read_A_32___P_N__q0;
  wire [63:0] read_A_32___edge_list_ch_32__q0;
  wire [63:0] edge_list_ch_32_read_addr__din;
  wire edge_list_ch_32_read_addr__full_n;
  wire edge_list_ch_32_read_addr__write;
  wire [255:0] edge_list_ch_32_read_data__dout;
  wire edge_list_ch_32_read_data__empty_n;
  wire edge_list_ch_32_read_data__read;
  wire [63:0] edge_list_ch_32_write_addr__din;
  wire edge_list_ch_32_write_addr__full_n;
  wire edge_list_ch_32_write_addr__write;
  wire [255:0] edge_list_ch_32_write_data__din;
  wire edge_list_ch_32_write_data__full_n;
  wire edge_list_ch_32_write_data__write;
  wire [7:0] edge_list_ch_32_write_resp__dout;
  wire edge_list_ch_32_write_resp__empty_n;
  wire edge_list_ch_32_write_resp__read;
  wire read_A_32__ap_start;
  wire read_A_32__ap_ready;
  wire read_A_32__ap_done;
  wire read_A_32__ap_idle;
  wire [31:0] read_A_33___NUM_A_LEN__q0;
  wire [31:0] read_A_33___P_N__q0;
  wire [63:0] read_A_33___edge_list_ch_33__q0;
  wire [63:0] edge_list_ch_33_read_addr__din;
  wire edge_list_ch_33_read_addr__full_n;
  wire edge_list_ch_33_read_addr__write;
  wire [255:0] edge_list_ch_33_read_data__dout;
  wire edge_list_ch_33_read_data__empty_n;
  wire edge_list_ch_33_read_data__read;
  wire [63:0] edge_list_ch_33_write_addr__din;
  wire edge_list_ch_33_write_addr__full_n;
  wire edge_list_ch_33_write_addr__write;
  wire [255:0] edge_list_ch_33_write_data__din;
  wire edge_list_ch_33_write_data__full_n;
  wire edge_list_ch_33_write_data__write;
  wire [7:0] edge_list_ch_33_write_resp__dout;
  wire edge_list_ch_33_write_resp__empty_n;
  wire edge_list_ch_33_write_resp__read;
  wire read_A_33__ap_start;
  wire read_A_33__ap_ready;
  wire read_A_33__ap_done;
  wire read_A_33__ap_idle;
  wire [31:0] read_A_34___NUM_A_LEN__q0;
  wire [31:0] read_A_34___P_N__q0;
  wire [63:0] read_A_34___edge_list_ch_34__q0;
  wire [63:0] edge_list_ch_34_read_addr__din;
  wire edge_list_ch_34_read_addr__full_n;
  wire edge_list_ch_34_read_addr__write;
  wire [255:0] edge_list_ch_34_read_data__dout;
  wire edge_list_ch_34_read_data__empty_n;
  wire edge_list_ch_34_read_data__read;
  wire [63:0] edge_list_ch_34_write_addr__din;
  wire edge_list_ch_34_write_addr__full_n;
  wire edge_list_ch_34_write_addr__write;
  wire [255:0] edge_list_ch_34_write_data__din;
  wire edge_list_ch_34_write_data__full_n;
  wire edge_list_ch_34_write_data__write;
  wire [7:0] edge_list_ch_34_write_resp__dout;
  wire edge_list_ch_34_write_resp__empty_n;
  wire edge_list_ch_34_write_resp__read;
  wire read_A_34__ap_start;
  wire read_A_34__ap_ready;
  wire read_A_34__ap_done;
  wire read_A_34__ap_idle;
  wire [31:0] read_A_35___NUM_A_LEN__q0;
  wire [31:0] read_A_35___P_N__q0;
  wire [63:0] read_A_35___edge_list_ch_35__q0;
  wire [63:0] edge_list_ch_35_read_addr__din;
  wire edge_list_ch_35_read_addr__full_n;
  wire edge_list_ch_35_read_addr__write;
  wire [255:0] edge_list_ch_35_read_data__dout;
  wire edge_list_ch_35_read_data__empty_n;
  wire edge_list_ch_35_read_data__read;
  wire [63:0] edge_list_ch_35_write_addr__din;
  wire edge_list_ch_35_write_addr__full_n;
  wire edge_list_ch_35_write_addr__write;
  wire [255:0] edge_list_ch_35_write_data__din;
  wire edge_list_ch_35_write_data__full_n;
  wire edge_list_ch_35_write_data__write;
  wire [7:0] edge_list_ch_35_write_resp__dout;
  wire edge_list_ch_35_write_resp__empty_n;
  wire edge_list_ch_35_write_resp__read;
  wire read_A_35__ap_start;
  wire read_A_35__ap_ready;
  wire read_A_35__ap_done;
  wire read_A_35__ap_idle;
  wire [31:0] read_A_36___NUM_A_LEN__q0;
  wire [31:0] read_A_36___P_N__q0;
  wire [63:0] read_A_36___edge_list_ch_36__q0;
  wire [63:0] edge_list_ch_36_read_addr__din;
  wire edge_list_ch_36_read_addr__full_n;
  wire edge_list_ch_36_read_addr__write;
  wire [255:0] edge_list_ch_36_read_data__dout;
  wire edge_list_ch_36_read_data__empty_n;
  wire edge_list_ch_36_read_data__read;
  wire [63:0] edge_list_ch_36_write_addr__din;
  wire edge_list_ch_36_write_addr__full_n;
  wire edge_list_ch_36_write_addr__write;
  wire [255:0] edge_list_ch_36_write_data__din;
  wire edge_list_ch_36_write_data__full_n;
  wire edge_list_ch_36_write_data__write;
  wire [7:0] edge_list_ch_36_write_resp__dout;
  wire edge_list_ch_36_write_resp__empty_n;
  wire edge_list_ch_36_write_resp__read;
  wire read_A_36__ap_start;
  wire read_A_36__ap_ready;
  wire read_A_36__ap_done;
  wire read_A_36__ap_idle;
  wire [31:0] read_A_37___NUM_A_LEN__q0;
  wire [31:0] read_A_37___P_N__q0;
  wire [63:0] read_A_37___edge_list_ch_37__q0;
  wire [63:0] edge_list_ch_37_read_addr__din;
  wire edge_list_ch_37_read_addr__full_n;
  wire edge_list_ch_37_read_addr__write;
  wire [255:0] edge_list_ch_37_read_data__dout;
  wire edge_list_ch_37_read_data__empty_n;
  wire edge_list_ch_37_read_data__read;
  wire [63:0] edge_list_ch_37_write_addr__din;
  wire edge_list_ch_37_write_addr__full_n;
  wire edge_list_ch_37_write_addr__write;
  wire [255:0] edge_list_ch_37_write_data__din;
  wire edge_list_ch_37_write_data__full_n;
  wire edge_list_ch_37_write_data__write;
  wire [7:0] edge_list_ch_37_write_resp__dout;
  wire edge_list_ch_37_write_resp__empty_n;
  wire edge_list_ch_37_write_resp__read;
  wire read_A_37__ap_start;
  wire read_A_37__ap_ready;
  wire read_A_37__ap_done;
  wire read_A_37__ap_idle;
  wire [31:0] read_A_38___NUM_A_LEN__q0;
  wire [31:0] read_A_38___P_N__q0;
  wire [63:0] read_A_38___edge_list_ch_38__q0;
  wire [63:0] edge_list_ch_38_read_addr__din;
  wire edge_list_ch_38_read_addr__full_n;
  wire edge_list_ch_38_read_addr__write;
  wire [255:0] edge_list_ch_38_read_data__dout;
  wire edge_list_ch_38_read_data__empty_n;
  wire edge_list_ch_38_read_data__read;
  wire [63:0] edge_list_ch_38_write_addr__din;
  wire edge_list_ch_38_write_addr__full_n;
  wire edge_list_ch_38_write_addr__write;
  wire [255:0] edge_list_ch_38_write_data__din;
  wire edge_list_ch_38_write_data__full_n;
  wire edge_list_ch_38_write_data__write;
  wire [7:0] edge_list_ch_38_write_resp__dout;
  wire edge_list_ch_38_write_resp__empty_n;
  wire edge_list_ch_38_write_resp__read;
  wire read_A_38__ap_start;
  wire read_A_38__ap_ready;
  wire read_A_38__ap_done;
  wire read_A_38__ap_idle;
  wire [31:0] read_A_39___NUM_A_LEN__q0;
  wire [31:0] read_A_39___P_N__q0;
  wire [63:0] read_A_39___edge_list_ch_39__q0;
  wire [63:0] edge_list_ch_39_read_addr__din;
  wire edge_list_ch_39_read_addr__full_n;
  wire edge_list_ch_39_read_addr__write;
  wire [255:0] edge_list_ch_39_read_data__dout;
  wire edge_list_ch_39_read_data__empty_n;
  wire edge_list_ch_39_read_data__read;
  wire [63:0] edge_list_ch_39_write_addr__din;
  wire edge_list_ch_39_write_addr__full_n;
  wire edge_list_ch_39_write_addr__write;
  wire [255:0] edge_list_ch_39_write_data__din;
  wire edge_list_ch_39_write_data__full_n;
  wire edge_list_ch_39_write_data__write;
  wire [7:0] edge_list_ch_39_write_resp__dout;
  wire edge_list_ch_39_write_resp__empty_n;
  wire edge_list_ch_39_write_resp__read;
  wire read_A_39__ap_start;
  wire read_A_39__ap_ready;
  wire read_A_39__ap_done;
  wire read_A_39__ap_idle;
  wire [31:0] read_A_40___NUM_A_LEN__q0;
  wire [31:0] read_A_40___P_N__q0;
  wire [63:0] read_A_40___edge_list_ch_40__q0;
  wire [63:0] edge_list_ch_40_read_addr__din;
  wire edge_list_ch_40_read_addr__full_n;
  wire edge_list_ch_40_read_addr__write;
  wire [255:0] edge_list_ch_40_read_data__dout;
  wire edge_list_ch_40_read_data__empty_n;
  wire edge_list_ch_40_read_data__read;
  wire [63:0] edge_list_ch_40_write_addr__din;
  wire edge_list_ch_40_write_addr__full_n;
  wire edge_list_ch_40_write_addr__write;
  wire [255:0] edge_list_ch_40_write_data__din;
  wire edge_list_ch_40_write_data__full_n;
  wire edge_list_ch_40_write_data__write;
  wire [7:0] edge_list_ch_40_write_resp__dout;
  wire edge_list_ch_40_write_resp__empty_n;
  wire edge_list_ch_40_write_resp__read;
  wire read_A_40__ap_start;
  wire read_A_40__ap_ready;
  wire read_A_40__ap_done;
  wire read_A_40__ap_idle;
  wire [31:0] read_A_41___NUM_A_LEN__q0;
  wire [31:0] read_A_41___P_N__q0;
  wire [63:0] read_A_41___edge_list_ch_41__q0;
  wire [63:0] edge_list_ch_41_read_addr__din;
  wire edge_list_ch_41_read_addr__full_n;
  wire edge_list_ch_41_read_addr__write;
  wire [255:0] edge_list_ch_41_read_data__dout;
  wire edge_list_ch_41_read_data__empty_n;
  wire edge_list_ch_41_read_data__read;
  wire [63:0] edge_list_ch_41_write_addr__din;
  wire edge_list_ch_41_write_addr__full_n;
  wire edge_list_ch_41_write_addr__write;
  wire [255:0] edge_list_ch_41_write_data__din;
  wire edge_list_ch_41_write_data__full_n;
  wire edge_list_ch_41_write_data__write;
  wire [7:0] edge_list_ch_41_write_resp__dout;
  wire edge_list_ch_41_write_resp__empty_n;
  wire edge_list_ch_41_write_resp__read;
  wire read_A_41__ap_start;
  wire read_A_41__ap_ready;
  wire read_A_41__ap_done;
  wire read_A_41__ap_idle;
  wire [31:0] read_A_42___NUM_A_LEN__q0;
  wire [31:0] read_A_42___P_N__q0;
  wire [63:0] read_A_42___edge_list_ch_42__q0;
  wire [63:0] edge_list_ch_42_read_addr__din;
  wire edge_list_ch_42_read_addr__full_n;
  wire edge_list_ch_42_read_addr__write;
  wire [255:0] edge_list_ch_42_read_data__dout;
  wire edge_list_ch_42_read_data__empty_n;
  wire edge_list_ch_42_read_data__read;
  wire [63:0] edge_list_ch_42_write_addr__din;
  wire edge_list_ch_42_write_addr__full_n;
  wire edge_list_ch_42_write_addr__write;
  wire [255:0] edge_list_ch_42_write_data__din;
  wire edge_list_ch_42_write_data__full_n;
  wire edge_list_ch_42_write_data__write;
  wire [7:0] edge_list_ch_42_write_resp__dout;
  wire edge_list_ch_42_write_resp__empty_n;
  wire edge_list_ch_42_write_resp__read;
  wire read_A_42__ap_start;
  wire read_A_42__ap_ready;
  wire read_A_42__ap_done;
  wire read_A_42__ap_idle;
  wire [31:0] read_A_43___NUM_A_LEN__q0;
  wire [31:0] read_A_43___P_N__q0;
  wire [63:0] read_A_43___edge_list_ch_43__q0;
  wire [63:0] edge_list_ch_43_read_addr__din;
  wire edge_list_ch_43_read_addr__full_n;
  wire edge_list_ch_43_read_addr__write;
  wire [255:0] edge_list_ch_43_read_data__dout;
  wire edge_list_ch_43_read_data__empty_n;
  wire edge_list_ch_43_read_data__read;
  wire [63:0] edge_list_ch_43_write_addr__din;
  wire edge_list_ch_43_write_addr__full_n;
  wire edge_list_ch_43_write_addr__write;
  wire [255:0] edge_list_ch_43_write_data__din;
  wire edge_list_ch_43_write_data__full_n;
  wire edge_list_ch_43_write_data__write;
  wire [7:0] edge_list_ch_43_write_resp__dout;
  wire edge_list_ch_43_write_resp__empty_n;
  wire edge_list_ch_43_write_resp__read;
  wire read_A_43__ap_start;
  wire read_A_43__ap_ready;
  wire read_A_43__ap_done;
  wire read_A_43__ap_idle;
  wire [31:0] read_A_44___NUM_A_LEN__q0;
  wire [31:0] read_A_44___P_N__q0;
  wire [63:0] read_A_44___edge_list_ch_44__q0;
  wire [63:0] edge_list_ch_44_read_addr__din;
  wire edge_list_ch_44_read_addr__full_n;
  wire edge_list_ch_44_read_addr__write;
  wire [255:0] edge_list_ch_44_read_data__dout;
  wire edge_list_ch_44_read_data__empty_n;
  wire edge_list_ch_44_read_data__read;
  wire [63:0] edge_list_ch_44_write_addr__din;
  wire edge_list_ch_44_write_addr__full_n;
  wire edge_list_ch_44_write_addr__write;
  wire [255:0] edge_list_ch_44_write_data__din;
  wire edge_list_ch_44_write_data__full_n;
  wire edge_list_ch_44_write_data__write;
  wire [7:0] edge_list_ch_44_write_resp__dout;
  wire edge_list_ch_44_write_resp__empty_n;
  wire edge_list_ch_44_write_resp__read;
  wire read_A_44__ap_start;
  wire read_A_44__ap_ready;
  wire read_A_44__ap_done;
  wire read_A_44__ap_idle;
  wire [31:0] read_A_45___NUM_A_LEN__q0;
  wire [31:0] read_A_45___P_N__q0;
  wire [63:0] read_A_45___edge_list_ch_45__q0;
  wire [63:0] edge_list_ch_45_read_addr__din;
  wire edge_list_ch_45_read_addr__full_n;
  wire edge_list_ch_45_read_addr__write;
  wire [255:0] edge_list_ch_45_read_data__dout;
  wire edge_list_ch_45_read_data__empty_n;
  wire edge_list_ch_45_read_data__read;
  wire [63:0] edge_list_ch_45_write_addr__din;
  wire edge_list_ch_45_write_addr__full_n;
  wire edge_list_ch_45_write_addr__write;
  wire [255:0] edge_list_ch_45_write_data__din;
  wire edge_list_ch_45_write_data__full_n;
  wire edge_list_ch_45_write_data__write;
  wire [7:0] edge_list_ch_45_write_resp__dout;
  wire edge_list_ch_45_write_resp__empty_n;
  wire edge_list_ch_45_write_resp__read;
  wire read_A_45__ap_start;
  wire read_A_45__ap_ready;
  wire read_A_45__ap_done;
  wire read_A_45__ap_idle;
  wire [31:0] read_A_46___NUM_A_LEN__q0;
  wire [31:0] read_A_46___P_N__q0;
  wire [63:0] read_A_46___edge_list_ch_46__q0;
  wire [63:0] edge_list_ch_46_read_addr__din;
  wire edge_list_ch_46_read_addr__full_n;
  wire edge_list_ch_46_read_addr__write;
  wire [255:0] edge_list_ch_46_read_data__dout;
  wire edge_list_ch_46_read_data__empty_n;
  wire edge_list_ch_46_read_data__read;
  wire [63:0] edge_list_ch_46_write_addr__din;
  wire edge_list_ch_46_write_addr__full_n;
  wire edge_list_ch_46_write_addr__write;
  wire [255:0] edge_list_ch_46_write_data__din;
  wire edge_list_ch_46_write_data__full_n;
  wire edge_list_ch_46_write_data__write;
  wire [7:0] edge_list_ch_46_write_resp__dout;
  wire edge_list_ch_46_write_resp__empty_n;
  wire edge_list_ch_46_write_resp__read;
  wire read_A_46__ap_start;
  wire read_A_46__ap_ready;
  wire read_A_46__ap_done;
  wire read_A_46__ap_idle;
  wire [31:0] read_A_47___NUM_A_LEN__q0;
  wire [31:0] read_A_47___P_N__q0;
  wire [63:0] read_A_47___edge_list_ch_47__q0;
  wire [63:0] edge_list_ch_47_read_addr__din;
  wire edge_list_ch_47_read_addr__full_n;
  wire edge_list_ch_47_read_addr__write;
  wire [255:0] edge_list_ch_47_read_data__dout;
  wire edge_list_ch_47_read_data__empty_n;
  wire edge_list_ch_47_read_data__read;
  wire [63:0] edge_list_ch_47_write_addr__din;
  wire edge_list_ch_47_write_addr__full_n;
  wire edge_list_ch_47_write_addr__write;
  wire [255:0] edge_list_ch_47_write_data__din;
  wire edge_list_ch_47_write_data__full_n;
  wire edge_list_ch_47_write_data__write;
  wire [7:0] edge_list_ch_47_write_resp__dout;
  wire edge_list_ch_47_write_resp__empty_n;
  wire edge_list_ch_47_write_resp__read;
  wire read_A_47__ap_start;
  wire read_A_47__ap_ready;
  wire read_A_47__ap_done;
  wire read_A_47__ap_idle;
  wire [31:0] read_X_0___K__q0;
  wire [31:0] read_X_0___P_N__q0;
  wire [63:0] read_X_0___vec_X__q0;
  wire [63:0] vec_X_read_addr__din;
  wire vec_X_read_addr__full_n;
  wire vec_X_read_addr__write;
  wire [255:0] vec_X_read_data__dout;
  wire vec_X_read_data__empty_n;
  wire vec_X_read_data__read;
  wire [63:0] vec_X_write_addr__din;
  wire vec_X_write_addr__full_n;
  wire vec_X_write_addr__write;
  wire [255:0] vec_X_write_data__din;
  wire vec_X_write_data__full_n;
  wire vec_X_write_data__write;
  wire [7:0] vec_X_write_resp__dout;
  wire vec_X_write_resp__empty_n;
  wire vec_X_write_resp__read;
  wire read_X_0__ap_start;
  wire read_X_0__ap_ready;
  wire read_X_0__ap_done;
  wire read_X_0__ap_idle;
  wire [31:0] read_Y_0___M__q0;
  wire [31:0] read_Y_0___P_N__q0;
  wire [63:0] read_Y_0___vec_Y__q0;
  wire [63:0] vec_Y_read_addr__din;
  wire vec_Y_read_addr__full_n;
  wire vec_Y_read_addr__write;
  wire [255:0] vec_Y_read_data__dout;
  wire vec_Y_read_data__empty_n;
  wire vec_Y_read_data__read;
  wire [63:0] vec_Y_write_addr__din;
  wire vec_Y_write_addr__full_n;
  wire vec_Y_write_addr__write;
  wire [255:0] vec_Y_write_data__din;
  wire vec_Y_write_data__full_n;
  wire vec_Y_write_data__write;
  wire [7:0] vec_Y_write_resp__dout;
  wire vec_Y_write_resp__empty_n;
  wire vec_Y_write_resp__read;
  wire read_Y_0__ap_start;
  wire read_Y_0__ap_ready;
  wire read_Y_0__ap_done;
  wire read_Y_0__ap_idle;
  wire [31:0] read_edge_list_ptr_0___K__q0;
  wire [31:0] read_edge_list_ptr_0___M__q0;
  wire [31:0] read_edge_list_ptr_0___NUM_ITE__q0;
  wire [31:0] read_edge_list_ptr_0___P_N__q0;
  wire [63:0] read_edge_list_ptr_0___edge_list_ptr__q0;
  wire [63:0] edge_list_ptr_read_addr__din;
  wire edge_list_ptr_read_addr__full_n;
  wire edge_list_ptr_read_addr__write;
  wire [31:0] edge_list_ptr_read_data__dout;
  wire edge_list_ptr_read_data__empty_n;
  wire edge_list_ptr_read_data__read;
  wire [63:0] edge_list_ptr_write_addr__din;
  wire edge_list_ptr_write_addr__full_n;
  wire edge_list_ptr_write_addr__write;
  wire [31:0] edge_list_ptr_write_data__din;
  wire edge_list_ptr_write_data__full_n;
  wire edge_list_ptr_write_data__write;
  wire [7:0] edge_list_ptr_write_resp__dout;
  wire edge_list_ptr_write_resp__empty_n;
  wire edge_list_ptr_write_resp__read;
  wire read_edge_list_ptr_0__ap_start;
  wire read_edge_list_ptr_0__ap_ready;
  wire read_edge_list_ptr_0__ap_done;
  wire read_edge_list_ptr_0__ap_idle;
  wire [31:0] write_Y_0___M__q0;
  wire [31:0] write_Y_0___P_N__q0;
  wire [63:0] write_Y_0___vec_Y_out__q0;
  wire [63:0] vec_Y_out_read_addr__din;
  wire vec_Y_out_read_addr__full_n;
  wire vec_Y_out_read_addr__write;
  wire [255:0] vec_Y_out_read_data__dout;
  wire vec_Y_out_read_data__empty_n;
  wire vec_Y_out_read_data__read;
  wire [63:0] vec_Y_out_write_addr__din;
  wire vec_Y_out_write_addr__full_n;
  wire vec_Y_out_write_addr__write;
  wire [255:0] vec_Y_out_write_data__din;
  wire vec_Y_out_write_data__full_n;
  wire vec_Y_out_write_data__write;
  wire [7:0] vec_Y_out_write_resp__dout;
  wire vec_Y_out_write_resp__empty_n;
  wire vec_Y_out_write_resp__read;
  wire write_Y_0__ap_start;
  wire write_Y_0__ap_ready;
  wire write_Y_0__ap_done;
  wire write_Y_0__ap_idle;
  wire ap_rst_n_inv;
  wire ap_done;
  wire ap_idle;
  wire ap_ready;
  assign ap_rst_n_inv = (~ap_rst_n);
  assign control_s_axi_U_ACLK = ap_clk;
  assign control_s_axi_U_ACLK_EN = 1'b1;
  assign control_s_axi_U_ARADDR = s_axi_control_ARADDR;
  assign control_s_axi_U_ARESET = ap_rst_n_inv;
  assign s_axi_control_ARREADY = control_s_axi_U_ARREADY;
  assign control_s_axi_U_ARVALID = s_axi_control_ARVALID;
  assign control_s_axi_U_AWADDR = s_axi_control_AWADDR;
  assign s_axi_control_AWREADY = control_s_axi_U_AWREADY;
  assign control_s_axi_U_AWVALID = s_axi_control_AWVALID;
  assign control_s_axi_U_BREADY = s_axi_control_BREADY;
  assign s_axi_control_BRESP = control_s_axi_U_BRESP;
  assign s_axi_control_BVALID = control_s_axi_U_BVALID;
  assign K = control_s_axi_U_K;
  assign M = control_s_axi_U_M;
  assign NUM_A_LEN = control_s_axi_U_NUM_A_LEN;
  assign NUM_ITE = control_s_axi_U_NUM_ITE;
  assign P_N = control_s_axi_U_P_N;
  assign s_axi_control_RDATA = control_s_axi_U_RDATA;
  assign control_s_axi_U_RREADY = s_axi_control_RREADY;
  assign s_axi_control_RRESP = control_s_axi_U_RRESP;
  assign s_axi_control_RVALID = control_s_axi_U_RVALID;
  assign control_s_axi_U_WDATA = s_axi_control_WDATA;
  assign s_axi_control_WREADY = control_s_axi_U_WREADY;
  assign control_s_axi_U_WSTRB = s_axi_control_WSTRB;
  assign control_s_axi_U_WVALID = s_axi_control_WVALID;
  assign alpha_u = control_s_axi_U_alpha_u;
  assign control_s_axi_U_ap_done = ap_done;
  assign control_s_axi_U_ap_idle = ap_idle;
  assign control_s_axi_U_ap_ready = ap_ready;
  assign ap_start = control_s_axi_U_ap_start;
  assign beta_u = control_s_axi_U_beta_u;
  assign edge_list_ch_0 = control_s_axi_U_edge_list_ch_0;
  assign edge_list_ch_1 = control_s_axi_U_edge_list_ch_1;
  assign edge_list_ch_10 = control_s_axi_U_edge_list_ch_10;
  assign edge_list_ch_11 = control_s_axi_U_edge_list_ch_11;
  assign edge_list_ch_12 = control_s_axi_U_edge_list_ch_12;
  assign edge_list_ch_13 = control_s_axi_U_edge_list_ch_13;
  assign edge_list_ch_14 = control_s_axi_U_edge_list_ch_14;
  assign edge_list_ch_15 = control_s_axi_U_edge_list_ch_15;
  assign edge_list_ch_16 = control_s_axi_U_edge_list_ch_16;
  assign edge_list_ch_17 = control_s_axi_U_edge_list_ch_17;
  assign edge_list_ch_18 = control_s_axi_U_edge_list_ch_18;
  assign edge_list_ch_19 = control_s_axi_U_edge_list_ch_19;
  assign edge_list_ch_2 = control_s_axi_U_edge_list_ch_2;
  assign edge_list_ch_20 = control_s_axi_U_edge_list_ch_20;
  assign edge_list_ch_21 = control_s_axi_U_edge_list_ch_21;
  assign edge_list_ch_22 = control_s_axi_U_edge_list_ch_22;
  assign edge_list_ch_23 = control_s_axi_U_edge_list_ch_23;
  assign edge_list_ch_24 = control_s_axi_U_edge_list_ch_24;
  assign edge_list_ch_25 = control_s_axi_U_edge_list_ch_25;
  assign edge_list_ch_26 = control_s_axi_U_edge_list_ch_26;
  assign edge_list_ch_27 = control_s_axi_U_edge_list_ch_27;
  assign edge_list_ch_28 = control_s_axi_U_edge_list_ch_28;
  assign edge_list_ch_29 = control_s_axi_U_edge_list_ch_29;
  assign edge_list_ch_3 = control_s_axi_U_edge_list_ch_3;
  assign edge_list_ch_30 = control_s_axi_U_edge_list_ch_30;
  assign edge_list_ch_31 = control_s_axi_U_edge_list_ch_31;
  assign edge_list_ch_32 = control_s_axi_U_edge_list_ch_32;
  assign edge_list_ch_33 = control_s_axi_U_edge_list_ch_33;
  assign edge_list_ch_34 = control_s_axi_U_edge_list_ch_34;
  assign edge_list_ch_35 = control_s_axi_U_edge_list_ch_35;
  assign edge_list_ch_36 = control_s_axi_U_edge_list_ch_36;
  assign edge_list_ch_37 = control_s_axi_U_edge_list_ch_37;
  assign edge_list_ch_38 = control_s_axi_U_edge_list_ch_38;
  assign edge_list_ch_39 = control_s_axi_U_edge_list_ch_39;
  assign edge_list_ch_4 = control_s_axi_U_edge_list_ch_4;
  assign edge_list_ch_40 = control_s_axi_U_edge_list_ch_40;
  assign edge_list_ch_41 = control_s_axi_U_edge_list_ch_41;
  assign edge_list_ch_42 = control_s_axi_U_edge_list_ch_42;
  assign edge_list_ch_43 = control_s_axi_U_edge_list_ch_43;
  assign edge_list_ch_44 = control_s_axi_U_edge_list_ch_44;
  assign edge_list_ch_45 = control_s_axi_U_edge_list_ch_45;
  assign edge_list_ch_46 = control_s_axi_U_edge_list_ch_46;
  assign edge_list_ch_47 = control_s_axi_U_edge_list_ch_47;
  assign edge_list_ch_5 = control_s_axi_U_edge_list_ch_5;
  assign edge_list_ch_6 = control_s_axi_U_edge_list_ch_6;
  assign edge_list_ch_7 = control_s_axi_U_edge_list_ch_7;
  assign edge_list_ch_8 = control_s_axi_U_edge_list_ch_8;
  assign edge_list_ch_9 = control_s_axi_U_edge_list_ch_9;
  assign edge_list_ptr = control_s_axi_U_edge_list_ptr;
  assign interrupt = control_s_axi_U_interrupt;
  assign vec_X = control_s_axi_U_vec_X;
  assign vec_Y = control_s_axi_U_vec_Y;
  assign vec_Y_out = control_s_axi_U_vec_Y_out;
  assign PE_inst_0_clk = ap_clk;
  assign PE_inst_0_if_din = PE_inst_0__din;
  assign PE_inst_0__dout = PE_inst_0_if_dout;
  assign PE_inst_0__empty_n = PE_inst_0_if_empty_n;
  assign PE_inst_0__full_n = PE_inst_0_if_full_n;
  assign PE_inst_0_if_read = PE_inst_0__read;
  assign PE_inst_0_if_read_ce = 1'b1;
  assign PE_inst_0_if_write = PE_inst_0__write;
  assign PE_inst_0_if_write_ce = 1'b1;
  assign PE_inst_0_reset = ~ ap_rst_n;
  assign PE_inst_10_clk = ap_clk;
  assign PE_inst_10_if_din = PE_inst_10__din;
  assign PE_inst_10__dout = PE_inst_10_if_dout;
  assign PE_inst_10__empty_n = PE_inst_10_if_empty_n;
  assign PE_inst_10__full_n = PE_inst_10_if_full_n;
  assign PE_inst_10_if_read = PE_inst_10__read;
  assign PE_inst_10_if_read_ce = 1'b1;
  assign PE_inst_10_if_write = PE_inst_10__write;
  assign PE_inst_10_if_write_ce = 1'b1;
  assign PE_inst_10_reset = ~ ap_rst_n;
  assign PE_inst_11_clk = ap_clk;
  assign PE_inst_11_if_din = PE_inst_11__din;
  assign PE_inst_11__dout = PE_inst_11_if_dout;
  assign PE_inst_11__empty_n = PE_inst_11_if_empty_n;
  assign PE_inst_11__full_n = PE_inst_11_if_full_n;
  assign PE_inst_11_if_read = PE_inst_11__read;
  assign PE_inst_11_if_read_ce = 1'b1;
  assign PE_inst_11_if_write = PE_inst_11__write;
  assign PE_inst_11_if_write_ce = 1'b1;
  assign PE_inst_11_reset = ~ ap_rst_n;
  assign PE_inst_12_clk = ap_clk;
  assign PE_inst_12_if_din = PE_inst_12__din;
  assign PE_inst_12__dout = PE_inst_12_if_dout;
  assign PE_inst_12__empty_n = PE_inst_12_if_empty_n;
  assign PE_inst_12__full_n = PE_inst_12_if_full_n;
  assign PE_inst_12_if_read = PE_inst_12__read;
  assign PE_inst_12_if_read_ce = 1'b1;
  assign PE_inst_12_if_write = PE_inst_12__write;
  assign PE_inst_12_if_write_ce = 1'b1;
  assign PE_inst_12_reset = ~ ap_rst_n;
  assign PE_inst_13_clk = ap_clk;
  assign PE_inst_13_if_din = PE_inst_13__din;
  assign PE_inst_13__dout = PE_inst_13_if_dout;
  assign PE_inst_13__empty_n = PE_inst_13_if_empty_n;
  assign PE_inst_13__full_n = PE_inst_13_if_full_n;
  assign PE_inst_13_if_read = PE_inst_13__read;
  assign PE_inst_13_if_read_ce = 1'b1;
  assign PE_inst_13_if_write = PE_inst_13__write;
  assign PE_inst_13_if_write_ce = 1'b1;
  assign PE_inst_13_reset = ~ ap_rst_n;
  assign PE_inst_14_clk = ap_clk;
  assign PE_inst_14_if_din = PE_inst_14__din;
  assign PE_inst_14__dout = PE_inst_14_if_dout;
  assign PE_inst_14__empty_n = PE_inst_14_if_empty_n;
  assign PE_inst_14__full_n = PE_inst_14_if_full_n;
  assign PE_inst_14_if_read = PE_inst_14__read;
  assign PE_inst_14_if_read_ce = 1'b1;
  assign PE_inst_14_if_write = PE_inst_14__write;
  assign PE_inst_14_if_write_ce = 1'b1;
  assign PE_inst_14_reset = ~ ap_rst_n;
  assign PE_inst_15_clk = ap_clk;
  assign PE_inst_15_if_din = PE_inst_15__din;
  assign PE_inst_15__dout = PE_inst_15_if_dout;
  assign PE_inst_15__empty_n = PE_inst_15_if_empty_n;
  assign PE_inst_15__full_n = PE_inst_15_if_full_n;
  assign PE_inst_15_if_read = PE_inst_15__read;
  assign PE_inst_15_if_read_ce = 1'b1;
  assign PE_inst_15_if_write = PE_inst_15__write;
  assign PE_inst_15_if_write_ce = 1'b1;
  assign PE_inst_15_reset = ~ ap_rst_n;
  assign PE_inst_16_clk = ap_clk;
  assign PE_inst_16_if_din = PE_inst_16__din;
  assign PE_inst_16__dout = PE_inst_16_if_dout;
  assign PE_inst_16__empty_n = PE_inst_16_if_empty_n;
  assign PE_inst_16__full_n = PE_inst_16_if_full_n;
  assign PE_inst_16_if_read = PE_inst_16__read;
  assign PE_inst_16_if_read_ce = 1'b1;
  assign PE_inst_16_if_write = PE_inst_16__write;
  assign PE_inst_16_if_write_ce = 1'b1;
  assign PE_inst_16_reset = ~ ap_rst_n;
  assign PE_inst_17_clk = ap_clk;
  assign PE_inst_17_if_din = PE_inst_17__din;
  assign PE_inst_17__dout = PE_inst_17_if_dout;
  assign PE_inst_17__empty_n = PE_inst_17_if_empty_n;
  assign PE_inst_17__full_n = PE_inst_17_if_full_n;
  assign PE_inst_17_if_read = PE_inst_17__read;
  assign PE_inst_17_if_read_ce = 1'b1;
  assign PE_inst_17_if_write = PE_inst_17__write;
  assign PE_inst_17_if_write_ce = 1'b1;
  assign PE_inst_17_reset = ~ ap_rst_n;
  assign PE_inst_18_clk = ap_clk;
  assign PE_inst_18_if_din = PE_inst_18__din;
  assign PE_inst_18__dout = PE_inst_18_if_dout;
  assign PE_inst_18__empty_n = PE_inst_18_if_empty_n;
  assign PE_inst_18__full_n = PE_inst_18_if_full_n;
  assign PE_inst_18_if_read = PE_inst_18__read;
  assign PE_inst_18_if_read_ce = 1'b1;
  assign PE_inst_18_if_write = PE_inst_18__write;
  assign PE_inst_18_if_write_ce = 1'b1;
  assign PE_inst_18_reset = ~ ap_rst_n;
  assign PE_inst_19_clk = ap_clk;
  assign PE_inst_19_if_din = PE_inst_19__din;
  assign PE_inst_19__dout = PE_inst_19_if_dout;
  assign PE_inst_19__empty_n = PE_inst_19_if_empty_n;
  assign PE_inst_19__full_n = PE_inst_19_if_full_n;
  assign PE_inst_19_if_read = PE_inst_19__read;
  assign PE_inst_19_if_read_ce = 1'b1;
  assign PE_inst_19_if_write = PE_inst_19__write;
  assign PE_inst_19_if_write_ce = 1'b1;
  assign PE_inst_19_reset = ~ ap_rst_n;
  assign PE_inst_1_clk = ap_clk;
  assign PE_inst_1_if_din = PE_inst_1__din;
  assign PE_inst_1__dout = PE_inst_1_if_dout;
  assign PE_inst_1__empty_n = PE_inst_1_if_empty_n;
  assign PE_inst_1__full_n = PE_inst_1_if_full_n;
  assign PE_inst_1_if_read = PE_inst_1__read;
  assign PE_inst_1_if_read_ce = 1'b1;
  assign PE_inst_1_if_write = PE_inst_1__write;
  assign PE_inst_1_if_write_ce = 1'b1;
  assign PE_inst_1_reset = ~ ap_rst_n;
  assign PE_inst_20_clk = ap_clk;
  assign PE_inst_20_if_din = PE_inst_20__din;
  assign PE_inst_20__dout = PE_inst_20_if_dout;
  assign PE_inst_20__empty_n = PE_inst_20_if_empty_n;
  assign PE_inst_20__full_n = PE_inst_20_if_full_n;
  assign PE_inst_20_if_read = PE_inst_20__read;
  assign PE_inst_20_if_read_ce = 1'b1;
  assign PE_inst_20_if_write = PE_inst_20__write;
  assign PE_inst_20_if_write_ce = 1'b1;
  assign PE_inst_20_reset = ~ ap_rst_n;
  assign PE_inst_21_clk = ap_clk;
  assign PE_inst_21_if_din = PE_inst_21__din;
  assign PE_inst_21__dout = PE_inst_21_if_dout;
  assign PE_inst_21__empty_n = PE_inst_21_if_empty_n;
  assign PE_inst_21__full_n = PE_inst_21_if_full_n;
  assign PE_inst_21_if_read = PE_inst_21__read;
  assign PE_inst_21_if_read_ce = 1'b1;
  assign PE_inst_21_if_write = PE_inst_21__write;
  assign PE_inst_21_if_write_ce = 1'b1;
  assign PE_inst_21_reset = ~ ap_rst_n;
  assign PE_inst_22_clk = ap_clk;
  assign PE_inst_22_if_din = PE_inst_22__din;
  assign PE_inst_22__dout = PE_inst_22_if_dout;
  assign PE_inst_22__empty_n = PE_inst_22_if_empty_n;
  assign PE_inst_22__full_n = PE_inst_22_if_full_n;
  assign PE_inst_22_if_read = PE_inst_22__read;
  assign PE_inst_22_if_read_ce = 1'b1;
  assign PE_inst_22_if_write = PE_inst_22__write;
  assign PE_inst_22_if_write_ce = 1'b1;
  assign PE_inst_22_reset = ~ ap_rst_n;
  assign PE_inst_23_clk = ap_clk;
  assign PE_inst_23_if_din = PE_inst_23__din;
  assign PE_inst_23__dout = PE_inst_23_if_dout;
  assign PE_inst_23__empty_n = PE_inst_23_if_empty_n;
  assign PE_inst_23__full_n = PE_inst_23_if_full_n;
  assign PE_inst_23_if_read = PE_inst_23__read;
  assign PE_inst_23_if_read_ce = 1'b1;
  assign PE_inst_23_if_write = PE_inst_23__write;
  assign PE_inst_23_if_write_ce = 1'b1;
  assign PE_inst_23_reset = ~ ap_rst_n;
  assign PE_inst_24_clk = ap_clk;
  assign PE_inst_24_if_din = PE_inst_24__din;
  assign PE_inst_24__dout = PE_inst_24_if_dout;
  assign PE_inst_24__empty_n = PE_inst_24_if_empty_n;
  assign PE_inst_24__full_n = PE_inst_24_if_full_n;
  assign PE_inst_24_if_read = PE_inst_24__read;
  assign PE_inst_24_if_read_ce = 1'b1;
  assign PE_inst_24_if_write = PE_inst_24__write;
  assign PE_inst_24_if_write_ce = 1'b1;
  assign PE_inst_24_reset = ~ ap_rst_n;
  assign PE_inst_25_clk = ap_clk;
  assign PE_inst_25_if_din = PE_inst_25__din;
  assign PE_inst_25__dout = PE_inst_25_if_dout;
  assign PE_inst_25__empty_n = PE_inst_25_if_empty_n;
  assign PE_inst_25__full_n = PE_inst_25_if_full_n;
  assign PE_inst_25_if_read = PE_inst_25__read;
  assign PE_inst_25_if_read_ce = 1'b1;
  assign PE_inst_25_if_write = PE_inst_25__write;
  assign PE_inst_25_if_write_ce = 1'b1;
  assign PE_inst_25_reset = ~ ap_rst_n;
  assign PE_inst_26_clk = ap_clk;
  assign PE_inst_26_if_din = PE_inst_26__din;
  assign PE_inst_26__dout = PE_inst_26_if_dout;
  assign PE_inst_26__empty_n = PE_inst_26_if_empty_n;
  assign PE_inst_26__full_n = PE_inst_26_if_full_n;
  assign PE_inst_26_if_read = PE_inst_26__read;
  assign PE_inst_26_if_read_ce = 1'b1;
  assign PE_inst_26_if_write = PE_inst_26__write;
  assign PE_inst_26_if_write_ce = 1'b1;
  assign PE_inst_26_reset = ~ ap_rst_n;
  assign PE_inst_27_clk = ap_clk;
  assign PE_inst_27_if_din = PE_inst_27__din;
  assign PE_inst_27__dout = PE_inst_27_if_dout;
  assign PE_inst_27__empty_n = PE_inst_27_if_empty_n;
  assign PE_inst_27__full_n = PE_inst_27_if_full_n;
  assign PE_inst_27_if_read = PE_inst_27__read;
  assign PE_inst_27_if_read_ce = 1'b1;
  assign PE_inst_27_if_write = PE_inst_27__write;
  assign PE_inst_27_if_write_ce = 1'b1;
  assign PE_inst_27_reset = ~ ap_rst_n;
  assign PE_inst_28_clk = ap_clk;
  assign PE_inst_28_if_din = PE_inst_28__din;
  assign PE_inst_28__dout = PE_inst_28_if_dout;
  assign PE_inst_28__empty_n = PE_inst_28_if_empty_n;
  assign PE_inst_28__full_n = PE_inst_28_if_full_n;
  assign PE_inst_28_if_read = PE_inst_28__read;
  assign PE_inst_28_if_read_ce = 1'b1;
  assign PE_inst_28_if_write = PE_inst_28__write;
  assign PE_inst_28_if_write_ce = 1'b1;
  assign PE_inst_28_reset = ~ ap_rst_n;
  assign PE_inst_29_clk = ap_clk;
  assign PE_inst_29_if_din = PE_inst_29__din;
  assign PE_inst_29__dout = PE_inst_29_if_dout;
  assign PE_inst_29__empty_n = PE_inst_29_if_empty_n;
  assign PE_inst_29__full_n = PE_inst_29_if_full_n;
  assign PE_inst_29_if_read = PE_inst_29__read;
  assign PE_inst_29_if_read_ce = 1'b1;
  assign PE_inst_29_if_write = PE_inst_29__write;
  assign PE_inst_29_if_write_ce = 1'b1;
  assign PE_inst_29_reset = ~ ap_rst_n;
  assign PE_inst_2_clk = ap_clk;
  assign PE_inst_2_if_din = PE_inst_2__din;
  assign PE_inst_2__dout = PE_inst_2_if_dout;
  assign PE_inst_2__empty_n = PE_inst_2_if_empty_n;
  assign PE_inst_2__full_n = PE_inst_2_if_full_n;
  assign PE_inst_2_if_read = PE_inst_2__read;
  assign PE_inst_2_if_read_ce = 1'b1;
  assign PE_inst_2_if_write = PE_inst_2__write;
  assign PE_inst_2_if_write_ce = 1'b1;
  assign PE_inst_2_reset = ~ ap_rst_n;
  assign PE_inst_30_clk = ap_clk;
  assign PE_inst_30_if_din = PE_inst_30__din;
  assign PE_inst_30__dout = PE_inst_30_if_dout;
  assign PE_inst_30__empty_n = PE_inst_30_if_empty_n;
  assign PE_inst_30__full_n = PE_inst_30_if_full_n;
  assign PE_inst_30_if_read = PE_inst_30__read;
  assign PE_inst_30_if_read_ce = 1'b1;
  assign PE_inst_30_if_write = PE_inst_30__write;
  assign PE_inst_30_if_write_ce = 1'b1;
  assign PE_inst_30_reset = ~ ap_rst_n;
  assign PE_inst_31_clk = ap_clk;
  assign PE_inst_31_if_din = PE_inst_31__din;
  assign PE_inst_31__dout = PE_inst_31_if_dout;
  assign PE_inst_31__empty_n = PE_inst_31_if_empty_n;
  assign PE_inst_31__full_n = PE_inst_31_if_full_n;
  assign PE_inst_31_if_read = PE_inst_31__read;
  assign PE_inst_31_if_read_ce = 1'b1;
  assign PE_inst_31_if_write = PE_inst_31__write;
  assign PE_inst_31_if_write_ce = 1'b1;
  assign PE_inst_31_reset = ~ ap_rst_n;
  assign PE_inst_32_clk = ap_clk;
  assign PE_inst_32_if_din = PE_inst_32__din;
  assign PE_inst_32__dout = PE_inst_32_if_dout;
  assign PE_inst_32__empty_n = PE_inst_32_if_empty_n;
  assign PE_inst_32__full_n = PE_inst_32_if_full_n;
  assign PE_inst_32_if_read = PE_inst_32__read;
  assign PE_inst_32_if_read_ce = 1'b1;
  assign PE_inst_32_if_write = PE_inst_32__write;
  assign PE_inst_32_if_write_ce = 1'b1;
  assign PE_inst_32_reset = ~ ap_rst_n;
  assign PE_inst_33_clk = ap_clk;
  assign PE_inst_33_if_din = PE_inst_33__din;
  assign PE_inst_33__dout = PE_inst_33_if_dout;
  assign PE_inst_33__empty_n = PE_inst_33_if_empty_n;
  assign PE_inst_33__full_n = PE_inst_33_if_full_n;
  assign PE_inst_33_if_read = PE_inst_33__read;
  assign PE_inst_33_if_read_ce = 1'b1;
  assign PE_inst_33_if_write = PE_inst_33__write;
  assign PE_inst_33_if_write_ce = 1'b1;
  assign PE_inst_33_reset = ~ ap_rst_n;
  assign PE_inst_34_clk = ap_clk;
  assign PE_inst_34_if_din = PE_inst_34__din;
  assign PE_inst_34__dout = PE_inst_34_if_dout;
  assign PE_inst_34__empty_n = PE_inst_34_if_empty_n;
  assign PE_inst_34__full_n = PE_inst_34_if_full_n;
  assign PE_inst_34_if_read = PE_inst_34__read;
  assign PE_inst_34_if_read_ce = 1'b1;
  assign PE_inst_34_if_write = PE_inst_34__write;
  assign PE_inst_34_if_write_ce = 1'b1;
  assign PE_inst_34_reset = ~ ap_rst_n;
  assign PE_inst_35_clk = ap_clk;
  assign PE_inst_35_if_din = PE_inst_35__din;
  assign PE_inst_35__dout = PE_inst_35_if_dout;
  assign PE_inst_35__empty_n = PE_inst_35_if_empty_n;
  assign PE_inst_35__full_n = PE_inst_35_if_full_n;
  assign PE_inst_35_if_read = PE_inst_35__read;
  assign PE_inst_35_if_read_ce = 1'b1;
  assign PE_inst_35_if_write = PE_inst_35__write;
  assign PE_inst_35_if_write_ce = 1'b1;
  assign PE_inst_35_reset = ~ ap_rst_n;
  assign PE_inst_36_clk = ap_clk;
  assign PE_inst_36_if_din = PE_inst_36__din;
  assign PE_inst_36__dout = PE_inst_36_if_dout;
  assign PE_inst_36__empty_n = PE_inst_36_if_empty_n;
  assign PE_inst_36__full_n = PE_inst_36_if_full_n;
  assign PE_inst_36_if_read = PE_inst_36__read;
  assign PE_inst_36_if_read_ce = 1'b1;
  assign PE_inst_36_if_write = PE_inst_36__write;
  assign PE_inst_36_if_write_ce = 1'b1;
  assign PE_inst_36_reset = ~ ap_rst_n;
  assign PE_inst_37_clk = ap_clk;
  assign PE_inst_37_if_din = PE_inst_37__din;
  assign PE_inst_37__dout = PE_inst_37_if_dout;
  assign PE_inst_37__empty_n = PE_inst_37_if_empty_n;
  assign PE_inst_37__full_n = PE_inst_37_if_full_n;
  assign PE_inst_37_if_read = PE_inst_37__read;
  assign PE_inst_37_if_read_ce = 1'b1;
  assign PE_inst_37_if_write = PE_inst_37__write;
  assign PE_inst_37_if_write_ce = 1'b1;
  assign PE_inst_37_reset = ~ ap_rst_n;
  assign PE_inst_38_clk = ap_clk;
  assign PE_inst_38_if_din = PE_inst_38__din;
  assign PE_inst_38__dout = PE_inst_38_if_dout;
  assign PE_inst_38__empty_n = PE_inst_38_if_empty_n;
  assign PE_inst_38__full_n = PE_inst_38_if_full_n;
  assign PE_inst_38_if_read = PE_inst_38__read;
  assign PE_inst_38_if_read_ce = 1'b1;
  assign PE_inst_38_if_write = PE_inst_38__write;
  assign PE_inst_38_if_write_ce = 1'b1;
  assign PE_inst_38_reset = ~ ap_rst_n;
  assign PE_inst_39_clk = ap_clk;
  assign PE_inst_39_if_din = PE_inst_39__din;
  assign PE_inst_39__dout = PE_inst_39_if_dout;
  assign PE_inst_39__empty_n = PE_inst_39_if_empty_n;
  assign PE_inst_39__full_n = PE_inst_39_if_full_n;
  assign PE_inst_39_if_read = PE_inst_39__read;
  assign PE_inst_39_if_read_ce = 1'b1;
  assign PE_inst_39_if_write = PE_inst_39__write;
  assign PE_inst_39_if_write_ce = 1'b1;
  assign PE_inst_39_reset = ~ ap_rst_n;
  assign PE_inst_3_clk = ap_clk;
  assign PE_inst_3_if_din = PE_inst_3__din;
  assign PE_inst_3__dout = PE_inst_3_if_dout;
  assign PE_inst_3__empty_n = PE_inst_3_if_empty_n;
  assign PE_inst_3__full_n = PE_inst_3_if_full_n;
  assign PE_inst_3_if_read = PE_inst_3__read;
  assign PE_inst_3_if_read_ce = 1'b1;
  assign PE_inst_3_if_write = PE_inst_3__write;
  assign PE_inst_3_if_write_ce = 1'b1;
  assign PE_inst_3_reset = ~ ap_rst_n;
  assign PE_inst_40_clk = ap_clk;
  assign PE_inst_40_if_din = PE_inst_40__din;
  assign PE_inst_40__dout = PE_inst_40_if_dout;
  assign PE_inst_40__empty_n = PE_inst_40_if_empty_n;
  assign PE_inst_40__full_n = PE_inst_40_if_full_n;
  assign PE_inst_40_if_read = PE_inst_40__read;
  assign PE_inst_40_if_read_ce = 1'b1;
  assign PE_inst_40_if_write = PE_inst_40__write;
  assign PE_inst_40_if_write_ce = 1'b1;
  assign PE_inst_40_reset = ~ ap_rst_n;
  assign PE_inst_41_clk = ap_clk;
  assign PE_inst_41_if_din = PE_inst_41__din;
  assign PE_inst_41__dout = PE_inst_41_if_dout;
  assign PE_inst_41__empty_n = PE_inst_41_if_empty_n;
  assign PE_inst_41__full_n = PE_inst_41_if_full_n;
  assign PE_inst_41_if_read = PE_inst_41__read;
  assign PE_inst_41_if_read_ce = 1'b1;
  assign PE_inst_41_if_write = PE_inst_41__write;
  assign PE_inst_41_if_write_ce = 1'b1;
  assign PE_inst_41_reset = ~ ap_rst_n;
  assign PE_inst_42_clk = ap_clk;
  assign PE_inst_42_if_din = PE_inst_42__din;
  assign PE_inst_42__dout = PE_inst_42_if_dout;
  assign PE_inst_42__empty_n = PE_inst_42_if_empty_n;
  assign PE_inst_42__full_n = PE_inst_42_if_full_n;
  assign PE_inst_42_if_read = PE_inst_42__read;
  assign PE_inst_42_if_read_ce = 1'b1;
  assign PE_inst_42_if_write = PE_inst_42__write;
  assign PE_inst_42_if_write_ce = 1'b1;
  assign PE_inst_42_reset = ~ ap_rst_n;
  assign PE_inst_43_clk = ap_clk;
  assign PE_inst_43_if_din = PE_inst_43__din;
  assign PE_inst_43__dout = PE_inst_43_if_dout;
  assign PE_inst_43__empty_n = PE_inst_43_if_empty_n;
  assign PE_inst_43__full_n = PE_inst_43_if_full_n;
  assign PE_inst_43_if_read = PE_inst_43__read;
  assign PE_inst_43_if_read_ce = 1'b1;
  assign PE_inst_43_if_write = PE_inst_43__write;
  assign PE_inst_43_if_write_ce = 1'b1;
  assign PE_inst_43_reset = ~ ap_rst_n;
  assign PE_inst_44_clk = ap_clk;
  assign PE_inst_44_if_din = PE_inst_44__din;
  assign PE_inst_44__dout = PE_inst_44_if_dout;
  assign PE_inst_44__empty_n = PE_inst_44_if_empty_n;
  assign PE_inst_44__full_n = PE_inst_44_if_full_n;
  assign PE_inst_44_if_read = PE_inst_44__read;
  assign PE_inst_44_if_read_ce = 1'b1;
  assign PE_inst_44_if_write = PE_inst_44__write;
  assign PE_inst_44_if_write_ce = 1'b1;
  assign PE_inst_44_reset = ~ ap_rst_n;
  assign PE_inst_45_clk = ap_clk;
  assign PE_inst_45_if_din = PE_inst_45__din;
  assign PE_inst_45__dout = PE_inst_45_if_dout;
  assign PE_inst_45__empty_n = PE_inst_45_if_empty_n;
  assign PE_inst_45__full_n = PE_inst_45_if_full_n;
  assign PE_inst_45_if_read = PE_inst_45__read;
  assign PE_inst_45_if_read_ce = 1'b1;
  assign PE_inst_45_if_write = PE_inst_45__write;
  assign PE_inst_45_if_write_ce = 1'b1;
  assign PE_inst_45_reset = ~ ap_rst_n;
  assign PE_inst_46_clk = ap_clk;
  assign PE_inst_46_if_din = PE_inst_46__din;
  assign PE_inst_46__dout = PE_inst_46_if_dout;
  assign PE_inst_46__empty_n = PE_inst_46_if_empty_n;
  assign PE_inst_46__full_n = PE_inst_46_if_full_n;
  assign PE_inst_46_if_read = PE_inst_46__read;
  assign PE_inst_46_if_read_ce = 1'b1;
  assign PE_inst_46_if_write = PE_inst_46__write;
  assign PE_inst_46_if_write_ce = 1'b1;
  assign PE_inst_46_reset = ~ ap_rst_n;
  assign PE_inst_47_clk = ap_clk;
  assign PE_inst_47_if_din = PE_inst_47__din;
  assign PE_inst_47__dout = PE_inst_47_if_dout;
  assign PE_inst_47__empty_n = PE_inst_47_if_empty_n;
  assign PE_inst_47__full_n = PE_inst_47_if_full_n;
  assign PE_inst_47_if_read = PE_inst_47__read;
  assign PE_inst_47_if_read_ce = 1'b1;
  assign PE_inst_47_if_write = PE_inst_47__write;
  assign PE_inst_47_if_write_ce = 1'b1;
  assign PE_inst_47_reset = ~ ap_rst_n;
  assign PE_inst_48_clk = ap_clk;
  assign PE_inst_48_if_din = PE_inst_48__din;
  assign PE_inst_48__dout = PE_inst_48_if_dout;
  assign PE_inst_48__empty_n = PE_inst_48_if_empty_n;
  assign PE_inst_48__full_n = PE_inst_48_if_full_n;
  assign PE_inst_48_if_read = PE_inst_48__read;
  assign PE_inst_48_if_read_ce = 1'b1;
  assign PE_inst_48_if_write = PE_inst_48__write;
  assign PE_inst_48_if_write_ce = 1'b1;
  assign PE_inst_48_reset = ~ ap_rst_n;
  assign PE_inst_4_clk = ap_clk;
  assign PE_inst_4_if_din = PE_inst_4__din;
  assign PE_inst_4__dout = PE_inst_4_if_dout;
  assign PE_inst_4__empty_n = PE_inst_4_if_empty_n;
  assign PE_inst_4__full_n = PE_inst_4_if_full_n;
  assign PE_inst_4_if_read = PE_inst_4__read;
  assign PE_inst_4_if_read_ce = 1'b1;
  assign PE_inst_4_if_write = PE_inst_4__write;
  assign PE_inst_4_if_write_ce = 1'b1;
  assign PE_inst_4_reset = ~ ap_rst_n;
  assign PE_inst_5_clk = ap_clk;
  assign PE_inst_5_if_din = PE_inst_5__din;
  assign PE_inst_5__dout = PE_inst_5_if_dout;
  assign PE_inst_5__empty_n = PE_inst_5_if_empty_n;
  assign PE_inst_5__full_n = PE_inst_5_if_full_n;
  assign PE_inst_5_if_read = PE_inst_5__read;
  assign PE_inst_5_if_read_ce = 1'b1;
  assign PE_inst_5_if_write = PE_inst_5__write;
  assign PE_inst_5_if_write_ce = 1'b1;
  assign PE_inst_5_reset = ~ ap_rst_n;
  assign PE_inst_6_clk = ap_clk;
  assign PE_inst_6_if_din = PE_inst_6__din;
  assign PE_inst_6__dout = PE_inst_6_if_dout;
  assign PE_inst_6__empty_n = PE_inst_6_if_empty_n;
  assign PE_inst_6__full_n = PE_inst_6_if_full_n;
  assign PE_inst_6_if_read = PE_inst_6__read;
  assign PE_inst_6_if_read_ce = 1'b1;
  assign PE_inst_6_if_write = PE_inst_6__write;
  assign PE_inst_6_if_write_ce = 1'b1;
  assign PE_inst_6_reset = ~ ap_rst_n;
  assign PE_inst_7_clk = ap_clk;
  assign PE_inst_7_if_din = PE_inst_7__din;
  assign PE_inst_7__dout = PE_inst_7_if_dout;
  assign PE_inst_7__empty_n = PE_inst_7_if_empty_n;
  assign PE_inst_7__full_n = PE_inst_7_if_full_n;
  assign PE_inst_7_if_read = PE_inst_7__read;
  assign PE_inst_7_if_read_ce = 1'b1;
  assign PE_inst_7_if_write = PE_inst_7__write;
  assign PE_inst_7_if_write_ce = 1'b1;
  assign PE_inst_7_reset = ~ ap_rst_n;
  assign PE_inst_8_clk = ap_clk;
  assign PE_inst_8_if_din = PE_inst_8__din;
  assign PE_inst_8__dout = PE_inst_8_if_dout;
  assign PE_inst_8__empty_n = PE_inst_8_if_empty_n;
  assign PE_inst_8__full_n = PE_inst_8_if_full_n;
  assign PE_inst_8_if_read = PE_inst_8__read;
  assign PE_inst_8_if_read_ce = 1'b1;
  assign PE_inst_8_if_write = PE_inst_8__write;
  assign PE_inst_8_if_write_ce = 1'b1;
  assign PE_inst_8_reset = ~ ap_rst_n;
  assign PE_inst_9_clk = ap_clk;
  assign PE_inst_9_if_din = PE_inst_9__din;
  assign PE_inst_9__dout = PE_inst_9_if_dout;
  assign PE_inst_9__empty_n = PE_inst_9_if_empty_n;
  assign PE_inst_9__full_n = PE_inst_9_if_full_n;
  assign PE_inst_9_if_read = PE_inst_9__read;
  assign PE_inst_9_if_read_ce = 1'b1;
  assign PE_inst_9_if_write = PE_inst_9__write;
  assign PE_inst_9_if_write_ce = 1'b1;
  assign PE_inst_9_reset = ~ ap_rst_n;
  assign Yvec_inst_0_clk = ap_clk;
  assign Yvec_inst_0_if_din = Yvec_inst_0__din;
  assign Yvec_inst_0__dout = Yvec_inst_0_if_dout;
  assign Yvec_inst_0__empty_n = Yvec_inst_0_if_empty_n;
  assign Yvec_inst_0__full_n = Yvec_inst_0_if_full_n;
  assign Yvec_inst_0_if_read = Yvec_inst_0__read;
  assign Yvec_inst_0_if_read_ce = 1'b1;
  assign Yvec_inst_0_if_write = Yvec_inst_0__write;
  assign Yvec_inst_0_if_write_ce = 1'b1;
  assign Yvec_inst_0_reset = ~ ap_rst_n;
  assign Yvec_inst_10_clk = ap_clk;
  assign Yvec_inst_10_if_din = Yvec_inst_10__din;
  assign Yvec_inst_10__dout = Yvec_inst_10_if_dout;
  assign Yvec_inst_10__empty_n = Yvec_inst_10_if_empty_n;
  assign Yvec_inst_10__full_n = Yvec_inst_10_if_full_n;
  assign Yvec_inst_10_if_read = Yvec_inst_10__read;
  assign Yvec_inst_10_if_read_ce = 1'b1;
  assign Yvec_inst_10_if_write = Yvec_inst_10__write;
  assign Yvec_inst_10_if_write_ce = 1'b1;
  assign Yvec_inst_10_reset = ~ ap_rst_n;
  assign Yvec_inst_11_clk = ap_clk;
  assign Yvec_inst_11_if_din = Yvec_inst_11__din;
  assign Yvec_inst_11__dout = Yvec_inst_11_if_dout;
  assign Yvec_inst_11__empty_n = Yvec_inst_11_if_empty_n;
  assign Yvec_inst_11__full_n = Yvec_inst_11_if_full_n;
  assign Yvec_inst_11_if_read = Yvec_inst_11__read;
  assign Yvec_inst_11_if_read_ce = 1'b1;
  assign Yvec_inst_11_if_write = Yvec_inst_11__write;
  assign Yvec_inst_11_if_write_ce = 1'b1;
  assign Yvec_inst_11_reset = ~ ap_rst_n;
  assign Yvec_inst_12_clk = ap_clk;
  assign Yvec_inst_12_if_din = Yvec_inst_12__din;
  assign Yvec_inst_12__dout = Yvec_inst_12_if_dout;
  assign Yvec_inst_12__empty_n = Yvec_inst_12_if_empty_n;
  assign Yvec_inst_12__full_n = Yvec_inst_12_if_full_n;
  assign Yvec_inst_12_if_read = Yvec_inst_12__read;
  assign Yvec_inst_12_if_read_ce = 1'b1;
  assign Yvec_inst_12_if_write = Yvec_inst_12__write;
  assign Yvec_inst_12_if_write_ce = 1'b1;
  assign Yvec_inst_12_reset = ~ ap_rst_n;
  assign Yvec_inst_13_clk = ap_clk;
  assign Yvec_inst_13_if_din = Yvec_inst_13__din;
  assign Yvec_inst_13__dout = Yvec_inst_13_if_dout;
  assign Yvec_inst_13__empty_n = Yvec_inst_13_if_empty_n;
  assign Yvec_inst_13__full_n = Yvec_inst_13_if_full_n;
  assign Yvec_inst_13_if_read = Yvec_inst_13__read;
  assign Yvec_inst_13_if_read_ce = 1'b1;
  assign Yvec_inst_13_if_write = Yvec_inst_13__write;
  assign Yvec_inst_13_if_write_ce = 1'b1;
  assign Yvec_inst_13_reset = ~ ap_rst_n;
  assign Yvec_inst_14_clk = ap_clk;
  assign Yvec_inst_14_if_din = Yvec_inst_14__din;
  assign Yvec_inst_14__dout = Yvec_inst_14_if_dout;
  assign Yvec_inst_14__empty_n = Yvec_inst_14_if_empty_n;
  assign Yvec_inst_14__full_n = Yvec_inst_14_if_full_n;
  assign Yvec_inst_14_if_read = Yvec_inst_14__read;
  assign Yvec_inst_14_if_read_ce = 1'b1;
  assign Yvec_inst_14_if_write = Yvec_inst_14__write;
  assign Yvec_inst_14_if_write_ce = 1'b1;
  assign Yvec_inst_14_reset = ~ ap_rst_n;
  assign Yvec_inst_15_clk = ap_clk;
  assign Yvec_inst_15_if_din = Yvec_inst_15__din;
  assign Yvec_inst_15__dout = Yvec_inst_15_if_dout;
  assign Yvec_inst_15__empty_n = Yvec_inst_15_if_empty_n;
  assign Yvec_inst_15__full_n = Yvec_inst_15_if_full_n;
  assign Yvec_inst_15_if_read = Yvec_inst_15__read;
  assign Yvec_inst_15_if_read_ce = 1'b1;
  assign Yvec_inst_15_if_write = Yvec_inst_15__write;
  assign Yvec_inst_15_if_write_ce = 1'b1;
  assign Yvec_inst_15_reset = ~ ap_rst_n;
  assign Yvec_inst_16_clk = ap_clk;
  assign Yvec_inst_16_if_din = Yvec_inst_16__din;
  assign Yvec_inst_16__dout = Yvec_inst_16_if_dout;
  assign Yvec_inst_16__empty_n = Yvec_inst_16_if_empty_n;
  assign Yvec_inst_16__full_n = Yvec_inst_16_if_full_n;
  assign Yvec_inst_16_if_read = Yvec_inst_16__read;
  assign Yvec_inst_16_if_read_ce = 1'b1;
  assign Yvec_inst_16_if_write = Yvec_inst_16__write;
  assign Yvec_inst_16_if_write_ce = 1'b1;
  assign Yvec_inst_16_reset = ~ ap_rst_n;
  assign Yvec_inst_17_clk = ap_clk;
  assign Yvec_inst_17_if_din = Yvec_inst_17__din;
  assign Yvec_inst_17__dout = Yvec_inst_17_if_dout;
  assign Yvec_inst_17__empty_n = Yvec_inst_17_if_empty_n;
  assign Yvec_inst_17__full_n = Yvec_inst_17_if_full_n;
  assign Yvec_inst_17_if_read = Yvec_inst_17__read;
  assign Yvec_inst_17_if_read_ce = 1'b1;
  assign Yvec_inst_17_if_write = Yvec_inst_17__write;
  assign Yvec_inst_17_if_write_ce = 1'b1;
  assign Yvec_inst_17_reset = ~ ap_rst_n;
  assign Yvec_inst_18_clk = ap_clk;
  assign Yvec_inst_18_if_din = Yvec_inst_18__din;
  assign Yvec_inst_18__dout = Yvec_inst_18_if_dout;
  assign Yvec_inst_18__empty_n = Yvec_inst_18_if_empty_n;
  assign Yvec_inst_18__full_n = Yvec_inst_18_if_full_n;
  assign Yvec_inst_18_if_read = Yvec_inst_18__read;
  assign Yvec_inst_18_if_read_ce = 1'b1;
  assign Yvec_inst_18_if_write = Yvec_inst_18__write;
  assign Yvec_inst_18_if_write_ce = 1'b1;
  assign Yvec_inst_18_reset = ~ ap_rst_n;
  assign Yvec_inst_19_clk = ap_clk;
  assign Yvec_inst_19_if_din = Yvec_inst_19__din;
  assign Yvec_inst_19__dout = Yvec_inst_19_if_dout;
  assign Yvec_inst_19__empty_n = Yvec_inst_19_if_empty_n;
  assign Yvec_inst_19__full_n = Yvec_inst_19_if_full_n;
  assign Yvec_inst_19_if_read = Yvec_inst_19__read;
  assign Yvec_inst_19_if_read_ce = 1'b1;
  assign Yvec_inst_19_if_write = Yvec_inst_19__write;
  assign Yvec_inst_19_if_write_ce = 1'b1;
  assign Yvec_inst_19_reset = ~ ap_rst_n;
  assign Yvec_inst_1_clk = ap_clk;
  assign Yvec_inst_1_if_din = Yvec_inst_1__din;
  assign Yvec_inst_1__dout = Yvec_inst_1_if_dout;
  assign Yvec_inst_1__empty_n = Yvec_inst_1_if_empty_n;
  assign Yvec_inst_1__full_n = Yvec_inst_1_if_full_n;
  assign Yvec_inst_1_if_read = Yvec_inst_1__read;
  assign Yvec_inst_1_if_read_ce = 1'b1;
  assign Yvec_inst_1_if_write = Yvec_inst_1__write;
  assign Yvec_inst_1_if_write_ce = 1'b1;
  assign Yvec_inst_1_reset = ~ ap_rst_n;
  assign Yvec_inst_20_clk = ap_clk;
  assign Yvec_inst_20_if_din = Yvec_inst_20__din;
  assign Yvec_inst_20__dout = Yvec_inst_20_if_dout;
  assign Yvec_inst_20__empty_n = Yvec_inst_20_if_empty_n;
  assign Yvec_inst_20__full_n = Yvec_inst_20_if_full_n;
  assign Yvec_inst_20_if_read = Yvec_inst_20__read;
  assign Yvec_inst_20_if_read_ce = 1'b1;
  assign Yvec_inst_20_if_write = Yvec_inst_20__write;
  assign Yvec_inst_20_if_write_ce = 1'b1;
  assign Yvec_inst_20_reset = ~ ap_rst_n;
  assign Yvec_inst_21_clk = ap_clk;
  assign Yvec_inst_21_if_din = Yvec_inst_21__din;
  assign Yvec_inst_21__dout = Yvec_inst_21_if_dout;
  assign Yvec_inst_21__empty_n = Yvec_inst_21_if_empty_n;
  assign Yvec_inst_21__full_n = Yvec_inst_21_if_full_n;
  assign Yvec_inst_21_if_read = Yvec_inst_21__read;
  assign Yvec_inst_21_if_read_ce = 1'b1;
  assign Yvec_inst_21_if_write = Yvec_inst_21__write;
  assign Yvec_inst_21_if_write_ce = 1'b1;
  assign Yvec_inst_21_reset = ~ ap_rst_n;
  assign Yvec_inst_22_clk = ap_clk;
  assign Yvec_inst_22_if_din = Yvec_inst_22__din;
  assign Yvec_inst_22__dout = Yvec_inst_22_if_dout;
  assign Yvec_inst_22__empty_n = Yvec_inst_22_if_empty_n;
  assign Yvec_inst_22__full_n = Yvec_inst_22_if_full_n;
  assign Yvec_inst_22_if_read = Yvec_inst_22__read;
  assign Yvec_inst_22_if_read_ce = 1'b1;
  assign Yvec_inst_22_if_write = Yvec_inst_22__write;
  assign Yvec_inst_22_if_write_ce = 1'b1;
  assign Yvec_inst_22_reset = ~ ap_rst_n;
  assign Yvec_inst_23_clk = ap_clk;
  assign Yvec_inst_23_if_din = Yvec_inst_23__din;
  assign Yvec_inst_23__dout = Yvec_inst_23_if_dout;
  assign Yvec_inst_23__empty_n = Yvec_inst_23_if_empty_n;
  assign Yvec_inst_23__full_n = Yvec_inst_23_if_full_n;
  assign Yvec_inst_23_if_read = Yvec_inst_23__read;
  assign Yvec_inst_23_if_read_ce = 1'b1;
  assign Yvec_inst_23_if_write = Yvec_inst_23__write;
  assign Yvec_inst_23_if_write_ce = 1'b1;
  assign Yvec_inst_23_reset = ~ ap_rst_n;
  assign Yvec_inst_24_clk = ap_clk;
  assign Yvec_inst_24_if_din = Yvec_inst_24__din;
  assign Yvec_inst_24__dout = Yvec_inst_24_if_dout;
  assign Yvec_inst_24__empty_n = Yvec_inst_24_if_empty_n;
  assign Yvec_inst_24__full_n = Yvec_inst_24_if_full_n;
  assign Yvec_inst_24_if_read = Yvec_inst_24__read;
  assign Yvec_inst_24_if_read_ce = 1'b1;
  assign Yvec_inst_24_if_write = Yvec_inst_24__write;
  assign Yvec_inst_24_if_write_ce = 1'b1;
  assign Yvec_inst_24_reset = ~ ap_rst_n;
  assign Yvec_inst_25_clk = ap_clk;
  assign Yvec_inst_25_if_din = Yvec_inst_25__din;
  assign Yvec_inst_25__dout = Yvec_inst_25_if_dout;
  assign Yvec_inst_25__empty_n = Yvec_inst_25_if_empty_n;
  assign Yvec_inst_25__full_n = Yvec_inst_25_if_full_n;
  assign Yvec_inst_25_if_read = Yvec_inst_25__read;
  assign Yvec_inst_25_if_read_ce = 1'b1;
  assign Yvec_inst_25_if_write = Yvec_inst_25__write;
  assign Yvec_inst_25_if_write_ce = 1'b1;
  assign Yvec_inst_25_reset = ~ ap_rst_n;
  assign Yvec_inst_26_clk = ap_clk;
  assign Yvec_inst_26_if_din = Yvec_inst_26__din;
  assign Yvec_inst_26__dout = Yvec_inst_26_if_dout;
  assign Yvec_inst_26__empty_n = Yvec_inst_26_if_empty_n;
  assign Yvec_inst_26__full_n = Yvec_inst_26_if_full_n;
  assign Yvec_inst_26_if_read = Yvec_inst_26__read;
  assign Yvec_inst_26_if_read_ce = 1'b1;
  assign Yvec_inst_26_if_write = Yvec_inst_26__write;
  assign Yvec_inst_26_if_write_ce = 1'b1;
  assign Yvec_inst_26_reset = ~ ap_rst_n;
  assign Yvec_inst_27_clk = ap_clk;
  assign Yvec_inst_27_if_din = Yvec_inst_27__din;
  assign Yvec_inst_27__dout = Yvec_inst_27_if_dout;
  assign Yvec_inst_27__empty_n = Yvec_inst_27_if_empty_n;
  assign Yvec_inst_27__full_n = Yvec_inst_27_if_full_n;
  assign Yvec_inst_27_if_read = Yvec_inst_27__read;
  assign Yvec_inst_27_if_read_ce = 1'b1;
  assign Yvec_inst_27_if_write = Yvec_inst_27__write;
  assign Yvec_inst_27_if_write_ce = 1'b1;
  assign Yvec_inst_27_reset = ~ ap_rst_n;
  assign Yvec_inst_28_clk = ap_clk;
  assign Yvec_inst_28_if_din = Yvec_inst_28__din;
  assign Yvec_inst_28__dout = Yvec_inst_28_if_dout;
  assign Yvec_inst_28__empty_n = Yvec_inst_28_if_empty_n;
  assign Yvec_inst_28__full_n = Yvec_inst_28_if_full_n;
  assign Yvec_inst_28_if_read = Yvec_inst_28__read;
  assign Yvec_inst_28_if_read_ce = 1'b1;
  assign Yvec_inst_28_if_write = Yvec_inst_28__write;
  assign Yvec_inst_28_if_write_ce = 1'b1;
  assign Yvec_inst_28_reset = ~ ap_rst_n;
  assign Yvec_inst_29_clk = ap_clk;
  assign Yvec_inst_29_if_din = Yvec_inst_29__din;
  assign Yvec_inst_29__dout = Yvec_inst_29_if_dout;
  assign Yvec_inst_29__empty_n = Yvec_inst_29_if_empty_n;
  assign Yvec_inst_29__full_n = Yvec_inst_29_if_full_n;
  assign Yvec_inst_29_if_read = Yvec_inst_29__read;
  assign Yvec_inst_29_if_read_ce = 1'b1;
  assign Yvec_inst_29_if_write = Yvec_inst_29__write;
  assign Yvec_inst_29_if_write_ce = 1'b1;
  assign Yvec_inst_29_reset = ~ ap_rst_n;
  assign Yvec_inst_2_clk = ap_clk;
  assign Yvec_inst_2_if_din = Yvec_inst_2__din;
  assign Yvec_inst_2__dout = Yvec_inst_2_if_dout;
  assign Yvec_inst_2__empty_n = Yvec_inst_2_if_empty_n;
  assign Yvec_inst_2__full_n = Yvec_inst_2_if_full_n;
  assign Yvec_inst_2_if_read = Yvec_inst_2__read;
  assign Yvec_inst_2_if_read_ce = 1'b1;
  assign Yvec_inst_2_if_write = Yvec_inst_2__write;
  assign Yvec_inst_2_if_write_ce = 1'b1;
  assign Yvec_inst_2_reset = ~ ap_rst_n;
  assign Yvec_inst_30_clk = ap_clk;
  assign Yvec_inst_30_if_din = Yvec_inst_30__din;
  assign Yvec_inst_30__dout = Yvec_inst_30_if_dout;
  assign Yvec_inst_30__empty_n = Yvec_inst_30_if_empty_n;
  assign Yvec_inst_30__full_n = Yvec_inst_30_if_full_n;
  assign Yvec_inst_30_if_read = Yvec_inst_30__read;
  assign Yvec_inst_30_if_read_ce = 1'b1;
  assign Yvec_inst_30_if_write = Yvec_inst_30__write;
  assign Yvec_inst_30_if_write_ce = 1'b1;
  assign Yvec_inst_30_reset = ~ ap_rst_n;
  assign Yvec_inst_31_clk = ap_clk;
  assign Yvec_inst_31_if_din = Yvec_inst_31__din;
  assign Yvec_inst_31__dout = Yvec_inst_31_if_dout;
  assign Yvec_inst_31__empty_n = Yvec_inst_31_if_empty_n;
  assign Yvec_inst_31__full_n = Yvec_inst_31_if_full_n;
  assign Yvec_inst_31_if_read = Yvec_inst_31__read;
  assign Yvec_inst_31_if_read_ce = 1'b1;
  assign Yvec_inst_31_if_write = Yvec_inst_31__write;
  assign Yvec_inst_31_if_write_ce = 1'b1;
  assign Yvec_inst_31_reset = ~ ap_rst_n;
  assign Yvec_inst_32_clk = ap_clk;
  assign Yvec_inst_32_if_din = Yvec_inst_32__din;
  assign Yvec_inst_32__dout = Yvec_inst_32_if_dout;
  assign Yvec_inst_32__empty_n = Yvec_inst_32_if_empty_n;
  assign Yvec_inst_32__full_n = Yvec_inst_32_if_full_n;
  assign Yvec_inst_32_if_read = Yvec_inst_32__read;
  assign Yvec_inst_32_if_read_ce = 1'b1;
  assign Yvec_inst_32_if_write = Yvec_inst_32__write;
  assign Yvec_inst_32_if_write_ce = 1'b1;
  assign Yvec_inst_32_reset = ~ ap_rst_n;
  assign Yvec_inst_33_clk = ap_clk;
  assign Yvec_inst_33_if_din = Yvec_inst_33__din;
  assign Yvec_inst_33__dout = Yvec_inst_33_if_dout;
  assign Yvec_inst_33__empty_n = Yvec_inst_33_if_empty_n;
  assign Yvec_inst_33__full_n = Yvec_inst_33_if_full_n;
  assign Yvec_inst_33_if_read = Yvec_inst_33__read;
  assign Yvec_inst_33_if_read_ce = 1'b1;
  assign Yvec_inst_33_if_write = Yvec_inst_33__write;
  assign Yvec_inst_33_if_write_ce = 1'b1;
  assign Yvec_inst_33_reset = ~ ap_rst_n;
  assign Yvec_inst_34_clk = ap_clk;
  assign Yvec_inst_34_if_din = Yvec_inst_34__din;
  assign Yvec_inst_34__dout = Yvec_inst_34_if_dout;
  assign Yvec_inst_34__empty_n = Yvec_inst_34_if_empty_n;
  assign Yvec_inst_34__full_n = Yvec_inst_34_if_full_n;
  assign Yvec_inst_34_if_read = Yvec_inst_34__read;
  assign Yvec_inst_34_if_read_ce = 1'b1;
  assign Yvec_inst_34_if_write = Yvec_inst_34__write;
  assign Yvec_inst_34_if_write_ce = 1'b1;
  assign Yvec_inst_34_reset = ~ ap_rst_n;
  assign Yvec_inst_35_clk = ap_clk;
  assign Yvec_inst_35_if_din = Yvec_inst_35__din;
  assign Yvec_inst_35__dout = Yvec_inst_35_if_dout;
  assign Yvec_inst_35__empty_n = Yvec_inst_35_if_empty_n;
  assign Yvec_inst_35__full_n = Yvec_inst_35_if_full_n;
  assign Yvec_inst_35_if_read = Yvec_inst_35__read;
  assign Yvec_inst_35_if_read_ce = 1'b1;
  assign Yvec_inst_35_if_write = Yvec_inst_35__write;
  assign Yvec_inst_35_if_write_ce = 1'b1;
  assign Yvec_inst_35_reset = ~ ap_rst_n;
  assign Yvec_inst_36_clk = ap_clk;
  assign Yvec_inst_36_if_din = Yvec_inst_36__din;
  assign Yvec_inst_36__dout = Yvec_inst_36_if_dout;
  assign Yvec_inst_36__empty_n = Yvec_inst_36_if_empty_n;
  assign Yvec_inst_36__full_n = Yvec_inst_36_if_full_n;
  assign Yvec_inst_36_if_read = Yvec_inst_36__read;
  assign Yvec_inst_36_if_read_ce = 1'b1;
  assign Yvec_inst_36_if_write = Yvec_inst_36__write;
  assign Yvec_inst_36_if_write_ce = 1'b1;
  assign Yvec_inst_36_reset = ~ ap_rst_n;
  assign Yvec_inst_37_clk = ap_clk;
  assign Yvec_inst_37_if_din = Yvec_inst_37__din;
  assign Yvec_inst_37__dout = Yvec_inst_37_if_dout;
  assign Yvec_inst_37__empty_n = Yvec_inst_37_if_empty_n;
  assign Yvec_inst_37__full_n = Yvec_inst_37_if_full_n;
  assign Yvec_inst_37_if_read = Yvec_inst_37__read;
  assign Yvec_inst_37_if_read_ce = 1'b1;
  assign Yvec_inst_37_if_write = Yvec_inst_37__write;
  assign Yvec_inst_37_if_write_ce = 1'b1;
  assign Yvec_inst_37_reset = ~ ap_rst_n;
  assign Yvec_inst_38_clk = ap_clk;
  assign Yvec_inst_38_if_din = Yvec_inst_38__din;
  assign Yvec_inst_38__dout = Yvec_inst_38_if_dout;
  assign Yvec_inst_38__empty_n = Yvec_inst_38_if_empty_n;
  assign Yvec_inst_38__full_n = Yvec_inst_38_if_full_n;
  assign Yvec_inst_38_if_read = Yvec_inst_38__read;
  assign Yvec_inst_38_if_read_ce = 1'b1;
  assign Yvec_inst_38_if_write = Yvec_inst_38__write;
  assign Yvec_inst_38_if_write_ce = 1'b1;
  assign Yvec_inst_38_reset = ~ ap_rst_n;
  assign Yvec_inst_39_clk = ap_clk;
  assign Yvec_inst_39_if_din = Yvec_inst_39__din;
  assign Yvec_inst_39__dout = Yvec_inst_39_if_dout;
  assign Yvec_inst_39__empty_n = Yvec_inst_39_if_empty_n;
  assign Yvec_inst_39__full_n = Yvec_inst_39_if_full_n;
  assign Yvec_inst_39_if_read = Yvec_inst_39__read;
  assign Yvec_inst_39_if_read_ce = 1'b1;
  assign Yvec_inst_39_if_write = Yvec_inst_39__write;
  assign Yvec_inst_39_if_write_ce = 1'b1;
  assign Yvec_inst_39_reset = ~ ap_rst_n;
  assign Yvec_inst_3_clk = ap_clk;
  assign Yvec_inst_3_if_din = Yvec_inst_3__din;
  assign Yvec_inst_3__dout = Yvec_inst_3_if_dout;
  assign Yvec_inst_3__empty_n = Yvec_inst_3_if_empty_n;
  assign Yvec_inst_3__full_n = Yvec_inst_3_if_full_n;
  assign Yvec_inst_3_if_read = Yvec_inst_3__read;
  assign Yvec_inst_3_if_read_ce = 1'b1;
  assign Yvec_inst_3_if_write = Yvec_inst_3__write;
  assign Yvec_inst_3_if_write_ce = 1'b1;
  assign Yvec_inst_3_reset = ~ ap_rst_n;
  assign Yvec_inst_40_clk = ap_clk;
  assign Yvec_inst_40_if_din = Yvec_inst_40__din;
  assign Yvec_inst_40__dout = Yvec_inst_40_if_dout;
  assign Yvec_inst_40__empty_n = Yvec_inst_40_if_empty_n;
  assign Yvec_inst_40__full_n = Yvec_inst_40_if_full_n;
  assign Yvec_inst_40_if_read = Yvec_inst_40__read;
  assign Yvec_inst_40_if_read_ce = 1'b1;
  assign Yvec_inst_40_if_write = Yvec_inst_40__write;
  assign Yvec_inst_40_if_write_ce = 1'b1;
  assign Yvec_inst_40_reset = ~ ap_rst_n;
  assign Yvec_inst_41_clk = ap_clk;
  assign Yvec_inst_41_if_din = Yvec_inst_41__din;
  assign Yvec_inst_41__dout = Yvec_inst_41_if_dout;
  assign Yvec_inst_41__empty_n = Yvec_inst_41_if_empty_n;
  assign Yvec_inst_41__full_n = Yvec_inst_41_if_full_n;
  assign Yvec_inst_41_if_read = Yvec_inst_41__read;
  assign Yvec_inst_41_if_read_ce = 1'b1;
  assign Yvec_inst_41_if_write = Yvec_inst_41__write;
  assign Yvec_inst_41_if_write_ce = 1'b1;
  assign Yvec_inst_41_reset = ~ ap_rst_n;
  assign Yvec_inst_42_clk = ap_clk;
  assign Yvec_inst_42_if_din = Yvec_inst_42__din;
  assign Yvec_inst_42__dout = Yvec_inst_42_if_dout;
  assign Yvec_inst_42__empty_n = Yvec_inst_42_if_empty_n;
  assign Yvec_inst_42__full_n = Yvec_inst_42_if_full_n;
  assign Yvec_inst_42_if_read = Yvec_inst_42__read;
  assign Yvec_inst_42_if_read_ce = 1'b1;
  assign Yvec_inst_42_if_write = Yvec_inst_42__write;
  assign Yvec_inst_42_if_write_ce = 1'b1;
  assign Yvec_inst_42_reset = ~ ap_rst_n;
  assign Yvec_inst_43_clk = ap_clk;
  assign Yvec_inst_43_if_din = Yvec_inst_43__din;
  assign Yvec_inst_43__dout = Yvec_inst_43_if_dout;
  assign Yvec_inst_43__empty_n = Yvec_inst_43_if_empty_n;
  assign Yvec_inst_43__full_n = Yvec_inst_43_if_full_n;
  assign Yvec_inst_43_if_read = Yvec_inst_43__read;
  assign Yvec_inst_43_if_read_ce = 1'b1;
  assign Yvec_inst_43_if_write = Yvec_inst_43__write;
  assign Yvec_inst_43_if_write_ce = 1'b1;
  assign Yvec_inst_43_reset = ~ ap_rst_n;
  assign Yvec_inst_44_clk = ap_clk;
  assign Yvec_inst_44_if_din = Yvec_inst_44__din;
  assign Yvec_inst_44__dout = Yvec_inst_44_if_dout;
  assign Yvec_inst_44__empty_n = Yvec_inst_44_if_empty_n;
  assign Yvec_inst_44__full_n = Yvec_inst_44_if_full_n;
  assign Yvec_inst_44_if_read = Yvec_inst_44__read;
  assign Yvec_inst_44_if_read_ce = 1'b1;
  assign Yvec_inst_44_if_write = Yvec_inst_44__write;
  assign Yvec_inst_44_if_write_ce = 1'b1;
  assign Yvec_inst_44_reset = ~ ap_rst_n;
  assign Yvec_inst_45_clk = ap_clk;
  assign Yvec_inst_45_if_din = Yvec_inst_45__din;
  assign Yvec_inst_45__dout = Yvec_inst_45_if_dout;
  assign Yvec_inst_45__empty_n = Yvec_inst_45_if_empty_n;
  assign Yvec_inst_45__full_n = Yvec_inst_45_if_full_n;
  assign Yvec_inst_45_if_read = Yvec_inst_45__read;
  assign Yvec_inst_45_if_read_ce = 1'b1;
  assign Yvec_inst_45_if_write = Yvec_inst_45__write;
  assign Yvec_inst_45_if_write_ce = 1'b1;
  assign Yvec_inst_45_reset = ~ ap_rst_n;
  assign Yvec_inst_46_clk = ap_clk;
  assign Yvec_inst_46_if_din = Yvec_inst_46__din;
  assign Yvec_inst_46__dout = Yvec_inst_46_if_dout;
  assign Yvec_inst_46__empty_n = Yvec_inst_46_if_empty_n;
  assign Yvec_inst_46__full_n = Yvec_inst_46_if_full_n;
  assign Yvec_inst_46_if_read = Yvec_inst_46__read;
  assign Yvec_inst_46_if_read_ce = 1'b1;
  assign Yvec_inst_46_if_write = Yvec_inst_46__write;
  assign Yvec_inst_46_if_write_ce = 1'b1;
  assign Yvec_inst_46_reset = ~ ap_rst_n;
  assign Yvec_inst_47_clk = ap_clk;
  assign Yvec_inst_47_if_din = Yvec_inst_47__din;
  assign Yvec_inst_47__dout = Yvec_inst_47_if_dout;
  assign Yvec_inst_47__empty_n = Yvec_inst_47_if_empty_n;
  assign Yvec_inst_47__full_n = Yvec_inst_47_if_full_n;
  assign Yvec_inst_47_if_read = Yvec_inst_47__read;
  assign Yvec_inst_47_if_read_ce = 1'b1;
  assign Yvec_inst_47_if_write = Yvec_inst_47__write;
  assign Yvec_inst_47_if_write_ce = 1'b1;
  assign Yvec_inst_47_reset = ~ ap_rst_n;
  assign Yvec_inst_4_clk = ap_clk;
  assign Yvec_inst_4_if_din = Yvec_inst_4__din;
  assign Yvec_inst_4__dout = Yvec_inst_4_if_dout;
  assign Yvec_inst_4__empty_n = Yvec_inst_4_if_empty_n;
  assign Yvec_inst_4__full_n = Yvec_inst_4_if_full_n;
  assign Yvec_inst_4_if_read = Yvec_inst_4__read;
  assign Yvec_inst_4_if_read_ce = 1'b1;
  assign Yvec_inst_4_if_write = Yvec_inst_4__write;
  assign Yvec_inst_4_if_write_ce = 1'b1;
  assign Yvec_inst_4_reset = ~ ap_rst_n;
  assign Yvec_inst_5_clk = ap_clk;
  assign Yvec_inst_5_if_din = Yvec_inst_5__din;
  assign Yvec_inst_5__dout = Yvec_inst_5_if_dout;
  assign Yvec_inst_5__empty_n = Yvec_inst_5_if_empty_n;
  assign Yvec_inst_5__full_n = Yvec_inst_5_if_full_n;
  assign Yvec_inst_5_if_read = Yvec_inst_5__read;
  assign Yvec_inst_5_if_read_ce = 1'b1;
  assign Yvec_inst_5_if_write = Yvec_inst_5__write;
  assign Yvec_inst_5_if_write_ce = 1'b1;
  assign Yvec_inst_5_reset = ~ ap_rst_n;
  assign Yvec_inst_6_clk = ap_clk;
  assign Yvec_inst_6_if_din = Yvec_inst_6__din;
  assign Yvec_inst_6__dout = Yvec_inst_6_if_dout;
  assign Yvec_inst_6__empty_n = Yvec_inst_6_if_empty_n;
  assign Yvec_inst_6__full_n = Yvec_inst_6_if_full_n;
  assign Yvec_inst_6_if_read = Yvec_inst_6__read;
  assign Yvec_inst_6_if_read_ce = 1'b1;
  assign Yvec_inst_6_if_write = Yvec_inst_6__write;
  assign Yvec_inst_6_if_write_ce = 1'b1;
  assign Yvec_inst_6_reset = ~ ap_rst_n;
  assign Yvec_inst_7_clk = ap_clk;
  assign Yvec_inst_7_if_din = Yvec_inst_7__din;
  assign Yvec_inst_7__dout = Yvec_inst_7_if_dout;
  assign Yvec_inst_7__empty_n = Yvec_inst_7_if_empty_n;
  assign Yvec_inst_7__full_n = Yvec_inst_7_if_full_n;
  assign Yvec_inst_7_if_read = Yvec_inst_7__read;
  assign Yvec_inst_7_if_read_ce = 1'b1;
  assign Yvec_inst_7_if_write = Yvec_inst_7__write;
  assign Yvec_inst_7_if_write_ce = 1'b1;
  assign Yvec_inst_7_reset = ~ ap_rst_n;
  assign Yvec_inst_8_clk = ap_clk;
  assign Yvec_inst_8_if_din = Yvec_inst_8__din;
  assign Yvec_inst_8__dout = Yvec_inst_8_if_dout;
  assign Yvec_inst_8__empty_n = Yvec_inst_8_if_empty_n;
  assign Yvec_inst_8__full_n = Yvec_inst_8_if_full_n;
  assign Yvec_inst_8_if_read = Yvec_inst_8__read;
  assign Yvec_inst_8_if_read_ce = 1'b1;
  assign Yvec_inst_8_if_write = Yvec_inst_8__write;
  assign Yvec_inst_8_if_write_ce = 1'b1;
  assign Yvec_inst_8_reset = ~ ap_rst_n;
  assign Yvec_inst_9_clk = ap_clk;
  assign Yvec_inst_9_if_din = Yvec_inst_9__din;
  assign Yvec_inst_9__dout = Yvec_inst_9_if_dout;
  assign Yvec_inst_9__empty_n = Yvec_inst_9_if_empty_n;
  assign Yvec_inst_9__full_n = Yvec_inst_9_if_full_n;
  assign Yvec_inst_9_if_read = Yvec_inst_9__read;
  assign Yvec_inst_9_if_read_ce = 1'b1;
  assign Yvec_inst_9_if_write = Yvec_inst_9__write;
  assign Yvec_inst_9_if_write_ce = 1'b1;
  assign Yvec_inst_9_reset = ~ ap_rst_n;
  assign fifo_A_0_clk = ap_clk;
  assign fifo_A_0_if_din = fifo_A_0__din;
  assign fifo_A_0__dout = fifo_A_0_if_dout;
  assign fifo_A_0__empty_n = fifo_A_0_if_empty_n;
  assign fifo_A_0__full_n = fifo_A_0_if_full_n;
  assign fifo_A_0_if_read = fifo_A_0__read;
  assign fifo_A_0_if_read_ce = 1'b1;
  assign fifo_A_0_if_write = fifo_A_0__write;
  assign fifo_A_0_if_write_ce = 1'b1;
  assign fifo_A_0_reset = ~ ap_rst_n;
  assign fifo_A_10_clk = ap_clk;
  assign fifo_A_10_if_din = fifo_A_10__din;
  assign fifo_A_10__dout = fifo_A_10_if_dout;
  assign fifo_A_10__empty_n = fifo_A_10_if_empty_n;
  assign fifo_A_10__full_n = fifo_A_10_if_full_n;
  assign fifo_A_10_if_read = fifo_A_10__read;
  assign fifo_A_10_if_read_ce = 1'b1;
  assign fifo_A_10_if_write = fifo_A_10__write;
  assign fifo_A_10_if_write_ce = 1'b1;
  assign fifo_A_10_reset = ~ ap_rst_n;
  assign fifo_A_11_clk = ap_clk;
  assign fifo_A_11_if_din = fifo_A_11__din;
  assign fifo_A_11__dout = fifo_A_11_if_dout;
  assign fifo_A_11__empty_n = fifo_A_11_if_empty_n;
  assign fifo_A_11__full_n = fifo_A_11_if_full_n;
  assign fifo_A_11_if_read = fifo_A_11__read;
  assign fifo_A_11_if_read_ce = 1'b1;
  assign fifo_A_11_if_write = fifo_A_11__write;
  assign fifo_A_11_if_write_ce = 1'b1;
  assign fifo_A_11_reset = ~ ap_rst_n;
  assign fifo_A_12_clk = ap_clk;
  assign fifo_A_12_if_din = fifo_A_12__din;
  assign fifo_A_12__dout = fifo_A_12_if_dout;
  assign fifo_A_12__empty_n = fifo_A_12_if_empty_n;
  assign fifo_A_12__full_n = fifo_A_12_if_full_n;
  assign fifo_A_12_if_read = fifo_A_12__read;
  assign fifo_A_12_if_read_ce = 1'b1;
  assign fifo_A_12_if_write = fifo_A_12__write;
  assign fifo_A_12_if_write_ce = 1'b1;
  assign fifo_A_12_reset = ~ ap_rst_n;
  assign fifo_A_13_clk = ap_clk;
  assign fifo_A_13_if_din = fifo_A_13__din;
  assign fifo_A_13__dout = fifo_A_13_if_dout;
  assign fifo_A_13__empty_n = fifo_A_13_if_empty_n;
  assign fifo_A_13__full_n = fifo_A_13_if_full_n;
  assign fifo_A_13_if_read = fifo_A_13__read;
  assign fifo_A_13_if_read_ce = 1'b1;
  assign fifo_A_13_if_write = fifo_A_13__write;
  assign fifo_A_13_if_write_ce = 1'b1;
  assign fifo_A_13_reset = ~ ap_rst_n;
  assign fifo_A_14_clk = ap_clk;
  assign fifo_A_14_if_din = fifo_A_14__din;
  assign fifo_A_14__dout = fifo_A_14_if_dout;
  assign fifo_A_14__empty_n = fifo_A_14_if_empty_n;
  assign fifo_A_14__full_n = fifo_A_14_if_full_n;
  assign fifo_A_14_if_read = fifo_A_14__read;
  assign fifo_A_14_if_read_ce = 1'b1;
  assign fifo_A_14_if_write = fifo_A_14__write;
  assign fifo_A_14_if_write_ce = 1'b1;
  assign fifo_A_14_reset = ~ ap_rst_n;
  assign fifo_A_15_clk = ap_clk;
  assign fifo_A_15_if_din = fifo_A_15__din;
  assign fifo_A_15__dout = fifo_A_15_if_dout;
  assign fifo_A_15__empty_n = fifo_A_15_if_empty_n;
  assign fifo_A_15__full_n = fifo_A_15_if_full_n;
  assign fifo_A_15_if_read = fifo_A_15__read;
  assign fifo_A_15_if_read_ce = 1'b1;
  assign fifo_A_15_if_write = fifo_A_15__write;
  assign fifo_A_15_if_write_ce = 1'b1;
  assign fifo_A_15_reset = ~ ap_rst_n;
  assign fifo_A_16_clk = ap_clk;
  assign fifo_A_16_if_din = fifo_A_16__din;
  assign fifo_A_16__dout = fifo_A_16_if_dout;
  assign fifo_A_16__empty_n = fifo_A_16_if_empty_n;
  assign fifo_A_16__full_n = fifo_A_16_if_full_n;
  assign fifo_A_16_if_read = fifo_A_16__read;
  assign fifo_A_16_if_read_ce = 1'b1;
  assign fifo_A_16_if_write = fifo_A_16__write;
  assign fifo_A_16_if_write_ce = 1'b1;
  assign fifo_A_16_reset = ~ ap_rst_n;
  assign fifo_A_17_clk = ap_clk;
  assign fifo_A_17_if_din = fifo_A_17__din;
  assign fifo_A_17__dout = fifo_A_17_if_dout;
  assign fifo_A_17__empty_n = fifo_A_17_if_empty_n;
  assign fifo_A_17__full_n = fifo_A_17_if_full_n;
  assign fifo_A_17_if_read = fifo_A_17__read;
  assign fifo_A_17_if_read_ce = 1'b1;
  assign fifo_A_17_if_write = fifo_A_17__write;
  assign fifo_A_17_if_write_ce = 1'b1;
  assign fifo_A_17_reset = ~ ap_rst_n;
  assign fifo_A_18_clk = ap_clk;
  assign fifo_A_18_if_din = fifo_A_18__din;
  assign fifo_A_18__dout = fifo_A_18_if_dout;
  assign fifo_A_18__empty_n = fifo_A_18_if_empty_n;
  assign fifo_A_18__full_n = fifo_A_18_if_full_n;
  assign fifo_A_18_if_read = fifo_A_18__read;
  assign fifo_A_18_if_read_ce = 1'b1;
  assign fifo_A_18_if_write = fifo_A_18__write;
  assign fifo_A_18_if_write_ce = 1'b1;
  assign fifo_A_18_reset = ~ ap_rst_n;
  assign fifo_A_19_clk = ap_clk;
  assign fifo_A_19_if_din = fifo_A_19__din;
  assign fifo_A_19__dout = fifo_A_19_if_dout;
  assign fifo_A_19__empty_n = fifo_A_19_if_empty_n;
  assign fifo_A_19__full_n = fifo_A_19_if_full_n;
  assign fifo_A_19_if_read = fifo_A_19__read;
  assign fifo_A_19_if_read_ce = 1'b1;
  assign fifo_A_19_if_write = fifo_A_19__write;
  assign fifo_A_19_if_write_ce = 1'b1;
  assign fifo_A_19_reset = ~ ap_rst_n;
  assign fifo_A_1_clk = ap_clk;
  assign fifo_A_1_if_din = fifo_A_1__din;
  assign fifo_A_1__dout = fifo_A_1_if_dout;
  assign fifo_A_1__empty_n = fifo_A_1_if_empty_n;
  assign fifo_A_1__full_n = fifo_A_1_if_full_n;
  assign fifo_A_1_if_read = fifo_A_1__read;
  assign fifo_A_1_if_read_ce = 1'b1;
  assign fifo_A_1_if_write = fifo_A_1__write;
  assign fifo_A_1_if_write_ce = 1'b1;
  assign fifo_A_1_reset = ~ ap_rst_n;
  assign fifo_A_20_clk = ap_clk;
  assign fifo_A_20_if_din = fifo_A_20__din;
  assign fifo_A_20__dout = fifo_A_20_if_dout;
  assign fifo_A_20__empty_n = fifo_A_20_if_empty_n;
  assign fifo_A_20__full_n = fifo_A_20_if_full_n;
  assign fifo_A_20_if_read = fifo_A_20__read;
  assign fifo_A_20_if_read_ce = 1'b1;
  assign fifo_A_20_if_write = fifo_A_20__write;
  assign fifo_A_20_if_write_ce = 1'b1;
  assign fifo_A_20_reset = ~ ap_rst_n;
  assign fifo_A_21_clk = ap_clk;
  assign fifo_A_21_if_din = fifo_A_21__din;
  assign fifo_A_21__dout = fifo_A_21_if_dout;
  assign fifo_A_21__empty_n = fifo_A_21_if_empty_n;
  assign fifo_A_21__full_n = fifo_A_21_if_full_n;
  assign fifo_A_21_if_read = fifo_A_21__read;
  assign fifo_A_21_if_read_ce = 1'b1;
  assign fifo_A_21_if_write = fifo_A_21__write;
  assign fifo_A_21_if_write_ce = 1'b1;
  assign fifo_A_21_reset = ~ ap_rst_n;
  assign fifo_A_22_clk = ap_clk;
  assign fifo_A_22_if_din = fifo_A_22__din;
  assign fifo_A_22__dout = fifo_A_22_if_dout;
  assign fifo_A_22__empty_n = fifo_A_22_if_empty_n;
  assign fifo_A_22__full_n = fifo_A_22_if_full_n;
  assign fifo_A_22_if_read = fifo_A_22__read;
  assign fifo_A_22_if_read_ce = 1'b1;
  assign fifo_A_22_if_write = fifo_A_22__write;
  assign fifo_A_22_if_write_ce = 1'b1;
  assign fifo_A_22_reset = ~ ap_rst_n;
  assign fifo_A_23_clk = ap_clk;
  assign fifo_A_23_if_din = fifo_A_23__din;
  assign fifo_A_23__dout = fifo_A_23_if_dout;
  assign fifo_A_23__empty_n = fifo_A_23_if_empty_n;
  assign fifo_A_23__full_n = fifo_A_23_if_full_n;
  assign fifo_A_23_if_read = fifo_A_23__read;
  assign fifo_A_23_if_read_ce = 1'b1;
  assign fifo_A_23_if_write = fifo_A_23__write;
  assign fifo_A_23_if_write_ce = 1'b1;
  assign fifo_A_23_reset = ~ ap_rst_n;
  assign fifo_A_24_clk = ap_clk;
  assign fifo_A_24_if_din = fifo_A_24__din;
  assign fifo_A_24__dout = fifo_A_24_if_dout;
  assign fifo_A_24__empty_n = fifo_A_24_if_empty_n;
  assign fifo_A_24__full_n = fifo_A_24_if_full_n;
  assign fifo_A_24_if_read = fifo_A_24__read;
  assign fifo_A_24_if_read_ce = 1'b1;
  assign fifo_A_24_if_write = fifo_A_24__write;
  assign fifo_A_24_if_write_ce = 1'b1;
  assign fifo_A_24_reset = ~ ap_rst_n;
  assign fifo_A_25_clk = ap_clk;
  assign fifo_A_25_if_din = fifo_A_25__din;
  assign fifo_A_25__dout = fifo_A_25_if_dout;
  assign fifo_A_25__empty_n = fifo_A_25_if_empty_n;
  assign fifo_A_25__full_n = fifo_A_25_if_full_n;
  assign fifo_A_25_if_read = fifo_A_25__read;
  assign fifo_A_25_if_read_ce = 1'b1;
  assign fifo_A_25_if_write = fifo_A_25__write;
  assign fifo_A_25_if_write_ce = 1'b1;
  assign fifo_A_25_reset = ~ ap_rst_n;
  assign fifo_A_26_clk = ap_clk;
  assign fifo_A_26_if_din = fifo_A_26__din;
  assign fifo_A_26__dout = fifo_A_26_if_dout;
  assign fifo_A_26__empty_n = fifo_A_26_if_empty_n;
  assign fifo_A_26__full_n = fifo_A_26_if_full_n;
  assign fifo_A_26_if_read = fifo_A_26__read;
  assign fifo_A_26_if_read_ce = 1'b1;
  assign fifo_A_26_if_write = fifo_A_26__write;
  assign fifo_A_26_if_write_ce = 1'b1;
  assign fifo_A_26_reset = ~ ap_rst_n;
  assign fifo_A_27_clk = ap_clk;
  assign fifo_A_27_if_din = fifo_A_27__din;
  assign fifo_A_27__dout = fifo_A_27_if_dout;
  assign fifo_A_27__empty_n = fifo_A_27_if_empty_n;
  assign fifo_A_27__full_n = fifo_A_27_if_full_n;
  assign fifo_A_27_if_read = fifo_A_27__read;
  assign fifo_A_27_if_read_ce = 1'b1;
  assign fifo_A_27_if_write = fifo_A_27__write;
  assign fifo_A_27_if_write_ce = 1'b1;
  assign fifo_A_27_reset = ~ ap_rst_n;
  assign fifo_A_28_clk = ap_clk;
  assign fifo_A_28_if_din = fifo_A_28__din;
  assign fifo_A_28__dout = fifo_A_28_if_dout;
  assign fifo_A_28__empty_n = fifo_A_28_if_empty_n;
  assign fifo_A_28__full_n = fifo_A_28_if_full_n;
  assign fifo_A_28_if_read = fifo_A_28__read;
  assign fifo_A_28_if_read_ce = 1'b1;
  assign fifo_A_28_if_write = fifo_A_28__write;
  assign fifo_A_28_if_write_ce = 1'b1;
  assign fifo_A_28_reset = ~ ap_rst_n;
  assign fifo_A_29_clk = ap_clk;
  assign fifo_A_29_if_din = fifo_A_29__din;
  assign fifo_A_29__dout = fifo_A_29_if_dout;
  assign fifo_A_29__empty_n = fifo_A_29_if_empty_n;
  assign fifo_A_29__full_n = fifo_A_29_if_full_n;
  assign fifo_A_29_if_read = fifo_A_29__read;
  assign fifo_A_29_if_read_ce = 1'b1;
  assign fifo_A_29_if_write = fifo_A_29__write;
  assign fifo_A_29_if_write_ce = 1'b1;
  assign fifo_A_29_reset = ~ ap_rst_n;
  assign fifo_A_2_clk = ap_clk;
  assign fifo_A_2_if_din = fifo_A_2__din;
  assign fifo_A_2__dout = fifo_A_2_if_dout;
  assign fifo_A_2__empty_n = fifo_A_2_if_empty_n;
  assign fifo_A_2__full_n = fifo_A_2_if_full_n;
  assign fifo_A_2_if_read = fifo_A_2__read;
  assign fifo_A_2_if_read_ce = 1'b1;
  assign fifo_A_2_if_write = fifo_A_2__write;
  assign fifo_A_2_if_write_ce = 1'b1;
  assign fifo_A_2_reset = ~ ap_rst_n;
  assign fifo_A_30_clk = ap_clk;
  assign fifo_A_30_if_din = fifo_A_30__din;
  assign fifo_A_30__dout = fifo_A_30_if_dout;
  assign fifo_A_30__empty_n = fifo_A_30_if_empty_n;
  assign fifo_A_30__full_n = fifo_A_30_if_full_n;
  assign fifo_A_30_if_read = fifo_A_30__read;
  assign fifo_A_30_if_read_ce = 1'b1;
  assign fifo_A_30_if_write = fifo_A_30__write;
  assign fifo_A_30_if_write_ce = 1'b1;
  assign fifo_A_30_reset = ~ ap_rst_n;
  assign fifo_A_31_clk = ap_clk;
  assign fifo_A_31_if_din = fifo_A_31__din;
  assign fifo_A_31__dout = fifo_A_31_if_dout;
  assign fifo_A_31__empty_n = fifo_A_31_if_empty_n;
  assign fifo_A_31__full_n = fifo_A_31_if_full_n;
  assign fifo_A_31_if_read = fifo_A_31__read;
  assign fifo_A_31_if_read_ce = 1'b1;
  assign fifo_A_31_if_write = fifo_A_31__write;
  assign fifo_A_31_if_write_ce = 1'b1;
  assign fifo_A_31_reset = ~ ap_rst_n;
  assign fifo_A_32_clk = ap_clk;
  assign fifo_A_32_if_din = fifo_A_32__din;
  assign fifo_A_32__dout = fifo_A_32_if_dout;
  assign fifo_A_32__empty_n = fifo_A_32_if_empty_n;
  assign fifo_A_32__full_n = fifo_A_32_if_full_n;
  assign fifo_A_32_if_read = fifo_A_32__read;
  assign fifo_A_32_if_read_ce = 1'b1;
  assign fifo_A_32_if_write = fifo_A_32__write;
  assign fifo_A_32_if_write_ce = 1'b1;
  assign fifo_A_32_reset = ~ ap_rst_n;
  assign fifo_A_33_clk = ap_clk;
  assign fifo_A_33_if_din = fifo_A_33__din;
  assign fifo_A_33__dout = fifo_A_33_if_dout;
  assign fifo_A_33__empty_n = fifo_A_33_if_empty_n;
  assign fifo_A_33__full_n = fifo_A_33_if_full_n;
  assign fifo_A_33_if_read = fifo_A_33__read;
  assign fifo_A_33_if_read_ce = 1'b1;
  assign fifo_A_33_if_write = fifo_A_33__write;
  assign fifo_A_33_if_write_ce = 1'b1;
  assign fifo_A_33_reset = ~ ap_rst_n;
  assign fifo_A_34_clk = ap_clk;
  assign fifo_A_34_if_din = fifo_A_34__din;
  assign fifo_A_34__dout = fifo_A_34_if_dout;
  assign fifo_A_34__empty_n = fifo_A_34_if_empty_n;
  assign fifo_A_34__full_n = fifo_A_34_if_full_n;
  assign fifo_A_34_if_read = fifo_A_34__read;
  assign fifo_A_34_if_read_ce = 1'b1;
  assign fifo_A_34_if_write = fifo_A_34__write;
  assign fifo_A_34_if_write_ce = 1'b1;
  assign fifo_A_34_reset = ~ ap_rst_n;
  assign fifo_A_35_clk = ap_clk;
  assign fifo_A_35_if_din = fifo_A_35__din;
  assign fifo_A_35__dout = fifo_A_35_if_dout;
  assign fifo_A_35__empty_n = fifo_A_35_if_empty_n;
  assign fifo_A_35__full_n = fifo_A_35_if_full_n;
  assign fifo_A_35_if_read = fifo_A_35__read;
  assign fifo_A_35_if_read_ce = 1'b1;
  assign fifo_A_35_if_write = fifo_A_35__write;
  assign fifo_A_35_if_write_ce = 1'b1;
  assign fifo_A_35_reset = ~ ap_rst_n;
  assign fifo_A_36_clk = ap_clk;
  assign fifo_A_36_if_din = fifo_A_36__din;
  assign fifo_A_36__dout = fifo_A_36_if_dout;
  assign fifo_A_36__empty_n = fifo_A_36_if_empty_n;
  assign fifo_A_36__full_n = fifo_A_36_if_full_n;
  assign fifo_A_36_if_read = fifo_A_36__read;
  assign fifo_A_36_if_read_ce = 1'b1;
  assign fifo_A_36_if_write = fifo_A_36__write;
  assign fifo_A_36_if_write_ce = 1'b1;
  assign fifo_A_36_reset = ~ ap_rst_n;
  assign fifo_A_37_clk = ap_clk;
  assign fifo_A_37_if_din = fifo_A_37__din;
  assign fifo_A_37__dout = fifo_A_37_if_dout;
  assign fifo_A_37__empty_n = fifo_A_37_if_empty_n;
  assign fifo_A_37__full_n = fifo_A_37_if_full_n;
  assign fifo_A_37_if_read = fifo_A_37__read;
  assign fifo_A_37_if_read_ce = 1'b1;
  assign fifo_A_37_if_write = fifo_A_37__write;
  assign fifo_A_37_if_write_ce = 1'b1;
  assign fifo_A_37_reset = ~ ap_rst_n;
  assign fifo_A_38_clk = ap_clk;
  assign fifo_A_38_if_din = fifo_A_38__din;
  assign fifo_A_38__dout = fifo_A_38_if_dout;
  assign fifo_A_38__empty_n = fifo_A_38_if_empty_n;
  assign fifo_A_38__full_n = fifo_A_38_if_full_n;
  assign fifo_A_38_if_read = fifo_A_38__read;
  assign fifo_A_38_if_read_ce = 1'b1;
  assign fifo_A_38_if_write = fifo_A_38__write;
  assign fifo_A_38_if_write_ce = 1'b1;
  assign fifo_A_38_reset = ~ ap_rst_n;
  assign fifo_A_39_clk = ap_clk;
  assign fifo_A_39_if_din = fifo_A_39__din;
  assign fifo_A_39__dout = fifo_A_39_if_dout;
  assign fifo_A_39__empty_n = fifo_A_39_if_empty_n;
  assign fifo_A_39__full_n = fifo_A_39_if_full_n;
  assign fifo_A_39_if_read = fifo_A_39__read;
  assign fifo_A_39_if_read_ce = 1'b1;
  assign fifo_A_39_if_write = fifo_A_39__write;
  assign fifo_A_39_if_write_ce = 1'b1;
  assign fifo_A_39_reset = ~ ap_rst_n;
  assign fifo_A_3_clk = ap_clk;
  assign fifo_A_3_if_din = fifo_A_3__din;
  assign fifo_A_3__dout = fifo_A_3_if_dout;
  assign fifo_A_3__empty_n = fifo_A_3_if_empty_n;
  assign fifo_A_3__full_n = fifo_A_3_if_full_n;
  assign fifo_A_3_if_read = fifo_A_3__read;
  assign fifo_A_3_if_read_ce = 1'b1;
  assign fifo_A_3_if_write = fifo_A_3__write;
  assign fifo_A_3_if_write_ce = 1'b1;
  assign fifo_A_3_reset = ~ ap_rst_n;
  assign fifo_A_40_clk = ap_clk;
  assign fifo_A_40_if_din = fifo_A_40__din;
  assign fifo_A_40__dout = fifo_A_40_if_dout;
  assign fifo_A_40__empty_n = fifo_A_40_if_empty_n;
  assign fifo_A_40__full_n = fifo_A_40_if_full_n;
  assign fifo_A_40_if_read = fifo_A_40__read;
  assign fifo_A_40_if_read_ce = 1'b1;
  assign fifo_A_40_if_write = fifo_A_40__write;
  assign fifo_A_40_if_write_ce = 1'b1;
  assign fifo_A_40_reset = ~ ap_rst_n;
  assign fifo_A_41_clk = ap_clk;
  assign fifo_A_41_if_din = fifo_A_41__din;
  assign fifo_A_41__dout = fifo_A_41_if_dout;
  assign fifo_A_41__empty_n = fifo_A_41_if_empty_n;
  assign fifo_A_41__full_n = fifo_A_41_if_full_n;
  assign fifo_A_41_if_read = fifo_A_41__read;
  assign fifo_A_41_if_read_ce = 1'b1;
  assign fifo_A_41_if_write = fifo_A_41__write;
  assign fifo_A_41_if_write_ce = 1'b1;
  assign fifo_A_41_reset = ~ ap_rst_n;
  assign fifo_A_42_clk = ap_clk;
  assign fifo_A_42_if_din = fifo_A_42__din;
  assign fifo_A_42__dout = fifo_A_42_if_dout;
  assign fifo_A_42__empty_n = fifo_A_42_if_empty_n;
  assign fifo_A_42__full_n = fifo_A_42_if_full_n;
  assign fifo_A_42_if_read = fifo_A_42__read;
  assign fifo_A_42_if_read_ce = 1'b1;
  assign fifo_A_42_if_write = fifo_A_42__write;
  assign fifo_A_42_if_write_ce = 1'b1;
  assign fifo_A_42_reset = ~ ap_rst_n;
  assign fifo_A_43_clk = ap_clk;
  assign fifo_A_43_if_din = fifo_A_43__din;
  assign fifo_A_43__dout = fifo_A_43_if_dout;
  assign fifo_A_43__empty_n = fifo_A_43_if_empty_n;
  assign fifo_A_43__full_n = fifo_A_43_if_full_n;
  assign fifo_A_43_if_read = fifo_A_43__read;
  assign fifo_A_43_if_read_ce = 1'b1;
  assign fifo_A_43_if_write = fifo_A_43__write;
  assign fifo_A_43_if_write_ce = 1'b1;
  assign fifo_A_43_reset = ~ ap_rst_n;
  assign fifo_A_44_clk = ap_clk;
  assign fifo_A_44_if_din = fifo_A_44__din;
  assign fifo_A_44__dout = fifo_A_44_if_dout;
  assign fifo_A_44__empty_n = fifo_A_44_if_empty_n;
  assign fifo_A_44__full_n = fifo_A_44_if_full_n;
  assign fifo_A_44_if_read = fifo_A_44__read;
  assign fifo_A_44_if_read_ce = 1'b1;
  assign fifo_A_44_if_write = fifo_A_44__write;
  assign fifo_A_44_if_write_ce = 1'b1;
  assign fifo_A_44_reset = ~ ap_rst_n;
  assign fifo_A_45_clk = ap_clk;
  assign fifo_A_45_if_din = fifo_A_45__din;
  assign fifo_A_45__dout = fifo_A_45_if_dout;
  assign fifo_A_45__empty_n = fifo_A_45_if_empty_n;
  assign fifo_A_45__full_n = fifo_A_45_if_full_n;
  assign fifo_A_45_if_read = fifo_A_45__read;
  assign fifo_A_45_if_read_ce = 1'b1;
  assign fifo_A_45_if_write = fifo_A_45__write;
  assign fifo_A_45_if_write_ce = 1'b1;
  assign fifo_A_45_reset = ~ ap_rst_n;
  assign fifo_A_46_clk = ap_clk;
  assign fifo_A_46_if_din = fifo_A_46__din;
  assign fifo_A_46__dout = fifo_A_46_if_dout;
  assign fifo_A_46__empty_n = fifo_A_46_if_empty_n;
  assign fifo_A_46__full_n = fifo_A_46_if_full_n;
  assign fifo_A_46_if_read = fifo_A_46__read;
  assign fifo_A_46_if_read_ce = 1'b1;
  assign fifo_A_46_if_write = fifo_A_46__write;
  assign fifo_A_46_if_write_ce = 1'b1;
  assign fifo_A_46_reset = ~ ap_rst_n;
  assign fifo_A_47_clk = ap_clk;
  assign fifo_A_47_if_din = fifo_A_47__din;
  assign fifo_A_47__dout = fifo_A_47_if_dout;
  assign fifo_A_47__empty_n = fifo_A_47_if_empty_n;
  assign fifo_A_47__full_n = fifo_A_47_if_full_n;
  assign fifo_A_47_if_read = fifo_A_47__read;
  assign fifo_A_47_if_read_ce = 1'b1;
  assign fifo_A_47_if_write = fifo_A_47__write;
  assign fifo_A_47_if_write_ce = 1'b1;
  assign fifo_A_47_reset = ~ ap_rst_n;
  assign fifo_A_4_clk = ap_clk;
  assign fifo_A_4_if_din = fifo_A_4__din;
  assign fifo_A_4__dout = fifo_A_4_if_dout;
  assign fifo_A_4__empty_n = fifo_A_4_if_empty_n;
  assign fifo_A_4__full_n = fifo_A_4_if_full_n;
  assign fifo_A_4_if_read = fifo_A_4__read;
  assign fifo_A_4_if_read_ce = 1'b1;
  assign fifo_A_4_if_write = fifo_A_4__write;
  assign fifo_A_4_if_write_ce = 1'b1;
  assign fifo_A_4_reset = ~ ap_rst_n;
  assign fifo_A_5_clk = ap_clk;
  assign fifo_A_5_if_din = fifo_A_5__din;
  assign fifo_A_5__dout = fifo_A_5_if_dout;
  assign fifo_A_5__empty_n = fifo_A_5_if_empty_n;
  assign fifo_A_5__full_n = fifo_A_5_if_full_n;
  assign fifo_A_5_if_read = fifo_A_5__read;
  assign fifo_A_5_if_read_ce = 1'b1;
  assign fifo_A_5_if_write = fifo_A_5__write;
  assign fifo_A_5_if_write_ce = 1'b1;
  assign fifo_A_5_reset = ~ ap_rst_n;
  assign fifo_A_6_clk = ap_clk;
  assign fifo_A_6_if_din = fifo_A_6__din;
  assign fifo_A_6__dout = fifo_A_6_if_dout;
  assign fifo_A_6__empty_n = fifo_A_6_if_empty_n;
  assign fifo_A_6__full_n = fifo_A_6_if_full_n;
  assign fifo_A_6_if_read = fifo_A_6__read;
  assign fifo_A_6_if_read_ce = 1'b1;
  assign fifo_A_6_if_write = fifo_A_6__write;
  assign fifo_A_6_if_write_ce = 1'b1;
  assign fifo_A_6_reset = ~ ap_rst_n;
  assign fifo_A_7_clk = ap_clk;
  assign fifo_A_7_if_din = fifo_A_7__din;
  assign fifo_A_7__dout = fifo_A_7_if_dout;
  assign fifo_A_7__empty_n = fifo_A_7_if_empty_n;
  assign fifo_A_7__full_n = fifo_A_7_if_full_n;
  assign fifo_A_7_if_read = fifo_A_7__read;
  assign fifo_A_7_if_read_ce = 1'b1;
  assign fifo_A_7_if_write = fifo_A_7__write;
  assign fifo_A_7_if_write_ce = 1'b1;
  assign fifo_A_7_reset = ~ ap_rst_n;
  assign fifo_A_8_clk = ap_clk;
  assign fifo_A_8_if_din = fifo_A_8__din;
  assign fifo_A_8__dout = fifo_A_8_if_dout;
  assign fifo_A_8__empty_n = fifo_A_8_if_empty_n;
  assign fifo_A_8__full_n = fifo_A_8_if_full_n;
  assign fifo_A_8_if_read = fifo_A_8__read;
  assign fifo_A_8_if_read_ce = 1'b1;
  assign fifo_A_8_if_write = fifo_A_8__write;
  assign fifo_A_8_if_write_ce = 1'b1;
  assign fifo_A_8_reset = ~ ap_rst_n;
  assign fifo_A_9_clk = ap_clk;
  assign fifo_A_9_if_din = fifo_A_9__din;
  assign fifo_A_9__dout = fifo_A_9_if_dout;
  assign fifo_A_9__empty_n = fifo_A_9_if_empty_n;
  assign fifo_A_9__full_n = fifo_A_9_if_full_n;
  assign fifo_A_9_if_read = fifo_A_9__read;
  assign fifo_A_9_if_read_ce = 1'b1;
  assign fifo_A_9_if_write = fifo_A_9__write;
  assign fifo_A_9_if_write_ce = 1'b1;
  assign fifo_A_9_reset = ~ ap_rst_n;
  assign fifo_X_pe_0_clk = ap_clk;
  assign fifo_X_pe_0_if_din = fifo_X_pe_0__din;
  assign fifo_X_pe_0__dout = fifo_X_pe_0_if_dout;
  assign fifo_X_pe_0__empty_n = fifo_X_pe_0_if_empty_n;
  assign fifo_X_pe_0__full_n = fifo_X_pe_0_if_full_n;
  assign fifo_X_pe_0_if_read = fifo_X_pe_0__read;
  assign fifo_X_pe_0_if_read_ce = 1'b1;
  assign fifo_X_pe_0_if_write = fifo_X_pe_0__write;
  assign fifo_X_pe_0_if_write_ce = 1'b1;
  assign fifo_X_pe_0_reset = ~ ap_rst_n;
  assign fifo_X_pe_10_clk = ap_clk;
  assign fifo_X_pe_10_if_din = fifo_X_pe_10__din;
  assign fifo_X_pe_10__dout = fifo_X_pe_10_if_dout;
  assign fifo_X_pe_10__empty_n = fifo_X_pe_10_if_empty_n;
  assign fifo_X_pe_10__full_n = fifo_X_pe_10_if_full_n;
  assign fifo_X_pe_10_if_read = fifo_X_pe_10__read;
  assign fifo_X_pe_10_if_read_ce = 1'b1;
  assign fifo_X_pe_10_if_write = fifo_X_pe_10__write;
  assign fifo_X_pe_10_if_write_ce = 1'b1;
  assign fifo_X_pe_10_reset = ~ ap_rst_n;
  assign fifo_X_pe_11_clk = ap_clk;
  assign fifo_X_pe_11_if_din = fifo_X_pe_11__din;
  assign fifo_X_pe_11__dout = fifo_X_pe_11_if_dout;
  assign fifo_X_pe_11__empty_n = fifo_X_pe_11_if_empty_n;
  assign fifo_X_pe_11__full_n = fifo_X_pe_11_if_full_n;
  assign fifo_X_pe_11_if_read = fifo_X_pe_11__read;
  assign fifo_X_pe_11_if_read_ce = 1'b1;
  assign fifo_X_pe_11_if_write = fifo_X_pe_11__write;
  assign fifo_X_pe_11_if_write_ce = 1'b1;
  assign fifo_X_pe_11_reset = ~ ap_rst_n;
  assign fifo_X_pe_12_clk = ap_clk;
  assign fifo_X_pe_12_if_din = fifo_X_pe_12__din;
  assign fifo_X_pe_12__dout = fifo_X_pe_12_if_dout;
  assign fifo_X_pe_12__empty_n = fifo_X_pe_12_if_empty_n;
  assign fifo_X_pe_12__full_n = fifo_X_pe_12_if_full_n;
  assign fifo_X_pe_12_if_read = fifo_X_pe_12__read;
  assign fifo_X_pe_12_if_read_ce = 1'b1;
  assign fifo_X_pe_12_if_write = fifo_X_pe_12__write;
  assign fifo_X_pe_12_if_write_ce = 1'b1;
  assign fifo_X_pe_12_reset = ~ ap_rst_n;
  assign fifo_X_pe_13_clk = ap_clk;
  assign fifo_X_pe_13_if_din = fifo_X_pe_13__din;
  assign fifo_X_pe_13__dout = fifo_X_pe_13_if_dout;
  assign fifo_X_pe_13__empty_n = fifo_X_pe_13_if_empty_n;
  assign fifo_X_pe_13__full_n = fifo_X_pe_13_if_full_n;
  assign fifo_X_pe_13_if_read = fifo_X_pe_13__read;
  assign fifo_X_pe_13_if_read_ce = 1'b1;
  assign fifo_X_pe_13_if_write = fifo_X_pe_13__write;
  assign fifo_X_pe_13_if_write_ce = 1'b1;
  assign fifo_X_pe_13_reset = ~ ap_rst_n;
  assign fifo_X_pe_14_clk = ap_clk;
  assign fifo_X_pe_14_if_din = fifo_X_pe_14__din;
  assign fifo_X_pe_14__dout = fifo_X_pe_14_if_dout;
  assign fifo_X_pe_14__empty_n = fifo_X_pe_14_if_empty_n;
  assign fifo_X_pe_14__full_n = fifo_X_pe_14_if_full_n;
  assign fifo_X_pe_14_if_read = fifo_X_pe_14__read;
  assign fifo_X_pe_14_if_read_ce = 1'b1;
  assign fifo_X_pe_14_if_write = fifo_X_pe_14__write;
  assign fifo_X_pe_14_if_write_ce = 1'b1;
  assign fifo_X_pe_14_reset = ~ ap_rst_n;
  assign fifo_X_pe_15_clk = ap_clk;
  assign fifo_X_pe_15_if_din = fifo_X_pe_15__din;
  assign fifo_X_pe_15__dout = fifo_X_pe_15_if_dout;
  assign fifo_X_pe_15__empty_n = fifo_X_pe_15_if_empty_n;
  assign fifo_X_pe_15__full_n = fifo_X_pe_15_if_full_n;
  assign fifo_X_pe_15_if_read = fifo_X_pe_15__read;
  assign fifo_X_pe_15_if_read_ce = 1'b1;
  assign fifo_X_pe_15_if_write = fifo_X_pe_15__write;
  assign fifo_X_pe_15_if_write_ce = 1'b1;
  assign fifo_X_pe_15_reset = ~ ap_rst_n;
  assign fifo_X_pe_16_clk = ap_clk;
  assign fifo_X_pe_16_if_din = fifo_X_pe_16__din;
  assign fifo_X_pe_16__dout = fifo_X_pe_16_if_dout;
  assign fifo_X_pe_16__empty_n = fifo_X_pe_16_if_empty_n;
  assign fifo_X_pe_16__full_n = fifo_X_pe_16_if_full_n;
  assign fifo_X_pe_16_if_read = fifo_X_pe_16__read;
  assign fifo_X_pe_16_if_read_ce = 1'b1;
  assign fifo_X_pe_16_if_write = fifo_X_pe_16__write;
  assign fifo_X_pe_16_if_write_ce = 1'b1;
  assign fifo_X_pe_16_reset = ~ ap_rst_n;
  assign fifo_X_pe_17_clk = ap_clk;
  assign fifo_X_pe_17_if_din = fifo_X_pe_17__din;
  assign fifo_X_pe_17__dout = fifo_X_pe_17_if_dout;
  assign fifo_X_pe_17__empty_n = fifo_X_pe_17_if_empty_n;
  assign fifo_X_pe_17__full_n = fifo_X_pe_17_if_full_n;
  assign fifo_X_pe_17_if_read = fifo_X_pe_17__read;
  assign fifo_X_pe_17_if_read_ce = 1'b1;
  assign fifo_X_pe_17_if_write = fifo_X_pe_17__write;
  assign fifo_X_pe_17_if_write_ce = 1'b1;
  assign fifo_X_pe_17_reset = ~ ap_rst_n;
  assign fifo_X_pe_18_clk = ap_clk;
  assign fifo_X_pe_18_if_din = fifo_X_pe_18__din;
  assign fifo_X_pe_18__dout = fifo_X_pe_18_if_dout;
  assign fifo_X_pe_18__empty_n = fifo_X_pe_18_if_empty_n;
  assign fifo_X_pe_18__full_n = fifo_X_pe_18_if_full_n;
  assign fifo_X_pe_18_if_read = fifo_X_pe_18__read;
  assign fifo_X_pe_18_if_read_ce = 1'b1;
  assign fifo_X_pe_18_if_write = fifo_X_pe_18__write;
  assign fifo_X_pe_18_if_write_ce = 1'b1;
  assign fifo_X_pe_18_reset = ~ ap_rst_n;
  assign fifo_X_pe_19_clk = ap_clk;
  assign fifo_X_pe_19_if_din = fifo_X_pe_19__din;
  assign fifo_X_pe_19__dout = fifo_X_pe_19_if_dout;
  assign fifo_X_pe_19__empty_n = fifo_X_pe_19_if_empty_n;
  assign fifo_X_pe_19__full_n = fifo_X_pe_19_if_full_n;
  assign fifo_X_pe_19_if_read = fifo_X_pe_19__read;
  assign fifo_X_pe_19_if_read_ce = 1'b1;
  assign fifo_X_pe_19_if_write = fifo_X_pe_19__write;
  assign fifo_X_pe_19_if_write_ce = 1'b1;
  assign fifo_X_pe_19_reset = ~ ap_rst_n;
  assign fifo_X_pe_1_clk = ap_clk;
  assign fifo_X_pe_1_if_din = fifo_X_pe_1__din;
  assign fifo_X_pe_1__dout = fifo_X_pe_1_if_dout;
  assign fifo_X_pe_1__empty_n = fifo_X_pe_1_if_empty_n;
  assign fifo_X_pe_1__full_n = fifo_X_pe_1_if_full_n;
  assign fifo_X_pe_1_if_read = fifo_X_pe_1__read;
  assign fifo_X_pe_1_if_read_ce = 1'b1;
  assign fifo_X_pe_1_if_write = fifo_X_pe_1__write;
  assign fifo_X_pe_1_if_write_ce = 1'b1;
  assign fifo_X_pe_1_reset = ~ ap_rst_n;
  assign fifo_X_pe_20_clk = ap_clk;
  assign fifo_X_pe_20_if_din = fifo_X_pe_20__din;
  assign fifo_X_pe_20__dout = fifo_X_pe_20_if_dout;
  assign fifo_X_pe_20__empty_n = fifo_X_pe_20_if_empty_n;
  assign fifo_X_pe_20__full_n = fifo_X_pe_20_if_full_n;
  assign fifo_X_pe_20_if_read = fifo_X_pe_20__read;
  assign fifo_X_pe_20_if_read_ce = 1'b1;
  assign fifo_X_pe_20_if_write = fifo_X_pe_20__write;
  assign fifo_X_pe_20_if_write_ce = 1'b1;
  assign fifo_X_pe_20_reset = ~ ap_rst_n;
  assign fifo_X_pe_21_clk = ap_clk;
  assign fifo_X_pe_21_if_din = fifo_X_pe_21__din;
  assign fifo_X_pe_21__dout = fifo_X_pe_21_if_dout;
  assign fifo_X_pe_21__empty_n = fifo_X_pe_21_if_empty_n;
  assign fifo_X_pe_21__full_n = fifo_X_pe_21_if_full_n;
  assign fifo_X_pe_21_if_read = fifo_X_pe_21__read;
  assign fifo_X_pe_21_if_read_ce = 1'b1;
  assign fifo_X_pe_21_if_write = fifo_X_pe_21__write;
  assign fifo_X_pe_21_if_write_ce = 1'b1;
  assign fifo_X_pe_21_reset = ~ ap_rst_n;
  assign fifo_X_pe_22_clk = ap_clk;
  assign fifo_X_pe_22_if_din = fifo_X_pe_22__din;
  assign fifo_X_pe_22__dout = fifo_X_pe_22_if_dout;
  assign fifo_X_pe_22__empty_n = fifo_X_pe_22_if_empty_n;
  assign fifo_X_pe_22__full_n = fifo_X_pe_22_if_full_n;
  assign fifo_X_pe_22_if_read = fifo_X_pe_22__read;
  assign fifo_X_pe_22_if_read_ce = 1'b1;
  assign fifo_X_pe_22_if_write = fifo_X_pe_22__write;
  assign fifo_X_pe_22_if_write_ce = 1'b1;
  assign fifo_X_pe_22_reset = ~ ap_rst_n;
  assign fifo_X_pe_23_clk = ap_clk;
  assign fifo_X_pe_23_if_din = fifo_X_pe_23__din;
  assign fifo_X_pe_23__dout = fifo_X_pe_23_if_dout;
  assign fifo_X_pe_23__empty_n = fifo_X_pe_23_if_empty_n;
  assign fifo_X_pe_23__full_n = fifo_X_pe_23_if_full_n;
  assign fifo_X_pe_23_if_read = fifo_X_pe_23__read;
  assign fifo_X_pe_23_if_read_ce = 1'b1;
  assign fifo_X_pe_23_if_write = fifo_X_pe_23__write;
  assign fifo_X_pe_23_if_write_ce = 1'b1;
  assign fifo_X_pe_23_reset = ~ ap_rst_n;
  assign fifo_X_pe_24_clk = ap_clk;
  assign fifo_X_pe_24_if_din = fifo_X_pe_24__din;
  assign fifo_X_pe_24__dout = fifo_X_pe_24_if_dout;
  assign fifo_X_pe_24__empty_n = fifo_X_pe_24_if_empty_n;
  assign fifo_X_pe_24__full_n = fifo_X_pe_24_if_full_n;
  assign fifo_X_pe_24_if_read = fifo_X_pe_24__read;
  assign fifo_X_pe_24_if_read_ce = 1'b1;
  assign fifo_X_pe_24_if_write = fifo_X_pe_24__write;
  assign fifo_X_pe_24_if_write_ce = 1'b1;
  assign fifo_X_pe_24_reset = ~ ap_rst_n;
  assign fifo_X_pe_25_clk = ap_clk;
  assign fifo_X_pe_25_if_din = fifo_X_pe_25__din;
  assign fifo_X_pe_25__dout = fifo_X_pe_25_if_dout;
  assign fifo_X_pe_25__empty_n = fifo_X_pe_25_if_empty_n;
  assign fifo_X_pe_25__full_n = fifo_X_pe_25_if_full_n;
  assign fifo_X_pe_25_if_read = fifo_X_pe_25__read;
  assign fifo_X_pe_25_if_read_ce = 1'b1;
  assign fifo_X_pe_25_if_write = fifo_X_pe_25__write;
  assign fifo_X_pe_25_if_write_ce = 1'b1;
  assign fifo_X_pe_25_reset = ~ ap_rst_n;
  assign fifo_X_pe_26_clk = ap_clk;
  assign fifo_X_pe_26_if_din = fifo_X_pe_26__din;
  assign fifo_X_pe_26__dout = fifo_X_pe_26_if_dout;
  assign fifo_X_pe_26__empty_n = fifo_X_pe_26_if_empty_n;
  assign fifo_X_pe_26__full_n = fifo_X_pe_26_if_full_n;
  assign fifo_X_pe_26_if_read = fifo_X_pe_26__read;
  assign fifo_X_pe_26_if_read_ce = 1'b1;
  assign fifo_X_pe_26_if_write = fifo_X_pe_26__write;
  assign fifo_X_pe_26_if_write_ce = 1'b1;
  assign fifo_X_pe_26_reset = ~ ap_rst_n;
  assign fifo_X_pe_27_clk = ap_clk;
  assign fifo_X_pe_27_if_din = fifo_X_pe_27__din;
  assign fifo_X_pe_27__dout = fifo_X_pe_27_if_dout;
  assign fifo_X_pe_27__empty_n = fifo_X_pe_27_if_empty_n;
  assign fifo_X_pe_27__full_n = fifo_X_pe_27_if_full_n;
  assign fifo_X_pe_27_if_read = fifo_X_pe_27__read;
  assign fifo_X_pe_27_if_read_ce = 1'b1;
  assign fifo_X_pe_27_if_write = fifo_X_pe_27__write;
  assign fifo_X_pe_27_if_write_ce = 1'b1;
  assign fifo_X_pe_27_reset = ~ ap_rst_n;
  assign fifo_X_pe_28_clk = ap_clk;
  assign fifo_X_pe_28_if_din = fifo_X_pe_28__din;
  assign fifo_X_pe_28__dout = fifo_X_pe_28_if_dout;
  assign fifo_X_pe_28__empty_n = fifo_X_pe_28_if_empty_n;
  assign fifo_X_pe_28__full_n = fifo_X_pe_28_if_full_n;
  assign fifo_X_pe_28_if_read = fifo_X_pe_28__read;
  assign fifo_X_pe_28_if_read_ce = 1'b1;
  assign fifo_X_pe_28_if_write = fifo_X_pe_28__write;
  assign fifo_X_pe_28_if_write_ce = 1'b1;
  assign fifo_X_pe_28_reset = ~ ap_rst_n;
  assign fifo_X_pe_29_clk = ap_clk;
  assign fifo_X_pe_29_if_din = fifo_X_pe_29__din;
  assign fifo_X_pe_29__dout = fifo_X_pe_29_if_dout;
  assign fifo_X_pe_29__empty_n = fifo_X_pe_29_if_empty_n;
  assign fifo_X_pe_29__full_n = fifo_X_pe_29_if_full_n;
  assign fifo_X_pe_29_if_read = fifo_X_pe_29__read;
  assign fifo_X_pe_29_if_read_ce = 1'b1;
  assign fifo_X_pe_29_if_write = fifo_X_pe_29__write;
  assign fifo_X_pe_29_if_write_ce = 1'b1;
  assign fifo_X_pe_29_reset = ~ ap_rst_n;
  assign fifo_X_pe_2_clk = ap_clk;
  assign fifo_X_pe_2_if_din = fifo_X_pe_2__din;
  assign fifo_X_pe_2__dout = fifo_X_pe_2_if_dout;
  assign fifo_X_pe_2__empty_n = fifo_X_pe_2_if_empty_n;
  assign fifo_X_pe_2__full_n = fifo_X_pe_2_if_full_n;
  assign fifo_X_pe_2_if_read = fifo_X_pe_2__read;
  assign fifo_X_pe_2_if_read_ce = 1'b1;
  assign fifo_X_pe_2_if_write = fifo_X_pe_2__write;
  assign fifo_X_pe_2_if_write_ce = 1'b1;
  assign fifo_X_pe_2_reset = ~ ap_rst_n;
  assign fifo_X_pe_30_clk = ap_clk;
  assign fifo_X_pe_30_if_din = fifo_X_pe_30__din;
  assign fifo_X_pe_30__dout = fifo_X_pe_30_if_dout;
  assign fifo_X_pe_30__empty_n = fifo_X_pe_30_if_empty_n;
  assign fifo_X_pe_30__full_n = fifo_X_pe_30_if_full_n;
  assign fifo_X_pe_30_if_read = fifo_X_pe_30__read;
  assign fifo_X_pe_30_if_read_ce = 1'b1;
  assign fifo_X_pe_30_if_write = fifo_X_pe_30__write;
  assign fifo_X_pe_30_if_write_ce = 1'b1;
  assign fifo_X_pe_30_reset = ~ ap_rst_n;
  assign fifo_X_pe_31_clk = ap_clk;
  assign fifo_X_pe_31_if_din = fifo_X_pe_31__din;
  assign fifo_X_pe_31__dout = fifo_X_pe_31_if_dout;
  assign fifo_X_pe_31__empty_n = fifo_X_pe_31_if_empty_n;
  assign fifo_X_pe_31__full_n = fifo_X_pe_31_if_full_n;
  assign fifo_X_pe_31_if_read = fifo_X_pe_31__read;
  assign fifo_X_pe_31_if_read_ce = 1'b1;
  assign fifo_X_pe_31_if_write = fifo_X_pe_31__write;
  assign fifo_X_pe_31_if_write_ce = 1'b1;
  assign fifo_X_pe_31_reset = ~ ap_rst_n;
  assign fifo_X_pe_32_clk = ap_clk;
  assign fifo_X_pe_32_if_din = fifo_X_pe_32__din;
  assign fifo_X_pe_32__dout = fifo_X_pe_32_if_dout;
  assign fifo_X_pe_32__empty_n = fifo_X_pe_32_if_empty_n;
  assign fifo_X_pe_32__full_n = fifo_X_pe_32_if_full_n;
  assign fifo_X_pe_32_if_read = fifo_X_pe_32__read;
  assign fifo_X_pe_32_if_read_ce = 1'b1;
  assign fifo_X_pe_32_if_write = fifo_X_pe_32__write;
  assign fifo_X_pe_32_if_write_ce = 1'b1;
  assign fifo_X_pe_32_reset = ~ ap_rst_n;
  assign fifo_X_pe_33_clk = ap_clk;
  assign fifo_X_pe_33_if_din = fifo_X_pe_33__din;
  assign fifo_X_pe_33__dout = fifo_X_pe_33_if_dout;
  assign fifo_X_pe_33__empty_n = fifo_X_pe_33_if_empty_n;
  assign fifo_X_pe_33__full_n = fifo_X_pe_33_if_full_n;
  assign fifo_X_pe_33_if_read = fifo_X_pe_33__read;
  assign fifo_X_pe_33_if_read_ce = 1'b1;
  assign fifo_X_pe_33_if_write = fifo_X_pe_33__write;
  assign fifo_X_pe_33_if_write_ce = 1'b1;
  assign fifo_X_pe_33_reset = ~ ap_rst_n;
  assign fifo_X_pe_34_clk = ap_clk;
  assign fifo_X_pe_34_if_din = fifo_X_pe_34__din;
  assign fifo_X_pe_34__dout = fifo_X_pe_34_if_dout;
  assign fifo_X_pe_34__empty_n = fifo_X_pe_34_if_empty_n;
  assign fifo_X_pe_34__full_n = fifo_X_pe_34_if_full_n;
  assign fifo_X_pe_34_if_read = fifo_X_pe_34__read;
  assign fifo_X_pe_34_if_read_ce = 1'b1;
  assign fifo_X_pe_34_if_write = fifo_X_pe_34__write;
  assign fifo_X_pe_34_if_write_ce = 1'b1;
  assign fifo_X_pe_34_reset = ~ ap_rst_n;
  assign fifo_X_pe_35_clk = ap_clk;
  assign fifo_X_pe_35_if_din = fifo_X_pe_35__din;
  assign fifo_X_pe_35__dout = fifo_X_pe_35_if_dout;
  assign fifo_X_pe_35__empty_n = fifo_X_pe_35_if_empty_n;
  assign fifo_X_pe_35__full_n = fifo_X_pe_35_if_full_n;
  assign fifo_X_pe_35_if_read = fifo_X_pe_35__read;
  assign fifo_X_pe_35_if_read_ce = 1'b1;
  assign fifo_X_pe_35_if_write = fifo_X_pe_35__write;
  assign fifo_X_pe_35_if_write_ce = 1'b1;
  assign fifo_X_pe_35_reset = ~ ap_rst_n;
  assign fifo_X_pe_36_clk = ap_clk;
  assign fifo_X_pe_36_if_din = fifo_X_pe_36__din;
  assign fifo_X_pe_36__dout = fifo_X_pe_36_if_dout;
  assign fifo_X_pe_36__empty_n = fifo_X_pe_36_if_empty_n;
  assign fifo_X_pe_36__full_n = fifo_X_pe_36_if_full_n;
  assign fifo_X_pe_36_if_read = fifo_X_pe_36__read;
  assign fifo_X_pe_36_if_read_ce = 1'b1;
  assign fifo_X_pe_36_if_write = fifo_X_pe_36__write;
  assign fifo_X_pe_36_if_write_ce = 1'b1;
  assign fifo_X_pe_36_reset = ~ ap_rst_n;
  assign fifo_X_pe_37_clk = ap_clk;
  assign fifo_X_pe_37_if_din = fifo_X_pe_37__din;
  assign fifo_X_pe_37__dout = fifo_X_pe_37_if_dout;
  assign fifo_X_pe_37__empty_n = fifo_X_pe_37_if_empty_n;
  assign fifo_X_pe_37__full_n = fifo_X_pe_37_if_full_n;
  assign fifo_X_pe_37_if_read = fifo_X_pe_37__read;
  assign fifo_X_pe_37_if_read_ce = 1'b1;
  assign fifo_X_pe_37_if_write = fifo_X_pe_37__write;
  assign fifo_X_pe_37_if_write_ce = 1'b1;
  assign fifo_X_pe_37_reset = ~ ap_rst_n;
  assign fifo_X_pe_38_clk = ap_clk;
  assign fifo_X_pe_38_if_din = fifo_X_pe_38__din;
  assign fifo_X_pe_38__dout = fifo_X_pe_38_if_dout;
  assign fifo_X_pe_38__empty_n = fifo_X_pe_38_if_empty_n;
  assign fifo_X_pe_38__full_n = fifo_X_pe_38_if_full_n;
  assign fifo_X_pe_38_if_read = fifo_X_pe_38__read;
  assign fifo_X_pe_38_if_read_ce = 1'b1;
  assign fifo_X_pe_38_if_write = fifo_X_pe_38__write;
  assign fifo_X_pe_38_if_write_ce = 1'b1;
  assign fifo_X_pe_38_reset = ~ ap_rst_n;
  assign fifo_X_pe_39_clk = ap_clk;
  assign fifo_X_pe_39_if_din = fifo_X_pe_39__din;
  assign fifo_X_pe_39__dout = fifo_X_pe_39_if_dout;
  assign fifo_X_pe_39__empty_n = fifo_X_pe_39_if_empty_n;
  assign fifo_X_pe_39__full_n = fifo_X_pe_39_if_full_n;
  assign fifo_X_pe_39_if_read = fifo_X_pe_39__read;
  assign fifo_X_pe_39_if_read_ce = 1'b1;
  assign fifo_X_pe_39_if_write = fifo_X_pe_39__write;
  assign fifo_X_pe_39_if_write_ce = 1'b1;
  assign fifo_X_pe_39_reset = ~ ap_rst_n;
  assign fifo_X_pe_3_clk = ap_clk;
  assign fifo_X_pe_3_if_din = fifo_X_pe_3__din;
  assign fifo_X_pe_3__dout = fifo_X_pe_3_if_dout;
  assign fifo_X_pe_3__empty_n = fifo_X_pe_3_if_empty_n;
  assign fifo_X_pe_3__full_n = fifo_X_pe_3_if_full_n;
  assign fifo_X_pe_3_if_read = fifo_X_pe_3__read;
  assign fifo_X_pe_3_if_read_ce = 1'b1;
  assign fifo_X_pe_3_if_write = fifo_X_pe_3__write;
  assign fifo_X_pe_3_if_write_ce = 1'b1;
  assign fifo_X_pe_3_reset = ~ ap_rst_n;
  assign fifo_X_pe_40_clk = ap_clk;
  assign fifo_X_pe_40_if_din = fifo_X_pe_40__din;
  assign fifo_X_pe_40__dout = fifo_X_pe_40_if_dout;
  assign fifo_X_pe_40__empty_n = fifo_X_pe_40_if_empty_n;
  assign fifo_X_pe_40__full_n = fifo_X_pe_40_if_full_n;
  assign fifo_X_pe_40_if_read = fifo_X_pe_40__read;
  assign fifo_X_pe_40_if_read_ce = 1'b1;
  assign fifo_X_pe_40_if_write = fifo_X_pe_40__write;
  assign fifo_X_pe_40_if_write_ce = 1'b1;
  assign fifo_X_pe_40_reset = ~ ap_rst_n;
  assign fifo_X_pe_41_clk = ap_clk;
  assign fifo_X_pe_41_if_din = fifo_X_pe_41__din;
  assign fifo_X_pe_41__dout = fifo_X_pe_41_if_dout;
  assign fifo_X_pe_41__empty_n = fifo_X_pe_41_if_empty_n;
  assign fifo_X_pe_41__full_n = fifo_X_pe_41_if_full_n;
  assign fifo_X_pe_41_if_read = fifo_X_pe_41__read;
  assign fifo_X_pe_41_if_read_ce = 1'b1;
  assign fifo_X_pe_41_if_write = fifo_X_pe_41__write;
  assign fifo_X_pe_41_if_write_ce = 1'b1;
  assign fifo_X_pe_41_reset = ~ ap_rst_n;
  assign fifo_X_pe_42_clk = ap_clk;
  assign fifo_X_pe_42_if_din = fifo_X_pe_42__din;
  assign fifo_X_pe_42__dout = fifo_X_pe_42_if_dout;
  assign fifo_X_pe_42__empty_n = fifo_X_pe_42_if_empty_n;
  assign fifo_X_pe_42__full_n = fifo_X_pe_42_if_full_n;
  assign fifo_X_pe_42_if_read = fifo_X_pe_42__read;
  assign fifo_X_pe_42_if_read_ce = 1'b1;
  assign fifo_X_pe_42_if_write = fifo_X_pe_42__write;
  assign fifo_X_pe_42_if_write_ce = 1'b1;
  assign fifo_X_pe_42_reset = ~ ap_rst_n;
  assign fifo_X_pe_43_clk = ap_clk;
  assign fifo_X_pe_43_if_din = fifo_X_pe_43__din;
  assign fifo_X_pe_43__dout = fifo_X_pe_43_if_dout;
  assign fifo_X_pe_43__empty_n = fifo_X_pe_43_if_empty_n;
  assign fifo_X_pe_43__full_n = fifo_X_pe_43_if_full_n;
  assign fifo_X_pe_43_if_read = fifo_X_pe_43__read;
  assign fifo_X_pe_43_if_read_ce = 1'b1;
  assign fifo_X_pe_43_if_write = fifo_X_pe_43__write;
  assign fifo_X_pe_43_if_write_ce = 1'b1;
  assign fifo_X_pe_43_reset = ~ ap_rst_n;
  assign fifo_X_pe_44_clk = ap_clk;
  assign fifo_X_pe_44_if_din = fifo_X_pe_44__din;
  assign fifo_X_pe_44__dout = fifo_X_pe_44_if_dout;
  assign fifo_X_pe_44__empty_n = fifo_X_pe_44_if_empty_n;
  assign fifo_X_pe_44__full_n = fifo_X_pe_44_if_full_n;
  assign fifo_X_pe_44_if_read = fifo_X_pe_44__read;
  assign fifo_X_pe_44_if_read_ce = 1'b1;
  assign fifo_X_pe_44_if_write = fifo_X_pe_44__write;
  assign fifo_X_pe_44_if_write_ce = 1'b1;
  assign fifo_X_pe_44_reset = ~ ap_rst_n;
  assign fifo_X_pe_45_clk = ap_clk;
  assign fifo_X_pe_45_if_din = fifo_X_pe_45__din;
  assign fifo_X_pe_45__dout = fifo_X_pe_45_if_dout;
  assign fifo_X_pe_45__empty_n = fifo_X_pe_45_if_empty_n;
  assign fifo_X_pe_45__full_n = fifo_X_pe_45_if_full_n;
  assign fifo_X_pe_45_if_read = fifo_X_pe_45__read;
  assign fifo_X_pe_45_if_read_ce = 1'b1;
  assign fifo_X_pe_45_if_write = fifo_X_pe_45__write;
  assign fifo_X_pe_45_if_write_ce = 1'b1;
  assign fifo_X_pe_45_reset = ~ ap_rst_n;
  assign fifo_X_pe_46_clk = ap_clk;
  assign fifo_X_pe_46_if_din = fifo_X_pe_46__din;
  assign fifo_X_pe_46__dout = fifo_X_pe_46_if_dout;
  assign fifo_X_pe_46__empty_n = fifo_X_pe_46_if_empty_n;
  assign fifo_X_pe_46__full_n = fifo_X_pe_46_if_full_n;
  assign fifo_X_pe_46_if_read = fifo_X_pe_46__read;
  assign fifo_X_pe_46_if_read_ce = 1'b1;
  assign fifo_X_pe_46_if_write = fifo_X_pe_46__write;
  assign fifo_X_pe_46_if_write_ce = 1'b1;
  assign fifo_X_pe_46_reset = ~ ap_rst_n;
  assign fifo_X_pe_47_clk = ap_clk;
  assign fifo_X_pe_47_if_din = fifo_X_pe_47__din;
  assign fifo_X_pe_47__dout = fifo_X_pe_47_if_dout;
  assign fifo_X_pe_47__empty_n = fifo_X_pe_47_if_empty_n;
  assign fifo_X_pe_47__full_n = fifo_X_pe_47_if_full_n;
  assign fifo_X_pe_47_if_read = fifo_X_pe_47__read;
  assign fifo_X_pe_47_if_read_ce = 1'b1;
  assign fifo_X_pe_47_if_write = fifo_X_pe_47__write;
  assign fifo_X_pe_47_if_write_ce = 1'b1;
  assign fifo_X_pe_47_reset = ~ ap_rst_n;
  assign fifo_X_pe_48_clk = ap_clk;
  assign fifo_X_pe_48_if_din = fifo_X_pe_48__din;
  assign fifo_X_pe_48__dout = fifo_X_pe_48_if_dout;
  assign fifo_X_pe_48__empty_n = fifo_X_pe_48_if_empty_n;
  assign fifo_X_pe_48__full_n = fifo_X_pe_48_if_full_n;
  assign fifo_X_pe_48_if_read = fifo_X_pe_48__read;
  assign fifo_X_pe_48_if_read_ce = 1'b1;
  assign fifo_X_pe_48_if_write = fifo_X_pe_48__write;
  assign fifo_X_pe_48_if_write_ce = 1'b1;
  assign fifo_X_pe_48_reset = ~ ap_rst_n;
  assign fifo_X_pe_4_clk = ap_clk;
  assign fifo_X_pe_4_if_din = fifo_X_pe_4__din;
  assign fifo_X_pe_4__dout = fifo_X_pe_4_if_dout;
  assign fifo_X_pe_4__empty_n = fifo_X_pe_4_if_empty_n;
  assign fifo_X_pe_4__full_n = fifo_X_pe_4_if_full_n;
  assign fifo_X_pe_4_if_read = fifo_X_pe_4__read;
  assign fifo_X_pe_4_if_read_ce = 1'b1;
  assign fifo_X_pe_4_if_write = fifo_X_pe_4__write;
  assign fifo_X_pe_4_if_write_ce = 1'b1;
  assign fifo_X_pe_4_reset = ~ ap_rst_n;
  assign fifo_X_pe_5_clk = ap_clk;
  assign fifo_X_pe_5_if_din = fifo_X_pe_5__din;
  assign fifo_X_pe_5__dout = fifo_X_pe_5_if_dout;
  assign fifo_X_pe_5__empty_n = fifo_X_pe_5_if_empty_n;
  assign fifo_X_pe_5__full_n = fifo_X_pe_5_if_full_n;
  assign fifo_X_pe_5_if_read = fifo_X_pe_5__read;
  assign fifo_X_pe_5_if_read_ce = 1'b1;
  assign fifo_X_pe_5_if_write = fifo_X_pe_5__write;
  assign fifo_X_pe_5_if_write_ce = 1'b1;
  assign fifo_X_pe_5_reset = ~ ap_rst_n;
  assign fifo_X_pe_6_clk = ap_clk;
  assign fifo_X_pe_6_if_din = fifo_X_pe_6__din;
  assign fifo_X_pe_6__dout = fifo_X_pe_6_if_dout;
  assign fifo_X_pe_6__empty_n = fifo_X_pe_6_if_empty_n;
  assign fifo_X_pe_6__full_n = fifo_X_pe_6_if_full_n;
  assign fifo_X_pe_6_if_read = fifo_X_pe_6__read;
  assign fifo_X_pe_6_if_read_ce = 1'b1;
  assign fifo_X_pe_6_if_write = fifo_X_pe_6__write;
  assign fifo_X_pe_6_if_write_ce = 1'b1;
  assign fifo_X_pe_6_reset = ~ ap_rst_n;
  assign fifo_X_pe_7_clk = ap_clk;
  assign fifo_X_pe_7_if_din = fifo_X_pe_7__din;
  assign fifo_X_pe_7__dout = fifo_X_pe_7_if_dout;
  assign fifo_X_pe_7__empty_n = fifo_X_pe_7_if_empty_n;
  assign fifo_X_pe_7__full_n = fifo_X_pe_7_if_full_n;
  assign fifo_X_pe_7_if_read = fifo_X_pe_7__read;
  assign fifo_X_pe_7_if_read_ce = 1'b1;
  assign fifo_X_pe_7_if_write = fifo_X_pe_7__write;
  assign fifo_X_pe_7_if_write_ce = 1'b1;
  assign fifo_X_pe_7_reset = ~ ap_rst_n;
  assign fifo_X_pe_8_clk = ap_clk;
  assign fifo_X_pe_8_if_din = fifo_X_pe_8__din;
  assign fifo_X_pe_8__dout = fifo_X_pe_8_if_dout;
  assign fifo_X_pe_8__empty_n = fifo_X_pe_8_if_empty_n;
  assign fifo_X_pe_8__full_n = fifo_X_pe_8_if_full_n;
  assign fifo_X_pe_8_if_read = fifo_X_pe_8__read;
  assign fifo_X_pe_8_if_read_ce = 1'b1;
  assign fifo_X_pe_8_if_write = fifo_X_pe_8__write;
  assign fifo_X_pe_8_if_write_ce = 1'b1;
  assign fifo_X_pe_8_reset = ~ ap_rst_n;
  assign fifo_X_pe_9_clk = ap_clk;
  assign fifo_X_pe_9_if_din = fifo_X_pe_9__din;
  assign fifo_X_pe_9__dout = fifo_X_pe_9_if_dout;
  assign fifo_X_pe_9__empty_n = fifo_X_pe_9_if_empty_n;
  assign fifo_X_pe_9__full_n = fifo_X_pe_9_if_full_n;
  assign fifo_X_pe_9_if_read = fifo_X_pe_9__read;
  assign fifo_X_pe_9_if_read_ce = 1'b1;
  assign fifo_X_pe_9_if_write = fifo_X_pe_9__write;
  assign fifo_X_pe_9_if_write_ce = 1'b1;
  assign fifo_X_pe_9_reset = ~ ap_rst_n;
  assign fifo_Y_AX_clk = ap_clk;
  assign fifo_Y_AX_if_din = fifo_Y_AX__din;
  assign fifo_Y_AX__dout = fifo_Y_AX_if_dout;
  assign fifo_Y_AX__empty_n = fifo_Y_AX_if_empty_n;
  assign fifo_Y_AX__full_n = fifo_Y_AX_if_full_n;
  assign fifo_Y_AX_if_read = fifo_Y_AX__read;
  assign fifo_Y_AX_if_read_ce = 1'b1;
  assign fifo_Y_AX_if_write = fifo_Y_AX__write;
  assign fifo_Y_AX_if_write_ce = 1'b1;
  assign fifo_Y_AX_reset = ~ ap_rst_n;
  assign fifo_Y_alpha_AX_clk = ap_clk;
  assign fifo_Y_alpha_AX_if_din = fifo_Y_alpha_AX__din;
  assign fifo_Y_alpha_AX__dout = fifo_Y_alpha_AX_if_dout;
  assign fifo_Y_alpha_AX__empty_n = fifo_Y_alpha_AX_if_empty_n;
  assign fifo_Y_alpha_AX__full_n = fifo_Y_alpha_AX_if_full_n;
  assign fifo_Y_alpha_AX_if_read = fifo_Y_alpha_AX__read;
  assign fifo_Y_alpha_AX_if_read_ce = 1'b1;
  assign fifo_Y_alpha_AX_if_write = fifo_Y_alpha_AX__write;
  assign fifo_Y_alpha_AX_if_write_ce = 1'b1;
  assign fifo_Y_alpha_AX_reset = ~ ap_rst_n;
  assign fifo_Y_in_clk = ap_clk;
  assign fifo_Y_in_if_din = fifo_Y_in__din;
  assign fifo_Y_in__dout = fifo_Y_in_if_dout;
  assign fifo_Y_in__empty_n = fifo_Y_in_if_empty_n;
  assign fifo_Y_in__full_n = fifo_Y_in_if_full_n;
  assign fifo_Y_in_if_read = fifo_Y_in__read;
  assign fifo_Y_in_if_read_ce = 1'b1;
  assign fifo_Y_in_if_write = fifo_Y_in__write;
  assign fifo_Y_in_if_write_ce = 1'b1;
  assign fifo_Y_in_reset = ~ ap_rst_n;
  assign fifo_Y_in_beta_clk = ap_clk;
  assign fifo_Y_in_beta_if_din = fifo_Y_in_beta__din;
  assign fifo_Y_in_beta__dout = fifo_Y_in_beta_if_dout;
  assign fifo_Y_in_beta__empty_n = fifo_Y_in_beta_if_empty_n;
  assign fifo_Y_in_beta__full_n = fifo_Y_in_beta_if_full_n;
  assign fifo_Y_in_beta_if_read = fifo_Y_in_beta__read;
  assign fifo_Y_in_beta_if_read_ce = 1'b1;
  assign fifo_Y_in_beta_if_write = fifo_Y_in_beta__write;
  assign fifo_Y_in_beta_if_write_ce = 1'b1;
  assign fifo_Y_in_beta_reset = ~ ap_rst_n;
  assign fifo_Y_out_clk = ap_clk;
  assign fifo_Y_out_if_din = fifo_Y_out__din;
  assign fifo_Y_out__dout = fifo_Y_out_if_dout;
  assign fifo_Y_out__empty_n = fifo_Y_out_if_empty_n;
  assign fifo_Y_out__full_n = fifo_Y_out_if_full_n;
  assign fifo_Y_out_if_read = fifo_Y_out__read;
  assign fifo_Y_out_if_read_ce = 1'b1;
  assign fifo_Y_out_if_write = fifo_Y_out__write;
  assign fifo_Y_out_if_write_ce = 1'b1;
  assign fifo_Y_out_reset = ~ ap_rst_n;
  assign fifo_Y_pe_0_clk = ap_clk;
  assign fifo_Y_pe_0_if_din = fifo_Y_pe_0__din;
  assign fifo_Y_pe_0__dout = fifo_Y_pe_0_if_dout;
  assign fifo_Y_pe_0__empty_n = fifo_Y_pe_0_if_empty_n;
  assign fifo_Y_pe_0__full_n = fifo_Y_pe_0_if_full_n;
  assign fifo_Y_pe_0_if_read = fifo_Y_pe_0__read;
  assign fifo_Y_pe_0_if_read_ce = 1'b1;
  assign fifo_Y_pe_0_if_write = fifo_Y_pe_0__write;
  assign fifo_Y_pe_0_if_write_ce = 1'b1;
  assign fifo_Y_pe_0_reset = ~ ap_rst_n;
  assign fifo_Y_pe_10_clk = ap_clk;
  assign fifo_Y_pe_10_if_din = fifo_Y_pe_10__din;
  assign fifo_Y_pe_10__dout = fifo_Y_pe_10_if_dout;
  assign fifo_Y_pe_10__empty_n = fifo_Y_pe_10_if_empty_n;
  assign fifo_Y_pe_10__full_n = fifo_Y_pe_10_if_full_n;
  assign fifo_Y_pe_10_if_read = fifo_Y_pe_10__read;
  assign fifo_Y_pe_10_if_read_ce = 1'b1;
  assign fifo_Y_pe_10_if_write = fifo_Y_pe_10__write;
  assign fifo_Y_pe_10_if_write_ce = 1'b1;
  assign fifo_Y_pe_10_reset = ~ ap_rst_n;
  assign fifo_Y_pe_11_clk = ap_clk;
  assign fifo_Y_pe_11_if_din = fifo_Y_pe_11__din;
  assign fifo_Y_pe_11__dout = fifo_Y_pe_11_if_dout;
  assign fifo_Y_pe_11__empty_n = fifo_Y_pe_11_if_empty_n;
  assign fifo_Y_pe_11__full_n = fifo_Y_pe_11_if_full_n;
  assign fifo_Y_pe_11_if_read = fifo_Y_pe_11__read;
  assign fifo_Y_pe_11_if_read_ce = 1'b1;
  assign fifo_Y_pe_11_if_write = fifo_Y_pe_11__write;
  assign fifo_Y_pe_11_if_write_ce = 1'b1;
  assign fifo_Y_pe_11_reset = ~ ap_rst_n;
  assign fifo_Y_pe_12_clk = ap_clk;
  assign fifo_Y_pe_12_if_din = fifo_Y_pe_12__din;
  assign fifo_Y_pe_12__dout = fifo_Y_pe_12_if_dout;
  assign fifo_Y_pe_12__empty_n = fifo_Y_pe_12_if_empty_n;
  assign fifo_Y_pe_12__full_n = fifo_Y_pe_12_if_full_n;
  assign fifo_Y_pe_12_if_read = fifo_Y_pe_12__read;
  assign fifo_Y_pe_12_if_read_ce = 1'b1;
  assign fifo_Y_pe_12_if_write = fifo_Y_pe_12__write;
  assign fifo_Y_pe_12_if_write_ce = 1'b1;
  assign fifo_Y_pe_12_reset = ~ ap_rst_n;
  assign fifo_Y_pe_13_clk = ap_clk;
  assign fifo_Y_pe_13_if_din = fifo_Y_pe_13__din;
  assign fifo_Y_pe_13__dout = fifo_Y_pe_13_if_dout;
  assign fifo_Y_pe_13__empty_n = fifo_Y_pe_13_if_empty_n;
  assign fifo_Y_pe_13__full_n = fifo_Y_pe_13_if_full_n;
  assign fifo_Y_pe_13_if_read = fifo_Y_pe_13__read;
  assign fifo_Y_pe_13_if_read_ce = 1'b1;
  assign fifo_Y_pe_13_if_write = fifo_Y_pe_13__write;
  assign fifo_Y_pe_13_if_write_ce = 1'b1;
  assign fifo_Y_pe_13_reset = ~ ap_rst_n;
  assign fifo_Y_pe_14_clk = ap_clk;
  assign fifo_Y_pe_14_if_din = fifo_Y_pe_14__din;
  assign fifo_Y_pe_14__dout = fifo_Y_pe_14_if_dout;
  assign fifo_Y_pe_14__empty_n = fifo_Y_pe_14_if_empty_n;
  assign fifo_Y_pe_14__full_n = fifo_Y_pe_14_if_full_n;
  assign fifo_Y_pe_14_if_read = fifo_Y_pe_14__read;
  assign fifo_Y_pe_14_if_read_ce = 1'b1;
  assign fifo_Y_pe_14_if_write = fifo_Y_pe_14__write;
  assign fifo_Y_pe_14_if_write_ce = 1'b1;
  assign fifo_Y_pe_14_reset = ~ ap_rst_n;
  assign fifo_Y_pe_15_clk = ap_clk;
  assign fifo_Y_pe_15_if_din = fifo_Y_pe_15__din;
  assign fifo_Y_pe_15__dout = fifo_Y_pe_15_if_dout;
  assign fifo_Y_pe_15__empty_n = fifo_Y_pe_15_if_empty_n;
  assign fifo_Y_pe_15__full_n = fifo_Y_pe_15_if_full_n;
  assign fifo_Y_pe_15_if_read = fifo_Y_pe_15__read;
  assign fifo_Y_pe_15_if_read_ce = 1'b1;
  assign fifo_Y_pe_15_if_write = fifo_Y_pe_15__write;
  assign fifo_Y_pe_15_if_write_ce = 1'b1;
  assign fifo_Y_pe_15_reset = ~ ap_rst_n;
  assign fifo_Y_pe_16_clk = ap_clk;
  assign fifo_Y_pe_16_if_din = fifo_Y_pe_16__din;
  assign fifo_Y_pe_16__dout = fifo_Y_pe_16_if_dout;
  assign fifo_Y_pe_16__empty_n = fifo_Y_pe_16_if_empty_n;
  assign fifo_Y_pe_16__full_n = fifo_Y_pe_16_if_full_n;
  assign fifo_Y_pe_16_if_read = fifo_Y_pe_16__read;
  assign fifo_Y_pe_16_if_read_ce = 1'b1;
  assign fifo_Y_pe_16_if_write = fifo_Y_pe_16__write;
  assign fifo_Y_pe_16_if_write_ce = 1'b1;
  assign fifo_Y_pe_16_reset = ~ ap_rst_n;
  assign fifo_Y_pe_17_clk = ap_clk;
  assign fifo_Y_pe_17_if_din = fifo_Y_pe_17__din;
  assign fifo_Y_pe_17__dout = fifo_Y_pe_17_if_dout;
  assign fifo_Y_pe_17__empty_n = fifo_Y_pe_17_if_empty_n;
  assign fifo_Y_pe_17__full_n = fifo_Y_pe_17_if_full_n;
  assign fifo_Y_pe_17_if_read = fifo_Y_pe_17__read;
  assign fifo_Y_pe_17_if_read_ce = 1'b1;
  assign fifo_Y_pe_17_if_write = fifo_Y_pe_17__write;
  assign fifo_Y_pe_17_if_write_ce = 1'b1;
  assign fifo_Y_pe_17_reset = ~ ap_rst_n;
  assign fifo_Y_pe_18_clk = ap_clk;
  assign fifo_Y_pe_18_if_din = fifo_Y_pe_18__din;
  assign fifo_Y_pe_18__dout = fifo_Y_pe_18_if_dout;
  assign fifo_Y_pe_18__empty_n = fifo_Y_pe_18_if_empty_n;
  assign fifo_Y_pe_18__full_n = fifo_Y_pe_18_if_full_n;
  assign fifo_Y_pe_18_if_read = fifo_Y_pe_18__read;
  assign fifo_Y_pe_18_if_read_ce = 1'b1;
  assign fifo_Y_pe_18_if_write = fifo_Y_pe_18__write;
  assign fifo_Y_pe_18_if_write_ce = 1'b1;
  assign fifo_Y_pe_18_reset = ~ ap_rst_n;
  assign fifo_Y_pe_19_clk = ap_clk;
  assign fifo_Y_pe_19_if_din = fifo_Y_pe_19__din;
  assign fifo_Y_pe_19__dout = fifo_Y_pe_19_if_dout;
  assign fifo_Y_pe_19__empty_n = fifo_Y_pe_19_if_empty_n;
  assign fifo_Y_pe_19__full_n = fifo_Y_pe_19_if_full_n;
  assign fifo_Y_pe_19_if_read = fifo_Y_pe_19__read;
  assign fifo_Y_pe_19_if_read_ce = 1'b1;
  assign fifo_Y_pe_19_if_write = fifo_Y_pe_19__write;
  assign fifo_Y_pe_19_if_write_ce = 1'b1;
  assign fifo_Y_pe_19_reset = ~ ap_rst_n;
  assign fifo_Y_pe_1_clk = ap_clk;
  assign fifo_Y_pe_1_if_din = fifo_Y_pe_1__din;
  assign fifo_Y_pe_1__dout = fifo_Y_pe_1_if_dout;
  assign fifo_Y_pe_1__empty_n = fifo_Y_pe_1_if_empty_n;
  assign fifo_Y_pe_1__full_n = fifo_Y_pe_1_if_full_n;
  assign fifo_Y_pe_1_if_read = fifo_Y_pe_1__read;
  assign fifo_Y_pe_1_if_read_ce = 1'b1;
  assign fifo_Y_pe_1_if_write = fifo_Y_pe_1__write;
  assign fifo_Y_pe_1_if_write_ce = 1'b1;
  assign fifo_Y_pe_1_reset = ~ ap_rst_n;
  assign fifo_Y_pe_20_clk = ap_clk;
  assign fifo_Y_pe_20_if_din = fifo_Y_pe_20__din;
  assign fifo_Y_pe_20__dout = fifo_Y_pe_20_if_dout;
  assign fifo_Y_pe_20__empty_n = fifo_Y_pe_20_if_empty_n;
  assign fifo_Y_pe_20__full_n = fifo_Y_pe_20_if_full_n;
  assign fifo_Y_pe_20_if_read = fifo_Y_pe_20__read;
  assign fifo_Y_pe_20_if_read_ce = 1'b1;
  assign fifo_Y_pe_20_if_write = fifo_Y_pe_20__write;
  assign fifo_Y_pe_20_if_write_ce = 1'b1;
  assign fifo_Y_pe_20_reset = ~ ap_rst_n;
  assign fifo_Y_pe_21_clk = ap_clk;
  assign fifo_Y_pe_21_if_din = fifo_Y_pe_21__din;
  assign fifo_Y_pe_21__dout = fifo_Y_pe_21_if_dout;
  assign fifo_Y_pe_21__empty_n = fifo_Y_pe_21_if_empty_n;
  assign fifo_Y_pe_21__full_n = fifo_Y_pe_21_if_full_n;
  assign fifo_Y_pe_21_if_read = fifo_Y_pe_21__read;
  assign fifo_Y_pe_21_if_read_ce = 1'b1;
  assign fifo_Y_pe_21_if_write = fifo_Y_pe_21__write;
  assign fifo_Y_pe_21_if_write_ce = 1'b1;
  assign fifo_Y_pe_21_reset = ~ ap_rst_n;
  assign fifo_Y_pe_22_clk = ap_clk;
  assign fifo_Y_pe_22_if_din = fifo_Y_pe_22__din;
  assign fifo_Y_pe_22__dout = fifo_Y_pe_22_if_dout;
  assign fifo_Y_pe_22__empty_n = fifo_Y_pe_22_if_empty_n;
  assign fifo_Y_pe_22__full_n = fifo_Y_pe_22_if_full_n;
  assign fifo_Y_pe_22_if_read = fifo_Y_pe_22__read;
  assign fifo_Y_pe_22_if_read_ce = 1'b1;
  assign fifo_Y_pe_22_if_write = fifo_Y_pe_22__write;
  assign fifo_Y_pe_22_if_write_ce = 1'b1;
  assign fifo_Y_pe_22_reset = ~ ap_rst_n;
  assign fifo_Y_pe_23_clk = ap_clk;
  assign fifo_Y_pe_23_if_din = fifo_Y_pe_23__din;
  assign fifo_Y_pe_23__dout = fifo_Y_pe_23_if_dout;
  assign fifo_Y_pe_23__empty_n = fifo_Y_pe_23_if_empty_n;
  assign fifo_Y_pe_23__full_n = fifo_Y_pe_23_if_full_n;
  assign fifo_Y_pe_23_if_read = fifo_Y_pe_23__read;
  assign fifo_Y_pe_23_if_read_ce = 1'b1;
  assign fifo_Y_pe_23_if_write = fifo_Y_pe_23__write;
  assign fifo_Y_pe_23_if_write_ce = 1'b1;
  assign fifo_Y_pe_23_reset = ~ ap_rst_n;
  assign fifo_Y_pe_24_clk = ap_clk;
  assign fifo_Y_pe_24_if_din = fifo_Y_pe_24__din;
  assign fifo_Y_pe_24__dout = fifo_Y_pe_24_if_dout;
  assign fifo_Y_pe_24__empty_n = fifo_Y_pe_24_if_empty_n;
  assign fifo_Y_pe_24__full_n = fifo_Y_pe_24_if_full_n;
  assign fifo_Y_pe_24_if_read = fifo_Y_pe_24__read;
  assign fifo_Y_pe_24_if_read_ce = 1'b1;
  assign fifo_Y_pe_24_if_write = fifo_Y_pe_24__write;
  assign fifo_Y_pe_24_if_write_ce = 1'b1;
  assign fifo_Y_pe_24_reset = ~ ap_rst_n;
  assign fifo_Y_pe_25_clk = ap_clk;
  assign fifo_Y_pe_25_if_din = fifo_Y_pe_25__din;
  assign fifo_Y_pe_25__dout = fifo_Y_pe_25_if_dout;
  assign fifo_Y_pe_25__empty_n = fifo_Y_pe_25_if_empty_n;
  assign fifo_Y_pe_25__full_n = fifo_Y_pe_25_if_full_n;
  assign fifo_Y_pe_25_if_read = fifo_Y_pe_25__read;
  assign fifo_Y_pe_25_if_read_ce = 1'b1;
  assign fifo_Y_pe_25_if_write = fifo_Y_pe_25__write;
  assign fifo_Y_pe_25_if_write_ce = 1'b1;
  assign fifo_Y_pe_25_reset = ~ ap_rst_n;
  assign fifo_Y_pe_26_clk = ap_clk;
  assign fifo_Y_pe_26_if_din = fifo_Y_pe_26__din;
  assign fifo_Y_pe_26__dout = fifo_Y_pe_26_if_dout;
  assign fifo_Y_pe_26__empty_n = fifo_Y_pe_26_if_empty_n;
  assign fifo_Y_pe_26__full_n = fifo_Y_pe_26_if_full_n;
  assign fifo_Y_pe_26_if_read = fifo_Y_pe_26__read;
  assign fifo_Y_pe_26_if_read_ce = 1'b1;
  assign fifo_Y_pe_26_if_write = fifo_Y_pe_26__write;
  assign fifo_Y_pe_26_if_write_ce = 1'b1;
  assign fifo_Y_pe_26_reset = ~ ap_rst_n;
  assign fifo_Y_pe_27_clk = ap_clk;
  assign fifo_Y_pe_27_if_din = fifo_Y_pe_27__din;
  assign fifo_Y_pe_27__dout = fifo_Y_pe_27_if_dout;
  assign fifo_Y_pe_27__empty_n = fifo_Y_pe_27_if_empty_n;
  assign fifo_Y_pe_27__full_n = fifo_Y_pe_27_if_full_n;
  assign fifo_Y_pe_27_if_read = fifo_Y_pe_27__read;
  assign fifo_Y_pe_27_if_read_ce = 1'b1;
  assign fifo_Y_pe_27_if_write = fifo_Y_pe_27__write;
  assign fifo_Y_pe_27_if_write_ce = 1'b1;
  assign fifo_Y_pe_27_reset = ~ ap_rst_n;
  assign fifo_Y_pe_28_clk = ap_clk;
  assign fifo_Y_pe_28_if_din = fifo_Y_pe_28__din;
  assign fifo_Y_pe_28__dout = fifo_Y_pe_28_if_dout;
  assign fifo_Y_pe_28__empty_n = fifo_Y_pe_28_if_empty_n;
  assign fifo_Y_pe_28__full_n = fifo_Y_pe_28_if_full_n;
  assign fifo_Y_pe_28_if_read = fifo_Y_pe_28__read;
  assign fifo_Y_pe_28_if_read_ce = 1'b1;
  assign fifo_Y_pe_28_if_write = fifo_Y_pe_28__write;
  assign fifo_Y_pe_28_if_write_ce = 1'b1;
  assign fifo_Y_pe_28_reset = ~ ap_rst_n;
  assign fifo_Y_pe_29_clk = ap_clk;
  assign fifo_Y_pe_29_if_din = fifo_Y_pe_29__din;
  assign fifo_Y_pe_29__dout = fifo_Y_pe_29_if_dout;
  assign fifo_Y_pe_29__empty_n = fifo_Y_pe_29_if_empty_n;
  assign fifo_Y_pe_29__full_n = fifo_Y_pe_29_if_full_n;
  assign fifo_Y_pe_29_if_read = fifo_Y_pe_29__read;
  assign fifo_Y_pe_29_if_read_ce = 1'b1;
  assign fifo_Y_pe_29_if_write = fifo_Y_pe_29__write;
  assign fifo_Y_pe_29_if_write_ce = 1'b1;
  assign fifo_Y_pe_29_reset = ~ ap_rst_n;
  assign fifo_Y_pe_2_clk = ap_clk;
  assign fifo_Y_pe_2_if_din = fifo_Y_pe_2__din;
  assign fifo_Y_pe_2__dout = fifo_Y_pe_2_if_dout;
  assign fifo_Y_pe_2__empty_n = fifo_Y_pe_2_if_empty_n;
  assign fifo_Y_pe_2__full_n = fifo_Y_pe_2_if_full_n;
  assign fifo_Y_pe_2_if_read = fifo_Y_pe_2__read;
  assign fifo_Y_pe_2_if_read_ce = 1'b1;
  assign fifo_Y_pe_2_if_write = fifo_Y_pe_2__write;
  assign fifo_Y_pe_2_if_write_ce = 1'b1;
  assign fifo_Y_pe_2_reset = ~ ap_rst_n;
  assign fifo_Y_pe_30_clk = ap_clk;
  assign fifo_Y_pe_30_if_din = fifo_Y_pe_30__din;
  assign fifo_Y_pe_30__dout = fifo_Y_pe_30_if_dout;
  assign fifo_Y_pe_30__empty_n = fifo_Y_pe_30_if_empty_n;
  assign fifo_Y_pe_30__full_n = fifo_Y_pe_30_if_full_n;
  assign fifo_Y_pe_30_if_read = fifo_Y_pe_30__read;
  assign fifo_Y_pe_30_if_read_ce = 1'b1;
  assign fifo_Y_pe_30_if_write = fifo_Y_pe_30__write;
  assign fifo_Y_pe_30_if_write_ce = 1'b1;
  assign fifo_Y_pe_30_reset = ~ ap_rst_n;
  assign fifo_Y_pe_31_clk = ap_clk;
  assign fifo_Y_pe_31_if_din = fifo_Y_pe_31__din;
  assign fifo_Y_pe_31__dout = fifo_Y_pe_31_if_dout;
  assign fifo_Y_pe_31__empty_n = fifo_Y_pe_31_if_empty_n;
  assign fifo_Y_pe_31__full_n = fifo_Y_pe_31_if_full_n;
  assign fifo_Y_pe_31_if_read = fifo_Y_pe_31__read;
  assign fifo_Y_pe_31_if_read_ce = 1'b1;
  assign fifo_Y_pe_31_if_write = fifo_Y_pe_31__write;
  assign fifo_Y_pe_31_if_write_ce = 1'b1;
  assign fifo_Y_pe_31_reset = ~ ap_rst_n;
  assign fifo_Y_pe_32_clk = ap_clk;
  assign fifo_Y_pe_32_if_din = fifo_Y_pe_32__din;
  assign fifo_Y_pe_32__dout = fifo_Y_pe_32_if_dout;
  assign fifo_Y_pe_32__empty_n = fifo_Y_pe_32_if_empty_n;
  assign fifo_Y_pe_32__full_n = fifo_Y_pe_32_if_full_n;
  assign fifo_Y_pe_32_if_read = fifo_Y_pe_32__read;
  assign fifo_Y_pe_32_if_read_ce = 1'b1;
  assign fifo_Y_pe_32_if_write = fifo_Y_pe_32__write;
  assign fifo_Y_pe_32_if_write_ce = 1'b1;
  assign fifo_Y_pe_32_reset = ~ ap_rst_n;
  assign fifo_Y_pe_33_clk = ap_clk;
  assign fifo_Y_pe_33_if_din = fifo_Y_pe_33__din;
  assign fifo_Y_pe_33__dout = fifo_Y_pe_33_if_dout;
  assign fifo_Y_pe_33__empty_n = fifo_Y_pe_33_if_empty_n;
  assign fifo_Y_pe_33__full_n = fifo_Y_pe_33_if_full_n;
  assign fifo_Y_pe_33_if_read = fifo_Y_pe_33__read;
  assign fifo_Y_pe_33_if_read_ce = 1'b1;
  assign fifo_Y_pe_33_if_write = fifo_Y_pe_33__write;
  assign fifo_Y_pe_33_if_write_ce = 1'b1;
  assign fifo_Y_pe_33_reset = ~ ap_rst_n;
  assign fifo_Y_pe_34_clk = ap_clk;
  assign fifo_Y_pe_34_if_din = fifo_Y_pe_34__din;
  assign fifo_Y_pe_34__dout = fifo_Y_pe_34_if_dout;
  assign fifo_Y_pe_34__empty_n = fifo_Y_pe_34_if_empty_n;
  assign fifo_Y_pe_34__full_n = fifo_Y_pe_34_if_full_n;
  assign fifo_Y_pe_34_if_read = fifo_Y_pe_34__read;
  assign fifo_Y_pe_34_if_read_ce = 1'b1;
  assign fifo_Y_pe_34_if_write = fifo_Y_pe_34__write;
  assign fifo_Y_pe_34_if_write_ce = 1'b1;
  assign fifo_Y_pe_34_reset = ~ ap_rst_n;
  assign fifo_Y_pe_35_clk = ap_clk;
  assign fifo_Y_pe_35_if_din = fifo_Y_pe_35__din;
  assign fifo_Y_pe_35__dout = fifo_Y_pe_35_if_dout;
  assign fifo_Y_pe_35__empty_n = fifo_Y_pe_35_if_empty_n;
  assign fifo_Y_pe_35__full_n = fifo_Y_pe_35_if_full_n;
  assign fifo_Y_pe_35_if_read = fifo_Y_pe_35__read;
  assign fifo_Y_pe_35_if_read_ce = 1'b1;
  assign fifo_Y_pe_35_if_write = fifo_Y_pe_35__write;
  assign fifo_Y_pe_35_if_write_ce = 1'b1;
  assign fifo_Y_pe_35_reset = ~ ap_rst_n;
  assign fifo_Y_pe_36_clk = ap_clk;
  assign fifo_Y_pe_36_if_din = fifo_Y_pe_36__din;
  assign fifo_Y_pe_36__dout = fifo_Y_pe_36_if_dout;
  assign fifo_Y_pe_36__empty_n = fifo_Y_pe_36_if_empty_n;
  assign fifo_Y_pe_36__full_n = fifo_Y_pe_36_if_full_n;
  assign fifo_Y_pe_36_if_read = fifo_Y_pe_36__read;
  assign fifo_Y_pe_36_if_read_ce = 1'b1;
  assign fifo_Y_pe_36_if_write = fifo_Y_pe_36__write;
  assign fifo_Y_pe_36_if_write_ce = 1'b1;
  assign fifo_Y_pe_36_reset = ~ ap_rst_n;
  assign fifo_Y_pe_37_clk = ap_clk;
  assign fifo_Y_pe_37_if_din = fifo_Y_pe_37__din;
  assign fifo_Y_pe_37__dout = fifo_Y_pe_37_if_dout;
  assign fifo_Y_pe_37__empty_n = fifo_Y_pe_37_if_empty_n;
  assign fifo_Y_pe_37__full_n = fifo_Y_pe_37_if_full_n;
  assign fifo_Y_pe_37_if_read = fifo_Y_pe_37__read;
  assign fifo_Y_pe_37_if_read_ce = 1'b1;
  assign fifo_Y_pe_37_if_write = fifo_Y_pe_37__write;
  assign fifo_Y_pe_37_if_write_ce = 1'b1;
  assign fifo_Y_pe_37_reset = ~ ap_rst_n;
  assign fifo_Y_pe_38_clk = ap_clk;
  assign fifo_Y_pe_38_if_din = fifo_Y_pe_38__din;
  assign fifo_Y_pe_38__dout = fifo_Y_pe_38_if_dout;
  assign fifo_Y_pe_38__empty_n = fifo_Y_pe_38_if_empty_n;
  assign fifo_Y_pe_38__full_n = fifo_Y_pe_38_if_full_n;
  assign fifo_Y_pe_38_if_read = fifo_Y_pe_38__read;
  assign fifo_Y_pe_38_if_read_ce = 1'b1;
  assign fifo_Y_pe_38_if_write = fifo_Y_pe_38__write;
  assign fifo_Y_pe_38_if_write_ce = 1'b1;
  assign fifo_Y_pe_38_reset = ~ ap_rst_n;
  assign fifo_Y_pe_39_clk = ap_clk;
  assign fifo_Y_pe_39_if_din = fifo_Y_pe_39__din;
  assign fifo_Y_pe_39__dout = fifo_Y_pe_39_if_dout;
  assign fifo_Y_pe_39__empty_n = fifo_Y_pe_39_if_empty_n;
  assign fifo_Y_pe_39__full_n = fifo_Y_pe_39_if_full_n;
  assign fifo_Y_pe_39_if_read = fifo_Y_pe_39__read;
  assign fifo_Y_pe_39_if_read_ce = 1'b1;
  assign fifo_Y_pe_39_if_write = fifo_Y_pe_39__write;
  assign fifo_Y_pe_39_if_write_ce = 1'b1;
  assign fifo_Y_pe_39_reset = ~ ap_rst_n;
  assign fifo_Y_pe_3_clk = ap_clk;
  assign fifo_Y_pe_3_if_din = fifo_Y_pe_3__din;
  assign fifo_Y_pe_3__dout = fifo_Y_pe_3_if_dout;
  assign fifo_Y_pe_3__empty_n = fifo_Y_pe_3_if_empty_n;
  assign fifo_Y_pe_3__full_n = fifo_Y_pe_3_if_full_n;
  assign fifo_Y_pe_3_if_read = fifo_Y_pe_3__read;
  assign fifo_Y_pe_3_if_read_ce = 1'b1;
  assign fifo_Y_pe_3_if_write = fifo_Y_pe_3__write;
  assign fifo_Y_pe_3_if_write_ce = 1'b1;
  assign fifo_Y_pe_3_reset = ~ ap_rst_n;
  assign fifo_Y_pe_40_clk = ap_clk;
  assign fifo_Y_pe_40_if_din = fifo_Y_pe_40__din;
  assign fifo_Y_pe_40__dout = fifo_Y_pe_40_if_dout;
  assign fifo_Y_pe_40__empty_n = fifo_Y_pe_40_if_empty_n;
  assign fifo_Y_pe_40__full_n = fifo_Y_pe_40_if_full_n;
  assign fifo_Y_pe_40_if_read = fifo_Y_pe_40__read;
  assign fifo_Y_pe_40_if_read_ce = 1'b1;
  assign fifo_Y_pe_40_if_write = fifo_Y_pe_40__write;
  assign fifo_Y_pe_40_if_write_ce = 1'b1;
  assign fifo_Y_pe_40_reset = ~ ap_rst_n;
  assign fifo_Y_pe_41_clk = ap_clk;
  assign fifo_Y_pe_41_if_din = fifo_Y_pe_41__din;
  assign fifo_Y_pe_41__dout = fifo_Y_pe_41_if_dout;
  assign fifo_Y_pe_41__empty_n = fifo_Y_pe_41_if_empty_n;
  assign fifo_Y_pe_41__full_n = fifo_Y_pe_41_if_full_n;
  assign fifo_Y_pe_41_if_read = fifo_Y_pe_41__read;
  assign fifo_Y_pe_41_if_read_ce = 1'b1;
  assign fifo_Y_pe_41_if_write = fifo_Y_pe_41__write;
  assign fifo_Y_pe_41_if_write_ce = 1'b1;
  assign fifo_Y_pe_41_reset = ~ ap_rst_n;
  assign fifo_Y_pe_42_clk = ap_clk;
  assign fifo_Y_pe_42_if_din = fifo_Y_pe_42__din;
  assign fifo_Y_pe_42__dout = fifo_Y_pe_42_if_dout;
  assign fifo_Y_pe_42__empty_n = fifo_Y_pe_42_if_empty_n;
  assign fifo_Y_pe_42__full_n = fifo_Y_pe_42_if_full_n;
  assign fifo_Y_pe_42_if_read = fifo_Y_pe_42__read;
  assign fifo_Y_pe_42_if_read_ce = 1'b1;
  assign fifo_Y_pe_42_if_write = fifo_Y_pe_42__write;
  assign fifo_Y_pe_42_if_write_ce = 1'b1;
  assign fifo_Y_pe_42_reset = ~ ap_rst_n;
  assign fifo_Y_pe_43_clk = ap_clk;
  assign fifo_Y_pe_43_if_din = fifo_Y_pe_43__din;
  assign fifo_Y_pe_43__dout = fifo_Y_pe_43_if_dout;
  assign fifo_Y_pe_43__empty_n = fifo_Y_pe_43_if_empty_n;
  assign fifo_Y_pe_43__full_n = fifo_Y_pe_43_if_full_n;
  assign fifo_Y_pe_43_if_read = fifo_Y_pe_43__read;
  assign fifo_Y_pe_43_if_read_ce = 1'b1;
  assign fifo_Y_pe_43_if_write = fifo_Y_pe_43__write;
  assign fifo_Y_pe_43_if_write_ce = 1'b1;
  assign fifo_Y_pe_43_reset = ~ ap_rst_n;
  assign fifo_Y_pe_44_clk = ap_clk;
  assign fifo_Y_pe_44_if_din = fifo_Y_pe_44__din;
  assign fifo_Y_pe_44__dout = fifo_Y_pe_44_if_dout;
  assign fifo_Y_pe_44__empty_n = fifo_Y_pe_44_if_empty_n;
  assign fifo_Y_pe_44__full_n = fifo_Y_pe_44_if_full_n;
  assign fifo_Y_pe_44_if_read = fifo_Y_pe_44__read;
  assign fifo_Y_pe_44_if_read_ce = 1'b1;
  assign fifo_Y_pe_44_if_write = fifo_Y_pe_44__write;
  assign fifo_Y_pe_44_if_write_ce = 1'b1;
  assign fifo_Y_pe_44_reset = ~ ap_rst_n;
  assign fifo_Y_pe_45_clk = ap_clk;
  assign fifo_Y_pe_45_if_din = fifo_Y_pe_45__din;
  assign fifo_Y_pe_45__dout = fifo_Y_pe_45_if_dout;
  assign fifo_Y_pe_45__empty_n = fifo_Y_pe_45_if_empty_n;
  assign fifo_Y_pe_45__full_n = fifo_Y_pe_45_if_full_n;
  assign fifo_Y_pe_45_if_read = fifo_Y_pe_45__read;
  assign fifo_Y_pe_45_if_read_ce = 1'b1;
  assign fifo_Y_pe_45_if_write = fifo_Y_pe_45__write;
  assign fifo_Y_pe_45_if_write_ce = 1'b1;
  assign fifo_Y_pe_45_reset = ~ ap_rst_n;
  assign fifo_Y_pe_46_clk = ap_clk;
  assign fifo_Y_pe_46_if_din = fifo_Y_pe_46__din;
  assign fifo_Y_pe_46__dout = fifo_Y_pe_46_if_dout;
  assign fifo_Y_pe_46__empty_n = fifo_Y_pe_46_if_empty_n;
  assign fifo_Y_pe_46__full_n = fifo_Y_pe_46_if_full_n;
  assign fifo_Y_pe_46_if_read = fifo_Y_pe_46__read;
  assign fifo_Y_pe_46_if_read_ce = 1'b1;
  assign fifo_Y_pe_46_if_write = fifo_Y_pe_46__write;
  assign fifo_Y_pe_46_if_write_ce = 1'b1;
  assign fifo_Y_pe_46_reset = ~ ap_rst_n;
  assign fifo_Y_pe_47_clk = ap_clk;
  assign fifo_Y_pe_47_if_din = fifo_Y_pe_47__din;
  assign fifo_Y_pe_47__dout = fifo_Y_pe_47_if_dout;
  assign fifo_Y_pe_47__empty_n = fifo_Y_pe_47_if_empty_n;
  assign fifo_Y_pe_47__full_n = fifo_Y_pe_47_if_full_n;
  assign fifo_Y_pe_47_if_read = fifo_Y_pe_47__read;
  assign fifo_Y_pe_47_if_read_ce = 1'b1;
  assign fifo_Y_pe_47_if_write = fifo_Y_pe_47__write;
  assign fifo_Y_pe_47_if_write_ce = 1'b1;
  assign fifo_Y_pe_47_reset = ~ ap_rst_n;
  assign fifo_Y_pe_4_clk = ap_clk;
  assign fifo_Y_pe_4_if_din = fifo_Y_pe_4__din;
  assign fifo_Y_pe_4__dout = fifo_Y_pe_4_if_dout;
  assign fifo_Y_pe_4__empty_n = fifo_Y_pe_4_if_empty_n;
  assign fifo_Y_pe_4__full_n = fifo_Y_pe_4_if_full_n;
  assign fifo_Y_pe_4_if_read = fifo_Y_pe_4__read;
  assign fifo_Y_pe_4_if_read_ce = 1'b1;
  assign fifo_Y_pe_4_if_write = fifo_Y_pe_4__write;
  assign fifo_Y_pe_4_if_write_ce = 1'b1;
  assign fifo_Y_pe_4_reset = ~ ap_rst_n;
  assign fifo_Y_pe_5_clk = ap_clk;
  assign fifo_Y_pe_5_if_din = fifo_Y_pe_5__din;
  assign fifo_Y_pe_5__dout = fifo_Y_pe_5_if_dout;
  assign fifo_Y_pe_5__empty_n = fifo_Y_pe_5_if_empty_n;
  assign fifo_Y_pe_5__full_n = fifo_Y_pe_5_if_full_n;
  assign fifo_Y_pe_5_if_read = fifo_Y_pe_5__read;
  assign fifo_Y_pe_5_if_read_ce = 1'b1;
  assign fifo_Y_pe_5_if_write = fifo_Y_pe_5__write;
  assign fifo_Y_pe_5_if_write_ce = 1'b1;
  assign fifo_Y_pe_5_reset = ~ ap_rst_n;
  assign fifo_Y_pe_6_clk = ap_clk;
  assign fifo_Y_pe_6_if_din = fifo_Y_pe_6__din;
  assign fifo_Y_pe_6__dout = fifo_Y_pe_6_if_dout;
  assign fifo_Y_pe_6__empty_n = fifo_Y_pe_6_if_empty_n;
  assign fifo_Y_pe_6__full_n = fifo_Y_pe_6_if_full_n;
  assign fifo_Y_pe_6_if_read = fifo_Y_pe_6__read;
  assign fifo_Y_pe_6_if_read_ce = 1'b1;
  assign fifo_Y_pe_6_if_write = fifo_Y_pe_6__write;
  assign fifo_Y_pe_6_if_write_ce = 1'b1;
  assign fifo_Y_pe_6_reset = ~ ap_rst_n;
  assign fifo_Y_pe_7_clk = ap_clk;
  assign fifo_Y_pe_7_if_din = fifo_Y_pe_7__din;
  assign fifo_Y_pe_7__dout = fifo_Y_pe_7_if_dout;
  assign fifo_Y_pe_7__empty_n = fifo_Y_pe_7_if_empty_n;
  assign fifo_Y_pe_7__full_n = fifo_Y_pe_7_if_full_n;
  assign fifo_Y_pe_7_if_read = fifo_Y_pe_7__read;
  assign fifo_Y_pe_7_if_read_ce = 1'b1;
  assign fifo_Y_pe_7_if_write = fifo_Y_pe_7__write;
  assign fifo_Y_pe_7_if_write_ce = 1'b1;
  assign fifo_Y_pe_7_reset = ~ ap_rst_n;
  assign fifo_Y_pe_8_clk = ap_clk;
  assign fifo_Y_pe_8_if_din = fifo_Y_pe_8__din;
  assign fifo_Y_pe_8__dout = fifo_Y_pe_8_if_dout;
  assign fifo_Y_pe_8__empty_n = fifo_Y_pe_8_if_empty_n;
  assign fifo_Y_pe_8__full_n = fifo_Y_pe_8_if_full_n;
  assign fifo_Y_pe_8_if_read = fifo_Y_pe_8__read;
  assign fifo_Y_pe_8_if_read_ce = 1'b1;
  assign fifo_Y_pe_8_if_write = fifo_Y_pe_8__write;
  assign fifo_Y_pe_8_if_write_ce = 1'b1;
  assign fifo_Y_pe_8_reset = ~ ap_rst_n;
  assign fifo_Y_pe_9_clk = ap_clk;
  assign fifo_Y_pe_9_if_din = fifo_Y_pe_9__din;
  assign fifo_Y_pe_9__dout = fifo_Y_pe_9_if_dout;
  assign fifo_Y_pe_9__empty_n = fifo_Y_pe_9_if_empty_n;
  assign fifo_Y_pe_9__full_n = fifo_Y_pe_9_if_full_n;
  assign fifo_Y_pe_9_if_read = fifo_Y_pe_9__read;
  assign fifo_Y_pe_9_if_read_ce = 1'b1;
  assign fifo_Y_pe_9_if_write = fifo_Y_pe_9__write;
  assign fifo_Y_pe_9_if_write_ce = 1'b1;
  assign fifo_Y_pe_9_reset = ~ ap_rst_n;
  assign fifo_Y_pe_abd_0_clk = ap_clk;
  assign fifo_Y_pe_abd_0_if_din = fifo_Y_pe_abd_0__din;
  assign fifo_Y_pe_abd_0__dout = fifo_Y_pe_abd_0_if_dout;
  assign fifo_Y_pe_abd_0__empty_n = fifo_Y_pe_abd_0_if_empty_n;
  assign fifo_Y_pe_abd_0__full_n = fifo_Y_pe_abd_0_if_full_n;
  assign fifo_Y_pe_abd_0_if_read = fifo_Y_pe_abd_0__read;
  assign fifo_Y_pe_abd_0_if_read_ce = 1'b1;
  assign fifo_Y_pe_abd_0_if_write = fifo_Y_pe_abd_0__write;
  assign fifo_Y_pe_abd_0_if_write_ce = 1'b1;
  assign fifo_Y_pe_abd_0_reset = ~ ap_rst_n;
  assign fifo_Y_pe_abd_1_clk = ap_clk;
  assign fifo_Y_pe_abd_1_if_din = fifo_Y_pe_abd_1__din;
  assign fifo_Y_pe_abd_1__dout = fifo_Y_pe_abd_1_if_dout;
  assign fifo_Y_pe_abd_1__empty_n = fifo_Y_pe_abd_1_if_empty_n;
  assign fifo_Y_pe_abd_1__full_n = fifo_Y_pe_abd_1_if_full_n;
  assign fifo_Y_pe_abd_1_if_read = fifo_Y_pe_abd_1__read;
  assign fifo_Y_pe_abd_1_if_read_ce = 1'b1;
  assign fifo_Y_pe_abd_1_if_write = fifo_Y_pe_abd_1__write;
  assign fifo_Y_pe_abd_1_if_write_ce = 1'b1;
  assign fifo_Y_pe_abd_1_reset = ~ ap_rst_n;
  assign fifo_Y_pe_abd_2_clk = ap_clk;
  assign fifo_Y_pe_abd_2_if_din = fifo_Y_pe_abd_2__din;
  assign fifo_Y_pe_abd_2__dout = fifo_Y_pe_abd_2_if_dout;
  assign fifo_Y_pe_abd_2__empty_n = fifo_Y_pe_abd_2_if_empty_n;
  assign fifo_Y_pe_abd_2__full_n = fifo_Y_pe_abd_2_if_full_n;
  assign fifo_Y_pe_abd_2_if_read = fifo_Y_pe_abd_2__read;
  assign fifo_Y_pe_abd_2_if_read_ce = 1'b1;
  assign fifo_Y_pe_abd_2_if_write = fifo_Y_pe_abd_2__write;
  assign fifo_Y_pe_abd_2_if_write_ce = 1'b1;
  assign fifo_Y_pe_abd_2_reset = ~ ap_rst_n;
  assign fifo_Y_pe_abd_3_clk = ap_clk;
  assign fifo_Y_pe_abd_3_if_din = fifo_Y_pe_abd_3__din;
  assign fifo_Y_pe_abd_3__dout = fifo_Y_pe_abd_3_if_dout;
  assign fifo_Y_pe_abd_3__empty_n = fifo_Y_pe_abd_3_if_empty_n;
  assign fifo_Y_pe_abd_3__full_n = fifo_Y_pe_abd_3_if_full_n;
  assign fifo_Y_pe_abd_3_if_read = fifo_Y_pe_abd_3__read;
  assign fifo_Y_pe_abd_3_if_read_ce = 1'b1;
  assign fifo_Y_pe_abd_3_if_write = fifo_Y_pe_abd_3__write;
  assign fifo_Y_pe_abd_3_if_write_ce = 1'b1;
  assign fifo_Y_pe_abd_3_reset = ~ ap_rst_n;
  assign fifo_Y_pe_abd_4_clk = ap_clk;
  assign fifo_Y_pe_abd_4_if_din = fifo_Y_pe_abd_4__din;
  assign fifo_Y_pe_abd_4__dout = fifo_Y_pe_abd_4_if_dout;
  assign fifo_Y_pe_abd_4__empty_n = fifo_Y_pe_abd_4_if_empty_n;
  assign fifo_Y_pe_abd_4__full_n = fifo_Y_pe_abd_4_if_full_n;
  assign fifo_Y_pe_abd_4_if_read = fifo_Y_pe_abd_4__read;
  assign fifo_Y_pe_abd_4_if_read_ce = 1'b1;
  assign fifo_Y_pe_abd_4_if_write = fifo_Y_pe_abd_4__write;
  assign fifo_Y_pe_abd_4_if_write_ce = 1'b1;
  assign fifo_Y_pe_abd_4_reset = ~ ap_rst_n;
  assign fifo_Y_pe_abd_5_clk = ap_clk;
  assign fifo_Y_pe_abd_5_if_din = fifo_Y_pe_abd_5__din;
  assign fifo_Y_pe_abd_5__dout = fifo_Y_pe_abd_5_if_dout;
  assign fifo_Y_pe_abd_5__empty_n = fifo_Y_pe_abd_5_if_empty_n;
  assign fifo_Y_pe_abd_5__full_n = fifo_Y_pe_abd_5_if_full_n;
  assign fifo_Y_pe_abd_5_if_read = fifo_Y_pe_abd_5__read;
  assign fifo_Y_pe_abd_5_if_read_ce = 1'b1;
  assign fifo_Y_pe_abd_5_if_write = fifo_Y_pe_abd_5__write;
  assign fifo_Y_pe_abd_5_if_write_ce = 1'b1;
  assign fifo_Y_pe_abd_5_reset = ~ ap_rst_n;
  assign fifo_Y_pe_abd_6_clk = ap_clk;
  assign fifo_Y_pe_abd_6_if_din = fifo_Y_pe_abd_6__din;
  assign fifo_Y_pe_abd_6__dout = fifo_Y_pe_abd_6_if_dout;
  assign fifo_Y_pe_abd_6__empty_n = fifo_Y_pe_abd_6_if_empty_n;
  assign fifo_Y_pe_abd_6__full_n = fifo_Y_pe_abd_6_if_full_n;
  assign fifo_Y_pe_abd_6_if_read = fifo_Y_pe_abd_6__read;
  assign fifo_Y_pe_abd_6_if_read_ce = 1'b1;
  assign fifo_Y_pe_abd_6_if_write = fifo_Y_pe_abd_6__write;
  assign fifo_Y_pe_abd_6_if_write_ce = 1'b1;
  assign fifo_Y_pe_abd_6_reset = ~ ap_rst_n;
  assign fifo_Y_pe_abd_7_clk = ap_clk;
  assign fifo_Y_pe_abd_7_if_din = fifo_Y_pe_abd_7__din;
  assign fifo_Y_pe_abd_7__dout = fifo_Y_pe_abd_7_if_dout;
  assign fifo_Y_pe_abd_7__empty_n = fifo_Y_pe_abd_7_if_empty_n;
  assign fifo_Y_pe_abd_7__full_n = fifo_Y_pe_abd_7_if_full_n;
  assign fifo_Y_pe_abd_7_if_read = fifo_Y_pe_abd_7__read;
  assign fifo_Y_pe_abd_7_if_read_ce = 1'b1;
  assign fifo_Y_pe_abd_7_if_write = fifo_Y_pe_abd_7__write;
  assign fifo_Y_pe_abd_7_if_write_ce = 1'b1;
  assign fifo_Y_pe_abd_7_reset = ~ ap_rst_n;
  assign fifo_aXvec_0_clk = ap_clk;
  assign fifo_aXvec_0_if_din = fifo_aXvec_0__din;
  assign fifo_aXvec_0__dout = fifo_aXvec_0_if_dout;
  assign fifo_aXvec_0__empty_n = fifo_aXvec_0_if_empty_n;
  assign fifo_aXvec_0__full_n = fifo_aXvec_0_if_full_n;
  assign fifo_aXvec_0_if_read = fifo_aXvec_0__read;
  assign fifo_aXvec_0_if_read_ce = 1'b1;
  assign fifo_aXvec_0_if_write = fifo_aXvec_0__write;
  assign fifo_aXvec_0_if_write_ce = 1'b1;
  assign fifo_aXvec_0_reset = ~ ap_rst_n;
  assign fifo_aXvec_10_clk = ap_clk;
  assign fifo_aXvec_10_if_din = fifo_aXvec_10__din;
  assign fifo_aXvec_10__dout = fifo_aXvec_10_if_dout;
  assign fifo_aXvec_10__empty_n = fifo_aXvec_10_if_empty_n;
  assign fifo_aXvec_10__full_n = fifo_aXvec_10_if_full_n;
  assign fifo_aXvec_10_if_read = fifo_aXvec_10__read;
  assign fifo_aXvec_10_if_read_ce = 1'b1;
  assign fifo_aXvec_10_if_write = fifo_aXvec_10__write;
  assign fifo_aXvec_10_if_write_ce = 1'b1;
  assign fifo_aXvec_10_reset = ~ ap_rst_n;
  assign fifo_aXvec_11_clk = ap_clk;
  assign fifo_aXvec_11_if_din = fifo_aXvec_11__din;
  assign fifo_aXvec_11__dout = fifo_aXvec_11_if_dout;
  assign fifo_aXvec_11__empty_n = fifo_aXvec_11_if_empty_n;
  assign fifo_aXvec_11__full_n = fifo_aXvec_11_if_full_n;
  assign fifo_aXvec_11_if_read = fifo_aXvec_11__read;
  assign fifo_aXvec_11_if_read_ce = 1'b1;
  assign fifo_aXvec_11_if_write = fifo_aXvec_11__write;
  assign fifo_aXvec_11_if_write_ce = 1'b1;
  assign fifo_aXvec_11_reset = ~ ap_rst_n;
  assign fifo_aXvec_12_clk = ap_clk;
  assign fifo_aXvec_12_if_din = fifo_aXvec_12__din;
  assign fifo_aXvec_12__dout = fifo_aXvec_12_if_dout;
  assign fifo_aXvec_12__empty_n = fifo_aXvec_12_if_empty_n;
  assign fifo_aXvec_12__full_n = fifo_aXvec_12_if_full_n;
  assign fifo_aXvec_12_if_read = fifo_aXvec_12__read;
  assign fifo_aXvec_12_if_read_ce = 1'b1;
  assign fifo_aXvec_12_if_write = fifo_aXvec_12__write;
  assign fifo_aXvec_12_if_write_ce = 1'b1;
  assign fifo_aXvec_12_reset = ~ ap_rst_n;
  assign fifo_aXvec_13_clk = ap_clk;
  assign fifo_aXvec_13_if_din = fifo_aXvec_13__din;
  assign fifo_aXvec_13__dout = fifo_aXvec_13_if_dout;
  assign fifo_aXvec_13__empty_n = fifo_aXvec_13_if_empty_n;
  assign fifo_aXvec_13__full_n = fifo_aXvec_13_if_full_n;
  assign fifo_aXvec_13_if_read = fifo_aXvec_13__read;
  assign fifo_aXvec_13_if_read_ce = 1'b1;
  assign fifo_aXvec_13_if_write = fifo_aXvec_13__write;
  assign fifo_aXvec_13_if_write_ce = 1'b1;
  assign fifo_aXvec_13_reset = ~ ap_rst_n;
  assign fifo_aXvec_14_clk = ap_clk;
  assign fifo_aXvec_14_if_din = fifo_aXvec_14__din;
  assign fifo_aXvec_14__dout = fifo_aXvec_14_if_dout;
  assign fifo_aXvec_14__empty_n = fifo_aXvec_14_if_empty_n;
  assign fifo_aXvec_14__full_n = fifo_aXvec_14_if_full_n;
  assign fifo_aXvec_14_if_read = fifo_aXvec_14__read;
  assign fifo_aXvec_14_if_read_ce = 1'b1;
  assign fifo_aXvec_14_if_write = fifo_aXvec_14__write;
  assign fifo_aXvec_14_if_write_ce = 1'b1;
  assign fifo_aXvec_14_reset = ~ ap_rst_n;
  assign fifo_aXvec_15_clk = ap_clk;
  assign fifo_aXvec_15_if_din = fifo_aXvec_15__din;
  assign fifo_aXvec_15__dout = fifo_aXvec_15_if_dout;
  assign fifo_aXvec_15__empty_n = fifo_aXvec_15_if_empty_n;
  assign fifo_aXvec_15__full_n = fifo_aXvec_15_if_full_n;
  assign fifo_aXvec_15_if_read = fifo_aXvec_15__read;
  assign fifo_aXvec_15_if_read_ce = 1'b1;
  assign fifo_aXvec_15_if_write = fifo_aXvec_15__write;
  assign fifo_aXvec_15_if_write_ce = 1'b1;
  assign fifo_aXvec_15_reset = ~ ap_rst_n;
  assign fifo_aXvec_16_clk = ap_clk;
  assign fifo_aXvec_16_if_din = fifo_aXvec_16__din;
  assign fifo_aXvec_16__dout = fifo_aXvec_16_if_dout;
  assign fifo_aXvec_16__empty_n = fifo_aXvec_16_if_empty_n;
  assign fifo_aXvec_16__full_n = fifo_aXvec_16_if_full_n;
  assign fifo_aXvec_16_if_read = fifo_aXvec_16__read;
  assign fifo_aXvec_16_if_read_ce = 1'b1;
  assign fifo_aXvec_16_if_write = fifo_aXvec_16__write;
  assign fifo_aXvec_16_if_write_ce = 1'b1;
  assign fifo_aXvec_16_reset = ~ ap_rst_n;
  assign fifo_aXvec_17_clk = ap_clk;
  assign fifo_aXvec_17_if_din = fifo_aXvec_17__din;
  assign fifo_aXvec_17__dout = fifo_aXvec_17_if_dout;
  assign fifo_aXvec_17__empty_n = fifo_aXvec_17_if_empty_n;
  assign fifo_aXvec_17__full_n = fifo_aXvec_17_if_full_n;
  assign fifo_aXvec_17_if_read = fifo_aXvec_17__read;
  assign fifo_aXvec_17_if_read_ce = 1'b1;
  assign fifo_aXvec_17_if_write = fifo_aXvec_17__write;
  assign fifo_aXvec_17_if_write_ce = 1'b1;
  assign fifo_aXvec_17_reset = ~ ap_rst_n;
  assign fifo_aXvec_18_clk = ap_clk;
  assign fifo_aXvec_18_if_din = fifo_aXvec_18__din;
  assign fifo_aXvec_18__dout = fifo_aXvec_18_if_dout;
  assign fifo_aXvec_18__empty_n = fifo_aXvec_18_if_empty_n;
  assign fifo_aXvec_18__full_n = fifo_aXvec_18_if_full_n;
  assign fifo_aXvec_18_if_read = fifo_aXvec_18__read;
  assign fifo_aXvec_18_if_read_ce = 1'b1;
  assign fifo_aXvec_18_if_write = fifo_aXvec_18__write;
  assign fifo_aXvec_18_if_write_ce = 1'b1;
  assign fifo_aXvec_18_reset = ~ ap_rst_n;
  assign fifo_aXvec_19_clk = ap_clk;
  assign fifo_aXvec_19_if_din = fifo_aXvec_19__din;
  assign fifo_aXvec_19__dout = fifo_aXvec_19_if_dout;
  assign fifo_aXvec_19__empty_n = fifo_aXvec_19_if_empty_n;
  assign fifo_aXvec_19__full_n = fifo_aXvec_19_if_full_n;
  assign fifo_aXvec_19_if_read = fifo_aXvec_19__read;
  assign fifo_aXvec_19_if_read_ce = 1'b1;
  assign fifo_aXvec_19_if_write = fifo_aXvec_19__write;
  assign fifo_aXvec_19_if_write_ce = 1'b1;
  assign fifo_aXvec_19_reset = ~ ap_rst_n;
  assign fifo_aXvec_1_clk = ap_clk;
  assign fifo_aXvec_1_if_din = fifo_aXvec_1__din;
  assign fifo_aXvec_1__dout = fifo_aXvec_1_if_dout;
  assign fifo_aXvec_1__empty_n = fifo_aXvec_1_if_empty_n;
  assign fifo_aXvec_1__full_n = fifo_aXvec_1_if_full_n;
  assign fifo_aXvec_1_if_read = fifo_aXvec_1__read;
  assign fifo_aXvec_1_if_read_ce = 1'b1;
  assign fifo_aXvec_1_if_write = fifo_aXvec_1__write;
  assign fifo_aXvec_1_if_write_ce = 1'b1;
  assign fifo_aXvec_1_reset = ~ ap_rst_n;
  assign fifo_aXvec_20_clk = ap_clk;
  assign fifo_aXvec_20_if_din = fifo_aXvec_20__din;
  assign fifo_aXvec_20__dout = fifo_aXvec_20_if_dout;
  assign fifo_aXvec_20__empty_n = fifo_aXvec_20_if_empty_n;
  assign fifo_aXvec_20__full_n = fifo_aXvec_20_if_full_n;
  assign fifo_aXvec_20_if_read = fifo_aXvec_20__read;
  assign fifo_aXvec_20_if_read_ce = 1'b1;
  assign fifo_aXvec_20_if_write = fifo_aXvec_20__write;
  assign fifo_aXvec_20_if_write_ce = 1'b1;
  assign fifo_aXvec_20_reset = ~ ap_rst_n;
  assign fifo_aXvec_21_clk = ap_clk;
  assign fifo_aXvec_21_if_din = fifo_aXvec_21__din;
  assign fifo_aXvec_21__dout = fifo_aXvec_21_if_dout;
  assign fifo_aXvec_21__empty_n = fifo_aXvec_21_if_empty_n;
  assign fifo_aXvec_21__full_n = fifo_aXvec_21_if_full_n;
  assign fifo_aXvec_21_if_read = fifo_aXvec_21__read;
  assign fifo_aXvec_21_if_read_ce = 1'b1;
  assign fifo_aXvec_21_if_write = fifo_aXvec_21__write;
  assign fifo_aXvec_21_if_write_ce = 1'b1;
  assign fifo_aXvec_21_reset = ~ ap_rst_n;
  assign fifo_aXvec_22_clk = ap_clk;
  assign fifo_aXvec_22_if_din = fifo_aXvec_22__din;
  assign fifo_aXvec_22__dout = fifo_aXvec_22_if_dout;
  assign fifo_aXvec_22__empty_n = fifo_aXvec_22_if_empty_n;
  assign fifo_aXvec_22__full_n = fifo_aXvec_22_if_full_n;
  assign fifo_aXvec_22_if_read = fifo_aXvec_22__read;
  assign fifo_aXvec_22_if_read_ce = 1'b1;
  assign fifo_aXvec_22_if_write = fifo_aXvec_22__write;
  assign fifo_aXvec_22_if_write_ce = 1'b1;
  assign fifo_aXvec_22_reset = ~ ap_rst_n;
  assign fifo_aXvec_23_clk = ap_clk;
  assign fifo_aXvec_23_if_din = fifo_aXvec_23__din;
  assign fifo_aXvec_23__dout = fifo_aXvec_23_if_dout;
  assign fifo_aXvec_23__empty_n = fifo_aXvec_23_if_empty_n;
  assign fifo_aXvec_23__full_n = fifo_aXvec_23_if_full_n;
  assign fifo_aXvec_23_if_read = fifo_aXvec_23__read;
  assign fifo_aXvec_23_if_read_ce = 1'b1;
  assign fifo_aXvec_23_if_write = fifo_aXvec_23__write;
  assign fifo_aXvec_23_if_write_ce = 1'b1;
  assign fifo_aXvec_23_reset = ~ ap_rst_n;
  assign fifo_aXvec_24_clk = ap_clk;
  assign fifo_aXvec_24_if_din = fifo_aXvec_24__din;
  assign fifo_aXvec_24__dout = fifo_aXvec_24_if_dout;
  assign fifo_aXvec_24__empty_n = fifo_aXvec_24_if_empty_n;
  assign fifo_aXvec_24__full_n = fifo_aXvec_24_if_full_n;
  assign fifo_aXvec_24_if_read = fifo_aXvec_24__read;
  assign fifo_aXvec_24_if_read_ce = 1'b1;
  assign fifo_aXvec_24_if_write = fifo_aXvec_24__write;
  assign fifo_aXvec_24_if_write_ce = 1'b1;
  assign fifo_aXvec_24_reset = ~ ap_rst_n;
  assign fifo_aXvec_25_clk = ap_clk;
  assign fifo_aXvec_25_if_din = fifo_aXvec_25__din;
  assign fifo_aXvec_25__dout = fifo_aXvec_25_if_dout;
  assign fifo_aXvec_25__empty_n = fifo_aXvec_25_if_empty_n;
  assign fifo_aXvec_25__full_n = fifo_aXvec_25_if_full_n;
  assign fifo_aXvec_25_if_read = fifo_aXvec_25__read;
  assign fifo_aXvec_25_if_read_ce = 1'b1;
  assign fifo_aXvec_25_if_write = fifo_aXvec_25__write;
  assign fifo_aXvec_25_if_write_ce = 1'b1;
  assign fifo_aXvec_25_reset = ~ ap_rst_n;
  assign fifo_aXvec_26_clk = ap_clk;
  assign fifo_aXvec_26_if_din = fifo_aXvec_26__din;
  assign fifo_aXvec_26__dout = fifo_aXvec_26_if_dout;
  assign fifo_aXvec_26__empty_n = fifo_aXvec_26_if_empty_n;
  assign fifo_aXvec_26__full_n = fifo_aXvec_26_if_full_n;
  assign fifo_aXvec_26_if_read = fifo_aXvec_26__read;
  assign fifo_aXvec_26_if_read_ce = 1'b1;
  assign fifo_aXvec_26_if_write = fifo_aXvec_26__write;
  assign fifo_aXvec_26_if_write_ce = 1'b1;
  assign fifo_aXvec_26_reset = ~ ap_rst_n;
  assign fifo_aXvec_27_clk = ap_clk;
  assign fifo_aXvec_27_if_din = fifo_aXvec_27__din;
  assign fifo_aXvec_27__dout = fifo_aXvec_27_if_dout;
  assign fifo_aXvec_27__empty_n = fifo_aXvec_27_if_empty_n;
  assign fifo_aXvec_27__full_n = fifo_aXvec_27_if_full_n;
  assign fifo_aXvec_27_if_read = fifo_aXvec_27__read;
  assign fifo_aXvec_27_if_read_ce = 1'b1;
  assign fifo_aXvec_27_if_write = fifo_aXvec_27__write;
  assign fifo_aXvec_27_if_write_ce = 1'b1;
  assign fifo_aXvec_27_reset = ~ ap_rst_n;
  assign fifo_aXvec_28_clk = ap_clk;
  assign fifo_aXvec_28_if_din = fifo_aXvec_28__din;
  assign fifo_aXvec_28__dout = fifo_aXvec_28_if_dout;
  assign fifo_aXvec_28__empty_n = fifo_aXvec_28_if_empty_n;
  assign fifo_aXvec_28__full_n = fifo_aXvec_28_if_full_n;
  assign fifo_aXvec_28_if_read = fifo_aXvec_28__read;
  assign fifo_aXvec_28_if_read_ce = 1'b1;
  assign fifo_aXvec_28_if_write = fifo_aXvec_28__write;
  assign fifo_aXvec_28_if_write_ce = 1'b1;
  assign fifo_aXvec_28_reset = ~ ap_rst_n;
  assign fifo_aXvec_29_clk = ap_clk;
  assign fifo_aXvec_29_if_din = fifo_aXvec_29__din;
  assign fifo_aXvec_29__dout = fifo_aXvec_29_if_dout;
  assign fifo_aXvec_29__empty_n = fifo_aXvec_29_if_empty_n;
  assign fifo_aXvec_29__full_n = fifo_aXvec_29_if_full_n;
  assign fifo_aXvec_29_if_read = fifo_aXvec_29__read;
  assign fifo_aXvec_29_if_read_ce = 1'b1;
  assign fifo_aXvec_29_if_write = fifo_aXvec_29__write;
  assign fifo_aXvec_29_if_write_ce = 1'b1;
  assign fifo_aXvec_29_reset = ~ ap_rst_n;
  assign fifo_aXvec_2_clk = ap_clk;
  assign fifo_aXvec_2_if_din = fifo_aXvec_2__din;
  assign fifo_aXvec_2__dout = fifo_aXvec_2_if_dout;
  assign fifo_aXvec_2__empty_n = fifo_aXvec_2_if_empty_n;
  assign fifo_aXvec_2__full_n = fifo_aXvec_2_if_full_n;
  assign fifo_aXvec_2_if_read = fifo_aXvec_2__read;
  assign fifo_aXvec_2_if_read_ce = 1'b1;
  assign fifo_aXvec_2_if_write = fifo_aXvec_2__write;
  assign fifo_aXvec_2_if_write_ce = 1'b1;
  assign fifo_aXvec_2_reset = ~ ap_rst_n;
  assign fifo_aXvec_30_clk = ap_clk;
  assign fifo_aXvec_30_if_din = fifo_aXvec_30__din;
  assign fifo_aXvec_30__dout = fifo_aXvec_30_if_dout;
  assign fifo_aXvec_30__empty_n = fifo_aXvec_30_if_empty_n;
  assign fifo_aXvec_30__full_n = fifo_aXvec_30_if_full_n;
  assign fifo_aXvec_30_if_read = fifo_aXvec_30__read;
  assign fifo_aXvec_30_if_read_ce = 1'b1;
  assign fifo_aXvec_30_if_write = fifo_aXvec_30__write;
  assign fifo_aXvec_30_if_write_ce = 1'b1;
  assign fifo_aXvec_30_reset = ~ ap_rst_n;
  assign fifo_aXvec_31_clk = ap_clk;
  assign fifo_aXvec_31_if_din = fifo_aXvec_31__din;
  assign fifo_aXvec_31__dout = fifo_aXvec_31_if_dout;
  assign fifo_aXvec_31__empty_n = fifo_aXvec_31_if_empty_n;
  assign fifo_aXvec_31__full_n = fifo_aXvec_31_if_full_n;
  assign fifo_aXvec_31_if_read = fifo_aXvec_31__read;
  assign fifo_aXvec_31_if_read_ce = 1'b1;
  assign fifo_aXvec_31_if_write = fifo_aXvec_31__write;
  assign fifo_aXvec_31_if_write_ce = 1'b1;
  assign fifo_aXvec_31_reset = ~ ap_rst_n;
  assign fifo_aXvec_32_clk = ap_clk;
  assign fifo_aXvec_32_if_din = fifo_aXvec_32__din;
  assign fifo_aXvec_32__dout = fifo_aXvec_32_if_dout;
  assign fifo_aXvec_32__empty_n = fifo_aXvec_32_if_empty_n;
  assign fifo_aXvec_32__full_n = fifo_aXvec_32_if_full_n;
  assign fifo_aXvec_32_if_read = fifo_aXvec_32__read;
  assign fifo_aXvec_32_if_read_ce = 1'b1;
  assign fifo_aXvec_32_if_write = fifo_aXvec_32__write;
  assign fifo_aXvec_32_if_write_ce = 1'b1;
  assign fifo_aXvec_32_reset = ~ ap_rst_n;
  assign fifo_aXvec_33_clk = ap_clk;
  assign fifo_aXvec_33_if_din = fifo_aXvec_33__din;
  assign fifo_aXvec_33__dout = fifo_aXvec_33_if_dout;
  assign fifo_aXvec_33__empty_n = fifo_aXvec_33_if_empty_n;
  assign fifo_aXvec_33__full_n = fifo_aXvec_33_if_full_n;
  assign fifo_aXvec_33_if_read = fifo_aXvec_33__read;
  assign fifo_aXvec_33_if_read_ce = 1'b1;
  assign fifo_aXvec_33_if_write = fifo_aXvec_33__write;
  assign fifo_aXvec_33_if_write_ce = 1'b1;
  assign fifo_aXvec_33_reset = ~ ap_rst_n;
  assign fifo_aXvec_34_clk = ap_clk;
  assign fifo_aXvec_34_if_din = fifo_aXvec_34__din;
  assign fifo_aXvec_34__dout = fifo_aXvec_34_if_dout;
  assign fifo_aXvec_34__empty_n = fifo_aXvec_34_if_empty_n;
  assign fifo_aXvec_34__full_n = fifo_aXvec_34_if_full_n;
  assign fifo_aXvec_34_if_read = fifo_aXvec_34__read;
  assign fifo_aXvec_34_if_read_ce = 1'b1;
  assign fifo_aXvec_34_if_write = fifo_aXvec_34__write;
  assign fifo_aXvec_34_if_write_ce = 1'b1;
  assign fifo_aXvec_34_reset = ~ ap_rst_n;
  assign fifo_aXvec_35_clk = ap_clk;
  assign fifo_aXvec_35_if_din = fifo_aXvec_35__din;
  assign fifo_aXvec_35__dout = fifo_aXvec_35_if_dout;
  assign fifo_aXvec_35__empty_n = fifo_aXvec_35_if_empty_n;
  assign fifo_aXvec_35__full_n = fifo_aXvec_35_if_full_n;
  assign fifo_aXvec_35_if_read = fifo_aXvec_35__read;
  assign fifo_aXvec_35_if_read_ce = 1'b1;
  assign fifo_aXvec_35_if_write = fifo_aXvec_35__write;
  assign fifo_aXvec_35_if_write_ce = 1'b1;
  assign fifo_aXvec_35_reset = ~ ap_rst_n;
  assign fifo_aXvec_36_clk = ap_clk;
  assign fifo_aXvec_36_if_din = fifo_aXvec_36__din;
  assign fifo_aXvec_36__dout = fifo_aXvec_36_if_dout;
  assign fifo_aXvec_36__empty_n = fifo_aXvec_36_if_empty_n;
  assign fifo_aXvec_36__full_n = fifo_aXvec_36_if_full_n;
  assign fifo_aXvec_36_if_read = fifo_aXvec_36__read;
  assign fifo_aXvec_36_if_read_ce = 1'b1;
  assign fifo_aXvec_36_if_write = fifo_aXvec_36__write;
  assign fifo_aXvec_36_if_write_ce = 1'b1;
  assign fifo_aXvec_36_reset = ~ ap_rst_n;
  assign fifo_aXvec_37_clk = ap_clk;
  assign fifo_aXvec_37_if_din = fifo_aXvec_37__din;
  assign fifo_aXvec_37__dout = fifo_aXvec_37_if_dout;
  assign fifo_aXvec_37__empty_n = fifo_aXvec_37_if_empty_n;
  assign fifo_aXvec_37__full_n = fifo_aXvec_37_if_full_n;
  assign fifo_aXvec_37_if_read = fifo_aXvec_37__read;
  assign fifo_aXvec_37_if_read_ce = 1'b1;
  assign fifo_aXvec_37_if_write = fifo_aXvec_37__write;
  assign fifo_aXvec_37_if_write_ce = 1'b1;
  assign fifo_aXvec_37_reset = ~ ap_rst_n;
  assign fifo_aXvec_38_clk = ap_clk;
  assign fifo_aXvec_38_if_din = fifo_aXvec_38__din;
  assign fifo_aXvec_38__dout = fifo_aXvec_38_if_dout;
  assign fifo_aXvec_38__empty_n = fifo_aXvec_38_if_empty_n;
  assign fifo_aXvec_38__full_n = fifo_aXvec_38_if_full_n;
  assign fifo_aXvec_38_if_read = fifo_aXvec_38__read;
  assign fifo_aXvec_38_if_read_ce = 1'b1;
  assign fifo_aXvec_38_if_write = fifo_aXvec_38__write;
  assign fifo_aXvec_38_if_write_ce = 1'b1;
  assign fifo_aXvec_38_reset = ~ ap_rst_n;
  assign fifo_aXvec_39_clk = ap_clk;
  assign fifo_aXvec_39_if_din = fifo_aXvec_39__din;
  assign fifo_aXvec_39__dout = fifo_aXvec_39_if_dout;
  assign fifo_aXvec_39__empty_n = fifo_aXvec_39_if_empty_n;
  assign fifo_aXvec_39__full_n = fifo_aXvec_39_if_full_n;
  assign fifo_aXvec_39_if_read = fifo_aXvec_39__read;
  assign fifo_aXvec_39_if_read_ce = 1'b1;
  assign fifo_aXvec_39_if_write = fifo_aXvec_39__write;
  assign fifo_aXvec_39_if_write_ce = 1'b1;
  assign fifo_aXvec_39_reset = ~ ap_rst_n;
  assign fifo_aXvec_3_clk = ap_clk;
  assign fifo_aXvec_3_if_din = fifo_aXvec_3__din;
  assign fifo_aXvec_3__dout = fifo_aXvec_3_if_dout;
  assign fifo_aXvec_3__empty_n = fifo_aXvec_3_if_empty_n;
  assign fifo_aXvec_3__full_n = fifo_aXvec_3_if_full_n;
  assign fifo_aXvec_3_if_read = fifo_aXvec_3__read;
  assign fifo_aXvec_3_if_read_ce = 1'b1;
  assign fifo_aXvec_3_if_write = fifo_aXvec_3__write;
  assign fifo_aXvec_3_if_write_ce = 1'b1;
  assign fifo_aXvec_3_reset = ~ ap_rst_n;
  assign fifo_aXvec_40_clk = ap_clk;
  assign fifo_aXvec_40_if_din = fifo_aXvec_40__din;
  assign fifo_aXvec_40__dout = fifo_aXvec_40_if_dout;
  assign fifo_aXvec_40__empty_n = fifo_aXvec_40_if_empty_n;
  assign fifo_aXvec_40__full_n = fifo_aXvec_40_if_full_n;
  assign fifo_aXvec_40_if_read = fifo_aXvec_40__read;
  assign fifo_aXvec_40_if_read_ce = 1'b1;
  assign fifo_aXvec_40_if_write = fifo_aXvec_40__write;
  assign fifo_aXvec_40_if_write_ce = 1'b1;
  assign fifo_aXvec_40_reset = ~ ap_rst_n;
  assign fifo_aXvec_41_clk = ap_clk;
  assign fifo_aXvec_41_if_din = fifo_aXvec_41__din;
  assign fifo_aXvec_41__dout = fifo_aXvec_41_if_dout;
  assign fifo_aXvec_41__empty_n = fifo_aXvec_41_if_empty_n;
  assign fifo_aXvec_41__full_n = fifo_aXvec_41_if_full_n;
  assign fifo_aXvec_41_if_read = fifo_aXvec_41__read;
  assign fifo_aXvec_41_if_read_ce = 1'b1;
  assign fifo_aXvec_41_if_write = fifo_aXvec_41__write;
  assign fifo_aXvec_41_if_write_ce = 1'b1;
  assign fifo_aXvec_41_reset = ~ ap_rst_n;
  assign fifo_aXvec_42_clk = ap_clk;
  assign fifo_aXvec_42_if_din = fifo_aXvec_42__din;
  assign fifo_aXvec_42__dout = fifo_aXvec_42_if_dout;
  assign fifo_aXvec_42__empty_n = fifo_aXvec_42_if_empty_n;
  assign fifo_aXvec_42__full_n = fifo_aXvec_42_if_full_n;
  assign fifo_aXvec_42_if_read = fifo_aXvec_42__read;
  assign fifo_aXvec_42_if_read_ce = 1'b1;
  assign fifo_aXvec_42_if_write = fifo_aXvec_42__write;
  assign fifo_aXvec_42_if_write_ce = 1'b1;
  assign fifo_aXvec_42_reset = ~ ap_rst_n;
  assign fifo_aXvec_43_clk = ap_clk;
  assign fifo_aXvec_43_if_din = fifo_aXvec_43__din;
  assign fifo_aXvec_43__dout = fifo_aXvec_43_if_dout;
  assign fifo_aXvec_43__empty_n = fifo_aXvec_43_if_empty_n;
  assign fifo_aXvec_43__full_n = fifo_aXvec_43_if_full_n;
  assign fifo_aXvec_43_if_read = fifo_aXvec_43__read;
  assign fifo_aXvec_43_if_read_ce = 1'b1;
  assign fifo_aXvec_43_if_write = fifo_aXvec_43__write;
  assign fifo_aXvec_43_if_write_ce = 1'b1;
  assign fifo_aXvec_43_reset = ~ ap_rst_n;
  assign fifo_aXvec_44_clk = ap_clk;
  assign fifo_aXvec_44_if_din = fifo_aXvec_44__din;
  assign fifo_aXvec_44__dout = fifo_aXvec_44_if_dout;
  assign fifo_aXvec_44__empty_n = fifo_aXvec_44_if_empty_n;
  assign fifo_aXvec_44__full_n = fifo_aXvec_44_if_full_n;
  assign fifo_aXvec_44_if_read = fifo_aXvec_44__read;
  assign fifo_aXvec_44_if_read_ce = 1'b1;
  assign fifo_aXvec_44_if_write = fifo_aXvec_44__write;
  assign fifo_aXvec_44_if_write_ce = 1'b1;
  assign fifo_aXvec_44_reset = ~ ap_rst_n;
  assign fifo_aXvec_45_clk = ap_clk;
  assign fifo_aXvec_45_if_din = fifo_aXvec_45__din;
  assign fifo_aXvec_45__dout = fifo_aXvec_45_if_dout;
  assign fifo_aXvec_45__empty_n = fifo_aXvec_45_if_empty_n;
  assign fifo_aXvec_45__full_n = fifo_aXvec_45_if_full_n;
  assign fifo_aXvec_45_if_read = fifo_aXvec_45__read;
  assign fifo_aXvec_45_if_read_ce = 1'b1;
  assign fifo_aXvec_45_if_write = fifo_aXvec_45__write;
  assign fifo_aXvec_45_if_write_ce = 1'b1;
  assign fifo_aXvec_45_reset = ~ ap_rst_n;
  assign fifo_aXvec_46_clk = ap_clk;
  assign fifo_aXvec_46_if_din = fifo_aXvec_46__din;
  assign fifo_aXvec_46__dout = fifo_aXvec_46_if_dout;
  assign fifo_aXvec_46__empty_n = fifo_aXvec_46_if_empty_n;
  assign fifo_aXvec_46__full_n = fifo_aXvec_46_if_full_n;
  assign fifo_aXvec_46_if_read = fifo_aXvec_46__read;
  assign fifo_aXvec_46_if_read_ce = 1'b1;
  assign fifo_aXvec_46_if_write = fifo_aXvec_46__write;
  assign fifo_aXvec_46_if_write_ce = 1'b1;
  assign fifo_aXvec_46_reset = ~ ap_rst_n;
  assign fifo_aXvec_47_clk = ap_clk;
  assign fifo_aXvec_47_if_din = fifo_aXvec_47__din;
  assign fifo_aXvec_47__dout = fifo_aXvec_47_if_dout;
  assign fifo_aXvec_47__empty_n = fifo_aXvec_47_if_empty_n;
  assign fifo_aXvec_47__full_n = fifo_aXvec_47_if_full_n;
  assign fifo_aXvec_47_if_read = fifo_aXvec_47__read;
  assign fifo_aXvec_47_if_read_ce = 1'b1;
  assign fifo_aXvec_47_if_write = fifo_aXvec_47__write;
  assign fifo_aXvec_47_if_write_ce = 1'b1;
  assign fifo_aXvec_47_reset = ~ ap_rst_n;
  assign fifo_aXvec_4_clk = ap_clk;
  assign fifo_aXvec_4_if_din = fifo_aXvec_4__din;
  assign fifo_aXvec_4__dout = fifo_aXvec_4_if_dout;
  assign fifo_aXvec_4__empty_n = fifo_aXvec_4_if_empty_n;
  assign fifo_aXvec_4__full_n = fifo_aXvec_4_if_full_n;
  assign fifo_aXvec_4_if_read = fifo_aXvec_4__read;
  assign fifo_aXvec_4_if_read_ce = 1'b1;
  assign fifo_aXvec_4_if_write = fifo_aXvec_4__write;
  assign fifo_aXvec_4_if_write_ce = 1'b1;
  assign fifo_aXvec_4_reset = ~ ap_rst_n;
  assign fifo_aXvec_5_clk = ap_clk;
  assign fifo_aXvec_5_if_din = fifo_aXvec_5__din;
  assign fifo_aXvec_5__dout = fifo_aXvec_5_if_dout;
  assign fifo_aXvec_5__empty_n = fifo_aXvec_5_if_empty_n;
  assign fifo_aXvec_5__full_n = fifo_aXvec_5_if_full_n;
  assign fifo_aXvec_5_if_read = fifo_aXvec_5__read;
  assign fifo_aXvec_5_if_read_ce = 1'b1;
  assign fifo_aXvec_5_if_write = fifo_aXvec_5__write;
  assign fifo_aXvec_5_if_write_ce = 1'b1;
  assign fifo_aXvec_5_reset = ~ ap_rst_n;
  assign fifo_aXvec_6_clk = ap_clk;
  assign fifo_aXvec_6_if_din = fifo_aXvec_6__din;
  assign fifo_aXvec_6__dout = fifo_aXvec_6_if_dout;
  assign fifo_aXvec_6__empty_n = fifo_aXvec_6_if_empty_n;
  assign fifo_aXvec_6__full_n = fifo_aXvec_6_if_full_n;
  assign fifo_aXvec_6_if_read = fifo_aXvec_6__read;
  assign fifo_aXvec_6_if_read_ce = 1'b1;
  assign fifo_aXvec_6_if_write = fifo_aXvec_6__write;
  assign fifo_aXvec_6_if_write_ce = 1'b1;
  assign fifo_aXvec_6_reset = ~ ap_rst_n;
  assign fifo_aXvec_7_clk = ap_clk;
  assign fifo_aXvec_7_if_din = fifo_aXvec_7__din;
  assign fifo_aXvec_7__dout = fifo_aXvec_7_if_dout;
  assign fifo_aXvec_7__empty_n = fifo_aXvec_7_if_empty_n;
  assign fifo_aXvec_7__full_n = fifo_aXvec_7_if_full_n;
  assign fifo_aXvec_7_if_read = fifo_aXvec_7__read;
  assign fifo_aXvec_7_if_read_ce = 1'b1;
  assign fifo_aXvec_7_if_write = fifo_aXvec_7__write;
  assign fifo_aXvec_7_if_write_ce = 1'b1;
  assign fifo_aXvec_7_reset = ~ ap_rst_n;
  assign fifo_aXvec_8_clk = ap_clk;
  assign fifo_aXvec_8_if_din = fifo_aXvec_8__din;
  assign fifo_aXvec_8__dout = fifo_aXvec_8_if_dout;
  assign fifo_aXvec_8__empty_n = fifo_aXvec_8_if_empty_n;
  assign fifo_aXvec_8__full_n = fifo_aXvec_8_if_full_n;
  assign fifo_aXvec_8_if_read = fifo_aXvec_8__read;
  assign fifo_aXvec_8_if_read_ce = 1'b1;
  assign fifo_aXvec_8_if_write = fifo_aXvec_8__write;
  assign fifo_aXvec_8_if_write_ce = 1'b1;
  assign fifo_aXvec_8_reset = ~ ap_rst_n;
  assign fifo_aXvec_9_clk = ap_clk;
  assign fifo_aXvec_9_if_din = fifo_aXvec_9__din;
  assign fifo_aXvec_9__dout = fifo_aXvec_9_if_dout;
  assign fifo_aXvec_9__empty_n = fifo_aXvec_9_if_empty_n;
  assign fifo_aXvec_9__full_n = fifo_aXvec_9_if_full_n;
  assign fifo_aXvec_9_if_read = fifo_aXvec_9__read;
  assign fifo_aXvec_9_if_read_ce = 1'b1;
  assign fifo_aXvec_9_if_write = fifo_aXvec_9__write;
  assign fifo_aXvec_9_if_write_ce = 1'b1;
  assign fifo_aXvec_9_reset = ~ ap_rst_n;
  assign Arbiter_Y_0_M = Arbiter_Y_0___M__q0;
  assign Arbiter_Y_0_P_N = Arbiter_Y_0___P_N__q0;
  assign Arbiter_Y_0_ap_clk = ap_clk;
  assign Arbiter_Y_0__ap_done = Arbiter_Y_0_ap_done;
  assign Arbiter_Y_0__ap_idle = Arbiter_Y_0_ap_idle;
  assign Arbiter_Y_0__ap_ready = Arbiter_Y_0_ap_ready;
  assign Arbiter_Y_0_ap_rst_n = ap_rst_n;
  assign Arbiter_Y_0_ap_start = Arbiter_Y_0__ap_start;
  assign Arbiter_Y_0_fifo_in_0_dout = fifo_Y_pe_0__dout;
  assign Arbiter_Y_0_fifo_in_0_empty_n = fifo_Y_pe_0__empty_n;
  assign fifo_Y_pe_0__read = Arbiter_Y_0_fifo_in_0_read;
  assign Arbiter_Y_0_fifo_in_1_dout = fifo_Y_pe_1__dout;
  assign Arbiter_Y_0_fifo_in_1_empty_n = fifo_Y_pe_1__empty_n;
  assign fifo_Y_pe_1__read = Arbiter_Y_0_fifo_in_1_read;
  assign Arbiter_Y_0_fifo_in_2_dout = fifo_Y_pe_2__dout;
  assign Arbiter_Y_0_fifo_in_2_empty_n = fifo_Y_pe_2__empty_n;
  assign fifo_Y_pe_2__read = Arbiter_Y_0_fifo_in_2_read;
  assign Arbiter_Y_0_fifo_in_3_dout = fifo_Y_pe_3__dout;
  assign Arbiter_Y_0_fifo_in_3_empty_n = fifo_Y_pe_3__empty_n;
  assign fifo_Y_pe_3__read = Arbiter_Y_0_fifo_in_3_read;
  assign Arbiter_Y_0_fifo_in_4_dout = fifo_Y_pe_4__dout;
  assign Arbiter_Y_0_fifo_in_4_empty_n = fifo_Y_pe_4__empty_n;
  assign fifo_Y_pe_4__read = Arbiter_Y_0_fifo_in_4_read;
  assign Arbiter_Y_0_fifo_in_5_dout = fifo_Y_pe_5__dout;
  assign Arbiter_Y_0_fifo_in_5_empty_n = fifo_Y_pe_5__empty_n;
  assign fifo_Y_pe_5__read = Arbiter_Y_0_fifo_in_5_read;
  assign Arbiter_Y_0_fifo_in_peek_0_dout = fifo_Y_pe_0__dout;
  assign Arbiter_Y_0_fifo_in_peek_0_empty_n = fifo_Y_pe_0__empty_n;
  assign Arbiter_Y_0_fifo_in_peek_1_dout = fifo_Y_pe_1__dout;
  assign Arbiter_Y_0_fifo_in_peek_1_empty_n = fifo_Y_pe_1__empty_n;
  assign Arbiter_Y_0_fifo_in_peek_2_dout = fifo_Y_pe_2__dout;
  assign Arbiter_Y_0_fifo_in_peek_2_empty_n = fifo_Y_pe_2__empty_n;
  assign Arbiter_Y_0_fifo_in_peek_3_dout = fifo_Y_pe_3__dout;
  assign Arbiter_Y_0_fifo_in_peek_3_empty_n = fifo_Y_pe_3__empty_n;
  assign Arbiter_Y_0_fifo_in_peek_4_dout = fifo_Y_pe_4__dout;
  assign Arbiter_Y_0_fifo_in_peek_4_empty_n = fifo_Y_pe_4__empty_n;
  assign Arbiter_Y_0_fifo_in_peek_5_dout = fifo_Y_pe_5__dout;
  assign Arbiter_Y_0_fifo_in_peek_5_empty_n = fifo_Y_pe_5__empty_n;
  assign fifo_Y_pe_abd_0__din = Arbiter_Y_0_fifo_out_din;
  assign Arbiter_Y_0_fifo_out_full_n = fifo_Y_pe_abd_0__full_n;
  assign fifo_Y_pe_abd_0__write = Arbiter_Y_0_fifo_out_write;
  assign Arbiter_Y_1_M = Arbiter_Y_1___M__q0;
  assign Arbiter_Y_1_P_N = Arbiter_Y_1___P_N__q0;
  assign Arbiter_Y_1_ap_clk = ap_clk;
  assign Arbiter_Y_1__ap_done = Arbiter_Y_1_ap_done;
  assign Arbiter_Y_1__ap_idle = Arbiter_Y_1_ap_idle;
  assign Arbiter_Y_1__ap_ready = Arbiter_Y_1_ap_ready;
  assign Arbiter_Y_1_ap_rst_n = ap_rst_n;
  assign Arbiter_Y_1_ap_start = Arbiter_Y_1__ap_start;
  assign Arbiter_Y_1_fifo_in_0_dout = fifo_Y_pe_6__dout;
  assign Arbiter_Y_1_fifo_in_0_empty_n = fifo_Y_pe_6__empty_n;
  assign fifo_Y_pe_6__read = Arbiter_Y_1_fifo_in_0_read;
  assign Arbiter_Y_1_fifo_in_1_dout = fifo_Y_pe_7__dout;
  assign Arbiter_Y_1_fifo_in_1_empty_n = fifo_Y_pe_7__empty_n;
  assign fifo_Y_pe_7__read = Arbiter_Y_1_fifo_in_1_read;
  assign Arbiter_Y_1_fifo_in_2_dout = fifo_Y_pe_8__dout;
  assign Arbiter_Y_1_fifo_in_2_empty_n = fifo_Y_pe_8__empty_n;
  assign fifo_Y_pe_8__read = Arbiter_Y_1_fifo_in_2_read;
  assign Arbiter_Y_1_fifo_in_3_dout = fifo_Y_pe_9__dout;
  assign Arbiter_Y_1_fifo_in_3_empty_n = fifo_Y_pe_9__empty_n;
  assign fifo_Y_pe_9__read = Arbiter_Y_1_fifo_in_3_read;
  assign Arbiter_Y_1_fifo_in_4_dout = fifo_Y_pe_10__dout;
  assign Arbiter_Y_1_fifo_in_4_empty_n = fifo_Y_pe_10__empty_n;
  assign fifo_Y_pe_10__read = Arbiter_Y_1_fifo_in_4_read;
  assign Arbiter_Y_1_fifo_in_5_dout = fifo_Y_pe_11__dout;
  assign Arbiter_Y_1_fifo_in_5_empty_n = fifo_Y_pe_11__empty_n;
  assign fifo_Y_pe_11__read = Arbiter_Y_1_fifo_in_5_read;
  assign Arbiter_Y_1_fifo_in_peek_0_dout = fifo_Y_pe_6__dout;
  assign Arbiter_Y_1_fifo_in_peek_0_empty_n = fifo_Y_pe_6__empty_n;
  assign Arbiter_Y_1_fifo_in_peek_1_dout = fifo_Y_pe_7__dout;
  assign Arbiter_Y_1_fifo_in_peek_1_empty_n = fifo_Y_pe_7__empty_n;
  assign Arbiter_Y_1_fifo_in_peek_2_dout = fifo_Y_pe_8__dout;
  assign Arbiter_Y_1_fifo_in_peek_2_empty_n = fifo_Y_pe_8__empty_n;
  assign Arbiter_Y_1_fifo_in_peek_3_dout = fifo_Y_pe_9__dout;
  assign Arbiter_Y_1_fifo_in_peek_3_empty_n = fifo_Y_pe_9__empty_n;
  assign Arbiter_Y_1_fifo_in_peek_4_dout = fifo_Y_pe_10__dout;
  assign Arbiter_Y_1_fifo_in_peek_4_empty_n = fifo_Y_pe_10__empty_n;
  assign Arbiter_Y_1_fifo_in_peek_5_dout = fifo_Y_pe_11__dout;
  assign Arbiter_Y_1_fifo_in_peek_5_empty_n = fifo_Y_pe_11__empty_n;
  assign fifo_Y_pe_abd_1__din = Arbiter_Y_1_fifo_out_din;
  assign Arbiter_Y_1_fifo_out_full_n = fifo_Y_pe_abd_1__full_n;
  assign fifo_Y_pe_abd_1__write = Arbiter_Y_1_fifo_out_write;
  assign Arbiter_Y_2_M = Arbiter_Y_2___M__q0;
  assign Arbiter_Y_2_P_N = Arbiter_Y_2___P_N__q0;
  assign Arbiter_Y_2_ap_clk = ap_clk;
  assign Arbiter_Y_2__ap_done = Arbiter_Y_2_ap_done;
  assign Arbiter_Y_2__ap_idle = Arbiter_Y_2_ap_idle;
  assign Arbiter_Y_2__ap_ready = Arbiter_Y_2_ap_ready;
  assign Arbiter_Y_2_ap_rst_n = ap_rst_n;
  assign Arbiter_Y_2_ap_start = Arbiter_Y_2__ap_start;
  assign Arbiter_Y_2_fifo_in_0_dout = fifo_Y_pe_12__dout;
  assign Arbiter_Y_2_fifo_in_0_empty_n = fifo_Y_pe_12__empty_n;
  assign fifo_Y_pe_12__read = Arbiter_Y_2_fifo_in_0_read;
  assign Arbiter_Y_2_fifo_in_1_dout = fifo_Y_pe_13__dout;
  assign Arbiter_Y_2_fifo_in_1_empty_n = fifo_Y_pe_13__empty_n;
  assign fifo_Y_pe_13__read = Arbiter_Y_2_fifo_in_1_read;
  assign Arbiter_Y_2_fifo_in_2_dout = fifo_Y_pe_14__dout;
  assign Arbiter_Y_2_fifo_in_2_empty_n = fifo_Y_pe_14__empty_n;
  assign fifo_Y_pe_14__read = Arbiter_Y_2_fifo_in_2_read;
  assign Arbiter_Y_2_fifo_in_3_dout = fifo_Y_pe_15__dout;
  assign Arbiter_Y_2_fifo_in_3_empty_n = fifo_Y_pe_15__empty_n;
  assign fifo_Y_pe_15__read = Arbiter_Y_2_fifo_in_3_read;
  assign Arbiter_Y_2_fifo_in_4_dout = fifo_Y_pe_16__dout;
  assign Arbiter_Y_2_fifo_in_4_empty_n = fifo_Y_pe_16__empty_n;
  assign fifo_Y_pe_16__read = Arbiter_Y_2_fifo_in_4_read;
  assign Arbiter_Y_2_fifo_in_5_dout = fifo_Y_pe_17__dout;
  assign Arbiter_Y_2_fifo_in_5_empty_n = fifo_Y_pe_17__empty_n;
  assign fifo_Y_pe_17__read = Arbiter_Y_2_fifo_in_5_read;
  assign Arbiter_Y_2_fifo_in_peek_0_dout = fifo_Y_pe_12__dout;
  assign Arbiter_Y_2_fifo_in_peek_0_empty_n = fifo_Y_pe_12__empty_n;
  assign Arbiter_Y_2_fifo_in_peek_1_dout = fifo_Y_pe_13__dout;
  assign Arbiter_Y_2_fifo_in_peek_1_empty_n = fifo_Y_pe_13__empty_n;
  assign Arbiter_Y_2_fifo_in_peek_2_dout = fifo_Y_pe_14__dout;
  assign Arbiter_Y_2_fifo_in_peek_2_empty_n = fifo_Y_pe_14__empty_n;
  assign Arbiter_Y_2_fifo_in_peek_3_dout = fifo_Y_pe_15__dout;
  assign Arbiter_Y_2_fifo_in_peek_3_empty_n = fifo_Y_pe_15__empty_n;
  assign Arbiter_Y_2_fifo_in_peek_4_dout = fifo_Y_pe_16__dout;
  assign Arbiter_Y_2_fifo_in_peek_4_empty_n = fifo_Y_pe_16__empty_n;
  assign Arbiter_Y_2_fifo_in_peek_5_dout = fifo_Y_pe_17__dout;
  assign Arbiter_Y_2_fifo_in_peek_5_empty_n = fifo_Y_pe_17__empty_n;
  assign fifo_Y_pe_abd_2__din = Arbiter_Y_2_fifo_out_din;
  assign Arbiter_Y_2_fifo_out_full_n = fifo_Y_pe_abd_2__full_n;
  assign fifo_Y_pe_abd_2__write = Arbiter_Y_2_fifo_out_write;
  assign Arbiter_Y_3_M = Arbiter_Y_3___M__q0;
  assign Arbiter_Y_3_P_N = Arbiter_Y_3___P_N__q0;
  assign Arbiter_Y_3_ap_clk = ap_clk;
  assign Arbiter_Y_3__ap_done = Arbiter_Y_3_ap_done;
  assign Arbiter_Y_3__ap_idle = Arbiter_Y_3_ap_idle;
  assign Arbiter_Y_3__ap_ready = Arbiter_Y_3_ap_ready;
  assign Arbiter_Y_3_ap_rst_n = ap_rst_n;
  assign Arbiter_Y_3_ap_start = Arbiter_Y_3__ap_start;
  assign Arbiter_Y_3_fifo_in_0_dout = fifo_Y_pe_18__dout;
  assign Arbiter_Y_3_fifo_in_0_empty_n = fifo_Y_pe_18__empty_n;
  assign fifo_Y_pe_18__read = Arbiter_Y_3_fifo_in_0_read;
  assign Arbiter_Y_3_fifo_in_1_dout = fifo_Y_pe_19__dout;
  assign Arbiter_Y_3_fifo_in_1_empty_n = fifo_Y_pe_19__empty_n;
  assign fifo_Y_pe_19__read = Arbiter_Y_3_fifo_in_1_read;
  assign Arbiter_Y_3_fifo_in_2_dout = fifo_Y_pe_20__dout;
  assign Arbiter_Y_3_fifo_in_2_empty_n = fifo_Y_pe_20__empty_n;
  assign fifo_Y_pe_20__read = Arbiter_Y_3_fifo_in_2_read;
  assign Arbiter_Y_3_fifo_in_3_dout = fifo_Y_pe_21__dout;
  assign Arbiter_Y_3_fifo_in_3_empty_n = fifo_Y_pe_21__empty_n;
  assign fifo_Y_pe_21__read = Arbiter_Y_3_fifo_in_3_read;
  assign Arbiter_Y_3_fifo_in_4_dout = fifo_Y_pe_22__dout;
  assign Arbiter_Y_3_fifo_in_4_empty_n = fifo_Y_pe_22__empty_n;
  assign fifo_Y_pe_22__read = Arbiter_Y_3_fifo_in_4_read;
  assign Arbiter_Y_3_fifo_in_5_dout = fifo_Y_pe_23__dout;
  assign Arbiter_Y_3_fifo_in_5_empty_n = fifo_Y_pe_23__empty_n;
  assign fifo_Y_pe_23__read = Arbiter_Y_3_fifo_in_5_read;
  assign Arbiter_Y_3_fifo_in_peek_0_dout = fifo_Y_pe_18__dout;
  assign Arbiter_Y_3_fifo_in_peek_0_empty_n = fifo_Y_pe_18__empty_n;
  assign Arbiter_Y_3_fifo_in_peek_1_dout = fifo_Y_pe_19__dout;
  assign Arbiter_Y_3_fifo_in_peek_1_empty_n = fifo_Y_pe_19__empty_n;
  assign Arbiter_Y_3_fifo_in_peek_2_dout = fifo_Y_pe_20__dout;
  assign Arbiter_Y_3_fifo_in_peek_2_empty_n = fifo_Y_pe_20__empty_n;
  assign Arbiter_Y_3_fifo_in_peek_3_dout = fifo_Y_pe_21__dout;
  assign Arbiter_Y_3_fifo_in_peek_3_empty_n = fifo_Y_pe_21__empty_n;
  assign Arbiter_Y_3_fifo_in_peek_4_dout = fifo_Y_pe_22__dout;
  assign Arbiter_Y_3_fifo_in_peek_4_empty_n = fifo_Y_pe_22__empty_n;
  assign Arbiter_Y_3_fifo_in_peek_5_dout = fifo_Y_pe_23__dout;
  assign Arbiter_Y_3_fifo_in_peek_5_empty_n = fifo_Y_pe_23__empty_n;
  assign fifo_Y_pe_abd_3__din = Arbiter_Y_3_fifo_out_din;
  assign Arbiter_Y_3_fifo_out_full_n = fifo_Y_pe_abd_3__full_n;
  assign fifo_Y_pe_abd_3__write = Arbiter_Y_3_fifo_out_write;
  assign Arbiter_Y_4_M = Arbiter_Y_4___M__q0;
  assign Arbiter_Y_4_P_N = Arbiter_Y_4___P_N__q0;
  assign Arbiter_Y_4_ap_clk = ap_clk;
  assign Arbiter_Y_4__ap_done = Arbiter_Y_4_ap_done;
  assign Arbiter_Y_4__ap_idle = Arbiter_Y_4_ap_idle;
  assign Arbiter_Y_4__ap_ready = Arbiter_Y_4_ap_ready;
  assign Arbiter_Y_4_ap_rst_n = ap_rst_n;
  assign Arbiter_Y_4_ap_start = Arbiter_Y_4__ap_start;
  assign Arbiter_Y_4_fifo_in_0_dout = fifo_Y_pe_24__dout;
  assign Arbiter_Y_4_fifo_in_0_empty_n = fifo_Y_pe_24__empty_n;
  assign fifo_Y_pe_24__read = Arbiter_Y_4_fifo_in_0_read;
  assign Arbiter_Y_4_fifo_in_1_dout = fifo_Y_pe_25__dout;
  assign Arbiter_Y_4_fifo_in_1_empty_n = fifo_Y_pe_25__empty_n;
  assign fifo_Y_pe_25__read = Arbiter_Y_4_fifo_in_1_read;
  assign Arbiter_Y_4_fifo_in_2_dout = fifo_Y_pe_26__dout;
  assign Arbiter_Y_4_fifo_in_2_empty_n = fifo_Y_pe_26__empty_n;
  assign fifo_Y_pe_26__read = Arbiter_Y_4_fifo_in_2_read;
  assign Arbiter_Y_4_fifo_in_3_dout = fifo_Y_pe_27__dout;
  assign Arbiter_Y_4_fifo_in_3_empty_n = fifo_Y_pe_27__empty_n;
  assign fifo_Y_pe_27__read = Arbiter_Y_4_fifo_in_3_read;
  assign Arbiter_Y_4_fifo_in_4_dout = fifo_Y_pe_28__dout;
  assign Arbiter_Y_4_fifo_in_4_empty_n = fifo_Y_pe_28__empty_n;
  assign fifo_Y_pe_28__read = Arbiter_Y_4_fifo_in_4_read;
  assign Arbiter_Y_4_fifo_in_5_dout = fifo_Y_pe_29__dout;
  assign Arbiter_Y_4_fifo_in_5_empty_n = fifo_Y_pe_29__empty_n;
  assign fifo_Y_pe_29__read = Arbiter_Y_4_fifo_in_5_read;
  assign Arbiter_Y_4_fifo_in_peek_0_dout = fifo_Y_pe_24__dout;
  assign Arbiter_Y_4_fifo_in_peek_0_empty_n = fifo_Y_pe_24__empty_n;
  assign Arbiter_Y_4_fifo_in_peek_1_dout = fifo_Y_pe_25__dout;
  assign Arbiter_Y_4_fifo_in_peek_1_empty_n = fifo_Y_pe_25__empty_n;
  assign Arbiter_Y_4_fifo_in_peek_2_dout = fifo_Y_pe_26__dout;
  assign Arbiter_Y_4_fifo_in_peek_2_empty_n = fifo_Y_pe_26__empty_n;
  assign Arbiter_Y_4_fifo_in_peek_3_dout = fifo_Y_pe_27__dout;
  assign Arbiter_Y_4_fifo_in_peek_3_empty_n = fifo_Y_pe_27__empty_n;
  assign Arbiter_Y_4_fifo_in_peek_4_dout = fifo_Y_pe_28__dout;
  assign Arbiter_Y_4_fifo_in_peek_4_empty_n = fifo_Y_pe_28__empty_n;
  assign Arbiter_Y_4_fifo_in_peek_5_dout = fifo_Y_pe_29__dout;
  assign Arbiter_Y_4_fifo_in_peek_5_empty_n = fifo_Y_pe_29__empty_n;
  assign fifo_Y_pe_abd_4__din = Arbiter_Y_4_fifo_out_din;
  assign Arbiter_Y_4_fifo_out_full_n = fifo_Y_pe_abd_4__full_n;
  assign fifo_Y_pe_abd_4__write = Arbiter_Y_4_fifo_out_write;
  assign Arbiter_Y_5_M = Arbiter_Y_5___M__q0;
  assign Arbiter_Y_5_P_N = Arbiter_Y_5___P_N__q0;
  assign Arbiter_Y_5_ap_clk = ap_clk;
  assign Arbiter_Y_5__ap_done = Arbiter_Y_5_ap_done;
  assign Arbiter_Y_5__ap_idle = Arbiter_Y_5_ap_idle;
  assign Arbiter_Y_5__ap_ready = Arbiter_Y_5_ap_ready;
  assign Arbiter_Y_5_ap_rst_n = ap_rst_n;
  assign Arbiter_Y_5_ap_start = Arbiter_Y_5__ap_start;
  assign Arbiter_Y_5_fifo_in_0_dout = fifo_Y_pe_30__dout;
  assign Arbiter_Y_5_fifo_in_0_empty_n = fifo_Y_pe_30__empty_n;
  assign fifo_Y_pe_30__read = Arbiter_Y_5_fifo_in_0_read;
  assign Arbiter_Y_5_fifo_in_1_dout = fifo_Y_pe_31__dout;
  assign Arbiter_Y_5_fifo_in_1_empty_n = fifo_Y_pe_31__empty_n;
  assign fifo_Y_pe_31__read = Arbiter_Y_5_fifo_in_1_read;
  assign Arbiter_Y_5_fifo_in_2_dout = fifo_Y_pe_32__dout;
  assign Arbiter_Y_5_fifo_in_2_empty_n = fifo_Y_pe_32__empty_n;
  assign fifo_Y_pe_32__read = Arbiter_Y_5_fifo_in_2_read;
  assign Arbiter_Y_5_fifo_in_3_dout = fifo_Y_pe_33__dout;
  assign Arbiter_Y_5_fifo_in_3_empty_n = fifo_Y_pe_33__empty_n;
  assign fifo_Y_pe_33__read = Arbiter_Y_5_fifo_in_3_read;
  assign Arbiter_Y_5_fifo_in_4_dout = fifo_Y_pe_34__dout;
  assign Arbiter_Y_5_fifo_in_4_empty_n = fifo_Y_pe_34__empty_n;
  assign fifo_Y_pe_34__read = Arbiter_Y_5_fifo_in_4_read;
  assign Arbiter_Y_5_fifo_in_5_dout = fifo_Y_pe_35__dout;
  assign Arbiter_Y_5_fifo_in_5_empty_n = fifo_Y_pe_35__empty_n;
  assign fifo_Y_pe_35__read = Arbiter_Y_5_fifo_in_5_read;
  assign Arbiter_Y_5_fifo_in_peek_0_dout = fifo_Y_pe_30__dout;
  assign Arbiter_Y_5_fifo_in_peek_0_empty_n = fifo_Y_pe_30__empty_n;
  assign Arbiter_Y_5_fifo_in_peek_1_dout = fifo_Y_pe_31__dout;
  assign Arbiter_Y_5_fifo_in_peek_1_empty_n = fifo_Y_pe_31__empty_n;
  assign Arbiter_Y_5_fifo_in_peek_2_dout = fifo_Y_pe_32__dout;
  assign Arbiter_Y_5_fifo_in_peek_2_empty_n = fifo_Y_pe_32__empty_n;
  assign Arbiter_Y_5_fifo_in_peek_3_dout = fifo_Y_pe_33__dout;
  assign Arbiter_Y_5_fifo_in_peek_3_empty_n = fifo_Y_pe_33__empty_n;
  assign Arbiter_Y_5_fifo_in_peek_4_dout = fifo_Y_pe_34__dout;
  assign Arbiter_Y_5_fifo_in_peek_4_empty_n = fifo_Y_pe_34__empty_n;
  assign Arbiter_Y_5_fifo_in_peek_5_dout = fifo_Y_pe_35__dout;
  assign Arbiter_Y_5_fifo_in_peek_5_empty_n = fifo_Y_pe_35__empty_n;
  assign fifo_Y_pe_abd_5__din = Arbiter_Y_5_fifo_out_din;
  assign Arbiter_Y_5_fifo_out_full_n = fifo_Y_pe_abd_5__full_n;
  assign fifo_Y_pe_abd_5__write = Arbiter_Y_5_fifo_out_write;
  assign Arbiter_Y_6_M = Arbiter_Y_6___M__q0;
  assign Arbiter_Y_6_P_N = Arbiter_Y_6___P_N__q0;
  assign Arbiter_Y_6_ap_clk = ap_clk;
  assign Arbiter_Y_6__ap_done = Arbiter_Y_6_ap_done;
  assign Arbiter_Y_6__ap_idle = Arbiter_Y_6_ap_idle;
  assign Arbiter_Y_6__ap_ready = Arbiter_Y_6_ap_ready;
  assign Arbiter_Y_6_ap_rst_n = ap_rst_n;
  assign Arbiter_Y_6_ap_start = Arbiter_Y_6__ap_start;
  assign Arbiter_Y_6_fifo_in_0_dout = fifo_Y_pe_36__dout;
  assign Arbiter_Y_6_fifo_in_0_empty_n = fifo_Y_pe_36__empty_n;
  assign fifo_Y_pe_36__read = Arbiter_Y_6_fifo_in_0_read;
  assign Arbiter_Y_6_fifo_in_1_dout = fifo_Y_pe_37__dout;
  assign Arbiter_Y_6_fifo_in_1_empty_n = fifo_Y_pe_37__empty_n;
  assign fifo_Y_pe_37__read = Arbiter_Y_6_fifo_in_1_read;
  assign Arbiter_Y_6_fifo_in_2_dout = fifo_Y_pe_38__dout;
  assign Arbiter_Y_6_fifo_in_2_empty_n = fifo_Y_pe_38__empty_n;
  assign fifo_Y_pe_38__read = Arbiter_Y_6_fifo_in_2_read;
  assign Arbiter_Y_6_fifo_in_3_dout = fifo_Y_pe_39__dout;
  assign Arbiter_Y_6_fifo_in_3_empty_n = fifo_Y_pe_39__empty_n;
  assign fifo_Y_pe_39__read = Arbiter_Y_6_fifo_in_3_read;
  assign Arbiter_Y_6_fifo_in_4_dout = fifo_Y_pe_40__dout;
  assign Arbiter_Y_6_fifo_in_4_empty_n = fifo_Y_pe_40__empty_n;
  assign fifo_Y_pe_40__read = Arbiter_Y_6_fifo_in_4_read;
  assign Arbiter_Y_6_fifo_in_5_dout = fifo_Y_pe_41__dout;
  assign Arbiter_Y_6_fifo_in_5_empty_n = fifo_Y_pe_41__empty_n;
  assign fifo_Y_pe_41__read = Arbiter_Y_6_fifo_in_5_read;
  assign Arbiter_Y_6_fifo_in_peek_0_dout = fifo_Y_pe_36__dout;
  assign Arbiter_Y_6_fifo_in_peek_0_empty_n = fifo_Y_pe_36__empty_n;
  assign Arbiter_Y_6_fifo_in_peek_1_dout = fifo_Y_pe_37__dout;
  assign Arbiter_Y_6_fifo_in_peek_1_empty_n = fifo_Y_pe_37__empty_n;
  assign Arbiter_Y_6_fifo_in_peek_2_dout = fifo_Y_pe_38__dout;
  assign Arbiter_Y_6_fifo_in_peek_2_empty_n = fifo_Y_pe_38__empty_n;
  assign Arbiter_Y_6_fifo_in_peek_3_dout = fifo_Y_pe_39__dout;
  assign Arbiter_Y_6_fifo_in_peek_3_empty_n = fifo_Y_pe_39__empty_n;
  assign Arbiter_Y_6_fifo_in_peek_4_dout = fifo_Y_pe_40__dout;
  assign Arbiter_Y_6_fifo_in_peek_4_empty_n = fifo_Y_pe_40__empty_n;
  assign Arbiter_Y_6_fifo_in_peek_5_dout = fifo_Y_pe_41__dout;
  assign Arbiter_Y_6_fifo_in_peek_5_empty_n = fifo_Y_pe_41__empty_n;
  assign fifo_Y_pe_abd_6__din = Arbiter_Y_6_fifo_out_din;
  assign Arbiter_Y_6_fifo_out_full_n = fifo_Y_pe_abd_6__full_n;
  assign fifo_Y_pe_abd_6__write = Arbiter_Y_6_fifo_out_write;
  assign Arbiter_Y_7_M = Arbiter_Y_7___M__q0;
  assign Arbiter_Y_7_P_N = Arbiter_Y_7___P_N__q0;
  assign Arbiter_Y_7_ap_clk = ap_clk;
  assign Arbiter_Y_7__ap_done = Arbiter_Y_7_ap_done;
  assign Arbiter_Y_7__ap_idle = Arbiter_Y_7_ap_idle;
  assign Arbiter_Y_7__ap_ready = Arbiter_Y_7_ap_ready;
  assign Arbiter_Y_7_ap_rst_n = ap_rst_n;
  assign Arbiter_Y_7_ap_start = Arbiter_Y_7__ap_start;
  assign Arbiter_Y_7_fifo_in_0_dout = fifo_Y_pe_42__dout;
  assign Arbiter_Y_7_fifo_in_0_empty_n = fifo_Y_pe_42__empty_n;
  assign fifo_Y_pe_42__read = Arbiter_Y_7_fifo_in_0_read;
  assign Arbiter_Y_7_fifo_in_1_dout = fifo_Y_pe_43__dout;
  assign Arbiter_Y_7_fifo_in_1_empty_n = fifo_Y_pe_43__empty_n;
  assign fifo_Y_pe_43__read = Arbiter_Y_7_fifo_in_1_read;
  assign Arbiter_Y_7_fifo_in_2_dout = fifo_Y_pe_44__dout;
  assign Arbiter_Y_7_fifo_in_2_empty_n = fifo_Y_pe_44__empty_n;
  assign fifo_Y_pe_44__read = Arbiter_Y_7_fifo_in_2_read;
  assign Arbiter_Y_7_fifo_in_3_dout = fifo_Y_pe_45__dout;
  assign Arbiter_Y_7_fifo_in_3_empty_n = fifo_Y_pe_45__empty_n;
  assign fifo_Y_pe_45__read = Arbiter_Y_7_fifo_in_3_read;
  assign Arbiter_Y_7_fifo_in_4_dout = fifo_Y_pe_46__dout;
  assign Arbiter_Y_7_fifo_in_4_empty_n = fifo_Y_pe_46__empty_n;
  assign fifo_Y_pe_46__read = Arbiter_Y_7_fifo_in_4_read;
  assign Arbiter_Y_7_fifo_in_5_dout = fifo_Y_pe_47__dout;
  assign Arbiter_Y_7_fifo_in_5_empty_n = fifo_Y_pe_47__empty_n;
  assign fifo_Y_pe_47__read = Arbiter_Y_7_fifo_in_5_read;
  assign Arbiter_Y_7_fifo_in_peek_0_dout = fifo_Y_pe_42__dout;
  assign Arbiter_Y_7_fifo_in_peek_0_empty_n = fifo_Y_pe_42__empty_n;
  assign Arbiter_Y_7_fifo_in_peek_1_dout = fifo_Y_pe_43__dout;
  assign Arbiter_Y_7_fifo_in_peek_1_empty_n = fifo_Y_pe_43__empty_n;
  assign Arbiter_Y_7_fifo_in_peek_2_dout = fifo_Y_pe_44__dout;
  assign Arbiter_Y_7_fifo_in_peek_2_empty_n = fifo_Y_pe_44__empty_n;
  assign Arbiter_Y_7_fifo_in_peek_3_dout = fifo_Y_pe_45__dout;
  assign Arbiter_Y_7_fifo_in_peek_3_empty_n = fifo_Y_pe_45__empty_n;
  assign Arbiter_Y_7_fifo_in_peek_4_dout = fifo_Y_pe_46__dout;
  assign Arbiter_Y_7_fifo_in_peek_4_empty_n = fifo_Y_pe_46__empty_n;
  assign Arbiter_Y_7_fifo_in_peek_5_dout = fifo_Y_pe_47__dout;
  assign Arbiter_Y_7_fifo_in_peek_5_empty_n = fifo_Y_pe_47__empty_n;
  assign fifo_Y_pe_abd_7__din = Arbiter_Y_7_fifo_out_din;
  assign Arbiter_Y_7_fifo_out_full_n = fifo_Y_pe_abd_7__full_n;
  assign fifo_Y_pe_abd_7__write = Arbiter_Y_7_fifo_out_write;
  assign FloatvAddFloatv_0_ap_clk = ap_clk;
  assign FloatvAddFloatv_0_ap_rst_n = ap_rst_n;
  assign FloatvAddFloatv_0_ap_start = FloatvAddFloatv_0__ap_start;
  assign FloatvAddFloatv_0_fifo_in0_peek_dout = fifo_Y_alpha_AX__dout;
  assign FloatvAddFloatv_0_fifo_in0_peek_empty_n = fifo_Y_alpha_AX__empty_n;
  assign FloatvAddFloatv_0_fifo_in0_s_dout = fifo_Y_alpha_AX__dout;
  assign FloatvAddFloatv_0_fifo_in0_s_empty_n = fifo_Y_alpha_AX__empty_n;
  assign fifo_Y_alpha_AX__read = FloatvAddFloatv_0_fifo_in0_s_read;
  assign FloatvAddFloatv_0_fifo_in1_peek_dout = fifo_Y_in_beta__dout;
  assign FloatvAddFloatv_0_fifo_in1_peek_empty_n = fifo_Y_in_beta__empty_n;
  assign FloatvAddFloatv_0_fifo_in1_s_dout = fifo_Y_in_beta__dout;
  assign FloatvAddFloatv_0_fifo_in1_s_empty_n = fifo_Y_in_beta__empty_n;
  assign fifo_Y_in_beta__read = FloatvAddFloatv_0_fifo_in1_s_read;
  assign fifo_Y_out__din = FloatvAddFloatv_0_fifo_out_din;
  assign FloatvAddFloatv_0_fifo_out_full_n = fifo_Y_out__full_n;
  assign fifo_Y_out__write = FloatvAddFloatv_0_fifo_out_write;
  assign FloatvMultConst_0_M = FloatvMultConst_0___M__q0;
  assign FloatvMultConst_0_P_N = FloatvMultConst_0___P_N__q0;
  assign FloatvMultConst_0_alpha_u = FloatvMultConst_0___alpha_u__q0;
  assign FloatvMultConst_0_ap_clk = ap_clk;
  assign FloatvMultConst_0__ap_done = FloatvMultConst_0_ap_done;
  assign FloatvMultConst_0__ap_idle = FloatvMultConst_0_ap_idle;
  assign FloatvMultConst_0__ap_ready = FloatvMultConst_0_ap_ready;
  assign FloatvMultConst_0_ap_rst_n = ap_rst_n;
  assign FloatvMultConst_0_ap_start = FloatvMultConst_0__ap_start;
  assign FloatvMultConst_0_fifo_in_peek_dout = fifo_Y_AX__dout;
  assign FloatvMultConst_0_fifo_in_peek_empty_n = fifo_Y_AX__empty_n;
  assign FloatvMultConst_0_fifo_in_s_dout = fifo_Y_AX__dout;
  assign FloatvMultConst_0_fifo_in_s_empty_n = fifo_Y_AX__empty_n;
  assign fifo_Y_AX__read = FloatvMultConst_0_fifo_in_s_read;
  assign fifo_Y_alpha_AX__din = FloatvMultConst_0_fifo_out_din;
  assign FloatvMultConst_0_fifo_out_full_n = fifo_Y_alpha_AX__full_n;
  assign fifo_Y_alpha_AX__write = FloatvMultConst_0_fifo_out_write;
  assign FloatvMultConst_1_M = FloatvMultConst_1___M__q0;
  assign FloatvMultConst_1_P_N = FloatvMultConst_1___P_N__q0;
  assign FloatvMultConst_1_alpha_u = FloatvMultConst_1___beta_u__q0;
  assign FloatvMultConst_1_ap_clk = ap_clk;
  assign FloatvMultConst_1__ap_done = FloatvMultConst_1_ap_done;
  assign FloatvMultConst_1__ap_idle = FloatvMultConst_1_ap_idle;
  assign FloatvMultConst_1__ap_ready = FloatvMultConst_1_ap_ready;
  assign FloatvMultConst_1_ap_rst_n = ap_rst_n;
  assign FloatvMultConst_1_ap_start = FloatvMultConst_1__ap_start;
  assign FloatvMultConst_1_fifo_in_peek_dout = fifo_Y_in__dout;
  assign FloatvMultConst_1_fifo_in_peek_empty_n = fifo_Y_in__empty_n;
  assign FloatvMultConst_1_fifo_in_s_dout = fifo_Y_in__dout;
  assign FloatvMultConst_1_fifo_in_s_empty_n = fifo_Y_in__empty_n;
  assign fifo_Y_in__read = FloatvMultConst_1_fifo_in_s_read;
  assign fifo_Y_in_beta__din = FloatvMultConst_1_fifo_out_din;
  assign FloatvMultConst_1_fifo_out_full_n = fifo_Y_in_beta__full_n;
  assign fifo_Y_in_beta__write = FloatvMultConst_1_fifo_out_write;
  assign Merger_Y_0_ap_clk = ap_clk;
  assign Merger_Y_0_ap_rst_n = ap_rst_n;
  assign Merger_Y_0_ap_start = Merger_Y_0__ap_start;
  assign Merger_Y_0_fifo_in_0_dout = fifo_Y_pe_abd_0__dout;
  assign Merger_Y_0_fifo_in_0_empty_n = fifo_Y_pe_abd_0__empty_n;
  assign fifo_Y_pe_abd_0__read = Merger_Y_0_fifo_in_0_read;
  assign Merger_Y_0_fifo_in_1_dout = fifo_Y_pe_abd_1__dout;
  assign Merger_Y_0_fifo_in_1_empty_n = fifo_Y_pe_abd_1__empty_n;
  assign fifo_Y_pe_abd_1__read = Merger_Y_0_fifo_in_1_read;
  assign Merger_Y_0_fifo_in_2_dout = fifo_Y_pe_abd_2__dout;
  assign Merger_Y_0_fifo_in_2_empty_n = fifo_Y_pe_abd_2__empty_n;
  assign fifo_Y_pe_abd_2__read = Merger_Y_0_fifo_in_2_read;
  assign Merger_Y_0_fifo_in_3_dout = fifo_Y_pe_abd_3__dout;
  assign Merger_Y_0_fifo_in_3_empty_n = fifo_Y_pe_abd_3__empty_n;
  assign fifo_Y_pe_abd_3__read = Merger_Y_0_fifo_in_3_read;
  assign Merger_Y_0_fifo_in_4_dout = fifo_Y_pe_abd_4__dout;
  assign Merger_Y_0_fifo_in_4_empty_n = fifo_Y_pe_abd_4__empty_n;
  assign fifo_Y_pe_abd_4__read = Merger_Y_0_fifo_in_4_read;
  assign Merger_Y_0_fifo_in_5_dout = fifo_Y_pe_abd_5__dout;
  assign Merger_Y_0_fifo_in_5_empty_n = fifo_Y_pe_abd_5__empty_n;
  assign fifo_Y_pe_abd_5__read = Merger_Y_0_fifo_in_5_read;
  assign Merger_Y_0_fifo_in_6_dout = fifo_Y_pe_abd_6__dout;
  assign Merger_Y_0_fifo_in_6_empty_n = fifo_Y_pe_abd_6__empty_n;
  assign fifo_Y_pe_abd_6__read = Merger_Y_0_fifo_in_6_read;
  assign Merger_Y_0_fifo_in_7_dout = fifo_Y_pe_abd_7__dout;
  assign Merger_Y_0_fifo_in_7_empty_n = fifo_Y_pe_abd_7__empty_n;
  assign fifo_Y_pe_abd_7__read = Merger_Y_0_fifo_in_7_read;
  assign Merger_Y_0_fifo_in_peek_0_dout = fifo_Y_pe_abd_0__dout;
  assign Merger_Y_0_fifo_in_peek_0_empty_n = fifo_Y_pe_abd_0__empty_n;
  assign Merger_Y_0_fifo_in_peek_1_dout = fifo_Y_pe_abd_1__dout;
  assign Merger_Y_0_fifo_in_peek_1_empty_n = fifo_Y_pe_abd_1__empty_n;
  assign Merger_Y_0_fifo_in_peek_2_dout = fifo_Y_pe_abd_2__dout;
  assign Merger_Y_0_fifo_in_peek_2_empty_n = fifo_Y_pe_abd_2__empty_n;
  assign Merger_Y_0_fifo_in_peek_3_dout = fifo_Y_pe_abd_3__dout;
  assign Merger_Y_0_fifo_in_peek_3_empty_n = fifo_Y_pe_abd_3__empty_n;
  assign Merger_Y_0_fifo_in_peek_4_dout = fifo_Y_pe_abd_4__dout;
  assign Merger_Y_0_fifo_in_peek_4_empty_n = fifo_Y_pe_abd_4__empty_n;
  assign Merger_Y_0_fifo_in_peek_5_dout = fifo_Y_pe_abd_5__dout;
  assign Merger_Y_0_fifo_in_peek_5_empty_n = fifo_Y_pe_abd_5__empty_n;
  assign Merger_Y_0_fifo_in_peek_6_dout = fifo_Y_pe_abd_6__dout;
  assign Merger_Y_0_fifo_in_peek_6_empty_n = fifo_Y_pe_abd_6__empty_n;
  assign Merger_Y_0_fifo_in_peek_7_dout = fifo_Y_pe_abd_7__dout;
  assign Merger_Y_0_fifo_in_peek_7_empty_n = fifo_Y_pe_abd_7__empty_n;
  assign fifo_Y_AX__din = Merger_Y_0_fifo_out_din;
  assign Merger_Y_0_fifo_out_full_n = fifo_Y_AX__full_n;
  assign fifo_Y_AX__write = Merger_Y_0_fifo_out_write;
  assign PEG_Xvec_0_ap_clk = ap_clk;
  assign PEG_Xvec_0__ap_done = PEG_Xvec_0_ap_done;
  assign PEG_Xvec_0__ap_idle = PEG_Xvec_0_ap_idle;
  assign PEG_Xvec_0__ap_ready = PEG_Xvec_0_ap_ready;
  assign PEG_Xvec_0_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_0_ap_start = PEG_Xvec_0__ap_start;
  assign PEG_Xvec_0_fifo_A_peek_dout = fifo_A_0__dout;
  assign PEG_Xvec_0_fifo_A_peek_empty_n = fifo_A_0__empty_n;
  assign PEG_Xvec_0_fifo_A_s_dout = fifo_A_0__dout;
  assign PEG_Xvec_0_fifo_A_s_empty_n = fifo_A_0__empty_n;
  assign fifo_A_0__read = PEG_Xvec_0_fifo_A_s_read;
  assign PEG_Xvec_0_fifo_X_in_peek_dout = fifo_X_pe_0__dout;
  assign PEG_Xvec_0_fifo_X_in_peek_empty_n = fifo_X_pe_0__empty_n;
  assign PEG_Xvec_0_fifo_X_in_s_dout = fifo_X_pe_0__dout;
  assign PEG_Xvec_0_fifo_X_in_s_empty_n = fifo_X_pe_0__empty_n;
  assign fifo_X_pe_0__read = PEG_Xvec_0_fifo_X_in_s_read;
  assign fifo_X_pe_1__din = PEG_Xvec_0_fifo_X_out_din;
  assign PEG_Xvec_0_fifo_X_out_full_n = fifo_X_pe_1__full_n;
  assign fifo_X_pe_1__write = PEG_Xvec_0_fifo_X_out_write;
  assign fifo_aXvec_0__din = PEG_Xvec_0_fifo_aXvec_din;
  assign PEG_Xvec_0_fifo_aXvec_full_n = fifo_aXvec_0__full_n;
  assign fifo_aXvec_0__write = PEG_Xvec_0_fifo_aXvec_write;
  assign PEG_Xvec_0_fifo_inst_in_peek_dout = PE_inst_0__dout;
  assign PEG_Xvec_0_fifo_inst_in_peek_empty_n = PE_inst_0__empty_n;
  assign PEG_Xvec_0_fifo_inst_in_s_dout = PE_inst_0__dout;
  assign PEG_Xvec_0_fifo_inst_in_s_empty_n = PE_inst_0__empty_n;
  assign PE_inst_0__read = PEG_Xvec_0_fifo_inst_in_s_read;
  assign PE_inst_1__din = PEG_Xvec_0_fifo_inst_out_din;
  assign PEG_Xvec_0_fifo_inst_out_full_n = PE_inst_1__full_n;
  assign Yvec_inst_0__din = PEG_Xvec_0_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_0_fifo_inst_out_to_Yvec_full_n = Yvec_inst_0__full_n;
  assign Yvec_inst_0__write = PEG_Xvec_0_fifo_inst_out_to_Yvec_write;
  assign PE_inst_1__write = PEG_Xvec_0_fifo_inst_out_write;
  assign PEG_Xvec_1_ap_clk = ap_clk;
  assign PEG_Xvec_1__ap_done = PEG_Xvec_1_ap_done;
  assign PEG_Xvec_1__ap_idle = PEG_Xvec_1_ap_idle;
  assign PEG_Xvec_1__ap_ready = PEG_Xvec_1_ap_ready;
  assign PEG_Xvec_1_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_1_ap_start = PEG_Xvec_1__ap_start;
  assign PEG_Xvec_1_fifo_A_peek_dout = fifo_A_1__dout;
  assign PEG_Xvec_1_fifo_A_peek_empty_n = fifo_A_1__empty_n;
  assign PEG_Xvec_1_fifo_A_s_dout = fifo_A_1__dout;
  assign PEG_Xvec_1_fifo_A_s_empty_n = fifo_A_1__empty_n;
  assign fifo_A_1__read = PEG_Xvec_1_fifo_A_s_read;
  assign PEG_Xvec_1_fifo_X_in_peek_dout = fifo_X_pe_1__dout;
  assign PEG_Xvec_1_fifo_X_in_peek_empty_n = fifo_X_pe_1__empty_n;
  assign PEG_Xvec_1_fifo_X_in_s_dout = fifo_X_pe_1__dout;
  assign PEG_Xvec_1_fifo_X_in_s_empty_n = fifo_X_pe_1__empty_n;
  assign fifo_X_pe_1__read = PEG_Xvec_1_fifo_X_in_s_read;
  assign fifo_X_pe_2__din = PEG_Xvec_1_fifo_X_out_din;
  assign PEG_Xvec_1_fifo_X_out_full_n = fifo_X_pe_2__full_n;
  assign fifo_X_pe_2__write = PEG_Xvec_1_fifo_X_out_write;
  assign fifo_aXvec_1__din = PEG_Xvec_1_fifo_aXvec_din;
  assign PEG_Xvec_1_fifo_aXvec_full_n = fifo_aXvec_1__full_n;
  assign fifo_aXvec_1__write = PEG_Xvec_1_fifo_aXvec_write;
  assign PEG_Xvec_1_fifo_inst_in_peek_dout = PE_inst_1__dout;
  assign PEG_Xvec_1_fifo_inst_in_peek_empty_n = PE_inst_1__empty_n;
  assign PEG_Xvec_1_fifo_inst_in_s_dout = PE_inst_1__dout;
  assign PEG_Xvec_1_fifo_inst_in_s_empty_n = PE_inst_1__empty_n;
  assign PE_inst_1__read = PEG_Xvec_1_fifo_inst_in_s_read;
  assign PE_inst_2__din = PEG_Xvec_1_fifo_inst_out_din;
  assign PEG_Xvec_1_fifo_inst_out_full_n = PE_inst_2__full_n;
  assign Yvec_inst_1__din = PEG_Xvec_1_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_1_fifo_inst_out_to_Yvec_full_n = Yvec_inst_1__full_n;
  assign Yvec_inst_1__write = PEG_Xvec_1_fifo_inst_out_to_Yvec_write;
  assign PE_inst_2__write = PEG_Xvec_1_fifo_inst_out_write;
  assign PEG_Xvec_2_ap_clk = ap_clk;
  assign PEG_Xvec_2__ap_done = PEG_Xvec_2_ap_done;
  assign PEG_Xvec_2__ap_idle = PEG_Xvec_2_ap_idle;
  assign PEG_Xvec_2__ap_ready = PEG_Xvec_2_ap_ready;
  assign PEG_Xvec_2_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_2_ap_start = PEG_Xvec_2__ap_start;
  assign PEG_Xvec_2_fifo_A_peek_dout = fifo_A_2__dout;
  assign PEG_Xvec_2_fifo_A_peek_empty_n = fifo_A_2__empty_n;
  assign PEG_Xvec_2_fifo_A_s_dout = fifo_A_2__dout;
  assign PEG_Xvec_2_fifo_A_s_empty_n = fifo_A_2__empty_n;
  assign fifo_A_2__read = PEG_Xvec_2_fifo_A_s_read;
  assign PEG_Xvec_2_fifo_X_in_peek_dout = fifo_X_pe_2__dout;
  assign PEG_Xvec_2_fifo_X_in_peek_empty_n = fifo_X_pe_2__empty_n;
  assign PEG_Xvec_2_fifo_X_in_s_dout = fifo_X_pe_2__dout;
  assign PEG_Xvec_2_fifo_X_in_s_empty_n = fifo_X_pe_2__empty_n;
  assign fifo_X_pe_2__read = PEG_Xvec_2_fifo_X_in_s_read;
  assign fifo_X_pe_3__din = PEG_Xvec_2_fifo_X_out_din;
  assign PEG_Xvec_2_fifo_X_out_full_n = fifo_X_pe_3__full_n;
  assign fifo_X_pe_3__write = PEG_Xvec_2_fifo_X_out_write;
  assign fifo_aXvec_2__din = PEG_Xvec_2_fifo_aXvec_din;
  assign PEG_Xvec_2_fifo_aXvec_full_n = fifo_aXvec_2__full_n;
  assign fifo_aXvec_2__write = PEG_Xvec_2_fifo_aXvec_write;
  assign PEG_Xvec_2_fifo_inst_in_peek_dout = PE_inst_2__dout;
  assign PEG_Xvec_2_fifo_inst_in_peek_empty_n = PE_inst_2__empty_n;
  assign PEG_Xvec_2_fifo_inst_in_s_dout = PE_inst_2__dout;
  assign PEG_Xvec_2_fifo_inst_in_s_empty_n = PE_inst_2__empty_n;
  assign PE_inst_2__read = PEG_Xvec_2_fifo_inst_in_s_read;
  assign PE_inst_3__din = PEG_Xvec_2_fifo_inst_out_din;
  assign PEG_Xvec_2_fifo_inst_out_full_n = PE_inst_3__full_n;
  assign Yvec_inst_2__din = PEG_Xvec_2_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_2_fifo_inst_out_to_Yvec_full_n = Yvec_inst_2__full_n;
  assign Yvec_inst_2__write = PEG_Xvec_2_fifo_inst_out_to_Yvec_write;
  assign PE_inst_3__write = PEG_Xvec_2_fifo_inst_out_write;
  assign PEG_Xvec_3_ap_clk = ap_clk;
  assign PEG_Xvec_3__ap_done = PEG_Xvec_3_ap_done;
  assign PEG_Xvec_3__ap_idle = PEG_Xvec_3_ap_idle;
  assign PEG_Xvec_3__ap_ready = PEG_Xvec_3_ap_ready;
  assign PEG_Xvec_3_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_3_ap_start = PEG_Xvec_3__ap_start;
  assign PEG_Xvec_3_fifo_A_peek_dout = fifo_A_3__dout;
  assign PEG_Xvec_3_fifo_A_peek_empty_n = fifo_A_3__empty_n;
  assign PEG_Xvec_3_fifo_A_s_dout = fifo_A_3__dout;
  assign PEG_Xvec_3_fifo_A_s_empty_n = fifo_A_3__empty_n;
  assign fifo_A_3__read = PEG_Xvec_3_fifo_A_s_read;
  assign PEG_Xvec_3_fifo_X_in_peek_dout = fifo_X_pe_3__dout;
  assign PEG_Xvec_3_fifo_X_in_peek_empty_n = fifo_X_pe_3__empty_n;
  assign PEG_Xvec_3_fifo_X_in_s_dout = fifo_X_pe_3__dout;
  assign PEG_Xvec_3_fifo_X_in_s_empty_n = fifo_X_pe_3__empty_n;
  assign fifo_X_pe_3__read = PEG_Xvec_3_fifo_X_in_s_read;
  assign fifo_X_pe_4__din = PEG_Xvec_3_fifo_X_out_din;
  assign PEG_Xvec_3_fifo_X_out_full_n = fifo_X_pe_4__full_n;
  assign fifo_X_pe_4__write = PEG_Xvec_3_fifo_X_out_write;
  assign fifo_aXvec_3__din = PEG_Xvec_3_fifo_aXvec_din;
  assign PEG_Xvec_3_fifo_aXvec_full_n = fifo_aXvec_3__full_n;
  assign fifo_aXvec_3__write = PEG_Xvec_3_fifo_aXvec_write;
  assign PEG_Xvec_3_fifo_inst_in_peek_dout = PE_inst_3__dout;
  assign PEG_Xvec_3_fifo_inst_in_peek_empty_n = PE_inst_3__empty_n;
  assign PEG_Xvec_3_fifo_inst_in_s_dout = PE_inst_3__dout;
  assign PEG_Xvec_3_fifo_inst_in_s_empty_n = PE_inst_3__empty_n;
  assign PE_inst_3__read = PEG_Xvec_3_fifo_inst_in_s_read;
  assign PE_inst_4__din = PEG_Xvec_3_fifo_inst_out_din;
  assign PEG_Xvec_3_fifo_inst_out_full_n = PE_inst_4__full_n;
  assign Yvec_inst_3__din = PEG_Xvec_3_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_3_fifo_inst_out_to_Yvec_full_n = Yvec_inst_3__full_n;
  assign Yvec_inst_3__write = PEG_Xvec_3_fifo_inst_out_to_Yvec_write;
  assign PE_inst_4__write = PEG_Xvec_3_fifo_inst_out_write;
  assign PEG_Xvec_4_ap_clk = ap_clk;
  assign PEG_Xvec_4__ap_done = PEG_Xvec_4_ap_done;
  assign PEG_Xvec_4__ap_idle = PEG_Xvec_4_ap_idle;
  assign PEG_Xvec_4__ap_ready = PEG_Xvec_4_ap_ready;
  assign PEG_Xvec_4_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_4_ap_start = PEG_Xvec_4__ap_start;
  assign PEG_Xvec_4_fifo_A_peek_dout = fifo_A_4__dout;
  assign PEG_Xvec_4_fifo_A_peek_empty_n = fifo_A_4__empty_n;
  assign PEG_Xvec_4_fifo_A_s_dout = fifo_A_4__dout;
  assign PEG_Xvec_4_fifo_A_s_empty_n = fifo_A_4__empty_n;
  assign fifo_A_4__read = PEG_Xvec_4_fifo_A_s_read;
  assign PEG_Xvec_4_fifo_X_in_peek_dout = fifo_X_pe_4__dout;
  assign PEG_Xvec_4_fifo_X_in_peek_empty_n = fifo_X_pe_4__empty_n;
  assign PEG_Xvec_4_fifo_X_in_s_dout = fifo_X_pe_4__dout;
  assign PEG_Xvec_4_fifo_X_in_s_empty_n = fifo_X_pe_4__empty_n;
  assign fifo_X_pe_4__read = PEG_Xvec_4_fifo_X_in_s_read;
  assign fifo_X_pe_5__din = PEG_Xvec_4_fifo_X_out_din;
  assign PEG_Xvec_4_fifo_X_out_full_n = fifo_X_pe_5__full_n;
  assign fifo_X_pe_5__write = PEG_Xvec_4_fifo_X_out_write;
  assign fifo_aXvec_4__din = PEG_Xvec_4_fifo_aXvec_din;
  assign PEG_Xvec_4_fifo_aXvec_full_n = fifo_aXvec_4__full_n;
  assign fifo_aXvec_4__write = PEG_Xvec_4_fifo_aXvec_write;
  assign PEG_Xvec_4_fifo_inst_in_peek_dout = PE_inst_4__dout;
  assign PEG_Xvec_4_fifo_inst_in_peek_empty_n = PE_inst_4__empty_n;
  assign PEG_Xvec_4_fifo_inst_in_s_dout = PE_inst_4__dout;
  assign PEG_Xvec_4_fifo_inst_in_s_empty_n = PE_inst_4__empty_n;
  assign PE_inst_4__read = PEG_Xvec_4_fifo_inst_in_s_read;
  assign PE_inst_5__din = PEG_Xvec_4_fifo_inst_out_din;
  assign PEG_Xvec_4_fifo_inst_out_full_n = PE_inst_5__full_n;
  assign Yvec_inst_4__din = PEG_Xvec_4_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_4_fifo_inst_out_to_Yvec_full_n = Yvec_inst_4__full_n;
  assign Yvec_inst_4__write = PEG_Xvec_4_fifo_inst_out_to_Yvec_write;
  assign PE_inst_5__write = PEG_Xvec_4_fifo_inst_out_write;
  assign PEG_Xvec_5_ap_clk = ap_clk;
  assign PEG_Xvec_5__ap_done = PEG_Xvec_5_ap_done;
  assign PEG_Xvec_5__ap_idle = PEG_Xvec_5_ap_idle;
  assign PEG_Xvec_5__ap_ready = PEG_Xvec_5_ap_ready;
  assign PEG_Xvec_5_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_5_ap_start = PEG_Xvec_5__ap_start;
  assign PEG_Xvec_5_fifo_A_peek_dout = fifo_A_5__dout;
  assign PEG_Xvec_5_fifo_A_peek_empty_n = fifo_A_5__empty_n;
  assign PEG_Xvec_5_fifo_A_s_dout = fifo_A_5__dout;
  assign PEG_Xvec_5_fifo_A_s_empty_n = fifo_A_5__empty_n;
  assign fifo_A_5__read = PEG_Xvec_5_fifo_A_s_read;
  assign PEG_Xvec_5_fifo_X_in_peek_dout = fifo_X_pe_5__dout;
  assign PEG_Xvec_5_fifo_X_in_peek_empty_n = fifo_X_pe_5__empty_n;
  assign PEG_Xvec_5_fifo_X_in_s_dout = fifo_X_pe_5__dout;
  assign PEG_Xvec_5_fifo_X_in_s_empty_n = fifo_X_pe_5__empty_n;
  assign fifo_X_pe_5__read = PEG_Xvec_5_fifo_X_in_s_read;
  assign fifo_X_pe_6__din = PEG_Xvec_5_fifo_X_out_din;
  assign PEG_Xvec_5_fifo_X_out_full_n = fifo_X_pe_6__full_n;
  assign fifo_X_pe_6__write = PEG_Xvec_5_fifo_X_out_write;
  assign fifo_aXvec_5__din = PEG_Xvec_5_fifo_aXvec_din;
  assign PEG_Xvec_5_fifo_aXvec_full_n = fifo_aXvec_5__full_n;
  assign fifo_aXvec_5__write = PEG_Xvec_5_fifo_aXvec_write;
  assign PEG_Xvec_5_fifo_inst_in_peek_dout = PE_inst_5__dout;
  assign PEG_Xvec_5_fifo_inst_in_peek_empty_n = PE_inst_5__empty_n;
  assign PEG_Xvec_5_fifo_inst_in_s_dout = PE_inst_5__dout;
  assign PEG_Xvec_5_fifo_inst_in_s_empty_n = PE_inst_5__empty_n;
  assign PE_inst_5__read = PEG_Xvec_5_fifo_inst_in_s_read;
  assign PE_inst_6__din = PEG_Xvec_5_fifo_inst_out_din;
  assign PEG_Xvec_5_fifo_inst_out_full_n = PE_inst_6__full_n;
  assign Yvec_inst_5__din = PEG_Xvec_5_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_5_fifo_inst_out_to_Yvec_full_n = Yvec_inst_5__full_n;
  assign Yvec_inst_5__write = PEG_Xvec_5_fifo_inst_out_to_Yvec_write;
  assign PE_inst_6__write = PEG_Xvec_5_fifo_inst_out_write;
  assign PEG_Xvec_6_ap_clk = ap_clk;
  assign PEG_Xvec_6__ap_done = PEG_Xvec_6_ap_done;
  assign PEG_Xvec_6__ap_idle = PEG_Xvec_6_ap_idle;
  assign PEG_Xvec_6__ap_ready = PEG_Xvec_6_ap_ready;
  assign PEG_Xvec_6_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_6_ap_start = PEG_Xvec_6__ap_start;
  assign PEG_Xvec_6_fifo_A_peek_dout = fifo_A_6__dout;
  assign PEG_Xvec_6_fifo_A_peek_empty_n = fifo_A_6__empty_n;
  assign PEG_Xvec_6_fifo_A_s_dout = fifo_A_6__dout;
  assign PEG_Xvec_6_fifo_A_s_empty_n = fifo_A_6__empty_n;
  assign fifo_A_6__read = PEG_Xvec_6_fifo_A_s_read;
  assign PEG_Xvec_6_fifo_X_in_peek_dout = fifo_X_pe_6__dout;
  assign PEG_Xvec_6_fifo_X_in_peek_empty_n = fifo_X_pe_6__empty_n;
  assign PEG_Xvec_6_fifo_X_in_s_dout = fifo_X_pe_6__dout;
  assign PEG_Xvec_6_fifo_X_in_s_empty_n = fifo_X_pe_6__empty_n;
  assign fifo_X_pe_6__read = PEG_Xvec_6_fifo_X_in_s_read;
  assign fifo_X_pe_7__din = PEG_Xvec_6_fifo_X_out_din;
  assign PEG_Xvec_6_fifo_X_out_full_n = fifo_X_pe_7__full_n;
  assign fifo_X_pe_7__write = PEG_Xvec_6_fifo_X_out_write;
  assign fifo_aXvec_6__din = PEG_Xvec_6_fifo_aXvec_din;
  assign PEG_Xvec_6_fifo_aXvec_full_n = fifo_aXvec_6__full_n;
  assign fifo_aXvec_6__write = PEG_Xvec_6_fifo_aXvec_write;
  assign PEG_Xvec_6_fifo_inst_in_peek_dout = PE_inst_6__dout;
  assign PEG_Xvec_6_fifo_inst_in_peek_empty_n = PE_inst_6__empty_n;
  assign PEG_Xvec_6_fifo_inst_in_s_dout = PE_inst_6__dout;
  assign PEG_Xvec_6_fifo_inst_in_s_empty_n = PE_inst_6__empty_n;
  assign PE_inst_6__read = PEG_Xvec_6_fifo_inst_in_s_read;
  assign PE_inst_7__din = PEG_Xvec_6_fifo_inst_out_din;
  assign PEG_Xvec_6_fifo_inst_out_full_n = PE_inst_7__full_n;
  assign Yvec_inst_6__din = PEG_Xvec_6_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_6_fifo_inst_out_to_Yvec_full_n = Yvec_inst_6__full_n;
  assign Yvec_inst_6__write = PEG_Xvec_6_fifo_inst_out_to_Yvec_write;
  assign PE_inst_7__write = PEG_Xvec_6_fifo_inst_out_write;
  assign PEG_Xvec_7_ap_clk = ap_clk;
  assign PEG_Xvec_7__ap_done = PEG_Xvec_7_ap_done;
  assign PEG_Xvec_7__ap_idle = PEG_Xvec_7_ap_idle;
  assign PEG_Xvec_7__ap_ready = PEG_Xvec_7_ap_ready;
  assign PEG_Xvec_7_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_7_ap_start = PEG_Xvec_7__ap_start;
  assign PEG_Xvec_7_fifo_A_peek_dout = fifo_A_7__dout;
  assign PEG_Xvec_7_fifo_A_peek_empty_n = fifo_A_7__empty_n;
  assign PEG_Xvec_7_fifo_A_s_dout = fifo_A_7__dout;
  assign PEG_Xvec_7_fifo_A_s_empty_n = fifo_A_7__empty_n;
  assign fifo_A_7__read = PEG_Xvec_7_fifo_A_s_read;
  assign PEG_Xvec_7_fifo_X_in_peek_dout = fifo_X_pe_7__dout;
  assign PEG_Xvec_7_fifo_X_in_peek_empty_n = fifo_X_pe_7__empty_n;
  assign PEG_Xvec_7_fifo_X_in_s_dout = fifo_X_pe_7__dout;
  assign PEG_Xvec_7_fifo_X_in_s_empty_n = fifo_X_pe_7__empty_n;
  assign fifo_X_pe_7__read = PEG_Xvec_7_fifo_X_in_s_read;
  assign fifo_X_pe_8__din = PEG_Xvec_7_fifo_X_out_din;
  assign PEG_Xvec_7_fifo_X_out_full_n = fifo_X_pe_8__full_n;
  assign fifo_X_pe_8__write = PEG_Xvec_7_fifo_X_out_write;
  assign fifo_aXvec_7__din = PEG_Xvec_7_fifo_aXvec_din;
  assign PEG_Xvec_7_fifo_aXvec_full_n = fifo_aXvec_7__full_n;
  assign fifo_aXvec_7__write = PEG_Xvec_7_fifo_aXvec_write;
  assign PEG_Xvec_7_fifo_inst_in_peek_dout = PE_inst_7__dout;
  assign PEG_Xvec_7_fifo_inst_in_peek_empty_n = PE_inst_7__empty_n;
  assign PEG_Xvec_7_fifo_inst_in_s_dout = PE_inst_7__dout;
  assign PEG_Xvec_7_fifo_inst_in_s_empty_n = PE_inst_7__empty_n;
  assign PE_inst_7__read = PEG_Xvec_7_fifo_inst_in_s_read;
  assign PE_inst_8__din = PEG_Xvec_7_fifo_inst_out_din;
  assign PEG_Xvec_7_fifo_inst_out_full_n = PE_inst_8__full_n;
  assign Yvec_inst_7__din = PEG_Xvec_7_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_7_fifo_inst_out_to_Yvec_full_n = Yvec_inst_7__full_n;
  assign Yvec_inst_7__write = PEG_Xvec_7_fifo_inst_out_to_Yvec_write;
  assign PE_inst_8__write = PEG_Xvec_7_fifo_inst_out_write;
  assign PEG_Xvec_8_ap_clk = ap_clk;
  assign PEG_Xvec_8__ap_done = PEG_Xvec_8_ap_done;
  assign PEG_Xvec_8__ap_idle = PEG_Xvec_8_ap_idle;
  assign PEG_Xvec_8__ap_ready = PEG_Xvec_8_ap_ready;
  assign PEG_Xvec_8_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_8_ap_start = PEG_Xvec_8__ap_start;
  assign PEG_Xvec_8_fifo_A_peek_dout = fifo_A_8__dout;
  assign PEG_Xvec_8_fifo_A_peek_empty_n = fifo_A_8__empty_n;
  assign PEG_Xvec_8_fifo_A_s_dout = fifo_A_8__dout;
  assign PEG_Xvec_8_fifo_A_s_empty_n = fifo_A_8__empty_n;
  assign fifo_A_8__read = PEG_Xvec_8_fifo_A_s_read;
  assign PEG_Xvec_8_fifo_X_in_peek_dout = fifo_X_pe_8__dout;
  assign PEG_Xvec_8_fifo_X_in_peek_empty_n = fifo_X_pe_8__empty_n;
  assign PEG_Xvec_8_fifo_X_in_s_dout = fifo_X_pe_8__dout;
  assign PEG_Xvec_8_fifo_X_in_s_empty_n = fifo_X_pe_8__empty_n;
  assign fifo_X_pe_8__read = PEG_Xvec_8_fifo_X_in_s_read;
  assign fifo_X_pe_9__din = PEG_Xvec_8_fifo_X_out_din;
  assign PEG_Xvec_8_fifo_X_out_full_n = fifo_X_pe_9__full_n;
  assign fifo_X_pe_9__write = PEG_Xvec_8_fifo_X_out_write;
  assign fifo_aXvec_8__din = PEG_Xvec_8_fifo_aXvec_din;
  assign PEG_Xvec_8_fifo_aXvec_full_n = fifo_aXvec_8__full_n;
  assign fifo_aXvec_8__write = PEG_Xvec_8_fifo_aXvec_write;
  assign PEG_Xvec_8_fifo_inst_in_peek_dout = PE_inst_8__dout;
  assign PEG_Xvec_8_fifo_inst_in_peek_empty_n = PE_inst_8__empty_n;
  assign PEG_Xvec_8_fifo_inst_in_s_dout = PE_inst_8__dout;
  assign PEG_Xvec_8_fifo_inst_in_s_empty_n = PE_inst_8__empty_n;
  assign PE_inst_8__read = PEG_Xvec_8_fifo_inst_in_s_read;
  assign PE_inst_9__din = PEG_Xvec_8_fifo_inst_out_din;
  assign PEG_Xvec_8_fifo_inst_out_full_n = PE_inst_9__full_n;
  assign Yvec_inst_8__din = PEG_Xvec_8_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_8_fifo_inst_out_to_Yvec_full_n = Yvec_inst_8__full_n;
  assign Yvec_inst_8__write = PEG_Xvec_8_fifo_inst_out_to_Yvec_write;
  assign PE_inst_9__write = PEG_Xvec_8_fifo_inst_out_write;
  assign PEG_Xvec_9_ap_clk = ap_clk;
  assign PEG_Xvec_9__ap_done = PEG_Xvec_9_ap_done;
  assign PEG_Xvec_9__ap_idle = PEG_Xvec_9_ap_idle;
  assign PEG_Xvec_9__ap_ready = PEG_Xvec_9_ap_ready;
  assign PEG_Xvec_9_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_9_ap_start = PEG_Xvec_9__ap_start;
  assign PEG_Xvec_9_fifo_A_peek_dout = fifo_A_9__dout;
  assign PEG_Xvec_9_fifo_A_peek_empty_n = fifo_A_9__empty_n;
  assign PEG_Xvec_9_fifo_A_s_dout = fifo_A_9__dout;
  assign PEG_Xvec_9_fifo_A_s_empty_n = fifo_A_9__empty_n;
  assign fifo_A_9__read = PEG_Xvec_9_fifo_A_s_read;
  assign PEG_Xvec_9_fifo_X_in_peek_dout = fifo_X_pe_9__dout;
  assign PEG_Xvec_9_fifo_X_in_peek_empty_n = fifo_X_pe_9__empty_n;
  assign PEG_Xvec_9_fifo_X_in_s_dout = fifo_X_pe_9__dout;
  assign PEG_Xvec_9_fifo_X_in_s_empty_n = fifo_X_pe_9__empty_n;
  assign fifo_X_pe_9__read = PEG_Xvec_9_fifo_X_in_s_read;
  assign fifo_X_pe_10__din = PEG_Xvec_9_fifo_X_out_din;
  assign PEG_Xvec_9_fifo_X_out_full_n = fifo_X_pe_10__full_n;
  assign fifo_X_pe_10__write = PEG_Xvec_9_fifo_X_out_write;
  assign fifo_aXvec_9__din = PEG_Xvec_9_fifo_aXvec_din;
  assign PEG_Xvec_9_fifo_aXvec_full_n = fifo_aXvec_9__full_n;
  assign fifo_aXvec_9__write = PEG_Xvec_9_fifo_aXvec_write;
  assign PEG_Xvec_9_fifo_inst_in_peek_dout = PE_inst_9__dout;
  assign PEG_Xvec_9_fifo_inst_in_peek_empty_n = PE_inst_9__empty_n;
  assign PEG_Xvec_9_fifo_inst_in_s_dout = PE_inst_9__dout;
  assign PEG_Xvec_9_fifo_inst_in_s_empty_n = PE_inst_9__empty_n;
  assign PE_inst_9__read = PEG_Xvec_9_fifo_inst_in_s_read;
  assign PE_inst_10__din = PEG_Xvec_9_fifo_inst_out_din;
  assign PEG_Xvec_9_fifo_inst_out_full_n = PE_inst_10__full_n;
  assign Yvec_inst_9__din = PEG_Xvec_9_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_9_fifo_inst_out_to_Yvec_full_n = Yvec_inst_9__full_n;
  assign Yvec_inst_9__write = PEG_Xvec_9_fifo_inst_out_to_Yvec_write;
  assign PE_inst_10__write = PEG_Xvec_9_fifo_inst_out_write;
  assign PEG_Xvec_10_ap_clk = ap_clk;
  assign PEG_Xvec_10__ap_done = PEG_Xvec_10_ap_done;
  assign PEG_Xvec_10__ap_idle = PEG_Xvec_10_ap_idle;
  assign PEG_Xvec_10__ap_ready = PEG_Xvec_10_ap_ready;
  assign PEG_Xvec_10_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_10_ap_start = PEG_Xvec_10__ap_start;
  assign PEG_Xvec_10_fifo_A_peek_dout = fifo_A_10__dout;
  assign PEG_Xvec_10_fifo_A_peek_empty_n = fifo_A_10__empty_n;
  assign PEG_Xvec_10_fifo_A_s_dout = fifo_A_10__dout;
  assign PEG_Xvec_10_fifo_A_s_empty_n = fifo_A_10__empty_n;
  assign fifo_A_10__read = PEG_Xvec_10_fifo_A_s_read;
  assign PEG_Xvec_10_fifo_X_in_peek_dout = fifo_X_pe_10__dout;
  assign PEG_Xvec_10_fifo_X_in_peek_empty_n = fifo_X_pe_10__empty_n;
  assign PEG_Xvec_10_fifo_X_in_s_dout = fifo_X_pe_10__dout;
  assign PEG_Xvec_10_fifo_X_in_s_empty_n = fifo_X_pe_10__empty_n;
  assign fifo_X_pe_10__read = PEG_Xvec_10_fifo_X_in_s_read;
  assign fifo_X_pe_11__din = PEG_Xvec_10_fifo_X_out_din;
  assign PEG_Xvec_10_fifo_X_out_full_n = fifo_X_pe_11__full_n;
  assign fifo_X_pe_11__write = PEG_Xvec_10_fifo_X_out_write;
  assign fifo_aXvec_10__din = PEG_Xvec_10_fifo_aXvec_din;
  assign PEG_Xvec_10_fifo_aXvec_full_n = fifo_aXvec_10__full_n;
  assign fifo_aXvec_10__write = PEG_Xvec_10_fifo_aXvec_write;
  assign PEG_Xvec_10_fifo_inst_in_peek_dout = PE_inst_10__dout;
  assign PEG_Xvec_10_fifo_inst_in_peek_empty_n = PE_inst_10__empty_n;
  assign PEG_Xvec_10_fifo_inst_in_s_dout = PE_inst_10__dout;
  assign PEG_Xvec_10_fifo_inst_in_s_empty_n = PE_inst_10__empty_n;
  assign PE_inst_10__read = PEG_Xvec_10_fifo_inst_in_s_read;
  assign PE_inst_11__din = PEG_Xvec_10_fifo_inst_out_din;
  assign PEG_Xvec_10_fifo_inst_out_full_n = PE_inst_11__full_n;
  assign Yvec_inst_10__din = PEG_Xvec_10_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_10_fifo_inst_out_to_Yvec_full_n = Yvec_inst_10__full_n;
  assign Yvec_inst_10__write = PEG_Xvec_10_fifo_inst_out_to_Yvec_write;
  assign PE_inst_11__write = PEG_Xvec_10_fifo_inst_out_write;
  assign PEG_Xvec_11_ap_clk = ap_clk;
  assign PEG_Xvec_11__ap_done = PEG_Xvec_11_ap_done;
  assign PEG_Xvec_11__ap_idle = PEG_Xvec_11_ap_idle;
  assign PEG_Xvec_11__ap_ready = PEG_Xvec_11_ap_ready;
  assign PEG_Xvec_11_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_11_ap_start = PEG_Xvec_11__ap_start;
  assign PEG_Xvec_11_fifo_A_peek_dout = fifo_A_11__dout;
  assign PEG_Xvec_11_fifo_A_peek_empty_n = fifo_A_11__empty_n;
  assign PEG_Xvec_11_fifo_A_s_dout = fifo_A_11__dout;
  assign PEG_Xvec_11_fifo_A_s_empty_n = fifo_A_11__empty_n;
  assign fifo_A_11__read = PEG_Xvec_11_fifo_A_s_read;
  assign PEG_Xvec_11_fifo_X_in_peek_dout = fifo_X_pe_11__dout;
  assign PEG_Xvec_11_fifo_X_in_peek_empty_n = fifo_X_pe_11__empty_n;
  assign PEG_Xvec_11_fifo_X_in_s_dout = fifo_X_pe_11__dout;
  assign PEG_Xvec_11_fifo_X_in_s_empty_n = fifo_X_pe_11__empty_n;
  assign fifo_X_pe_11__read = PEG_Xvec_11_fifo_X_in_s_read;
  assign fifo_X_pe_12__din = PEG_Xvec_11_fifo_X_out_din;
  assign PEG_Xvec_11_fifo_X_out_full_n = fifo_X_pe_12__full_n;
  assign fifo_X_pe_12__write = PEG_Xvec_11_fifo_X_out_write;
  assign fifo_aXvec_11__din = PEG_Xvec_11_fifo_aXvec_din;
  assign PEG_Xvec_11_fifo_aXvec_full_n = fifo_aXvec_11__full_n;
  assign fifo_aXvec_11__write = PEG_Xvec_11_fifo_aXvec_write;
  assign PEG_Xvec_11_fifo_inst_in_peek_dout = PE_inst_11__dout;
  assign PEG_Xvec_11_fifo_inst_in_peek_empty_n = PE_inst_11__empty_n;
  assign PEG_Xvec_11_fifo_inst_in_s_dout = PE_inst_11__dout;
  assign PEG_Xvec_11_fifo_inst_in_s_empty_n = PE_inst_11__empty_n;
  assign PE_inst_11__read = PEG_Xvec_11_fifo_inst_in_s_read;
  assign PE_inst_12__din = PEG_Xvec_11_fifo_inst_out_din;
  assign PEG_Xvec_11_fifo_inst_out_full_n = PE_inst_12__full_n;
  assign Yvec_inst_11__din = PEG_Xvec_11_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_11_fifo_inst_out_to_Yvec_full_n = Yvec_inst_11__full_n;
  assign Yvec_inst_11__write = PEG_Xvec_11_fifo_inst_out_to_Yvec_write;
  assign PE_inst_12__write = PEG_Xvec_11_fifo_inst_out_write;
  assign PEG_Xvec_12_ap_clk = ap_clk;
  assign PEG_Xvec_12__ap_done = PEG_Xvec_12_ap_done;
  assign PEG_Xvec_12__ap_idle = PEG_Xvec_12_ap_idle;
  assign PEG_Xvec_12__ap_ready = PEG_Xvec_12_ap_ready;
  assign PEG_Xvec_12_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_12_ap_start = PEG_Xvec_12__ap_start;
  assign PEG_Xvec_12_fifo_A_peek_dout = fifo_A_12__dout;
  assign PEG_Xvec_12_fifo_A_peek_empty_n = fifo_A_12__empty_n;
  assign PEG_Xvec_12_fifo_A_s_dout = fifo_A_12__dout;
  assign PEG_Xvec_12_fifo_A_s_empty_n = fifo_A_12__empty_n;
  assign fifo_A_12__read = PEG_Xvec_12_fifo_A_s_read;
  assign PEG_Xvec_12_fifo_X_in_peek_dout = fifo_X_pe_12__dout;
  assign PEG_Xvec_12_fifo_X_in_peek_empty_n = fifo_X_pe_12__empty_n;
  assign PEG_Xvec_12_fifo_X_in_s_dout = fifo_X_pe_12__dout;
  assign PEG_Xvec_12_fifo_X_in_s_empty_n = fifo_X_pe_12__empty_n;
  assign fifo_X_pe_12__read = PEG_Xvec_12_fifo_X_in_s_read;
  assign fifo_X_pe_13__din = PEG_Xvec_12_fifo_X_out_din;
  assign PEG_Xvec_12_fifo_X_out_full_n = fifo_X_pe_13__full_n;
  assign fifo_X_pe_13__write = PEG_Xvec_12_fifo_X_out_write;
  assign fifo_aXvec_12__din = PEG_Xvec_12_fifo_aXvec_din;
  assign PEG_Xvec_12_fifo_aXvec_full_n = fifo_aXvec_12__full_n;
  assign fifo_aXvec_12__write = PEG_Xvec_12_fifo_aXvec_write;
  assign PEG_Xvec_12_fifo_inst_in_peek_dout = PE_inst_12__dout;
  assign PEG_Xvec_12_fifo_inst_in_peek_empty_n = PE_inst_12__empty_n;
  assign PEG_Xvec_12_fifo_inst_in_s_dout = PE_inst_12__dout;
  assign PEG_Xvec_12_fifo_inst_in_s_empty_n = PE_inst_12__empty_n;
  assign PE_inst_12__read = PEG_Xvec_12_fifo_inst_in_s_read;
  assign PE_inst_13__din = PEG_Xvec_12_fifo_inst_out_din;
  assign PEG_Xvec_12_fifo_inst_out_full_n = PE_inst_13__full_n;
  assign Yvec_inst_12__din = PEG_Xvec_12_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_12_fifo_inst_out_to_Yvec_full_n = Yvec_inst_12__full_n;
  assign Yvec_inst_12__write = PEG_Xvec_12_fifo_inst_out_to_Yvec_write;
  assign PE_inst_13__write = PEG_Xvec_12_fifo_inst_out_write;
  assign PEG_Xvec_13_ap_clk = ap_clk;
  assign PEG_Xvec_13__ap_done = PEG_Xvec_13_ap_done;
  assign PEG_Xvec_13__ap_idle = PEG_Xvec_13_ap_idle;
  assign PEG_Xvec_13__ap_ready = PEG_Xvec_13_ap_ready;
  assign PEG_Xvec_13_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_13_ap_start = PEG_Xvec_13__ap_start;
  assign PEG_Xvec_13_fifo_A_peek_dout = fifo_A_13__dout;
  assign PEG_Xvec_13_fifo_A_peek_empty_n = fifo_A_13__empty_n;
  assign PEG_Xvec_13_fifo_A_s_dout = fifo_A_13__dout;
  assign PEG_Xvec_13_fifo_A_s_empty_n = fifo_A_13__empty_n;
  assign fifo_A_13__read = PEG_Xvec_13_fifo_A_s_read;
  assign PEG_Xvec_13_fifo_X_in_peek_dout = fifo_X_pe_13__dout;
  assign PEG_Xvec_13_fifo_X_in_peek_empty_n = fifo_X_pe_13__empty_n;
  assign PEG_Xvec_13_fifo_X_in_s_dout = fifo_X_pe_13__dout;
  assign PEG_Xvec_13_fifo_X_in_s_empty_n = fifo_X_pe_13__empty_n;
  assign fifo_X_pe_13__read = PEG_Xvec_13_fifo_X_in_s_read;
  assign fifo_X_pe_14__din = PEG_Xvec_13_fifo_X_out_din;
  assign PEG_Xvec_13_fifo_X_out_full_n = fifo_X_pe_14__full_n;
  assign fifo_X_pe_14__write = PEG_Xvec_13_fifo_X_out_write;
  assign fifo_aXvec_13__din = PEG_Xvec_13_fifo_aXvec_din;
  assign PEG_Xvec_13_fifo_aXvec_full_n = fifo_aXvec_13__full_n;
  assign fifo_aXvec_13__write = PEG_Xvec_13_fifo_aXvec_write;
  assign PEG_Xvec_13_fifo_inst_in_peek_dout = PE_inst_13__dout;
  assign PEG_Xvec_13_fifo_inst_in_peek_empty_n = PE_inst_13__empty_n;
  assign PEG_Xvec_13_fifo_inst_in_s_dout = PE_inst_13__dout;
  assign PEG_Xvec_13_fifo_inst_in_s_empty_n = PE_inst_13__empty_n;
  assign PE_inst_13__read = PEG_Xvec_13_fifo_inst_in_s_read;
  assign PE_inst_14__din = PEG_Xvec_13_fifo_inst_out_din;
  assign PEG_Xvec_13_fifo_inst_out_full_n = PE_inst_14__full_n;
  assign Yvec_inst_13__din = PEG_Xvec_13_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_13_fifo_inst_out_to_Yvec_full_n = Yvec_inst_13__full_n;
  assign Yvec_inst_13__write = PEG_Xvec_13_fifo_inst_out_to_Yvec_write;
  assign PE_inst_14__write = PEG_Xvec_13_fifo_inst_out_write;
  assign PEG_Xvec_14_ap_clk = ap_clk;
  assign PEG_Xvec_14__ap_done = PEG_Xvec_14_ap_done;
  assign PEG_Xvec_14__ap_idle = PEG_Xvec_14_ap_idle;
  assign PEG_Xvec_14__ap_ready = PEG_Xvec_14_ap_ready;
  assign PEG_Xvec_14_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_14_ap_start = PEG_Xvec_14__ap_start;
  assign PEG_Xvec_14_fifo_A_peek_dout = fifo_A_14__dout;
  assign PEG_Xvec_14_fifo_A_peek_empty_n = fifo_A_14__empty_n;
  assign PEG_Xvec_14_fifo_A_s_dout = fifo_A_14__dout;
  assign PEG_Xvec_14_fifo_A_s_empty_n = fifo_A_14__empty_n;
  assign fifo_A_14__read = PEG_Xvec_14_fifo_A_s_read;
  assign PEG_Xvec_14_fifo_X_in_peek_dout = fifo_X_pe_14__dout;
  assign PEG_Xvec_14_fifo_X_in_peek_empty_n = fifo_X_pe_14__empty_n;
  assign PEG_Xvec_14_fifo_X_in_s_dout = fifo_X_pe_14__dout;
  assign PEG_Xvec_14_fifo_X_in_s_empty_n = fifo_X_pe_14__empty_n;
  assign fifo_X_pe_14__read = PEG_Xvec_14_fifo_X_in_s_read;
  assign fifo_X_pe_15__din = PEG_Xvec_14_fifo_X_out_din;
  assign PEG_Xvec_14_fifo_X_out_full_n = fifo_X_pe_15__full_n;
  assign fifo_X_pe_15__write = PEG_Xvec_14_fifo_X_out_write;
  assign fifo_aXvec_14__din = PEG_Xvec_14_fifo_aXvec_din;
  assign PEG_Xvec_14_fifo_aXvec_full_n = fifo_aXvec_14__full_n;
  assign fifo_aXvec_14__write = PEG_Xvec_14_fifo_aXvec_write;
  assign PEG_Xvec_14_fifo_inst_in_peek_dout = PE_inst_14__dout;
  assign PEG_Xvec_14_fifo_inst_in_peek_empty_n = PE_inst_14__empty_n;
  assign PEG_Xvec_14_fifo_inst_in_s_dout = PE_inst_14__dout;
  assign PEG_Xvec_14_fifo_inst_in_s_empty_n = PE_inst_14__empty_n;
  assign PE_inst_14__read = PEG_Xvec_14_fifo_inst_in_s_read;
  assign PE_inst_15__din = PEG_Xvec_14_fifo_inst_out_din;
  assign PEG_Xvec_14_fifo_inst_out_full_n = PE_inst_15__full_n;
  assign Yvec_inst_14__din = PEG_Xvec_14_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_14_fifo_inst_out_to_Yvec_full_n = Yvec_inst_14__full_n;
  assign Yvec_inst_14__write = PEG_Xvec_14_fifo_inst_out_to_Yvec_write;
  assign PE_inst_15__write = PEG_Xvec_14_fifo_inst_out_write;
  assign PEG_Xvec_15_ap_clk = ap_clk;
  assign PEG_Xvec_15__ap_done = PEG_Xvec_15_ap_done;
  assign PEG_Xvec_15__ap_idle = PEG_Xvec_15_ap_idle;
  assign PEG_Xvec_15__ap_ready = PEG_Xvec_15_ap_ready;
  assign PEG_Xvec_15_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_15_ap_start = PEG_Xvec_15__ap_start;
  assign PEG_Xvec_15_fifo_A_peek_dout = fifo_A_15__dout;
  assign PEG_Xvec_15_fifo_A_peek_empty_n = fifo_A_15__empty_n;
  assign PEG_Xvec_15_fifo_A_s_dout = fifo_A_15__dout;
  assign PEG_Xvec_15_fifo_A_s_empty_n = fifo_A_15__empty_n;
  assign fifo_A_15__read = PEG_Xvec_15_fifo_A_s_read;
  assign PEG_Xvec_15_fifo_X_in_peek_dout = fifo_X_pe_15__dout;
  assign PEG_Xvec_15_fifo_X_in_peek_empty_n = fifo_X_pe_15__empty_n;
  assign PEG_Xvec_15_fifo_X_in_s_dout = fifo_X_pe_15__dout;
  assign PEG_Xvec_15_fifo_X_in_s_empty_n = fifo_X_pe_15__empty_n;
  assign fifo_X_pe_15__read = PEG_Xvec_15_fifo_X_in_s_read;
  assign fifo_X_pe_16__din = PEG_Xvec_15_fifo_X_out_din;
  assign PEG_Xvec_15_fifo_X_out_full_n = fifo_X_pe_16__full_n;
  assign fifo_X_pe_16__write = PEG_Xvec_15_fifo_X_out_write;
  assign fifo_aXvec_15__din = PEG_Xvec_15_fifo_aXvec_din;
  assign PEG_Xvec_15_fifo_aXvec_full_n = fifo_aXvec_15__full_n;
  assign fifo_aXvec_15__write = PEG_Xvec_15_fifo_aXvec_write;
  assign PEG_Xvec_15_fifo_inst_in_peek_dout = PE_inst_15__dout;
  assign PEG_Xvec_15_fifo_inst_in_peek_empty_n = PE_inst_15__empty_n;
  assign PEG_Xvec_15_fifo_inst_in_s_dout = PE_inst_15__dout;
  assign PEG_Xvec_15_fifo_inst_in_s_empty_n = PE_inst_15__empty_n;
  assign PE_inst_15__read = PEG_Xvec_15_fifo_inst_in_s_read;
  assign PE_inst_16__din = PEG_Xvec_15_fifo_inst_out_din;
  assign PEG_Xvec_15_fifo_inst_out_full_n = PE_inst_16__full_n;
  assign Yvec_inst_15__din = PEG_Xvec_15_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_15_fifo_inst_out_to_Yvec_full_n = Yvec_inst_15__full_n;
  assign Yvec_inst_15__write = PEG_Xvec_15_fifo_inst_out_to_Yvec_write;
  assign PE_inst_16__write = PEG_Xvec_15_fifo_inst_out_write;
  assign PEG_Xvec_16_ap_clk = ap_clk;
  assign PEG_Xvec_16__ap_done = PEG_Xvec_16_ap_done;
  assign PEG_Xvec_16__ap_idle = PEG_Xvec_16_ap_idle;
  assign PEG_Xvec_16__ap_ready = PEG_Xvec_16_ap_ready;
  assign PEG_Xvec_16_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_16_ap_start = PEG_Xvec_16__ap_start;
  assign PEG_Xvec_16_fifo_A_peek_dout = fifo_A_16__dout;
  assign PEG_Xvec_16_fifo_A_peek_empty_n = fifo_A_16__empty_n;
  assign PEG_Xvec_16_fifo_A_s_dout = fifo_A_16__dout;
  assign PEG_Xvec_16_fifo_A_s_empty_n = fifo_A_16__empty_n;
  assign fifo_A_16__read = PEG_Xvec_16_fifo_A_s_read;
  assign PEG_Xvec_16_fifo_X_in_peek_dout = fifo_X_pe_16__dout;
  assign PEG_Xvec_16_fifo_X_in_peek_empty_n = fifo_X_pe_16__empty_n;
  assign PEG_Xvec_16_fifo_X_in_s_dout = fifo_X_pe_16__dout;
  assign PEG_Xvec_16_fifo_X_in_s_empty_n = fifo_X_pe_16__empty_n;
  assign fifo_X_pe_16__read = PEG_Xvec_16_fifo_X_in_s_read;
  assign fifo_X_pe_17__din = PEG_Xvec_16_fifo_X_out_din;
  assign PEG_Xvec_16_fifo_X_out_full_n = fifo_X_pe_17__full_n;
  assign fifo_X_pe_17__write = PEG_Xvec_16_fifo_X_out_write;
  assign fifo_aXvec_16__din = PEG_Xvec_16_fifo_aXvec_din;
  assign PEG_Xvec_16_fifo_aXvec_full_n = fifo_aXvec_16__full_n;
  assign fifo_aXvec_16__write = PEG_Xvec_16_fifo_aXvec_write;
  assign PEG_Xvec_16_fifo_inst_in_peek_dout = PE_inst_16__dout;
  assign PEG_Xvec_16_fifo_inst_in_peek_empty_n = PE_inst_16__empty_n;
  assign PEG_Xvec_16_fifo_inst_in_s_dout = PE_inst_16__dout;
  assign PEG_Xvec_16_fifo_inst_in_s_empty_n = PE_inst_16__empty_n;
  assign PE_inst_16__read = PEG_Xvec_16_fifo_inst_in_s_read;
  assign PE_inst_17__din = PEG_Xvec_16_fifo_inst_out_din;
  assign PEG_Xvec_16_fifo_inst_out_full_n = PE_inst_17__full_n;
  assign Yvec_inst_16__din = PEG_Xvec_16_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_16_fifo_inst_out_to_Yvec_full_n = Yvec_inst_16__full_n;
  assign Yvec_inst_16__write = PEG_Xvec_16_fifo_inst_out_to_Yvec_write;
  assign PE_inst_17__write = PEG_Xvec_16_fifo_inst_out_write;
  assign PEG_Xvec_17_ap_clk = ap_clk;
  assign PEG_Xvec_17__ap_done = PEG_Xvec_17_ap_done;
  assign PEG_Xvec_17__ap_idle = PEG_Xvec_17_ap_idle;
  assign PEG_Xvec_17__ap_ready = PEG_Xvec_17_ap_ready;
  assign PEG_Xvec_17_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_17_ap_start = PEG_Xvec_17__ap_start;
  assign PEG_Xvec_17_fifo_A_peek_dout = fifo_A_17__dout;
  assign PEG_Xvec_17_fifo_A_peek_empty_n = fifo_A_17__empty_n;
  assign PEG_Xvec_17_fifo_A_s_dout = fifo_A_17__dout;
  assign PEG_Xvec_17_fifo_A_s_empty_n = fifo_A_17__empty_n;
  assign fifo_A_17__read = PEG_Xvec_17_fifo_A_s_read;
  assign PEG_Xvec_17_fifo_X_in_peek_dout = fifo_X_pe_17__dout;
  assign PEG_Xvec_17_fifo_X_in_peek_empty_n = fifo_X_pe_17__empty_n;
  assign PEG_Xvec_17_fifo_X_in_s_dout = fifo_X_pe_17__dout;
  assign PEG_Xvec_17_fifo_X_in_s_empty_n = fifo_X_pe_17__empty_n;
  assign fifo_X_pe_17__read = PEG_Xvec_17_fifo_X_in_s_read;
  assign fifo_X_pe_18__din = PEG_Xvec_17_fifo_X_out_din;
  assign PEG_Xvec_17_fifo_X_out_full_n = fifo_X_pe_18__full_n;
  assign fifo_X_pe_18__write = PEG_Xvec_17_fifo_X_out_write;
  assign fifo_aXvec_17__din = PEG_Xvec_17_fifo_aXvec_din;
  assign PEG_Xvec_17_fifo_aXvec_full_n = fifo_aXvec_17__full_n;
  assign fifo_aXvec_17__write = PEG_Xvec_17_fifo_aXvec_write;
  assign PEG_Xvec_17_fifo_inst_in_peek_dout = PE_inst_17__dout;
  assign PEG_Xvec_17_fifo_inst_in_peek_empty_n = PE_inst_17__empty_n;
  assign PEG_Xvec_17_fifo_inst_in_s_dout = PE_inst_17__dout;
  assign PEG_Xvec_17_fifo_inst_in_s_empty_n = PE_inst_17__empty_n;
  assign PE_inst_17__read = PEG_Xvec_17_fifo_inst_in_s_read;
  assign PE_inst_18__din = PEG_Xvec_17_fifo_inst_out_din;
  assign PEG_Xvec_17_fifo_inst_out_full_n = PE_inst_18__full_n;
  assign Yvec_inst_17__din = PEG_Xvec_17_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_17_fifo_inst_out_to_Yvec_full_n = Yvec_inst_17__full_n;
  assign Yvec_inst_17__write = PEG_Xvec_17_fifo_inst_out_to_Yvec_write;
  assign PE_inst_18__write = PEG_Xvec_17_fifo_inst_out_write;
  assign PEG_Xvec_18_ap_clk = ap_clk;
  assign PEG_Xvec_18__ap_done = PEG_Xvec_18_ap_done;
  assign PEG_Xvec_18__ap_idle = PEG_Xvec_18_ap_idle;
  assign PEG_Xvec_18__ap_ready = PEG_Xvec_18_ap_ready;
  assign PEG_Xvec_18_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_18_ap_start = PEG_Xvec_18__ap_start;
  assign PEG_Xvec_18_fifo_A_peek_dout = fifo_A_18__dout;
  assign PEG_Xvec_18_fifo_A_peek_empty_n = fifo_A_18__empty_n;
  assign PEG_Xvec_18_fifo_A_s_dout = fifo_A_18__dout;
  assign PEG_Xvec_18_fifo_A_s_empty_n = fifo_A_18__empty_n;
  assign fifo_A_18__read = PEG_Xvec_18_fifo_A_s_read;
  assign PEG_Xvec_18_fifo_X_in_peek_dout = fifo_X_pe_18__dout;
  assign PEG_Xvec_18_fifo_X_in_peek_empty_n = fifo_X_pe_18__empty_n;
  assign PEG_Xvec_18_fifo_X_in_s_dout = fifo_X_pe_18__dout;
  assign PEG_Xvec_18_fifo_X_in_s_empty_n = fifo_X_pe_18__empty_n;
  assign fifo_X_pe_18__read = PEG_Xvec_18_fifo_X_in_s_read;
  assign fifo_X_pe_19__din = PEG_Xvec_18_fifo_X_out_din;
  assign PEG_Xvec_18_fifo_X_out_full_n = fifo_X_pe_19__full_n;
  assign fifo_X_pe_19__write = PEG_Xvec_18_fifo_X_out_write;
  assign fifo_aXvec_18__din = PEG_Xvec_18_fifo_aXvec_din;
  assign PEG_Xvec_18_fifo_aXvec_full_n = fifo_aXvec_18__full_n;
  assign fifo_aXvec_18__write = PEG_Xvec_18_fifo_aXvec_write;
  assign PEG_Xvec_18_fifo_inst_in_peek_dout = PE_inst_18__dout;
  assign PEG_Xvec_18_fifo_inst_in_peek_empty_n = PE_inst_18__empty_n;
  assign PEG_Xvec_18_fifo_inst_in_s_dout = PE_inst_18__dout;
  assign PEG_Xvec_18_fifo_inst_in_s_empty_n = PE_inst_18__empty_n;
  assign PE_inst_18__read = PEG_Xvec_18_fifo_inst_in_s_read;
  assign PE_inst_19__din = PEG_Xvec_18_fifo_inst_out_din;
  assign PEG_Xvec_18_fifo_inst_out_full_n = PE_inst_19__full_n;
  assign Yvec_inst_18__din = PEG_Xvec_18_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_18_fifo_inst_out_to_Yvec_full_n = Yvec_inst_18__full_n;
  assign Yvec_inst_18__write = PEG_Xvec_18_fifo_inst_out_to_Yvec_write;
  assign PE_inst_19__write = PEG_Xvec_18_fifo_inst_out_write;
  assign PEG_Xvec_19_ap_clk = ap_clk;
  assign PEG_Xvec_19__ap_done = PEG_Xvec_19_ap_done;
  assign PEG_Xvec_19__ap_idle = PEG_Xvec_19_ap_idle;
  assign PEG_Xvec_19__ap_ready = PEG_Xvec_19_ap_ready;
  assign PEG_Xvec_19_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_19_ap_start = PEG_Xvec_19__ap_start;
  assign PEG_Xvec_19_fifo_A_peek_dout = fifo_A_19__dout;
  assign PEG_Xvec_19_fifo_A_peek_empty_n = fifo_A_19__empty_n;
  assign PEG_Xvec_19_fifo_A_s_dout = fifo_A_19__dout;
  assign PEG_Xvec_19_fifo_A_s_empty_n = fifo_A_19__empty_n;
  assign fifo_A_19__read = PEG_Xvec_19_fifo_A_s_read;
  assign PEG_Xvec_19_fifo_X_in_peek_dout = fifo_X_pe_19__dout;
  assign PEG_Xvec_19_fifo_X_in_peek_empty_n = fifo_X_pe_19__empty_n;
  assign PEG_Xvec_19_fifo_X_in_s_dout = fifo_X_pe_19__dout;
  assign PEG_Xvec_19_fifo_X_in_s_empty_n = fifo_X_pe_19__empty_n;
  assign fifo_X_pe_19__read = PEG_Xvec_19_fifo_X_in_s_read;
  assign fifo_X_pe_20__din = PEG_Xvec_19_fifo_X_out_din;
  assign PEG_Xvec_19_fifo_X_out_full_n = fifo_X_pe_20__full_n;
  assign fifo_X_pe_20__write = PEG_Xvec_19_fifo_X_out_write;
  assign fifo_aXvec_19__din = PEG_Xvec_19_fifo_aXvec_din;
  assign PEG_Xvec_19_fifo_aXvec_full_n = fifo_aXvec_19__full_n;
  assign fifo_aXvec_19__write = PEG_Xvec_19_fifo_aXvec_write;
  assign PEG_Xvec_19_fifo_inst_in_peek_dout = PE_inst_19__dout;
  assign PEG_Xvec_19_fifo_inst_in_peek_empty_n = PE_inst_19__empty_n;
  assign PEG_Xvec_19_fifo_inst_in_s_dout = PE_inst_19__dout;
  assign PEG_Xvec_19_fifo_inst_in_s_empty_n = PE_inst_19__empty_n;
  assign PE_inst_19__read = PEG_Xvec_19_fifo_inst_in_s_read;
  assign PE_inst_20__din = PEG_Xvec_19_fifo_inst_out_din;
  assign PEG_Xvec_19_fifo_inst_out_full_n = PE_inst_20__full_n;
  assign Yvec_inst_19__din = PEG_Xvec_19_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_19_fifo_inst_out_to_Yvec_full_n = Yvec_inst_19__full_n;
  assign Yvec_inst_19__write = PEG_Xvec_19_fifo_inst_out_to_Yvec_write;
  assign PE_inst_20__write = PEG_Xvec_19_fifo_inst_out_write;
  assign PEG_Xvec_20_ap_clk = ap_clk;
  assign PEG_Xvec_20__ap_done = PEG_Xvec_20_ap_done;
  assign PEG_Xvec_20__ap_idle = PEG_Xvec_20_ap_idle;
  assign PEG_Xvec_20__ap_ready = PEG_Xvec_20_ap_ready;
  assign PEG_Xvec_20_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_20_ap_start = PEG_Xvec_20__ap_start;
  assign PEG_Xvec_20_fifo_A_peek_dout = fifo_A_20__dout;
  assign PEG_Xvec_20_fifo_A_peek_empty_n = fifo_A_20__empty_n;
  assign PEG_Xvec_20_fifo_A_s_dout = fifo_A_20__dout;
  assign PEG_Xvec_20_fifo_A_s_empty_n = fifo_A_20__empty_n;
  assign fifo_A_20__read = PEG_Xvec_20_fifo_A_s_read;
  assign PEG_Xvec_20_fifo_X_in_peek_dout = fifo_X_pe_20__dout;
  assign PEG_Xvec_20_fifo_X_in_peek_empty_n = fifo_X_pe_20__empty_n;
  assign PEG_Xvec_20_fifo_X_in_s_dout = fifo_X_pe_20__dout;
  assign PEG_Xvec_20_fifo_X_in_s_empty_n = fifo_X_pe_20__empty_n;
  assign fifo_X_pe_20__read = PEG_Xvec_20_fifo_X_in_s_read;
  assign fifo_X_pe_21__din = PEG_Xvec_20_fifo_X_out_din;
  assign PEG_Xvec_20_fifo_X_out_full_n = fifo_X_pe_21__full_n;
  assign fifo_X_pe_21__write = PEG_Xvec_20_fifo_X_out_write;
  assign fifo_aXvec_20__din = PEG_Xvec_20_fifo_aXvec_din;
  assign PEG_Xvec_20_fifo_aXvec_full_n = fifo_aXvec_20__full_n;
  assign fifo_aXvec_20__write = PEG_Xvec_20_fifo_aXvec_write;
  assign PEG_Xvec_20_fifo_inst_in_peek_dout = PE_inst_20__dout;
  assign PEG_Xvec_20_fifo_inst_in_peek_empty_n = PE_inst_20__empty_n;
  assign PEG_Xvec_20_fifo_inst_in_s_dout = PE_inst_20__dout;
  assign PEG_Xvec_20_fifo_inst_in_s_empty_n = PE_inst_20__empty_n;
  assign PE_inst_20__read = PEG_Xvec_20_fifo_inst_in_s_read;
  assign PE_inst_21__din = PEG_Xvec_20_fifo_inst_out_din;
  assign PEG_Xvec_20_fifo_inst_out_full_n = PE_inst_21__full_n;
  assign Yvec_inst_20__din = PEG_Xvec_20_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_20_fifo_inst_out_to_Yvec_full_n = Yvec_inst_20__full_n;
  assign Yvec_inst_20__write = PEG_Xvec_20_fifo_inst_out_to_Yvec_write;
  assign PE_inst_21__write = PEG_Xvec_20_fifo_inst_out_write;
  assign PEG_Xvec_21_ap_clk = ap_clk;
  assign PEG_Xvec_21__ap_done = PEG_Xvec_21_ap_done;
  assign PEG_Xvec_21__ap_idle = PEG_Xvec_21_ap_idle;
  assign PEG_Xvec_21__ap_ready = PEG_Xvec_21_ap_ready;
  assign PEG_Xvec_21_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_21_ap_start = PEG_Xvec_21__ap_start;
  assign PEG_Xvec_21_fifo_A_peek_dout = fifo_A_21__dout;
  assign PEG_Xvec_21_fifo_A_peek_empty_n = fifo_A_21__empty_n;
  assign PEG_Xvec_21_fifo_A_s_dout = fifo_A_21__dout;
  assign PEG_Xvec_21_fifo_A_s_empty_n = fifo_A_21__empty_n;
  assign fifo_A_21__read = PEG_Xvec_21_fifo_A_s_read;
  assign PEG_Xvec_21_fifo_X_in_peek_dout = fifo_X_pe_21__dout;
  assign PEG_Xvec_21_fifo_X_in_peek_empty_n = fifo_X_pe_21__empty_n;
  assign PEG_Xvec_21_fifo_X_in_s_dout = fifo_X_pe_21__dout;
  assign PEG_Xvec_21_fifo_X_in_s_empty_n = fifo_X_pe_21__empty_n;
  assign fifo_X_pe_21__read = PEG_Xvec_21_fifo_X_in_s_read;
  assign fifo_X_pe_22__din = PEG_Xvec_21_fifo_X_out_din;
  assign PEG_Xvec_21_fifo_X_out_full_n = fifo_X_pe_22__full_n;
  assign fifo_X_pe_22__write = PEG_Xvec_21_fifo_X_out_write;
  assign fifo_aXvec_21__din = PEG_Xvec_21_fifo_aXvec_din;
  assign PEG_Xvec_21_fifo_aXvec_full_n = fifo_aXvec_21__full_n;
  assign fifo_aXvec_21__write = PEG_Xvec_21_fifo_aXvec_write;
  assign PEG_Xvec_21_fifo_inst_in_peek_dout = PE_inst_21__dout;
  assign PEG_Xvec_21_fifo_inst_in_peek_empty_n = PE_inst_21__empty_n;
  assign PEG_Xvec_21_fifo_inst_in_s_dout = PE_inst_21__dout;
  assign PEG_Xvec_21_fifo_inst_in_s_empty_n = PE_inst_21__empty_n;
  assign PE_inst_21__read = PEG_Xvec_21_fifo_inst_in_s_read;
  assign PE_inst_22__din = PEG_Xvec_21_fifo_inst_out_din;
  assign PEG_Xvec_21_fifo_inst_out_full_n = PE_inst_22__full_n;
  assign Yvec_inst_21__din = PEG_Xvec_21_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_21_fifo_inst_out_to_Yvec_full_n = Yvec_inst_21__full_n;
  assign Yvec_inst_21__write = PEG_Xvec_21_fifo_inst_out_to_Yvec_write;
  assign PE_inst_22__write = PEG_Xvec_21_fifo_inst_out_write;
  assign PEG_Xvec_22_ap_clk = ap_clk;
  assign PEG_Xvec_22__ap_done = PEG_Xvec_22_ap_done;
  assign PEG_Xvec_22__ap_idle = PEG_Xvec_22_ap_idle;
  assign PEG_Xvec_22__ap_ready = PEG_Xvec_22_ap_ready;
  assign PEG_Xvec_22_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_22_ap_start = PEG_Xvec_22__ap_start;
  assign PEG_Xvec_22_fifo_A_peek_dout = fifo_A_22__dout;
  assign PEG_Xvec_22_fifo_A_peek_empty_n = fifo_A_22__empty_n;
  assign PEG_Xvec_22_fifo_A_s_dout = fifo_A_22__dout;
  assign PEG_Xvec_22_fifo_A_s_empty_n = fifo_A_22__empty_n;
  assign fifo_A_22__read = PEG_Xvec_22_fifo_A_s_read;
  assign PEG_Xvec_22_fifo_X_in_peek_dout = fifo_X_pe_22__dout;
  assign PEG_Xvec_22_fifo_X_in_peek_empty_n = fifo_X_pe_22__empty_n;
  assign PEG_Xvec_22_fifo_X_in_s_dout = fifo_X_pe_22__dout;
  assign PEG_Xvec_22_fifo_X_in_s_empty_n = fifo_X_pe_22__empty_n;
  assign fifo_X_pe_22__read = PEG_Xvec_22_fifo_X_in_s_read;
  assign fifo_X_pe_23__din = PEG_Xvec_22_fifo_X_out_din;
  assign PEG_Xvec_22_fifo_X_out_full_n = fifo_X_pe_23__full_n;
  assign fifo_X_pe_23__write = PEG_Xvec_22_fifo_X_out_write;
  assign fifo_aXvec_22__din = PEG_Xvec_22_fifo_aXvec_din;
  assign PEG_Xvec_22_fifo_aXvec_full_n = fifo_aXvec_22__full_n;
  assign fifo_aXvec_22__write = PEG_Xvec_22_fifo_aXvec_write;
  assign PEG_Xvec_22_fifo_inst_in_peek_dout = PE_inst_22__dout;
  assign PEG_Xvec_22_fifo_inst_in_peek_empty_n = PE_inst_22__empty_n;
  assign PEG_Xvec_22_fifo_inst_in_s_dout = PE_inst_22__dout;
  assign PEG_Xvec_22_fifo_inst_in_s_empty_n = PE_inst_22__empty_n;
  assign PE_inst_22__read = PEG_Xvec_22_fifo_inst_in_s_read;
  assign PE_inst_23__din = PEG_Xvec_22_fifo_inst_out_din;
  assign PEG_Xvec_22_fifo_inst_out_full_n = PE_inst_23__full_n;
  assign Yvec_inst_22__din = PEG_Xvec_22_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_22_fifo_inst_out_to_Yvec_full_n = Yvec_inst_22__full_n;
  assign Yvec_inst_22__write = PEG_Xvec_22_fifo_inst_out_to_Yvec_write;
  assign PE_inst_23__write = PEG_Xvec_22_fifo_inst_out_write;
  assign PEG_Xvec_23_ap_clk = ap_clk;
  assign PEG_Xvec_23__ap_done = PEG_Xvec_23_ap_done;
  assign PEG_Xvec_23__ap_idle = PEG_Xvec_23_ap_idle;
  assign PEG_Xvec_23__ap_ready = PEG_Xvec_23_ap_ready;
  assign PEG_Xvec_23_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_23_ap_start = PEG_Xvec_23__ap_start;
  assign PEG_Xvec_23_fifo_A_peek_dout = fifo_A_23__dout;
  assign PEG_Xvec_23_fifo_A_peek_empty_n = fifo_A_23__empty_n;
  assign PEG_Xvec_23_fifo_A_s_dout = fifo_A_23__dout;
  assign PEG_Xvec_23_fifo_A_s_empty_n = fifo_A_23__empty_n;
  assign fifo_A_23__read = PEG_Xvec_23_fifo_A_s_read;
  assign PEG_Xvec_23_fifo_X_in_peek_dout = fifo_X_pe_23__dout;
  assign PEG_Xvec_23_fifo_X_in_peek_empty_n = fifo_X_pe_23__empty_n;
  assign PEG_Xvec_23_fifo_X_in_s_dout = fifo_X_pe_23__dout;
  assign PEG_Xvec_23_fifo_X_in_s_empty_n = fifo_X_pe_23__empty_n;
  assign fifo_X_pe_23__read = PEG_Xvec_23_fifo_X_in_s_read;
  assign fifo_X_pe_24__din = PEG_Xvec_23_fifo_X_out_din;
  assign PEG_Xvec_23_fifo_X_out_full_n = fifo_X_pe_24__full_n;
  assign fifo_X_pe_24__write = PEG_Xvec_23_fifo_X_out_write;
  assign fifo_aXvec_23__din = PEG_Xvec_23_fifo_aXvec_din;
  assign PEG_Xvec_23_fifo_aXvec_full_n = fifo_aXvec_23__full_n;
  assign fifo_aXvec_23__write = PEG_Xvec_23_fifo_aXvec_write;
  assign PEG_Xvec_23_fifo_inst_in_peek_dout = PE_inst_23__dout;
  assign PEG_Xvec_23_fifo_inst_in_peek_empty_n = PE_inst_23__empty_n;
  assign PEG_Xvec_23_fifo_inst_in_s_dout = PE_inst_23__dout;
  assign PEG_Xvec_23_fifo_inst_in_s_empty_n = PE_inst_23__empty_n;
  assign PE_inst_23__read = PEG_Xvec_23_fifo_inst_in_s_read;
  assign PE_inst_24__din = PEG_Xvec_23_fifo_inst_out_din;
  assign PEG_Xvec_23_fifo_inst_out_full_n = PE_inst_24__full_n;
  assign Yvec_inst_23__din = PEG_Xvec_23_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_23_fifo_inst_out_to_Yvec_full_n = Yvec_inst_23__full_n;
  assign Yvec_inst_23__write = PEG_Xvec_23_fifo_inst_out_to_Yvec_write;
  assign PE_inst_24__write = PEG_Xvec_23_fifo_inst_out_write;
  assign PEG_Xvec_24_ap_clk = ap_clk;
  assign PEG_Xvec_24__ap_done = PEG_Xvec_24_ap_done;
  assign PEG_Xvec_24__ap_idle = PEG_Xvec_24_ap_idle;
  assign PEG_Xvec_24__ap_ready = PEG_Xvec_24_ap_ready;
  assign PEG_Xvec_24_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_24_ap_start = PEG_Xvec_24__ap_start;
  assign PEG_Xvec_24_fifo_A_peek_dout = fifo_A_24__dout;
  assign PEG_Xvec_24_fifo_A_peek_empty_n = fifo_A_24__empty_n;
  assign PEG_Xvec_24_fifo_A_s_dout = fifo_A_24__dout;
  assign PEG_Xvec_24_fifo_A_s_empty_n = fifo_A_24__empty_n;
  assign fifo_A_24__read = PEG_Xvec_24_fifo_A_s_read;
  assign PEG_Xvec_24_fifo_X_in_peek_dout = fifo_X_pe_24__dout;
  assign PEG_Xvec_24_fifo_X_in_peek_empty_n = fifo_X_pe_24__empty_n;
  assign PEG_Xvec_24_fifo_X_in_s_dout = fifo_X_pe_24__dout;
  assign PEG_Xvec_24_fifo_X_in_s_empty_n = fifo_X_pe_24__empty_n;
  assign fifo_X_pe_24__read = PEG_Xvec_24_fifo_X_in_s_read;
  assign fifo_X_pe_25__din = PEG_Xvec_24_fifo_X_out_din;
  assign PEG_Xvec_24_fifo_X_out_full_n = fifo_X_pe_25__full_n;
  assign fifo_X_pe_25__write = PEG_Xvec_24_fifo_X_out_write;
  assign fifo_aXvec_24__din = PEG_Xvec_24_fifo_aXvec_din;
  assign PEG_Xvec_24_fifo_aXvec_full_n = fifo_aXvec_24__full_n;
  assign fifo_aXvec_24__write = PEG_Xvec_24_fifo_aXvec_write;
  assign PEG_Xvec_24_fifo_inst_in_peek_dout = PE_inst_24__dout;
  assign PEG_Xvec_24_fifo_inst_in_peek_empty_n = PE_inst_24__empty_n;
  assign PEG_Xvec_24_fifo_inst_in_s_dout = PE_inst_24__dout;
  assign PEG_Xvec_24_fifo_inst_in_s_empty_n = PE_inst_24__empty_n;
  assign PE_inst_24__read = PEG_Xvec_24_fifo_inst_in_s_read;
  assign PE_inst_25__din = PEG_Xvec_24_fifo_inst_out_din;
  assign PEG_Xvec_24_fifo_inst_out_full_n = PE_inst_25__full_n;
  assign Yvec_inst_24__din = PEG_Xvec_24_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_24_fifo_inst_out_to_Yvec_full_n = Yvec_inst_24__full_n;
  assign Yvec_inst_24__write = PEG_Xvec_24_fifo_inst_out_to_Yvec_write;
  assign PE_inst_25__write = PEG_Xvec_24_fifo_inst_out_write;
  assign PEG_Xvec_25_ap_clk = ap_clk;
  assign PEG_Xvec_25__ap_done = PEG_Xvec_25_ap_done;
  assign PEG_Xvec_25__ap_idle = PEG_Xvec_25_ap_idle;
  assign PEG_Xvec_25__ap_ready = PEG_Xvec_25_ap_ready;
  assign PEG_Xvec_25_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_25_ap_start = PEG_Xvec_25__ap_start;
  assign PEG_Xvec_25_fifo_A_peek_dout = fifo_A_25__dout;
  assign PEG_Xvec_25_fifo_A_peek_empty_n = fifo_A_25__empty_n;
  assign PEG_Xvec_25_fifo_A_s_dout = fifo_A_25__dout;
  assign PEG_Xvec_25_fifo_A_s_empty_n = fifo_A_25__empty_n;
  assign fifo_A_25__read = PEG_Xvec_25_fifo_A_s_read;
  assign PEG_Xvec_25_fifo_X_in_peek_dout = fifo_X_pe_25__dout;
  assign PEG_Xvec_25_fifo_X_in_peek_empty_n = fifo_X_pe_25__empty_n;
  assign PEG_Xvec_25_fifo_X_in_s_dout = fifo_X_pe_25__dout;
  assign PEG_Xvec_25_fifo_X_in_s_empty_n = fifo_X_pe_25__empty_n;
  assign fifo_X_pe_25__read = PEG_Xvec_25_fifo_X_in_s_read;
  assign fifo_X_pe_26__din = PEG_Xvec_25_fifo_X_out_din;
  assign PEG_Xvec_25_fifo_X_out_full_n = fifo_X_pe_26__full_n;
  assign fifo_X_pe_26__write = PEG_Xvec_25_fifo_X_out_write;
  assign fifo_aXvec_25__din = PEG_Xvec_25_fifo_aXvec_din;
  assign PEG_Xvec_25_fifo_aXvec_full_n = fifo_aXvec_25__full_n;
  assign fifo_aXvec_25__write = PEG_Xvec_25_fifo_aXvec_write;
  assign PEG_Xvec_25_fifo_inst_in_peek_dout = PE_inst_25__dout;
  assign PEG_Xvec_25_fifo_inst_in_peek_empty_n = PE_inst_25__empty_n;
  assign PEG_Xvec_25_fifo_inst_in_s_dout = PE_inst_25__dout;
  assign PEG_Xvec_25_fifo_inst_in_s_empty_n = PE_inst_25__empty_n;
  assign PE_inst_25__read = PEG_Xvec_25_fifo_inst_in_s_read;
  assign PE_inst_26__din = PEG_Xvec_25_fifo_inst_out_din;
  assign PEG_Xvec_25_fifo_inst_out_full_n = PE_inst_26__full_n;
  assign Yvec_inst_25__din = PEG_Xvec_25_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_25_fifo_inst_out_to_Yvec_full_n = Yvec_inst_25__full_n;
  assign Yvec_inst_25__write = PEG_Xvec_25_fifo_inst_out_to_Yvec_write;
  assign PE_inst_26__write = PEG_Xvec_25_fifo_inst_out_write;
  assign PEG_Xvec_26_ap_clk = ap_clk;
  assign PEG_Xvec_26__ap_done = PEG_Xvec_26_ap_done;
  assign PEG_Xvec_26__ap_idle = PEG_Xvec_26_ap_idle;
  assign PEG_Xvec_26__ap_ready = PEG_Xvec_26_ap_ready;
  assign PEG_Xvec_26_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_26_ap_start = PEG_Xvec_26__ap_start;
  assign PEG_Xvec_26_fifo_A_peek_dout = fifo_A_26__dout;
  assign PEG_Xvec_26_fifo_A_peek_empty_n = fifo_A_26__empty_n;
  assign PEG_Xvec_26_fifo_A_s_dout = fifo_A_26__dout;
  assign PEG_Xvec_26_fifo_A_s_empty_n = fifo_A_26__empty_n;
  assign fifo_A_26__read = PEG_Xvec_26_fifo_A_s_read;
  assign PEG_Xvec_26_fifo_X_in_peek_dout = fifo_X_pe_26__dout;
  assign PEG_Xvec_26_fifo_X_in_peek_empty_n = fifo_X_pe_26__empty_n;
  assign PEG_Xvec_26_fifo_X_in_s_dout = fifo_X_pe_26__dout;
  assign PEG_Xvec_26_fifo_X_in_s_empty_n = fifo_X_pe_26__empty_n;
  assign fifo_X_pe_26__read = PEG_Xvec_26_fifo_X_in_s_read;
  assign fifo_X_pe_27__din = PEG_Xvec_26_fifo_X_out_din;
  assign PEG_Xvec_26_fifo_X_out_full_n = fifo_X_pe_27__full_n;
  assign fifo_X_pe_27__write = PEG_Xvec_26_fifo_X_out_write;
  assign fifo_aXvec_26__din = PEG_Xvec_26_fifo_aXvec_din;
  assign PEG_Xvec_26_fifo_aXvec_full_n = fifo_aXvec_26__full_n;
  assign fifo_aXvec_26__write = PEG_Xvec_26_fifo_aXvec_write;
  assign PEG_Xvec_26_fifo_inst_in_peek_dout = PE_inst_26__dout;
  assign PEG_Xvec_26_fifo_inst_in_peek_empty_n = PE_inst_26__empty_n;
  assign PEG_Xvec_26_fifo_inst_in_s_dout = PE_inst_26__dout;
  assign PEG_Xvec_26_fifo_inst_in_s_empty_n = PE_inst_26__empty_n;
  assign PE_inst_26__read = PEG_Xvec_26_fifo_inst_in_s_read;
  assign PE_inst_27__din = PEG_Xvec_26_fifo_inst_out_din;
  assign PEG_Xvec_26_fifo_inst_out_full_n = PE_inst_27__full_n;
  assign Yvec_inst_26__din = PEG_Xvec_26_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_26_fifo_inst_out_to_Yvec_full_n = Yvec_inst_26__full_n;
  assign Yvec_inst_26__write = PEG_Xvec_26_fifo_inst_out_to_Yvec_write;
  assign PE_inst_27__write = PEG_Xvec_26_fifo_inst_out_write;
  assign PEG_Xvec_27_ap_clk = ap_clk;
  assign PEG_Xvec_27__ap_done = PEG_Xvec_27_ap_done;
  assign PEG_Xvec_27__ap_idle = PEG_Xvec_27_ap_idle;
  assign PEG_Xvec_27__ap_ready = PEG_Xvec_27_ap_ready;
  assign PEG_Xvec_27_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_27_ap_start = PEG_Xvec_27__ap_start;
  assign PEG_Xvec_27_fifo_A_peek_dout = fifo_A_27__dout;
  assign PEG_Xvec_27_fifo_A_peek_empty_n = fifo_A_27__empty_n;
  assign PEG_Xvec_27_fifo_A_s_dout = fifo_A_27__dout;
  assign PEG_Xvec_27_fifo_A_s_empty_n = fifo_A_27__empty_n;
  assign fifo_A_27__read = PEG_Xvec_27_fifo_A_s_read;
  assign PEG_Xvec_27_fifo_X_in_peek_dout = fifo_X_pe_27__dout;
  assign PEG_Xvec_27_fifo_X_in_peek_empty_n = fifo_X_pe_27__empty_n;
  assign PEG_Xvec_27_fifo_X_in_s_dout = fifo_X_pe_27__dout;
  assign PEG_Xvec_27_fifo_X_in_s_empty_n = fifo_X_pe_27__empty_n;
  assign fifo_X_pe_27__read = PEG_Xvec_27_fifo_X_in_s_read;
  assign fifo_X_pe_28__din = PEG_Xvec_27_fifo_X_out_din;
  assign PEG_Xvec_27_fifo_X_out_full_n = fifo_X_pe_28__full_n;
  assign fifo_X_pe_28__write = PEG_Xvec_27_fifo_X_out_write;
  assign fifo_aXvec_27__din = PEG_Xvec_27_fifo_aXvec_din;
  assign PEG_Xvec_27_fifo_aXvec_full_n = fifo_aXvec_27__full_n;
  assign fifo_aXvec_27__write = PEG_Xvec_27_fifo_aXvec_write;
  assign PEG_Xvec_27_fifo_inst_in_peek_dout = PE_inst_27__dout;
  assign PEG_Xvec_27_fifo_inst_in_peek_empty_n = PE_inst_27__empty_n;
  assign PEG_Xvec_27_fifo_inst_in_s_dout = PE_inst_27__dout;
  assign PEG_Xvec_27_fifo_inst_in_s_empty_n = PE_inst_27__empty_n;
  assign PE_inst_27__read = PEG_Xvec_27_fifo_inst_in_s_read;
  assign PE_inst_28__din = PEG_Xvec_27_fifo_inst_out_din;
  assign PEG_Xvec_27_fifo_inst_out_full_n = PE_inst_28__full_n;
  assign Yvec_inst_27__din = PEG_Xvec_27_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_27_fifo_inst_out_to_Yvec_full_n = Yvec_inst_27__full_n;
  assign Yvec_inst_27__write = PEG_Xvec_27_fifo_inst_out_to_Yvec_write;
  assign PE_inst_28__write = PEG_Xvec_27_fifo_inst_out_write;
  assign PEG_Xvec_28_ap_clk = ap_clk;
  assign PEG_Xvec_28__ap_done = PEG_Xvec_28_ap_done;
  assign PEG_Xvec_28__ap_idle = PEG_Xvec_28_ap_idle;
  assign PEG_Xvec_28__ap_ready = PEG_Xvec_28_ap_ready;
  assign PEG_Xvec_28_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_28_ap_start = PEG_Xvec_28__ap_start;
  assign PEG_Xvec_28_fifo_A_peek_dout = fifo_A_28__dout;
  assign PEG_Xvec_28_fifo_A_peek_empty_n = fifo_A_28__empty_n;
  assign PEG_Xvec_28_fifo_A_s_dout = fifo_A_28__dout;
  assign PEG_Xvec_28_fifo_A_s_empty_n = fifo_A_28__empty_n;
  assign fifo_A_28__read = PEG_Xvec_28_fifo_A_s_read;
  assign PEG_Xvec_28_fifo_X_in_peek_dout = fifo_X_pe_28__dout;
  assign PEG_Xvec_28_fifo_X_in_peek_empty_n = fifo_X_pe_28__empty_n;
  assign PEG_Xvec_28_fifo_X_in_s_dout = fifo_X_pe_28__dout;
  assign PEG_Xvec_28_fifo_X_in_s_empty_n = fifo_X_pe_28__empty_n;
  assign fifo_X_pe_28__read = PEG_Xvec_28_fifo_X_in_s_read;
  assign fifo_X_pe_29__din = PEG_Xvec_28_fifo_X_out_din;
  assign PEG_Xvec_28_fifo_X_out_full_n = fifo_X_pe_29__full_n;
  assign fifo_X_pe_29__write = PEG_Xvec_28_fifo_X_out_write;
  assign fifo_aXvec_28__din = PEG_Xvec_28_fifo_aXvec_din;
  assign PEG_Xvec_28_fifo_aXvec_full_n = fifo_aXvec_28__full_n;
  assign fifo_aXvec_28__write = PEG_Xvec_28_fifo_aXvec_write;
  assign PEG_Xvec_28_fifo_inst_in_peek_dout = PE_inst_28__dout;
  assign PEG_Xvec_28_fifo_inst_in_peek_empty_n = PE_inst_28__empty_n;
  assign PEG_Xvec_28_fifo_inst_in_s_dout = PE_inst_28__dout;
  assign PEG_Xvec_28_fifo_inst_in_s_empty_n = PE_inst_28__empty_n;
  assign PE_inst_28__read = PEG_Xvec_28_fifo_inst_in_s_read;
  assign PE_inst_29__din = PEG_Xvec_28_fifo_inst_out_din;
  assign PEG_Xvec_28_fifo_inst_out_full_n = PE_inst_29__full_n;
  assign Yvec_inst_28__din = PEG_Xvec_28_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_28_fifo_inst_out_to_Yvec_full_n = Yvec_inst_28__full_n;
  assign Yvec_inst_28__write = PEG_Xvec_28_fifo_inst_out_to_Yvec_write;
  assign PE_inst_29__write = PEG_Xvec_28_fifo_inst_out_write;
  assign PEG_Xvec_29_ap_clk = ap_clk;
  assign PEG_Xvec_29__ap_done = PEG_Xvec_29_ap_done;
  assign PEG_Xvec_29__ap_idle = PEG_Xvec_29_ap_idle;
  assign PEG_Xvec_29__ap_ready = PEG_Xvec_29_ap_ready;
  assign PEG_Xvec_29_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_29_ap_start = PEG_Xvec_29__ap_start;
  assign PEG_Xvec_29_fifo_A_peek_dout = fifo_A_29__dout;
  assign PEG_Xvec_29_fifo_A_peek_empty_n = fifo_A_29__empty_n;
  assign PEG_Xvec_29_fifo_A_s_dout = fifo_A_29__dout;
  assign PEG_Xvec_29_fifo_A_s_empty_n = fifo_A_29__empty_n;
  assign fifo_A_29__read = PEG_Xvec_29_fifo_A_s_read;
  assign PEG_Xvec_29_fifo_X_in_peek_dout = fifo_X_pe_29__dout;
  assign PEG_Xvec_29_fifo_X_in_peek_empty_n = fifo_X_pe_29__empty_n;
  assign PEG_Xvec_29_fifo_X_in_s_dout = fifo_X_pe_29__dout;
  assign PEG_Xvec_29_fifo_X_in_s_empty_n = fifo_X_pe_29__empty_n;
  assign fifo_X_pe_29__read = PEG_Xvec_29_fifo_X_in_s_read;
  assign fifo_X_pe_30__din = PEG_Xvec_29_fifo_X_out_din;
  assign PEG_Xvec_29_fifo_X_out_full_n = fifo_X_pe_30__full_n;
  assign fifo_X_pe_30__write = PEG_Xvec_29_fifo_X_out_write;
  assign fifo_aXvec_29__din = PEG_Xvec_29_fifo_aXvec_din;
  assign PEG_Xvec_29_fifo_aXvec_full_n = fifo_aXvec_29__full_n;
  assign fifo_aXvec_29__write = PEG_Xvec_29_fifo_aXvec_write;
  assign PEG_Xvec_29_fifo_inst_in_peek_dout = PE_inst_29__dout;
  assign PEG_Xvec_29_fifo_inst_in_peek_empty_n = PE_inst_29__empty_n;
  assign PEG_Xvec_29_fifo_inst_in_s_dout = PE_inst_29__dout;
  assign PEG_Xvec_29_fifo_inst_in_s_empty_n = PE_inst_29__empty_n;
  assign PE_inst_29__read = PEG_Xvec_29_fifo_inst_in_s_read;
  assign PE_inst_30__din = PEG_Xvec_29_fifo_inst_out_din;
  assign PEG_Xvec_29_fifo_inst_out_full_n = PE_inst_30__full_n;
  assign Yvec_inst_29__din = PEG_Xvec_29_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_29_fifo_inst_out_to_Yvec_full_n = Yvec_inst_29__full_n;
  assign Yvec_inst_29__write = PEG_Xvec_29_fifo_inst_out_to_Yvec_write;
  assign PE_inst_30__write = PEG_Xvec_29_fifo_inst_out_write;
  assign PEG_Xvec_30_ap_clk = ap_clk;
  assign PEG_Xvec_30__ap_done = PEG_Xvec_30_ap_done;
  assign PEG_Xvec_30__ap_idle = PEG_Xvec_30_ap_idle;
  assign PEG_Xvec_30__ap_ready = PEG_Xvec_30_ap_ready;
  assign PEG_Xvec_30_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_30_ap_start = PEG_Xvec_30__ap_start;
  assign PEG_Xvec_30_fifo_A_peek_dout = fifo_A_30__dout;
  assign PEG_Xvec_30_fifo_A_peek_empty_n = fifo_A_30__empty_n;
  assign PEG_Xvec_30_fifo_A_s_dout = fifo_A_30__dout;
  assign PEG_Xvec_30_fifo_A_s_empty_n = fifo_A_30__empty_n;
  assign fifo_A_30__read = PEG_Xvec_30_fifo_A_s_read;
  assign PEG_Xvec_30_fifo_X_in_peek_dout = fifo_X_pe_30__dout;
  assign PEG_Xvec_30_fifo_X_in_peek_empty_n = fifo_X_pe_30__empty_n;
  assign PEG_Xvec_30_fifo_X_in_s_dout = fifo_X_pe_30__dout;
  assign PEG_Xvec_30_fifo_X_in_s_empty_n = fifo_X_pe_30__empty_n;
  assign fifo_X_pe_30__read = PEG_Xvec_30_fifo_X_in_s_read;
  assign fifo_X_pe_31__din = PEG_Xvec_30_fifo_X_out_din;
  assign PEG_Xvec_30_fifo_X_out_full_n = fifo_X_pe_31__full_n;
  assign fifo_X_pe_31__write = PEG_Xvec_30_fifo_X_out_write;
  assign fifo_aXvec_30__din = PEG_Xvec_30_fifo_aXvec_din;
  assign PEG_Xvec_30_fifo_aXvec_full_n = fifo_aXvec_30__full_n;
  assign fifo_aXvec_30__write = PEG_Xvec_30_fifo_aXvec_write;
  assign PEG_Xvec_30_fifo_inst_in_peek_dout = PE_inst_30__dout;
  assign PEG_Xvec_30_fifo_inst_in_peek_empty_n = PE_inst_30__empty_n;
  assign PEG_Xvec_30_fifo_inst_in_s_dout = PE_inst_30__dout;
  assign PEG_Xvec_30_fifo_inst_in_s_empty_n = PE_inst_30__empty_n;
  assign PE_inst_30__read = PEG_Xvec_30_fifo_inst_in_s_read;
  assign PE_inst_31__din = PEG_Xvec_30_fifo_inst_out_din;
  assign PEG_Xvec_30_fifo_inst_out_full_n = PE_inst_31__full_n;
  assign Yvec_inst_30__din = PEG_Xvec_30_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_30_fifo_inst_out_to_Yvec_full_n = Yvec_inst_30__full_n;
  assign Yvec_inst_30__write = PEG_Xvec_30_fifo_inst_out_to_Yvec_write;
  assign PE_inst_31__write = PEG_Xvec_30_fifo_inst_out_write;
  assign PEG_Xvec_31_ap_clk = ap_clk;
  assign PEG_Xvec_31__ap_done = PEG_Xvec_31_ap_done;
  assign PEG_Xvec_31__ap_idle = PEG_Xvec_31_ap_idle;
  assign PEG_Xvec_31__ap_ready = PEG_Xvec_31_ap_ready;
  assign PEG_Xvec_31_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_31_ap_start = PEG_Xvec_31__ap_start;
  assign PEG_Xvec_31_fifo_A_peek_dout = fifo_A_31__dout;
  assign PEG_Xvec_31_fifo_A_peek_empty_n = fifo_A_31__empty_n;
  assign PEG_Xvec_31_fifo_A_s_dout = fifo_A_31__dout;
  assign PEG_Xvec_31_fifo_A_s_empty_n = fifo_A_31__empty_n;
  assign fifo_A_31__read = PEG_Xvec_31_fifo_A_s_read;
  assign PEG_Xvec_31_fifo_X_in_peek_dout = fifo_X_pe_31__dout;
  assign PEG_Xvec_31_fifo_X_in_peek_empty_n = fifo_X_pe_31__empty_n;
  assign PEG_Xvec_31_fifo_X_in_s_dout = fifo_X_pe_31__dout;
  assign PEG_Xvec_31_fifo_X_in_s_empty_n = fifo_X_pe_31__empty_n;
  assign fifo_X_pe_31__read = PEG_Xvec_31_fifo_X_in_s_read;
  assign fifo_X_pe_32__din = PEG_Xvec_31_fifo_X_out_din;
  assign PEG_Xvec_31_fifo_X_out_full_n = fifo_X_pe_32__full_n;
  assign fifo_X_pe_32__write = PEG_Xvec_31_fifo_X_out_write;
  assign fifo_aXvec_31__din = PEG_Xvec_31_fifo_aXvec_din;
  assign PEG_Xvec_31_fifo_aXvec_full_n = fifo_aXvec_31__full_n;
  assign fifo_aXvec_31__write = PEG_Xvec_31_fifo_aXvec_write;
  assign PEG_Xvec_31_fifo_inst_in_peek_dout = PE_inst_31__dout;
  assign PEG_Xvec_31_fifo_inst_in_peek_empty_n = PE_inst_31__empty_n;
  assign PEG_Xvec_31_fifo_inst_in_s_dout = PE_inst_31__dout;
  assign PEG_Xvec_31_fifo_inst_in_s_empty_n = PE_inst_31__empty_n;
  assign PE_inst_31__read = PEG_Xvec_31_fifo_inst_in_s_read;
  assign PE_inst_32__din = PEG_Xvec_31_fifo_inst_out_din;
  assign PEG_Xvec_31_fifo_inst_out_full_n = PE_inst_32__full_n;
  assign Yvec_inst_31__din = PEG_Xvec_31_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_31_fifo_inst_out_to_Yvec_full_n = Yvec_inst_31__full_n;
  assign Yvec_inst_31__write = PEG_Xvec_31_fifo_inst_out_to_Yvec_write;
  assign PE_inst_32__write = PEG_Xvec_31_fifo_inst_out_write;
  assign PEG_Xvec_32_ap_clk = ap_clk;
  assign PEG_Xvec_32__ap_done = PEG_Xvec_32_ap_done;
  assign PEG_Xvec_32__ap_idle = PEG_Xvec_32_ap_idle;
  assign PEG_Xvec_32__ap_ready = PEG_Xvec_32_ap_ready;
  assign PEG_Xvec_32_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_32_ap_start = PEG_Xvec_32__ap_start;
  assign PEG_Xvec_32_fifo_A_peek_dout = fifo_A_32__dout;
  assign PEG_Xvec_32_fifo_A_peek_empty_n = fifo_A_32__empty_n;
  assign PEG_Xvec_32_fifo_A_s_dout = fifo_A_32__dout;
  assign PEG_Xvec_32_fifo_A_s_empty_n = fifo_A_32__empty_n;
  assign fifo_A_32__read = PEG_Xvec_32_fifo_A_s_read;
  assign PEG_Xvec_32_fifo_X_in_peek_dout = fifo_X_pe_32__dout;
  assign PEG_Xvec_32_fifo_X_in_peek_empty_n = fifo_X_pe_32__empty_n;
  assign PEG_Xvec_32_fifo_X_in_s_dout = fifo_X_pe_32__dout;
  assign PEG_Xvec_32_fifo_X_in_s_empty_n = fifo_X_pe_32__empty_n;
  assign fifo_X_pe_32__read = PEG_Xvec_32_fifo_X_in_s_read;
  assign fifo_X_pe_33__din = PEG_Xvec_32_fifo_X_out_din;
  assign PEG_Xvec_32_fifo_X_out_full_n = fifo_X_pe_33__full_n;
  assign fifo_X_pe_33__write = PEG_Xvec_32_fifo_X_out_write;
  assign fifo_aXvec_32__din = PEG_Xvec_32_fifo_aXvec_din;
  assign PEG_Xvec_32_fifo_aXvec_full_n = fifo_aXvec_32__full_n;
  assign fifo_aXvec_32__write = PEG_Xvec_32_fifo_aXvec_write;
  assign PEG_Xvec_32_fifo_inst_in_peek_dout = PE_inst_32__dout;
  assign PEG_Xvec_32_fifo_inst_in_peek_empty_n = PE_inst_32__empty_n;
  assign PEG_Xvec_32_fifo_inst_in_s_dout = PE_inst_32__dout;
  assign PEG_Xvec_32_fifo_inst_in_s_empty_n = PE_inst_32__empty_n;
  assign PE_inst_32__read = PEG_Xvec_32_fifo_inst_in_s_read;
  assign PE_inst_33__din = PEG_Xvec_32_fifo_inst_out_din;
  assign PEG_Xvec_32_fifo_inst_out_full_n = PE_inst_33__full_n;
  assign Yvec_inst_32__din = PEG_Xvec_32_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_32_fifo_inst_out_to_Yvec_full_n = Yvec_inst_32__full_n;
  assign Yvec_inst_32__write = PEG_Xvec_32_fifo_inst_out_to_Yvec_write;
  assign PE_inst_33__write = PEG_Xvec_32_fifo_inst_out_write;
  assign PEG_Xvec_33_ap_clk = ap_clk;
  assign PEG_Xvec_33__ap_done = PEG_Xvec_33_ap_done;
  assign PEG_Xvec_33__ap_idle = PEG_Xvec_33_ap_idle;
  assign PEG_Xvec_33__ap_ready = PEG_Xvec_33_ap_ready;
  assign PEG_Xvec_33_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_33_ap_start = PEG_Xvec_33__ap_start;
  assign PEG_Xvec_33_fifo_A_peek_dout = fifo_A_33__dout;
  assign PEG_Xvec_33_fifo_A_peek_empty_n = fifo_A_33__empty_n;
  assign PEG_Xvec_33_fifo_A_s_dout = fifo_A_33__dout;
  assign PEG_Xvec_33_fifo_A_s_empty_n = fifo_A_33__empty_n;
  assign fifo_A_33__read = PEG_Xvec_33_fifo_A_s_read;
  assign PEG_Xvec_33_fifo_X_in_peek_dout = fifo_X_pe_33__dout;
  assign PEG_Xvec_33_fifo_X_in_peek_empty_n = fifo_X_pe_33__empty_n;
  assign PEG_Xvec_33_fifo_X_in_s_dout = fifo_X_pe_33__dout;
  assign PEG_Xvec_33_fifo_X_in_s_empty_n = fifo_X_pe_33__empty_n;
  assign fifo_X_pe_33__read = PEG_Xvec_33_fifo_X_in_s_read;
  assign fifo_X_pe_34__din = PEG_Xvec_33_fifo_X_out_din;
  assign PEG_Xvec_33_fifo_X_out_full_n = fifo_X_pe_34__full_n;
  assign fifo_X_pe_34__write = PEG_Xvec_33_fifo_X_out_write;
  assign fifo_aXvec_33__din = PEG_Xvec_33_fifo_aXvec_din;
  assign PEG_Xvec_33_fifo_aXvec_full_n = fifo_aXvec_33__full_n;
  assign fifo_aXvec_33__write = PEG_Xvec_33_fifo_aXvec_write;
  assign PEG_Xvec_33_fifo_inst_in_peek_dout = PE_inst_33__dout;
  assign PEG_Xvec_33_fifo_inst_in_peek_empty_n = PE_inst_33__empty_n;
  assign PEG_Xvec_33_fifo_inst_in_s_dout = PE_inst_33__dout;
  assign PEG_Xvec_33_fifo_inst_in_s_empty_n = PE_inst_33__empty_n;
  assign PE_inst_33__read = PEG_Xvec_33_fifo_inst_in_s_read;
  assign PE_inst_34__din = PEG_Xvec_33_fifo_inst_out_din;
  assign PEG_Xvec_33_fifo_inst_out_full_n = PE_inst_34__full_n;
  assign Yvec_inst_33__din = PEG_Xvec_33_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_33_fifo_inst_out_to_Yvec_full_n = Yvec_inst_33__full_n;
  assign Yvec_inst_33__write = PEG_Xvec_33_fifo_inst_out_to_Yvec_write;
  assign PE_inst_34__write = PEG_Xvec_33_fifo_inst_out_write;
  assign PEG_Xvec_34_ap_clk = ap_clk;
  assign PEG_Xvec_34__ap_done = PEG_Xvec_34_ap_done;
  assign PEG_Xvec_34__ap_idle = PEG_Xvec_34_ap_idle;
  assign PEG_Xvec_34__ap_ready = PEG_Xvec_34_ap_ready;
  assign PEG_Xvec_34_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_34_ap_start = PEG_Xvec_34__ap_start;
  assign PEG_Xvec_34_fifo_A_peek_dout = fifo_A_34__dout;
  assign PEG_Xvec_34_fifo_A_peek_empty_n = fifo_A_34__empty_n;
  assign PEG_Xvec_34_fifo_A_s_dout = fifo_A_34__dout;
  assign PEG_Xvec_34_fifo_A_s_empty_n = fifo_A_34__empty_n;
  assign fifo_A_34__read = PEG_Xvec_34_fifo_A_s_read;
  assign PEG_Xvec_34_fifo_X_in_peek_dout = fifo_X_pe_34__dout;
  assign PEG_Xvec_34_fifo_X_in_peek_empty_n = fifo_X_pe_34__empty_n;
  assign PEG_Xvec_34_fifo_X_in_s_dout = fifo_X_pe_34__dout;
  assign PEG_Xvec_34_fifo_X_in_s_empty_n = fifo_X_pe_34__empty_n;
  assign fifo_X_pe_34__read = PEG_Xvec_34_fifo_X_in_s_read;
  assign fifo_X_pe_35__din = PEG_Xvec_34_fifo_X_out_din;
  assign PEG_Xvec_34_fifo_X_out_full_n = fifo_X_pe_35__full_n;
  assign fifo_X_pe_35__write = PEG_Xvec_34_fifo_X_out_write;
  assign fifo_aXvec_34__din = PEG_Xvec_34_fifo_aXvec_din;
  assign PEG_Xvec_34_fifo_aXvec_full_n = fifo_aXvec_34__full_n;
  assign fifo_aXvec_34__write = PEG_Xvec_34_fifo_aXvec_write;
  assign PEG_Xvec_34_fifo_inst_in_peek_dout = PE_inst_34__dout;
  assign PEG_Xvec_34_fifo_inst_in_peek_empty_n = PE_inst_34__empty_n;
  assign PEG_Xvec_34_fifo_inst_in_s_dout = PE_inst_34__dout;
  assign PEG_Xvec_34_fifo_inst_in_s_empty_n = PE_inst_34__empty_n;
  assign PE_inst_34__read = PEG_Xvec_34_fifo_inst_in_s_read;
  assign PE_inst_35__din = PEG_Xvec_34_fifo_inst_out_din;
  assign PEG_Xvec_34_fifo_inst_out_full_n = PE_inst_35__full_n;
  assign Yvec_inst_34__din = PEG_Xvec_34_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_34_fifo_inst_out_to_Yvec_full_n = Yvec_inst_34__full_n;
  assign Yvec_inst_34__write = PEG_Xvec_34_fifo_inst_out_to_Yvec_write;
  assign PE_inst_35__write = PEG_Xvec_34_fifo_inst_out_write;
  assign PEG_Xvec_35_ap_clk = ap_clk;
  assign PEG_Xvec_35__ap_done = PEG_Xvec_35_ap_done;
  assign PEG_Xvec_35__ap_idle = PEG_Xvec_35_ap_idle;
  assign PEG_Xvec_35__ap_ready = PEG_Xvec_35_ap_ready;
  assign PEG_Xvec_35_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_35_ap_start = PEG_Xvec_35__ap_start;
  assign PEG_Xvec_35_fifo_A_peek_dout = fifo_A_35__dout;
  assign PEG_Xvec_35_fifo_A_peek_empty_n = fifo_A_35__empty_n;
  assign PEG_Xvec_35_fifo_A_s_dout = fifo_A_35__dout;
  assign PEG_Xvec_35_fifo_A_s_empty_n = fifo_A_35__empty_n;
  assign fifo_A_35__read = PEG_Xvec_35_fifo_A_s_read;
  assign PEG_Xvec_35_fifo_X_in_peek_dout = fifo_X_pe_35__dout;
  assign PEG_Xvec_35_fifo_X_in_peek_empty_n = fifo_X_pe_35__empty_n;
  assign PEG_Xvec_35_fifo_X_in_s_dout = fifo_X_pe_35__dout;
  assign PEG_Xvec_35_fifo_X_in_s_empty_n = fifo_X_pe_35__empty_n;
  assign fifo_X_pe_35__read = PEG_Xvec_35_fifo_X_in_s_read;
  assign fifo_X_pe_36__din = PEG_Xvec_35_fifo_X_out_din;
  assign PEG_Xvec_35_fifo_X_out_full_n = fifo_X_pe_36__full_n;
  assign fifo_X_pe_36__write = PEG_Xvec_35_fifo_X_out_write;
  assign fifo_aXvec_35__din = PEG_Xvec_35_fifo_aXvec_din;
  assign PEG_Xvec_35_fifo_aXvec_full_n = fifo_aXvec_35__full_n;
  assign fifo_aXvec_35__write = PEG_Xvec_35_fifo_aXvec_write;
  assign PEG_Xvec_35_fifo_inst_in_peek_dout = PE_inst_35__dout;
  assign PEG_Xvec_35_fifo_inst_in_peek_empty_n = PE_inst_35__empty_n;
  assign PEG_Xvec_35_fifo_inst_in_s_dout = PE_inst_35__dout;
  assign PEG_Xvec_35_fifo_inst_in_s_empty_n = PE_inst_35__empty_n;
  assign PE_inst_35__read = PEG_Xvec_35_fifo_inst_in_s_read;
  assign PE_inst_36__din = PEG_Xvec_35_fifo_inst_out_din;
  assign PEG_Xvec_35_fifo_inst_out_full_n = PE_inst_36__full_n;
  assign Yvec_inst_35__din = PEG_Xvec_35_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_35_fifo_inst_out_to_Yvec_full_n = Yvec_inst_35__full_n;
  assign Yvec_inst_35__write = PEG_Xvec_35_fifo_inst_out_to_Yvec_write;
  assign PE_inst_36__write = PEG_Xvec_35_fifo_inst_out_write;
  assign PEG_Xvec_36_ap_clk = ap_clk;
  assign PEG_Xvec_36__ap_done = PEG_Xvec_36_ap_done;
  assign PEG_Xvec_36__ap_idle = PEG_Xvec_36_ap_idle;
  assign PEG_Xvec_36__ap_ready = PEG_Xvec_36_ap_ready;
  assign PEG_Xvec_36_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_36_ap_start = PEG_Xvec_36__ap_start;
  assign PEG_Xvec_36_fifo_A_peek_dout = fifo_A_36__dout;
  assign PEG_Xvec_36_fifo_A_peek_empty_n = fifo_A_36__empty_n;
  assign PEG_Xvec_36_fifo_A_s_dout = fifo_A_36__dout;
  assign PEG_Xvec_36_fifo_A_s_empty_n = fifo_A_36__empty_n;
  assign fifo_A_36__read = PEG_Xvec_36_fifo_A_s_read;
  assign PEG_Xvec_36_fifo_X_in_peek_dout = fifo_X_pe_36__dout;
  assign PEG_Xvec_36_fifo_X_in_peek_empty_n = fifo_X_pe_36__empty_n;
  assign PEG_Xvec_36_fifo_X_in_s_dout = fifo_X_pe_36__dout;
  assign PEG_Xvec_36_fifo_X_in_s_empty_n = fifo_X_pe_36__empty_n;
  assign fifo_X_pe_36__read = PEG_Xvec_36_fifo_X_in_s_read;
  assign fifo_X_pe_37__din = PEG_Xvec_36_fifo_X_out_din;
  assign PEG_Xvec_36_fifo_X_out_full_n = fifo_X_pe_37__full_n;
  assign fifo_X_pe_37__write = PEG_Xvec_36_fifo_X_out_write;
  assign fifo_aXvec_36__din = PEG_Xvec_36_fifo_aXvec_din;
  assign PEG_Xvec_36_fifo_aXvec_full_n = fifo_aXvec_36__full_n;
  assign fifo_aXvec_36__write = PEG_Xvec_36_fifo_aXvec_write;
  assign PEG_Xvec_36_fifo_inst_in_peek_dout = PE_inst_36__dout;
  assign PEG_Xvec_36_fifo_inst_in_peek_empty_n = PE_inst_36__empty_n;
  assign PEG_Xvec_36_fifo_inst_in_s_dout = PE_inst_36__dout;
  assign PEG_Xvec_36_fifo_inst_in_s_empty_n = PE_inst_36__empty_n;
  assign PE_inst_36__read = PEG_Xvec_36_fifo_inst_in_s_read;
  assign PE_inst_37__din = PEG_Xvec_36_fifo_inst_out_din;
  assign PEG_Xvec_36_fifo_inst_out_full_n = PE_inst_37__full_n;
  assign Yvec_inst_36__din = PEG_Xvec_36_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_36_fifo_inst_out_to_Yvec_full_n = Yvec_inst_36__full_n;
  assign Yvec_inst_36__write = PEG_Xvec_36_fifo_inst_out_to_Yvec_write;
  assign PE_inst_37__write = PEG_Xvec_36_fifo_inst_out_write;
  assign PEG_Xvec_37_ap_clk = ap_clk;
  assign PEG_Xvec_37__ap_done = PEG_Xvec_37_ap_done;
  assign PEG_Xvec_37__ap_idle = PEG_Xvec_37_ap_idle;
  assign PEG_Xvec_37__ap_ready = PEG_Xvec_37_ap_ready;
  assign PEG_Xvec_37_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_37_ap_start = PEG_Xvec_37__ap_start;
  assign PEG_Xvec_37_fifo_A_peek_dout = fifo_A_37__dout;
  assign PEG_Xvec_37_fifo_A_peek_empty_n = fifo_A_37__empty_n;
  assign PEG_Xvec_37_fifo_A_s_dout = fifo_A_37__dout;
  assign PEG_Xvec_37_fifo_A_s_empty_n = fifo_A_37__empty_n;
  assign fifo_A_37__read = PEG_Xvec_37_fifo_A_s_read;
  assign PEG_Xvec_37_fifo_X_in_peek_dout = fifo_X_pe_37__dout;
  assign PEG_Xvec_37_fifo_X_in_peek_empty_n = fifo_X_pe_37__empty_n;
  assign PEG_Xvec_37_fifo_X_in_s_dout = fifo_X_pe_37__dout;
  assign PEG_Xvec_37_fifo_X_in_s_empty_n = fifo_X_pe_37__empty_n;
  assign fifo_X_pe_37__read = PEG_Xvec_37_fifo_X_in_s_read;
  assign fifo_X_pe_38__din = PEG_Xvec_37_fifo_X_out_din;
  assign PEG_Xvec_37_fifo_X_out_full_n = fifo_X_pe_38__full_n;
  assign fifo_X_pe_38__write = PEG_Xvec_37_fifo_X_out_write;
  assign fifo_aXvec_37__din = PEG_Xvec_37_fifo_aXvec_din;
  assign PEG_Xvec_37_fifo_aXvec_full_n = fifo_aXvec_37__full_n;
  assign fifo_aXvec_37__write = PEG_Xvec_37_fifo_aXvec_write;
  assign PEG_Xvec_37_fifo_inst_in_peek_dout = PE_inst_37__dout;
  assign PEG_Xvec_37_fifo_inst_in_peek_empty_n = PE_inst_37__empty_n;
  assign PEG_Xvec_37_fifo_inst_in_s_dout = PE_inst_37__dout;
  assign PEG_Xvec_37_fifo_inst_in_s_empty_n = PE_inst_37__empty_n;
  assign PE_inst_37__read = PEG_Xvec_37_fifo_inst_in_s_read;
  assign PE_inst_38__din = PEG_Xvec_37_fifo_inst_out_din;
  assign PEG_Xvec_37_fifo_inst_out_full_n = PE_inst_38__full_n;
  assign Yvec_inst_37__din = PEG_Xvec_37_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_37_fifo_inst_out_to_Yvec_full_n = Yvec_inst_37__full_n;
  assign Yvec_inst_37__write = PEG_Xvec_37_fifo_inst_out_to_Yvec_write;
  assign PE_inst_38__write = PEG_Xvec_37_fifo_inst_out_write;
  assign PEG_Xvec_38_ap_clk = ap_clk;
  assign PEG_Xvec_38__ap_done = PEG_Xvec_38_ap_done;
  assign PEG_Xvec_38__ap_idle = PEG_Xvec_38_ap_idle;
  assign PEG_Xvec_38__ap_ready = PEG_Xvec_38_ap_ready;
  assign PEG_Xvec_38_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_38_ap_start = PEG_Xvec_38__ap_start;
  assign PEG_Xvec_38_fifo_A_peek_dout = fifo_A_38__dout;
  assign PEG_Xvec_38_fifo_A_peek_empty_n = fifo_A_38__empty_n;
  assign PEG_Xvec_38_fifo_A_s_dout = fifo_A_38__dout;
  assign PEG_Xvec_38_fifo_A_s_empty_n = fifo_A_38__empty_n;
  assign fifo_A_38__read = PEG_Xvec_38_fifo_A_s_read;
  assign PEG_Xvec_38_fifo_X_in_peek_dout = fifo_X_pe_38__dout;
  assign PEG_Xvec_38_fifo_X_in_peek_empty_n = fifo_X_pe_38__empty_n;
  assign PEG_Xvec_38_fifo_X_in_s_dout = fifo_X_pe_38__dout;
  assign PEG_Xvec_38_fifo_X_in_s_empty_n = fifo_X_pe_38__empty_n;
  assign fifo_X_pe_38__read = PEG_Xvec_38_fifo_X_in_s_read;
  assign fifo_X_pe_39__din = PEG_Xvec_38_fifo_X_out_din;
  assign PEG_Xvec_38_fifo_X_out_full_n = fifo_X_pe_39__full_n;
  assign fifo_X_pe_39__write = PEG_Xvec_38_fifo_X_out_write;
  assign fifo_aXvec_38__din = PEG_Xvec_38_fifo_aXvec_din;
  assign PEG_Xvec_38_fifo_aXvec_full_n = fifo_aXvec_38__full_n;
  assign fifo_aXvec_38__write = PEG_Xvec_38_fifo_aXvec_write;
  assign PEG_Xvec_38_fifo_inst_in_peek_dout = PE_inst_38__dout;
  assign PEG_Xvec_38_fifo_inst_in_peek_empty_n = PE_inst_38__empty_n;
  assign PEG_Xvec_38_fifo_inst_in_s_dout = PE_inst_38__dout;
  assign PEG_Xvec_38_fifo_inst_in_s_empty_n = PE_inst_38__empty_n;
  assign PE_inst_38__read = PEG_Xvec_38_fifo_inst_in_s_read;
  assign PE_inst_39__din = PEG_Xvec_38_fifo_inst_out_din;
  assign PEG_Xvec_38_fifo_inst_out_full_n = PE_inst_39__full_n;
  assign Yvec_inst_38__din = PEG_Xvec_38_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_38_fifo_inst_out_to_Yvec_full_n = Yvec_inst_38__full_n;
  assign Yvec_inst_38__write = PEG_Xvec_38_fifo_inst_out_to_Yvec_write;
  assign PE_inst_39__write = PEG_Xvec_38_fifo_inst_out_write;
  assign PEG_Xvec_39_ap_clk = ap_clk;
  assign PEG_Xvec_39__ap_done = PEG_Xvec_39_ap_done;
  assign PEG_Xvec_39__ap_idle = PEG_Xvec_39_ap_idle;
  assign PEG_Xvec_39__ap_ready = PEG_Xvec_39_ap_ready;
  assign PEG_Xvec_39_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_39_ap_start = PEG_Xvec_39__ap_start;
  assign PEG_Xvec_39_fifo_A_peek_dout = fifo_A_39__dout;
  assign PEG_Xvec_39_fifo_A_peek_empty_n = fifo_A_39__empty_n;
  assign PEG_Xvec_39_fifo_A_s_dout = fifo_A_39__dout;
  assign PEG_Xvec_39_fifo_A_s_empty_n = fifo_A_39__empty_n;
  assign fifo_A_39__read = PEG_Xvec_39_fifo_A_s_read;
  assign PEG_Xvec_39_fifo_X_in_peek_dout = fifo_X_pe_39__dout;
  assign PEG_Xvec_39_fifo_X_in_peek_empty_n = fifo_X_pe_39__empty_n;
  assign PEG_Xvec_39_fifo_X_in_s_dout = fifo_X_pe_39__dout;
  assign PEG_Xvec_39_fifo_X_in_s_empty_n = fifo_X_pe_39__empty_n;
  assign fifo_X_pe_39__read = PEG_Xvec_39_fifo_X_in_s_read;
  assign fifo_X_pe_40__din = PEG_Xvec_39_fifo_X_out_din;
  assign PEG_Xvec_39_fifo_X_out_full_n = fifo_X_pe_40__full_n;
  assign fifo_X_pe_40__write = PEG_Xvec_39_fifo_X_out_write;
  assign fifo_aXvec_39__din = PEG_Xvec_39_fifo_aXvec_din;
  assign PEG_Xvec_39_fifo_aXvec_full_n = fifo_aXvec_39__full_n;
  assign fifo_aXvec_39__write = PEG_Xvec_39_fifo_aXvec_write;
  assign PEG_Xvec_39_fifo_inst_in_peek_dout = PE_inst_39__dout;
  assign PEG_Xvec_39_fifo_inst_in_peek_empty_n = PE_inst_39__empty_n;
  assign PEG_Xvec_39_fifo_inst_in_s_dout = PE_inst_39__dout;
  assign PEG_Xvec_39_fifo_inst_in_s_empty_n = PE_inst_39__empty_n;
  assign PE_inst_39__read = PEG_Xvec_39_fifo_inst_in_s_read;
  assign PE_inst_40__din = PEG_Xvec_39_fifo_inst_out_din;
  assign PEG_Xvec_39_fifo_inst_out_full_n = PE_inst_40__full_n;
  assign Yvec_inst_39__din = PEG_Xvec_39_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_39_fifo_inst_out_to_Yvec_full_n = Yvec_inst_39__full_n;
  assign Yvec_inst_39__write = PEG_Xvec_39_fifo_inst_out_to_Yvec_write;
  assign PE_inst_40__write = PEG_Xvec_39_fifo_inst_out_write;
  assign PEG_Xvec_40_ap_clk = ap_clk;
  assign PEG_Xvec_40__ap_done = PEG_Xvec_40_ap_done;
  assign PEG_Xvec_40__ap_idle = PEG_Xvec_40_ap_idle;
  assign PEG_Xvec_40__ap_ready = PEG_Xvec_40_ap_ready;
  assign PEG_Xvec_40_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_40_ap_start = PEG_Xvec_40__ap_start;
  assign PEG_Xvec_40_fifo_A_peek_dout = fifo_A_40__dout;
  assign PEG_Xvec_40_fifo_A_peek_empty_n = fifo_A_40__empty_n;
  assign PEG_Xvec_40_fifo_A_s_dout = fifo_A_40__dout;
  assign PEG_Xvec_40_fifo_A_s_empty_n = fifo_A_40__empty_n;
  assign fifo_A_40__read = PEG_Xvec_40_fifo_A_s_read;
  assign PEG_Xvec_40_fifo_X_in_peek_dout = fifo_X_pe_40__dout;
  assign PEG_Xvec_40_fifo_X_in_peek_empty_n = fifo_X_pe_40__empty_n;
  assign PEG_Xvec_40_fifo_X_in_s_dout = fifo_X_pe_40__dout;
  assign PEG_Xvec_40_fifo_X_in_s_empty_n = fifo_X_pe_40__empty_n;
  assign fifo_X_pe_40__read = PEG_Xvec_40_fifo_X_in_s_read;
  assign fifo_X_pe_41__din = PEG_Xvec_40_fifo_X_out_din;
  assign PEG_Xvec_40_fifo_X_out_full_n = fifo_X_pe_41__full_n;
  assign fifo_X_pe_41__write = PEG_Xvec_40_fifo_X_out_write;
  assign fifo_aXvec_40__din = PEG_Xvec_40_fifo_aXvec_din;
  assign PEG_Xvec_40_fifo_aXvec_full_n = fifo_aXvec_40__full_n;
  assign fifo_aXvec_40__write = PEG_Xvec_40_fifo_aXvec_write;
  assign PEG_Xvec_40_fifo_inst_in_peek_dout = PE_inst_40__dout;
  assign PEG_Xvec_40_fifo_inst_in_peek_empty_n = PE_inst_40__empty_n;
  assign PEG_Xvec_40_fifo_inst_in_s_dout = PE_inst_40__dout;
  assign PEG_Xvec_40_fifo_inst_in_s_empty_n = PE_inst_40__empty_n;
  assign PE_inst_40__read = PEG_Xvec_40_fifo_inst_in_s_read;
  assign PE_inst_41__din = PEG_Xvec_40_fifo_inst_out_din;
  assign PEG_Xvec_40_fifo_inst_out_full_n = PE_inst_41__full_n;
  assign Yvec_inst_40__din = PEG_Xvec_40_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_40_fifo_inst_out_to_Yvec_full_n = Yvec_inst_40__full_n;
  assign Yvec_inst_40__write = PEG_Xvec_40_fifo_inst_out_to_Yvec_write;
  assign PE_inst_41__write = PEG_Xvec_40_fifo_inst_out_write;
  assign PEG_Xvec_41_ap_clk = ap_clk;
  assign PEG_Xvec_41__ap_done = PEG_Xvec_41_ap_done;
  assign PEG_Xvec_41__ap_idle = PEG_Xvec_41_ap_idle;
  assign PEG_Xvec_41__ap_ready = PEG_Xvec_41_ap_ready;
  assign PEG_Xvec_41_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_41_ap_start = PEG_Xvec_41__ap_start;
  assign PEG_Xvec_41_fifo_A_peek_dout = fifo_A_41__dout;
  assign PEG_Xvec_41_fifo_A_peek_empty_n = fifo_A_41__empty_n;
  assign PEG_Xvec_41_fifo_A_s_dout = fifo_A_41__dout;
  assign PEG_Xvec_41_fifo_A_s_empty_n = fifo_A_41__empty_n;
  assign fifo_A_41__read = PEG_Xvec_41_fifo_A_s_read;
  assign PEG_Xvec_41_fifo_X_in_peek_dout = fifo_X_pe_41__dout;
  assign PEG_Xvec_41_fifo_X_in_peek_empty_n = fifo_X_pe_41__empty_n;
  assign PEG_Xvec_41_fifo_X_in_s_dout = fifo_X_pe_41__dout;
  assign PEG_Xvec_41_fifo_X_in_s_empty_n = fifo_X_pe_41__empty_n;
  assign fifo_X_pe_41__read = PEG_Xvec_41_fifo_X_in_s_read;
  assign fifo_X_pe_42__din = PEG_Xvec_41_fifo_X_out_din;
  assign PEG_Xvec_41_fifo_X_out_full_n = fifo_X_pe_42__full_n;
  assign fifo_X_pe_42__write = PEG_Xvec_41_fifo_X_out_write;
  assign fifo_aXvec_41__din = PEG_Xvec_41_fifo_aXvec_din;
  assign PEG_Xvec_41_fifo_aXvec_full_n = fifo_aXvec_41__full_n;
  assign fifo_aXvec_41__write = PEG_Xvec_41_fifo_aXvec_write;
  assign PEG_Xvec_41_fifo_inst_in_peek_dout = PE_inst_41__dout;
  assign PEG_Xvec_41_fifo_inst_in_peek_empty_n = PE_inst_41__empty_n;
  assign PEG_Xvec_41_fifo_inst_in_s_dout = PE_inst_41__dout;
  assign PEG_Xvec_41_fifo_inst_in_s_empty_n = PE_inst_41__empty_n;
  assign PE_inst_41__read = PEG_Xvec_41_fifo_inst_in_s_read;
  assign PE_inst_42__din = PEG_Xvec_41_fifo_inst_out_din;
  assign PEG_Xvec_41_fifo_inst_out_full_n = PE_inst_42__full_n;
  assign Yvec_inst_41__din = PEG_Xvec_41_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_41_fifo_inst_out_to_Yvec_full_n = Yvec_inst_41__full_n;
  assign Yvec_inst_41__write = PEG_Xvec_41_fifo_inst_out_to_Yvec_write;
  assign PE_inst_42__write = PEG_Xvec_41_fifo_inst_out_write;
  assign PEG_Xvec_42_ap_clk = ap_clk;
  assign PEG_Xvec_42__ap_done = PEG_Xvec_42_ap_done;
  assign PEG_Xvec_42__ap_idle = PEG_Xvec_42_ap_idle;
  assign PEG_Xvec_42__ap_ready = PEG_Xvec_42_ap_ready;
  assign PEG_Xvec_42_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_42_ap_start = PEG_Xvec_42__ap_start;
  assign PEG_Xvec_42_fifo_A_peek_dout = fifo_A_42__dout;
  assign PEG_Xvec_42_fifo_A_peek_empty_n = fifo_A_42__empty_n;
  assign PEG_Xvec_42_fifo_A_s_dout = fifo_A_42__dout;
  assign PEG_Xvec_42_fifo_A_s_empty_n = fifo_A_42__empty_n;
  assign fifo_A_42__read = PEG_Xvec_42_fifo_A_s_read;
  assign PEG_Xvec_42_fifo_X_in_peek_dout = fifo_X_pe_42__dout;
  assign PEG_Xvec_42_fifo_X_in_peek_empty_n = fifo_X_pe_42__empty_n;
  assign PEG_Xvec_42_fifo_X_in_s_dout = fifo_X_pe_42__dout;
  assign PEG_Xvec_42_fifo_X_in_s_empty_n = fifo_X_pe_42__empty_n;
  assign fifo_X_pe_42__read = PEG_Xvec_42_fifo_X_in_s_read;
  assign fifo_X_pe_43__din = PEG_Xvec_42_fifo_X_out_din;
  assign PEG_Xvec_42_fifo_X_out_full_n = fifo_X_pe_43__full_n;
  assign fifo_X_pe_43__write = PEG_Xvec_42_fifo_X_out_write;
  assign fifo_aXvec_42__din = PEG_Xvec_42_fifo_aXvec_din;
  assign PEG_Xvec_42_fifo_aXvec_full_n = fifo_aXvec_42__full_n;
  assign fifo_aXvec_42__write = PEG_Xvec_42_fifo_aXvec_write;
  assign PEG_Xvec_42_fifo_inst_in_peek_dout = PE_inst_42__dout;
  assign PEG_Xvec_42_fifo_inst_in_peek_empty_n = PE_inst_42__empty_n;
  assign PEG_Xvec_42_fifo_inst_in_s_dout = PE_inst_42__dout;
  assign PEG_Xvec_42_fifo_inst_in_s_empty_n = PE_inst_42__empty_n;
  assign PE_inst_42__read = PEG_Xvec_42_fifo_inst_in_s_read;
  assign PE_inst_43__din = PEG_Xvec_42_fifo_inst_out_din;
  assign PEG_Xvec_42_fifo_inst_out_full_n = PE_inst_43__full_n;
  assign Yvec_inst_42__din = PEG_Xvec_42_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_42_fifo_inst_out_to_Yvec_full_n = Yvec_inst_42__full_n;
  assign Yvec_inst_42__write = PEG_Xvec_42_fifo_inst_out_to_Yvec_write;
  assign PE_inst_43__write = PEG_Xvec_42_fifo_inst_out_write;
  assign PEG_Xvec_43_ap_clk = ap_clk;
  assign PEG_Xvec_43__ap_done = PEG_Xvec_43_ap_done;
  assign PEG_Xvec_43__ap_idle = PEG_Xvec_43_ap_idle;
  assign PEG_Xvec_43__ap_ready = PEG_Xvec_43_ap_ready;
  assign PEG_Xvec_43_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_43_ap_start = PEG_Xvec_43__ap_start;
  assign PEG_Xvec_43_fifo_A_peek_dout = fifo_A_43__dout;
  assign PEG_Xvec_43_fifo_A_peek_empty_n = fifo_A_43__empty_n;
  assign PEG_Xvec_43_fifo_A_s_dout = fifo_A_43__dout;
  assign PEG_Xvec_43_fifo_A_s_empty_n = fifo_A_43__empty_n;
  assign fifo_A_43__read = PEG_Xvec_43_fifo_A_s_read;
  assign PEG_Xvec_43_fifo_X_in_peek_dout = fifo_X_pe_43__dout;
  assign PEG_Xvec_43_fifo_X_in_peek_empty_n = fifo_X_pe_43__empty_n;
  assign PEG_Xvec_43_fifo_X_in_s_dout = fifo_X_pe_43__dout;
  assign PEG_Xvec_43_fifo_X_in_s_empty_n = fifo_X_pe_43__empty_n;
  assign fifo_X_pe_43__read = PEG_Xvec_43_fifo_X_in_s_read;
  assign fifo_X_pe_44__din = PEG_Xvec_43_fifo_X_out_din;
  assign PEG_Xvec_43_fifo_X_out_full_n = fifo_X_pe_44__full_n;
  assign fifo_X_pe_44__write = PEG_Xvec_43_fifo_X_out_write;
  assign fifo_aXvec_43__din = PEG_Xvec_43_fifo_aXvec_din;
  assign PEG_Xvec_43_fifo_aXvec_full_n = fifo_aXvec_43__full_n;
  assign fifo_aXvec_43__write = PEG_Xvec_43_fifo_aXvec_write;
  assign PEG_Xvec_43_fifo_inst_in_peek_dout = PE_inst_43__dout;
  assign PEG_Xvec_43_fifo_inst_in_peek_empty_n = PE_inst_43__empty_n;
  assign PEG_Xvec_43_fifo_inst_in_s_dout = PE_inst_43__dout;
  assign PEG_Xvec_43_fifo_inst_in_s_empty_n = PE_inst_43__empty_n;
  assign PE_inst_43__read = PEG_Xvec_43_fifo_inst_in_s_read;
  assign PE_inst_44__din = PEG_Xvec_43_fifo_inst_out_din;
  assign PEG_Xvec_43_fifo_inst_out_full_n = PE_inst_44__full_n;
  assign Yvec_inst_43__din = PEG_Xvec_43_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_43_fifo_inst_out_to_Yvec_full_n = Yvec_inst_43__full_n;
  assign Yvec_inst_43__write = PEG_Xvec_43_fifo_inst_out_to_Yvec_write;
  assign PE_inst_44__write = PEG_Xvec_43_fifo_inst_out_write;
  assign PEG_Xvec_44_ap_clk = ap_clk;
  assign PEG_Xvec_44__ap_done = PEG_Xvec_44_ap_done;
  assign PEG_Xvec_44__ap_idle = PEG_Xvec_44_ap_idle;
  assign PEG_Xvec_44__ap_ready = PEG_Xvec_44_ap_ready;
  assign PEG_Xvec_44_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_44_ap_start = PEG_Xvec_44__ap_start;
  assign PEG_Xvec_44_fifo_A_peek_dout = fifo_A_44__dout;
  assign PEG_Xvec_44_fifo_A_peek_empty_n = fifo_A_44__empty_n;
  assign PEG_Xvec_44_fifo_A_s_dout = fifo_A_44__dout;
  assign PEG_Xvec_44_fifo_A_s_empty_n = fifo_A_44__empty_n;
  assign fifo_A_44__read = PEG_Xvec_44_fifo_A_s_read;
  assign PEG_Xvec_44_fifo_X_in_peek_dout = fifo_X_pe_44__dout;
  assign PEG_Xvec_44_fifo_X_in_peek_empty_n = fifo_X_pe_44__empty_n;
  assign PEG_Xvec_44_fifo_X_in_s_dout = fifo_X_pe_44__dout;
  assign PEG_Xvec_44_fifo_X_in_s_empty_n = fifo_X_pe_44__empty_n;
  assign fifo_X_pe_44__read = PEG_Xvec_44_fifo_X_in_s_read;
  assign fifo_X_pe_45__din = PEG_Xvec_44_fifo_X_out_din;
  assign PEG_Xvec_44_fifo_X_out_full_n = fifo_X_pe_45__full_n;
  assign fifo_X_pe_45__write = PEG_Xvec_44_fifo_X_out_write;
  assign fifo_aXvec_44__din = PEG_Xvec_44_fifo_aXvec_din;
  assign PEG_Xvec_44_fifo_aXvec_full_n = fifo_aXvec_44__full_n;
  assign fifo_aXvec_44__write = PEG_Xvec_44_fifo_aXvec_write;
  assign PEG_Xvec_44_fifo_inst_in_peek_dout = PE_inst_44__dout;
  assign PEG_Xvec_44_fifo_inst_in_peek_empty_n = PE_inst_44__empty_n;
  assign PEG_Xvec_44_fifo_inst_in_s_dout = PE_inst_44__dout;
  assign PEG_Xvec_44_fifo_inst_in_s_empty_n = PE_inst_44__empty_n;
  assign PE_inst_44__read = PEG_Xvec_44_fifo_inst_in_s_read;
  assign PE_inst_45__din = PEG_Xvec_44_fifo_inst_out_din;
  assign PEG_Xvec_44_fifo_inst_out_full_n = PE_inst_45__full_n;
  assign Yvec_inst_44__din = PEG_Xvec_44_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_44_fifo_inst_out_to_Yvec_full_n = Yvec_inst_44__full_n;
  assign Yvec_inst_44__write = PEG_Xvec_44_fifo_inst_out_to_Yvec_write;
  assign PE_inst_45__write = PEG_Xvec_44_fifo_inst_out_write;
  assign PEG_Xvec_45_ap_clk = ap_clk;
  assign PEG_Xvec_45__ap_done = PEG_Xvec_45_ap_done;
  assign PEG_Xvec_45__ap_idle = PEG_Xvec_45_ap_idle;
  assign PEG_Xvec_45__ap_ready = PEG_Xvec_45_ap_ready;
  assign PEG_Xvec_45_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_45_ap_start = PEG_Xvec_45__ap_start;
  assign PEG_Xvec_45_fifo_A_peek_dout = fifo_A_45__dout;
  assign PEG_Xvec_45_fifo_A_peek_empty_n = fifo_A_45__empty_n;
  assign PEG_Xvec_45_fifo_A_s_dout = fifo_A_45__dout;
  assign PEG_Xvec_45_fifo_A_s_empty_n = fifo_A_45__empty_n;
  assign fifo_A_45__read = PEG_Xvec_45_fifo_A_s_read;
  assign PEG_Xvec_45_fifo_X_in_peek_dout = fifo_X_pe_45__dout;
  assign PEG_Xvec_45_fifo_X_in_peek_empty_n = fifo_X_pe_45__empty_n;
  assign PEG_Xvec_45_fifo_X_in_s_dout = fifo_X_pe_45__dout;
  assign PEG_Xvec_45_fifo_X_in_s_empty_n = fifo_X_pe_45__empty_n;
  assign fifo_X_pe_45__read = PEG_Xvec_45_fifo_X_in_s_read;
  assign fifo_X_pe_46__din = PEG_Xvec_45_fifo_X_out_din;
  assign PEG_Xvec_45_fifo_X_out_full_n = fifo_X_pe_46__full_n;
  assign fifo_X_pe_46__write = PEG_Xvec_45_fifo_X_out_write;
  assign fifo_aXvec_45__din = PEG_Xvec_45_fifo_aXvec_din;
  assign PEG_Xvec_45_fifo_aXvec_full_n = fifo_aXvec_45__full_n;
  assign fifo_aXvec_45__write = PEG_Xvec_45_fifo_aXvec_write;
  assign PEG_Xvec_45_fifo_inst_in_peek_dout = PE_inst_45__dout;
  assign PEG_Xvec_45_fifo_inst_in_peek_empty_n = PE_inst_45__empty_n;
  assign PEG_Xvec_45_fifo_inst_in_s_dout = PE_inst_45__dout;
  assign PEG_Xvec_45_fifo_inst_in_s_empty_n = PE_inst_45__empty_n;
  assign PE_inst_45__read = PEG_Xvec_45_fifo_inst_in_s_read;
  assign PE_inst_46__din = PEG_Xvec_45_fifo_inst_out_din;
  assign PEG_Xvec_45_fifo_inst_out_full_n = PE_inst_46__full_n;
  assign Yvec_inst_45__din = PEG_Xvec_45_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_45_fifo_inst_out_to_Yvec_full_n = Yvec_inst_45__full_n;
  assign Yvec_inst_45__write = PEG_Xvec_45_fifo_inst_out_to_Yvec_write;
  assign PE_inst_46__write = PEG_Xvec_45_fifo_inst_out_write;
  assign PEG_Xvec_46_ap_clk = ap_clk;
  assign PEG_Xvec_46__ap_done = PEG_Xvec_46_ap_done;
  assign PEG_Xvec_46__ap_idle = PEG_Xvec_46_ap_idle;
  assign PEG_Xvec_46__ap_ready = PEG_Xvec_46_ap_ready;
  assign PEG_Xvec_46_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_46_ap_start = PEG_Xvec_46__ap_start;
  assign PEG_Xvec_46_fifo_A_peek_dout = fifo_A_46__dout;
  assign PEG_Xvec_46_fifo_A_peek_empty_n = fifo_A_46__empty_n;
  assign PEG_Xvec_46_fifo_A_s_dout = fifo_A_46__dout;
  assign PEG_Xvec_46_fifo_A_s_empty_n = fifo_A_46__empty_n;
  assign fifo_A_46__read = PEG_Xvec_46_fifo_A_s_read;
  assign PEG_Xvec_46_fifo_X_in_peek_dout = fifo_X_pe_46__dout;
  assign PEG_Xvec_46_fifo_X_in_peek_empty_n = fifo_X_pe_46__empty_n;
  assign PEG_Xvec_46_fifo_X_in_s_dout = fifo_X_pe_46__dout;
  assign PEG_Xvec_46_fifo_X_in_s_empty_n = fifo_X_pe_46__empty_n;
  assign fifo_X_pe_46__read = PEG_Xvec_46_fifo_X_in_s_read;
  assign fifo_X_pe_47__din = PEG_Xvec_46_fifo_X_out_din;
  assign PEG_Xvec_46_fifo_X_out_full_n = fifo_X_pe_47__full_n;
  assign fifo_X_pe_47__write = PEG_Xvec_46_fifo_X_out_write;
  assign fifo_aXvec_46__din = PEG_Xvec_46_fifo_aXvec_din;
  assign PEG_Xvec_46_fifo_aXvec_full_n = fifo_aXvec_46__full_n;
  assign fifo_aXvec_46__write = PEG_Xvec_46_fifo_aXvec_write;
  assign PEG_Xvec_46_fifo_inst_in_peek_dout = PE_inst_46__dout;
  assign PEG_Xvec_46_fifo_inst_in_peek_empty_n = PE_inst_46__empty_n;
  assign PEG_Xvec_46_fifo_inst_in_s_dout = PE_inst_46__dout;
  assign PEG_Xvec_46_fifo_inst_in_s_empty_n = PE_inst_46__empty_n;
  assign PE_inst_46__read = PEG_Xvec_46_fifo_inst_in_s_read;
  assign PE_inst_47__din = PEG_Xvec_46_fifo_inst_out_din;
  assign PEG_Xvec_46_fifo_inst_out_full_n = PE_inst_47__full_n;
  assign Yvec_inst_46__din = PEG_Xvec_46_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_46_fifo_inst_out_to_Yvec_full_n = Yvec_inst_46__full_n;
  assign Yvec_inst_46__write = PEG_Xvec_46_fifo_inst_out_to_Yvec_write;
  assign PE_inst_47__write = PEG_Xvec_46_fifo_inst_out_write;
  assign PEG_Xvec_47_ap_clk = ap_clk;
  assign PEG_Xvec_47__ap_done = PEG_Xvec_47_ap_done;
  assign PEG_Xvec_47__ap_idle = PEG_Xvec_47_ap_idle;
  assign PEG_Xvec_47__ap_ready = PEG_Xvec_47_ap_ready;
  assign PEG_Xvec_47_ap_rst_n = ap_rst_n;
  assign PEG_Xvec_47_ap_start = PEG_Xvec_47__ap_start;
  assign PEG_Xvec_47_fifo_A_peek_dout = fifo_A_47__dout;
  assign PEG_Xvec_47_fifo_A_peek_empty_n = fifo_A_47__empty_n;
  assign PEG_Xvec_47_fifo_A_s_dout = fifo_A_47__dout;
  assign PEG_Xvec_47_fifo_A_s_empty_n = fifo_A_47__empty_n;
  assign fifo_A_47__read = PEG_Xvec_47_fifo_A_s_read;
  assign PEG_Xvec_47_fifo_X_in_peek_dout = fifo_X_pe_47__dout;
  assign PEG_Xvec_47_fifo_X_in_peek_empty_n = fifo_X_pe_47__empty_n;
  assign PEG_Xvec_47_fifo_X_in_s_dout = fifo_X_pe_47__dout;
  assign PEG_Xvec_47_fifo_X_in_s_empty_n = fifo_X_pe_47__empty_n;
  assign fifo_X_pe_47__read = PEG_Xvec_47_fifo_X_in_s_read;
  assign fifo_X_pe_48__din = PEG_Xvec_47_fifo_X_out_din;
  assign PEG_Xvec_47_fifo_X_out_full_n = fifo_X_pe_48__full_n;
  assign fifo_X_pe_48__write = PEG_Xvec_47_fifo_X_out_write;
  assign fifo_aXvec_47__din = PEG_Xvec_47_fifo_aXvec_din;
  assign PEG_Xvec_47_fifo_aXvec_full_n = fifo_aXvec_47__full_n;
  assign fifo_aXvec_47__write = PEG_Xvec_47_fifo_aXvec_write;
  assign PEG_Xvec_47_fifo_inst_in_peek_dout = PE_inst_47__dout;
  assign PEG_Xvec_47_fifo_inst_in_peek_empty_n = PE_inst_47__empty_n;
  assign PEG_Xvec_47_fifo_inst_in_s_dout = PE_inst_47__dout;
  assign PEG_Xvec_47_fifo_inst_in_s_empty_n = PE_inst_47__empty_n;
  assign PE_inst_47__read = PEG_Xvec_47_fifo_inst_in_s_read;
  assign PE_inst_48__din = PEG_Xvec_47_fifo_inst_out_din;
  assign PEG_Xvec_47_fifo_inst_out_full_n = PE_inst_48__full_n;
  assign Yvec_inst_47__din = PEG_Xvec_47_fifo_inst_out_to_Yvec_din;
  assign PEG_Xvec_47_fifo_inst_out_to_Yvec_full_n = Yvec_inst_47__full_n;
  assign Yvec_inst_47__write = PEG_Xvec_47_fifo_inst_out_to_Yvec_write;
  assign PE_inst_48__write = PEG_Xvec_47_fifo_inst_out_write;
  assign PEG_Yvec_0_ap_clk = ap_clk;
  assign PEG_Yvec_0__ap_done = PEG_Yvec_0_ap_done;
  assign PEG_Yvec_0__ap_idle = PEG_Yvec_0_ap_idle;
  assign PEG_Yvec_0__ap_ready = PEG_Yvec_0_ap_ready;
  assign PEG_Yvec_0_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_0_ap_start = PEG_Yvec_0__ap_start;
  assign fifo_Y_pe_0__din = PEG_Yvec_0_fifo_Y_out_din;
  assign PEG_Yvec_0_fifo_Y_out_full_n = fifo_Y_pe_0__full_n;
  assign fifo_Y_pe_0__write = PEG_Yvec_0_fifo_Y_out_write;
  assign PEG_Yvec_0_fifo_aXvec_peek_dout = fifo_aXvec_0__dout;
  assign PEG_Yvec_0_fifo_aXvec_peek_empty_n = fifo_aXvec_0__empty_n;
  assign PEG_Yvec_0_fifo_aXvec_s_dout = fifo_aXvec_0__dout;
  assign PEG_Yvec_0_fifo_aXvec_s_empty_n = fifo_aXvec_0__empty_n;
  assign fifo_aXvec_0__read = PEG_Yvec_0_fifo_aXvec_s_read;
  assign PEG_Yvec_0_fifo_inst_in_peek_dout = Yvec_inst_0__dout;
  assign PEG_Yvec_0_fifo_inst_in_peek_empty_n = Yvec_inst_0__empty_n;
  assign PEG_Yvec_0_fifo_inst_in_s_dout = Yvec_inst_0__dout;
  assign PEG_Yvec_0_fifo_inst_in_s_empty_n = Yvec_inst_0__empty_n;
  assign Yvec_inst_0__read = PEG_Yvec_0_fifo_inst_in_s_read;
  assign PEG_Yvec_1_ap_clk = ap_clk;
  assign PEG_Yvec_1__ap_done = PEG_Yvec_1_ap_done;
  assign PEG_Yvec_1__ap_idle = PEG_Yvec_1_ap_idle;
  assign PEG_Yvec_1__ap_ready = PEG_Yvec_1_ap_ready;
  assign PEG_Yvec_1_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_1_ap_start = PEG_Yvec_1__ap_start;
  assign fifo_Y_pe_1__din = PEG_Yvec_1_fifo_Y_out_din;
  assign PEG_Yvec_1_fifo_Y_out_full_n = fifo_Y_pe_1__full_n;
  assign fifo_Y_pe_1__write = PEG_Yvec_1_fifo_Y_out_write;
  assign PEG_Yvec_1_fifo_aXvec_peek_dout = fifo_aXvec_1__dout;
  assign PEG_Yvec_1_fifo_aXvec_peek_empty_n = fifo_aXvec_1__empty_n;
  assign PEG_Yvec_1_fifo_aXvec_s_dout = fifo_aXvec_1__dout;
  assign PEG_Yvec_1_fifo_aXvec_s_empty_n = fifo_aXvec_1__empty_n;
  assign fifo_aXvec_1__read = PEG_Yvec_1_fifo_aXvec_s_read;
  assign PEG_Yvec_1_fifo_inst_in_peek_dout = Yvec_inst_1__dout;
  assign PEG_Yvec_1_fifo_inst_in_peek_empty_n = Yvec_inst_1__empty_n;
  assign PEG_Yvec_1_fifo_inst_in_s_dout = Yvec_inst_1__dout;
  assign PEG_Yvec_1_fifo_inst_in_s_empty_n = Yvec_inst_1__empty_n;
  assign Yvec_inst_1__read = PEG_Yvec_1_fifo_inst_in_s_read;
  assign PEG_Yvec_2_ap_clk = ap_clk;
  assign PEG_Yvec_2__ap_done = PEG_Yvec_2_ap_done;
  assign PEG_Yvec_2__ap_idle = PEG_Yvec_2_ap_idle;
  assign PEG_Yvec_2__ap_ready = PEG_Yvec_2_ap_ready;
  assign PEG_Yvec_2_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_2_ap_start = PEG_Yvec_2__ap_start;
  assign fifo_Y_pe_2__din = PEG_Yvec_2_fifo_Y_out_din;
  assign PEG_Yvec_2_fifo_Y_out_full_n = fifo_Y_pe_2__full_n;
  assign fifo_Y_pe_2__write = PEG_Yvec_2_fifo_Y_out_write;
  assign PEG_Yvec_2_fifo_aXvec_peek_dout = fifo_aXvec_2__dout;
  assign PEG_Yvec_2_fifo_aXvec_peek_empty_n = fifo_aXvec_2__empty_n;
  assign PEG_Yvec_2_fifo_aXvec_s_dout = fifo_aXvec_2__dout;
  assign PEG_Yvec_2_fifo_aXvec_s_empty_n = fifo_aXvec_2__empty_n;
  assign fifo_aXvec_2__read = PEG_Yvec_2_fifo_aXvec_s_read;
  assign PEG_Yvec_2_fifo_inst_in_peek_dout = Yvec_inst_2__dout;
  assign PEG_Yvec_2_fifo_inst_in_peek_empty_n = Yvec_inst_2__empty_n;
  assign PEG_Yvec_2_fifo_inst_in_s_dout = Yvec_inst_2__dout;
  assign PEG_Yvec_2_fifo_inst_in_s_empty_n = Yvec_inst_2__empty_n;
  assign Yvec_inst_2__read = PEG_Yvec_2_fifo_inst_in_s_read;
  assign PEG_Yvec_3_ap_clk = ap_clk;
  assign PEG_Yvec_3__ap_done = PEG_Yvec_3_ap_done;
  assign PEG_Yvec_3__ap_idle = PEG_Yvec_3_ap_idle;
  assign PEG_Yvec_3__ap_ready = PEG_Yvec_3_ap_ready;
  assign PEG_Yvec_3_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_3_ap_start = PEG_Yvec_3__ap_start;
  assign fifo_Y_pe_3__din = PEG_Yvec_3_fifo_Y_out_din;
  assign PEG_Yvec_3_fifo_Y_out_full_n = fifo_Y_pe_3__full_n;
  assign fifo_Y_pe_3__write = PEG_Yvec_3_fifo_Y_out_write;
  assign PEG_Yvec_3_fifo_aXvec_peek_dout = fifo_aXvec_3__dout;
  assign PEG_Yvec_3_fifo_aXvec_peek_empty_n = fifo_aXvec_3__empty_n;
  assign PEG_Yvec_3_fifo_aXvec_s_dout = fifo_aXvec_3__dout;
  assign PEG_Yvec_3_fifo_aXvec_s_empty_n = fifo_aXvec_3__empty_n;
  assign fifo_aXvec_3__read = PEG_Yvec_3_fifo_aXvec_s_read;
  assign PEG_Yvec_3_fifo_inst_in_peek_dout = Yvec_inst_3__dout;
  assign PEG_Yvec_3_fifo_inst_in_peek_empty_n = Yvec_inst_3__empty_n;
  assign PEG_Yvec_3_fifo_inst_in_s_dout = Yvec_inst_3__dout;
  assign PEG_Yvec_3_fifo_inst_in_s_empty_n = Yvec_inst_3__empty_n;
  assign Yvec_inst_3__read = PEG_Yvec_3_fifo_inst_in_s_read;
  assign PEG_Yvec_4_ap_clk = ap_clk;
  assign PEG_Yvec_4__ap_done = PEG_Yvec_4_ap_done;
  assign PEG_Yvec_4__ap_idle = PEG_Yvec_4_ap_idle;
  assign PEG_Yvec_4__ap_ready = PEG_Yvec_4_ap_ready;
  assign PEG_Yvec_4_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_4_ap_start = PEG_Yvec_4__ap_start;
  assign fifo_Y_pe_4__din = PEG_Yvec_4_fifo_Y_out_din;
  assign PEG_Yvec_4_fifo_Y_out_full_n = fifo_Y_pe_4__full_n;
  assign fifo_Y_pe_4__write = PEG_Yvec_4_fifo_Y_out_write;
  assign PEG_Yvec_4_fifo_aXvec_peek_dout = fifo_aXvec_4__dout;
  assign PEG_Yvec_4_fifo_aXvec_peek_empty_n = fifo_aXvec_4__empty_n;
  assign PEG_Yvec_4_fifo_aXvec_s_dout = fifo_aXvec_4__dout;
  assign PEG_Yvec_4_fifo_aXvec_s_empty_n = fifo_aXvec_4__empty_n;
  assign fifo_aXvec_4__read = PEG_Yvec_4_fifo_aXvec_s_read;
  assign PEG_Yvec_4_fifo_inst_in_peek_dout = Yvec_inst_4__dout;
  assign PEG_Yvec_4_fifo_inst_in_peek_empty_n = Yvec_inst_4__empty_n;
  assign PEG_Yvec_4_fifo_inst_in_s_dout = Yvec_inst_4__dout;
  assign PEG_Yvec_4_fifo_inst_in_s_empty_n = Yvec_inst_4__empty_n;
  assign Yvec_inst_4__read = PEG_Yvec_4_fifo_inst_in_s_read;
  assign PEG_Yvec_5_ap_clk = ap_clk;
  assign PEG_Yvec_5__ap_done = PEG_Yvec_5_ap_done;
  assign PEG_Yvec_5__ap_idle = PEG_Yvec_5_ap_idle;
  assign PEG_Yvec_5__ap_ready = PEG_Yvec_5_ap_ready;
  assign PEG_Yvec_5_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_5_ap_start = PEG_Yvec_5__ap_start;
  assign fifo_Y_pe_5__din = PEG_Yvec_5_fifo_Y_out_din;
  assign PEG_Yvec_5_fifo_Y_out_full_n = fifo_Y_pe_5__full_n;
  assign fifo_Y_pe_5__write = PEG_Yvec_5_fifo_Y_out_write;
  assign PEG_Yvec_5_fifo_aXvec_peek_dout = fifo_aXvec_5__dout;
  assign PEG_Yvec_5_fifo_aXvec_peek_empty_n = fifo_aXvec_5__empty_n;
  assign PEG_Yvec_5_fifo_aXvec_s_dout = fifo_aXvec_5__dout;
  assign PEG_Yvec_5_fifo_aXvec_s_empty_n = fifo_aXvec_5__empty_n;
  assign fifo_aXvec_5__read = PEG_Yvec_5_fifo_aXvec_s_read;
  assign PEG_Yvec_5_fifo_inst_in_peek_dout = Yvec_inst_5__dout;
  assign PEG_Yvec_5_fifo_inst_in_peek_empty_n = Yvec_inst_5__empty_n;
  assign PEG_Yvec_5_fifo_inst_in_s_dout = Yvec_inst_5__dout;
  assign PEG_Yvec_5_fifo_inst_in_s_empty_n = Yvec_inst_5__empty_n;
  assign Yvec_inst_5__read = PEG_Yvec_5_fifo_inst_in_s_read;
  assign PEG_Yvec_6_ap_clk = ap_clk;
  assign PEG_Yvec_6__ap_done = PEG_Yvec_6_ap_done;
  assign PEG_Yvec_6__ap_idle = PEG_Yvec_6_ap_idle;
  assign PEG_Yvec_6__ap_ready = PEG_Yvec_6_ap_ready;
  assign PEG_Yvec_6_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_6_ap_start = PEG_Yvec_6__ap_start;
  assign fifo_Y_pe_6__din = PEG_Yvec_6_fifo_Y_out_din;
  assign PEG_Yvec_6_fifo_Y_out_full_n = fifo_Y_pe_6__full_n;
  assign fifo_Y_pe_6__write = PEG_Yvec_6_fifo_Y_out_write;
  assign PEG_Yvec_6_fifo_aXvec_peek_dout = fifo_aXvec_6__dout;
  assign PEG_Yvec_6_fifo_aXvec_peek_empty_n = fifo_aXvec_6__empty_n;
  assign PEG_Yvec_6_fifo_aXvec_s_dout = fifo_aXvec_6__dout;
  assign PEG_Yvec_6_fifo_aXvec_s_empty_n = fifo_aXvec_6__empty_n;
  assign fifo_aXvec_6__read = PEG_Yvec_6_fifo_aXvec_s_read;
  assign PEG_Yvec_6_fifo_inst_in_peek_dout = Yvec_inst_6__dout;
  assign PEG_Yvec_6_fifo_inst_in_peek_empty_n = Yvec_inst_6__empty_n;
  assign PEG_Yvec_6_fifo_inst_in_s_dout = Yvec_inst_6__dout;
  assign PEG_Yvec_6_fifo_inst_in_s_empty_n = Yvec_inst_6__empty_n;
  assign Yvec_inst_6__read = PEG_Yvec_6_fifo_inst_in_s_read;
  assign PEG_Yvec_7_ap_clk = ap_clk;
  assign PEG_Yvec_7__ap_done = PEG_Yvec_7_ap_done;
  assign PEG_Yvec_7__ap_idle = PEG_Yvec_7_ap_idle;
  assign PEG_Yvec_7__ap_ready = PEG_Yvec_7_ap_ready;
  assign PEG_Yvec_7_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_7_ap_start = PEG_Yvec_7__ap_start;
  assign fifo_Y_pe_7__din = PEG_Yvec_7_fifo_Y_out_din;
  assign PEG_Yvec_7_fifo_Y_out_full_n = fifo_Y_pe_7__full_n;
  assign fifo_Y_pe_7__write = PEG_Yvec_7_fifo_Y_out_write;
  assign PEG_Yvec_7_fifo_aXvec_peek_dout = fifo_aXvec_7__dout;
  assign PEG_Yvec_7_fifo_aXvec_peek_empty_n = fifo_aXvec_7__empty_n;
  assign PEG_Yvec_7_fifo_aXvec_s_dout = fifo_aXvec_7__dout;
  assign PEG_Yvec_7_fifo_aXvec_s_empty_n = fifo_aXvec_7__empty_n;
  assign fifo_aXvec_7__read = PEG_Yvec_7_fifo_aXvec_s_read;
  assign PEG_Yvec_7_fifo_inst_in_peek_dout = Yvec_inst_7__dout;
  assign PEG_Yvec_7_fifo_inst_in_peek_empty_n = Yvec_inst_7__empty_n;
  assign PEG_Yvec_7_fifo_inst_in_s_dout = Yvec_inst_7__dout;
  assign PEG_Yvec_7_fifo_inst_in_s_empty_n = Yvec_inst_7__empty_n;
  assign Yvec_inst_7__read = PEG_Yvec_7_fifo_inst_in_s_read;
  assign PEG_Yvec_8_ap_clk = ap_clk;
  assign PEG_Yvec_8__ap_done = PEG_Yvec_8_ap_done;
  assign PEG_Yvec_8__ap_idle = PEG_Yvec_8_ap_idle;
  assign PEG_Yvec_8__ap_ready = PEG_Yvec_8_ap_ready;
  assign PEG_Yvec_8_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_8_ap_start = PEG_Yvec_8__ap_start;
  assign fifo_Y_pe_8__din = PEG_Yvec_8_fifo_Y_out_din;
  assign PEG_Yvec_8_fifo_Y_out_full_n = fifo_Y_pe_8__full_n;
  assign fifo_Y_pe_8__write = PEG_Yvec_8_fifo_Y_out_write;
  assign PEG_Yvec_8_fifo_aXvec_peek_dout = fifo_aXvec_8__dout;
  assign PEG_Yvec_8_fifo_aXvec_peek_empty_n = fifo_aXvec_8__empty_n;
  assign PEG_Yvec_8_fifo_aXvec_s_dout = fifo_aXvec_8__dout;
  assign PEG_Yvec_8_fifo_aXvec_s_empty_n = fifo_aXvec_8__empty_n;
  assign fifo_aXvec_8__read = PEG_Yvec_8_fifo_aXvec_s_read;
  assign PEG_Yvec_8_fifo_inst_in_peek_dout = Yvec_inst_8__dout;
  assign PEG_Yvec_8_fifo_inst_in_peek_empty_n = Yvec_inst_8__empty_n;
  assign PEG_Yvec_8_fifo_inst_in_s_dout = Yvec_inst_8__dout;
  assign PEG_Yvec_8_fifo_inst_in_s_empty_n = Yvec_inst_8__empty_n;
  assign Yvec_inst_8__read = PEG_Yvec_8_fifo_inst_in_s_read;
  assign PEG_Yvec_9_ap_clk = ap_clk;
  assign PEG_Yvec_9__ap_done = PEG_Yvec_9_ap_done;
  assign PEG_Yvec_9__ap_idle = PEG_Yvec_9_ap_idle;
  assign PEG_Yvec_9__ap_ready = PEG_Yvec_9_ap_ready;
  assign PEG_Yvec_9_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_9_ap_start = PEG_Yvec_9__ap_start;
  assign fifo_Y_pe_9__din = PEG_Yvec_9_fifo_Y_out_din;
  assign PEG_Yvec_9_fifo_Y_out_full_n = fifo_Y_pe_9__full_n;
  assign fifo_Y_pe_9__write = PEG_Yvec_9_fifo_Y_out_write;
  assign PEG_Yvec_9_fifo_aXvec_peek_dout = fifo_aXvec_9__dout;
  assign PEG_Yvec_9_fifo_aXvec_peek_empty_n = fifo_aXvec_9__empty_n;
  assign PEG_Yvec_9_fifo_aXvec_s_dout = fifo_aXvec_9__dout;
  assign PEG_Yvec_9_fifo_aXvec_s_empty_n = fifo_aXvec_9__empty_n;
  assign fifo_aXvec_9__read = PEG_Yvec_9_fifo_aXvec_s_read;
  assign PEG_Yvec_9_fifo_inst_in_peek_dout = Yvec_inst_9__dout;
  assign PEG_Yvec_9_fifo_inst_in_peek_empty_n = Yvec_inst_9__empty_n;
  assign PEG_Yvec_9_fifo_inst_in_s_dout = Yvec_inst_9__dout;
  assign PEG_Yvec_9_fifo_inst_in_s_empty_n = Yvec_inst_9__empty_n;
  assign Yvec_inst_9__read = PEG_Yvec_9_fifo_inst_in_s_read;
  assign PEG_Yvec_10_ap_clk = ap_clk;
  assign PEG_Yvec_10__ap_done = PEG_Yvec_10_ap_done;
  assign PEG_Yvec_10__ap_idle = PEG_Yvec_10_ap_idle;
  assign PEG_Yvec_10__ap_ready = PEG_Yvec_10_ap_ready;
  assign PEG_Yvec_10_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_10_ap_start = PEG_Yvec_10__ap_start;
  assign fifo_Y_pe_10__din = PEG_Yvec_10_fifo_Y_out_din;
  assign PEG_Yvec_10_fifo_Y_out_full_n = fifo_Y_pe_10__full_n;
  assign fifo_Y_pe_10__write = PEG_Yvec_10_fifo_Y_out_write;
  assign PEG_Yvec_10_fifo_aXvec_peek_dout = fifo_aXvec_10__dout;
  assign PEG_Yvec_10_fifo_aXvec_peek_empty_n = fifo_aXvec_10__empty_n;
  assign PEG_Yvec_10_fifo_aXvec_s_dout = fifo_aXvec_10__dout;
  assign PEG_Yvec_10_fifo_aXvec_s_empty_n = fifo_aXvec_10__empty_n;
  assign fifo_aXvec_10__read = PEG_Yvec_10_fifo_aXvec_s_read;
  assign PEG_Yvec_10_fifo_inst_in_peek_dout = Yvec_inst_10__dout;
  assign PEG_Yvec_10_fifo_inst_in_peek_empty_n = Yvec_inst_10__empty_n;
  assign PEG_Yvec_10_fifo_inst_in_s_dout = Yvec_inst_10__dout;
  assign PEG_Yvec_10_fifo_inst_in_s_empty_n = Yvec_inst_10__empty_n;
  assign Yvec_inst_10__read = PEG_Yvec_10_fifo_inst_in_s_read;
  assign PEG_Yvec_11_ap_clk = ap_clk;
  assign PEG_Yvec_11__ap_done = PEG_Yvec_11_ap_done;
  assign PEG_Yvec_11__ap_idle = PEG_Yvec_11_ap_idle;
  assign PEG_Yvec_11__ap_ready = PEG_Yvec_11_ap_ready;
  assign PEG_Yvec_11_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_11_ap_start = PEG_Yvec_11__ap_start;
  assign fifo_Y_pe_11__din = PEG_Yvec_11_fifo_Y_out_din;
  assign PEG_Yvec_11_fifo_Y_out_full_n = fifo_Y_pe_11__full_n;
  assign fifo_Y_pe_11__write = PEG_Yvec_11_fifo_Y_out_write;
  assign PEG_Yvec_11_fifo_aXvec_peek_dout = fifo_aXvec_11__dout;
  assign PEG_Yvec_11_fifo_aXvec_peek_empty_n = fifo_aXvec_11__empty_n;
  assign PEG_Yvec_11_fifo_aXvec_s_dout = fifo_aXvec_11__dout;
  assign PEG_Yvec_11_fifo_aXvec_s_empty_n = fifo_aXvec_11__empty_n;
  assign fifo_aXvec_11__read = PEG_Yvec_11_fifo_aXvec_s_read;
  assign PEG_Yvec_11_fifo_inst_in_peek_dout = Yvec_inst_11__dout;
  assign PEG_Yvec_11_fifo_inst_in_peek_empty_n = Yvec_inst_11__empty_n;
  assign PEG_Yvec_11_fifo_inst_in_s_dout = Yvec_inst_11__dout;
  assign PEG_Yvec_11_fifo_inst_in_s_empty_n = Yvec_inst_11__empty_n;
  assign Yvec_inst_11__read = PEG_Yvec_11_fifo_inst_in_s_read;
  assign PEG_Yvec_12_ap_clk = ap_clk;
  assign PEG_Yvec_12__ap_done = PEG_Yvec_12_ap_done;
  assign PEG_Yvec_12__ap_idle = PEG_Yvec_12_ap_idle;
  assign PEG_Yvec_12__ap_ready = PEG_Yvec_12_ap_ready;
  assign PEG_Yvec_12_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_12_ap_start = PEG_Yvec_12__ap_start;
  assign fifo_Y_pe_12__din = PEG_Yvec_12_fifo_Y_out_din;
  assign PEG_Yvec_12_fifo_Y_out_full_n = fifo_Y_pe_12__full_n;
  assign fifo_Y_pe_12__write = PEG_Yvec_12_fifo_Y_out_write;
  assign PEG_Yvec_12_fifo_aXvec_peek_dout = fifo_aXvec_12__dout;
  assign PEG_Yvec_12_fifo_aXvec_peek_empty_n = fifo_aXvec_12__empty_n;
  assign PEG_Yvec_12_fifo_aXvec_s_dout = fifo_aXvec_12__dout;
  assign PEG_Yvec_12_fifo_aXvec_s_empty_n = fifo_aXvec_12__empty_n;
  assign fifo_aXvec_12__read = PEG_Yvec_12_fifo_aXvec_s_read;
  assign PEG_Yvec_12_fifo_inst_in_peek_dout = Yvec_inst_12__dout;
  assign PEG_Yvec_12_fifo_inst_in_peek_empty_n = Yvec_inst_12__empty_n;
  assign PEG_Yvec_12_fifo_inst_in_s_dout = Yvec_inst_12__dout;
  assign PEG_Yvec_12_fifo_inst_in_s_empty_n = Yvec_inst_12__empty_n;
  assign Yvec_inst_12__read = PEG_Yvec_12_fifo_inst_in_s_read;
  assign PEG_Yvec_13_ap_clk = ap_clk;
  assign PEG_Yvec_13__ap_done = PEG_Yvec_13_ap_done;
  assign PEG_Yvec_13__ap_idle = PEG_Yvec_13_ap_idle;
  assign PEG_Yvec_13__ap_ready = PEG_Yvec_13_ap_ready;
  assign PEG_Yvec_13_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_13_ap_start = PEG_Yvec_13__ap_start;
  assign fifo_Y_pe_13__din = PEG_Yvec_13_fifo_Y_out_din;
  assign PEG_Yvec_13_fifo_Y_out_full_n = fifo_Y_pe_13__full_n;
  assign fifo_Y_pe_13__write = PEG_Yvec_13_fifo_Y_out_write;
  assign PEG_Yvec_13_fifo_aXvec_peek_dout = fifo_aXvec_13__dout;
  assign PEG_Yvec_13_fifo_aXvec_peek_empty_n = fifo_aXvec_13__empty_n;
  assign PEG_Yvec_13_fifo_aXvec_s_dout = fifo_aXvec_13__dout;
  assign PEG_Yvec_13_fifo_aXvec_s_empty_n = fifo_aXvec_13__empty_n;
  assign fifo_aXvec_13__read = PEG_Yvec_13_fifo_aXvec_s_read;
  assign PEG_Yvec_13_fifo_inst_in_peek_dout = Yvec_inst_13__dout;
  assign PEG_Yvec_13_fifo_inst_in_peek_empty_n = Yvec_inst_13__empty_n;
  assign PEG_Yvec_13_fifo_inst_in_s_dout = Yvec_inst_13__dout;
  assign PEG_Yvec_13_fifo_inst_in_s_empty_n = Yvec_inst_13__empty_n;
  assign Yvec_inst_13__read = PEG_Yvec_13_fifo_inst_in_s_read;
  assign PEG_Yvec_14_ap_clk = ap_clk;
  assign PEG_Yvec_14__ap_done = PEG_Yvec_14_ap_done;
  assign PEG_Yvec_14__ap_idle = PEG_Yvec_14_ap_idle;
  assign PEG_Yvec_14__ap_ready = PEG_Yvec_14_ap_ready;
  assign PEG_Yvec_14_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_14_ap_start = PEG_Yvec_14__ap_start;
  assign fifo_Y_pe_14__din = PEG_Yvec_14_fifo_Y_out_din;
  assign PEG_Yvec_14_fifo_Y_out_full_n = fifo_Y_pe_14__full_n;
  assign fifo_Y_pe_14__write = PEG_Yvec_14_fifo_Y_out_write;
  assign PEG_Yvec_14_fifo_aXvec_peek_dout = fifo_aXvec_14__dout;
  assign PEG_Yvec_14_fifo_aXvec_peek_empty_n = fifo_aXvec_14__empty_n;
  assign PEG_Yvec_14_fifo_aXvec_s_dout = fifo_aXvec_14__dout;
  assign PEG_Yvec_14_fifo_aXvec_s_empty_n = fifo_aXvec_14__empty_n;
  assign fifo_aXvec_14__read = PEG_Yvec_14_fifo_aXvec_s_read;
  assign PEG_Yvec_14_fifo_inst_in_peek_dout = Yvec_inst_14__dout;
  assign PEG_Yvec_14_fifo_inst_in_peek_empty_n = Yvec_inst_14__empty_n;
  assign PEG_Yvec_14_fifo_inst_in_s_dout = Yvec_inst_14__dout;
  assign PEG_Yvec_14_fifo_inst_in_s_empty_n = Yvec_inst_14__empty_n;
  assign Yvec_inst_14__read = PEG_Yvec_14_fifo_inst_in_s_read;
  assign PEG_Yvec_15_ap_clk = ap_clk;
  assign PEG_Yvec_15__ap_done = PEG_Yvec_15_ap_done;
  assign PEG_Yvec_15__ap_idle = PEG_Yvec_15_ap_idle;
  assign PEG_Yvec_15__ap_ready = PEG_Yvec_15_ap_ready;
  assign PEG_Yvec_15_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_15_ap_start = PEG_Yvec_15__ap_start;
  assign fifo_Y_pe_15__din = PEG_Yvec_15_fifo_Y_out_din;
  assign PEG_Yvec_15_fifo_Y_out_full_n = fifo_Y_pe_15__full_n;
  assign fifo_Y_pe_15__write = PEG_Yvec_15_fifo_Y_out_write;
  assign PEG_Yvec_15_fifo_aXvec_peek_dout = fifo_aXvec_15__dout;
  assign PEG_Yvec_15_fifo_aXvec_peek_empty_n = fifo_aXvec_15__empty_n;
  assign PEG_Yvec_15_fifo_aXvec_s_dout = fifo_aXvec_15__dout;
  assign PEG_Yvec_15_fifo_aXvec_s_empty_n = fifo_aXvec_15__empty_n;
  assign fifo_aXvec_15__read = PEG_Yvec_15_fifo_aXvec_s_read;
  assign PEG_Yvec_15_fifo_inst_in_peek_dout = Yvec_inst_15__dout;
  assign PEG_Yvec_15_fifo_inst_in_peek_empty_n = Yvec_inst_15__empty_n;
  assign PEG_Yvec_15_fifo_inst_in_s_dout = Yvec_inst_15__dout;
  assign PEG_Yvec_15_fifo_inst_in_s_empty_n = Yvec_inst_15__empty_n;
  assign Yvec_inst_15__read = PEG_Yvec_15_fifo_inst_in_s_read;
  assign PEG_Yvec_16_ap_clk = ap_clk;
  assign PEG_Yvec_16__ap_done = PEG_Yvec_16_ap_done;
  assign PEG_Yvec_16__ap_idle = PEG_Yvec_16_ap_idle;
  assign PEG_Yvec_16__ap_ready = PEG_Yvec_16_ap_ready;
  assign PEG_Yvec_16_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_16_ap_start = PEG_Yvec_16__ap_start;
  assign fifo_Y_pe_16__din = PEG_Yvec_16_fifo_Y_out_din;
  assign PEG_Yvec_16_fifo_Y_out_full_n = fifo_Y_pe_16__full_n;
  assign fifo_Y_pe_16__write = PEG_Yvec_16_fifo_Y_out_write;
  assign PEG_Yvec_16_fifo_aXvec_peek_dout = fifo_aXvec_16__dout;
  assign PEG_Yvec_16_fifo_aXvec_peek_empty_n = fifo_aXvec_16__empty_n;
  assign PEG_Yvec_16_fifo_aXvec_s_dout = fifo_aXvec_16__dout;
  assign PEG_Yvec_16_fifo_aXvec_s_empty_n = fifo_aXvec_16__empty_n;
  assign fifo_aXvec_16__read = PEG_Yvec_16_fifo_aXvec_s_read;
  assign PEG_Yvec_16_fifo_inst_in_peek_dout = Yvec_inst_16__dout;
  assign PEG_Yvec_16_fifo_inst_in_peek_empty_n = Yvec_inst_16__empty_n;
  assign PEG_Yvec_16_fifo_inst_in_s_dout = Yvec_inst_16__dout;
  assign PEG_Yvec_16_fifo_inst_in_s_empty_n = Yvec_inst_16__empty_n;
  assign Yvec_inst_16__read = PEG_Yvec_16_fifo_inst_in_s_read;
  assign PEG_Yvec_17_ap_clk = ap_clk;
  assign PEG_Yvec_17__ap_done = PEG_Yvec_17_ap_done;
  assign PEG_Yvec_17__ap_idle = PEG_Yvec_17_ap_idle;
  assign PEG_Yvec_17__ap_ready = PEG_Yvec_17_ap_ready;
  assign PEG_Yvec_17_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_17_ap_start = PEG_Yvec_17__ap_start;
  assign fifo_Y_pe_17__din = PEG_Yvec_17_fifo_Y_out_din;
  assign PEG_Yvec_17_fifo_Y_out_full_n = fifo_Y_pe_17__full_n;
  assign fifo_Y_pe_17__write = PEG_Yvec_17_fifo_Y_out_write;
  assign PEG_Yvec_17_fifo_aXvec_peek_dout = fifo_aXvec_17__dout;
  assign PEG_Yvec_17_fifo_aXvec_peek_empty_n = fifo_aXvec_17__empty_n;
  assign PEG_Yvec_17_fifo_aXvec_s_dout = fifo_aXvec_17__dout;
  assign PEG_Yvec_17_fifo_aXvec_s_empty_n = fifo_aXvec_17__empty_n;
  assign fifo_aXvec_17__read = PEG_Yvec_17_fifo_aXvec_s_read;
  assign PEG_Yvec_17_fifo_inst_in_peek_dout = Yvec_inst_17__dout;
  assign PEG_Yvec_17_fifo_inst_in_peek_empty_n = Yvec_inst_17__empty_n;
  assign PEG_Yvec_17_fifo_inst_in_s_dout = Yvec_inst_17__dout;
  assign PEG_Yvec_17_fifo_inst_in_s_empty_n = Yvec_inst_17__empty_n;
  assign Yvec_inst_17__read = PEG_Yvec_17_fifo_inst_in_s_read;
  assign PEG_Yvec_18_ap_clk = ap_clk;
  assign PEG_Yvec_18__ap_done = PEG_Yvec_18_ap_done;
  assign PEG_Yvec_18__ap_idle = PEG_Yvec_18_ap_idle;
  assign PEG_Yvec_18__ap_ready = PEG_Yvec_18_ap_ready;
  assign PEG_Yvec_18_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_18_ap_start = PEG_Yvec_18__ap_start;
  assign fifo_Y_pe_18__din = PEG_Yvec_18_fifo_Y_out_din;
  assign PEG_Yvec_18_fifo_Y_out_full_n = fifo_Y_pe_18__full_n;
  assign fifo_Y_pe_18__write = PEG_Yvec_18_fifo_Y_out_write;
  assign PEG_Yvec_18_fifo_aXvec_peek_dout = fifo_aXvec_18__dout;
  assign PEG_Yvec_18_fifo_aXvec_peek_empty_n = fifo_aXvec_18__empty_n;
  assign PEG_Yvec_18_fifo_aXvec_s_dout = fifo_aXvec_18__dout;
  assign PEG_Yvec_18_fifo_aXvec_s_empty_n = fifo_aXvec_18__empty_n;
  assign fifo_aXvec_18__read = PEG_Yvec_18_fifo_aXvec_s_read;
  assign PEG_Yvec_18_fifo_inst_in_peek_dout = Yvec_inst_18__dout;
  assign PEG_Yvec_18_fifo_inst_in_peek_empty_n = Yvec_inst_18__empty_n;
  assign PEG_Yvec_18_fifo_inst_in_s_dout = Yvec_inst_18__dout;
  assign PEG_Yvec_18_fifo_inst_in_s_empty_n = Yvec_inst_18__empty_n;
  assign Yvec_inst_18__read = PEG_Yvec_18_fifo_inst_in_s_read;
  assign PEG_Yvec_19_ap_clk = ap_clk;
  assign PEG_Yvec_19__ap_done = PEG_Yvec_19_ap_done;
  assign PEG_Yvec_19__ap_idle = PEG_Yvec_19_ap_idle;
  assign PEG_Yvec_19__ap_ready = PEG_Yvec_19_ap_ready;
  assign PEG_Yvec_19_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_19_ap_start = PEG_Yvec_19__ap_start;
  assign fifo_Y_pe_19__din = PEG_Yvec_19_fifo_Y_out_din;
  assign PEG_Yvec_19_fifo_Y_out_full_n = fifo_Y_pe_19__full_n;
  assign fifo_Y_pe_19__write = PEG_Yvec_19_fifo_Y_out_write;
  assign PEG_Yvec_19_fifo_aXvec_peek_dout = fifo_aXvec_19__dout;
  assign PEG_Yvec_19_fifo_aXvec_peek_empty_n = fifo_aXvec_19__empty_n;
  assign PEG_Yvec_19_fifo_aXvec_s_dout = fifo_aXvec_19__dout;
  assign PEG_Yvec_19_fifo_aXvec_s_empty_n = fifo_aXvec_19__empty_n;
  assign fifo_aXvec_19__read = PEG_Yvec_19_fifo_aXvec_s_read;
  assign PEG_Yvec_19_fifo_inst_in_peek_dout = Yvec_inst_19__dout;
  assign PEG_Yvec_19_fifo_inst_in_peek_empty_n = Yvec_inst_19__empty_n;
  assign PEG_Yvec_19_fifo_inst_in_s_dout = Yvec_inst_19__dout;
  assign PEG_Yvec_19_fifo_inst_in_s_empty_n = Yvec_inst_19__empty_n;
  assign Yvec_inst_19__read = PEG_Yvec_19_fifo_inst_in_s_read;
  assign PEG_Yvec_20_ap_clk = ap_clk;
  assign PEG_Yvec_20__ap_done = PEG_Yvec_20_ap_done;
  assign PEG_Yvec_20__ap_idle = PEG_Yvec_20_ap_idle;
  assign PEG_Yvec_20__ap_ready = PEG_Yvec_20_ap_ready;
  assign PEG_Yvec_20_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_20_ap_start = PEG_Yvec_20__ap_start;
  assign fifo_Y_pe_20__din = PEG_Yvec_20_fifo_Y_out_din;
  assign PEG_Yvec_20_fifo_Y_out_full_n = fifo_Y_pe_20__full_n;
  assign fifo_Y_pe_20__write = PEG_Yvec_20_fifo_Y_out_write;
  assign PEG_Yvec_20_fifo_aXvec_peek_dout = fifo_aXvec_20__dout;
  assign PEG_Yvec_20_fifo_aXvec_peek_empty_n = fifo_aXvec_20__empty_n;
  assign PEG_Yvec_20_fifo_aXvec_s_dout = fifo_aXvec_20__dout;
  assign PEG_Yvec_20_fifo_aXvec_s_empty_n = fifo_aXvec_20__empty_n;
  assign fifo_aXvec_20__read = PEG_Yvec_20_fifo_aXvec_s_read;
  assign PEG_Yvec_20_fifo_inst_in_peek_dout = Yvec_inst_20__dout;
  assign PEG_Yvec_20_fifo_inst_in_peek_empty_n = Yvec_inst_20__empty_n;
  assign PEG_Yvec_20_fifo_inst_in_s_dout = Yvec_inst_20__dout;
  assign PEG_Yvec_20_fifo_inst_in_s_empty_n = Yvec_inst_20__empty_n;
  assign Yvec_inst_20__read = PEG_Yvec_20_fifo_inst_in_s_read;
  assign PEG_Yvec_21_ap_clk = ap_clk;
  assign PEG_Yvec_21__ap_done = PEG_Yvec_21_ap_done;
  assign PEG_Yvec_21__ap_idle = PEG_Yvec_21_ap_idle;
  assign PEG_Yvec_21__ap_ready = PEG_Yvec_21_ap_ready;
  assign PEG_Yvec_21_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_21_ap_start = PEG_Yvec_21__ap_start;
  assign fifo_Y_pe_21__din = PEG_Yvec_21_fifo_Y_out_din;
  assign PEG_Yvec_21_fifo_Y_out_full_n = fifo_Y_pe_21__full_n;
  assign fifo_Y_pe_21__write = PEG_Yvec_21_fifo_Y_out_write;
  assign PEG_Yvec_21_fifo_aXvec_peek_dout = fifo_aXvec_21__dout;
  assign PEG_Yvec_21_fifo_aXvec_peek_empty_n = fifo_aXvec_21__empty_n;
  assign PEG_Yvec_21_fifo_aXvec_s_dout = fifo_aXvec_21__dout;
  assign PEG_Yvec_21_fifo_aXvec_s_empty_n = fifo_aXvec_21__empty_n;
  assign fifo_aXvec_21__read = PEG_Yvec_21_fifo_aXvec_s_read;
  assign PEG_Yvec_21_fifo_inst_in_peek_dout = Yvec_inst_21__dout;
  assign PEG_Yvec_21_fifo_inst_in_peek_empty_n = Yvec_inst_21__empty_n;
  assign PEG_Yvec_21_fifo_inst_in_s_dout = Yvec_inst_21__dout;
  assign PEG_Yvec_21_fifo_inst_in_s_empty_n = Yvec_inst_21__empty_n;
  assign Yvec_inst_21__read = PEG_Yvec_21_fifo_inst_in_s_read;
  assign PEG_Yvec_22_ap_clk = ap_clk;
  assign PEG_Yvec_22__ap_done = PEG_Yvec_22_ap_done;
  assign PEG_Yvec_22__ap_idle = PEG_Yvec_22_ap_idle;
  assign PEG_Yvec_22__ap_ready = PEG_Yvec_22_ap_ready;
  assign PEG_Yvec_22_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_22_ap_start = PEG_Yvec_22__ap_start;
  assign fifo_Y_pe_22__din = PEG_Yvec_22_fifo_Y_out_din;
  assign PEG_Yvec_22_fifo_Y_out_full_n = fifo_Y_pe_22__full_n;
  assign fifo_Y_pe_22__write = PEG_Yvec_22_fifo_Y_out_write;
  assign PEG_Yvec_22_fifo_aXvec_peek_dout = fifo_aXvec_22__dout;
  assign PEG_Yvec_22_fifo_aXvec_peek_empty_n = fifo_aXvec_22__empty_n;
  assign PEG_Yvec_22_fifo_aXvec_s_dout = fifo_aXvec_22__dout;
  assign PEG_Yvec_22_fifo_aXvec_s_empty_n = fifo_aXvec_22__empty_n;
  assign fifo_aXvec_22__read = PEG_Yvec_22_fifo_aXvec_s_read;
  assign PEG_Yvec_22_fifo_inst_in_peek_dout = Yvec_inst_22__dout;
  assign PEG_Yvec_22_fifo_inst_in_peek_empty_n = Yvec_inst_22__empty_n;
  assign PEG_Yvec_22_fifo_inst_in_s_dout = Yvec_inst_22__dout;
  assign PEG_Yvec_22_fifo_inst_in_s_empty_n = Yvec_inst_22__empty_n;
  assign Yvec_inst_22__read = PEG_Yvec_22_fifo_inst_in_s_read;
  assign PEG_Yvec_23_ap_clk = ap_clk;
  assign PEG_Yvec_23__ap_done = PEG_Yvec_23_ap_done;
  assign PEG_Yvec_23__ap_idle = PEG_Yvec_23_ap_idle;
  assign PEG_Yvec_23__ap_ready = PEG_Yvec_23_ap_ready;
  assign PEG_Yvec_23_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_23_ap_start = PEG_Yvec_23__ap_start;
  assign fifo_Y_pe_23__din = PEG_Yvec_23_fifo_Y_out_din;
  assign PEG_Yvec_23_fifo_Y_out_full_n = fifo_Y_pe_23__full_n;
  assign fifo_Y_pe_23__write = PEG_Yvec_23_fifo_Y_out_write;
  assign PEG_Yvec_23_fifo_aXvec_peek_dout = fifo_aXvec_23__dout;
  assign PEG_Yvec_23_fifo_aXvec_peek_empty_n = fifo_aXvec_23__empty_n;
  assign PEG_Yvec_23_fifo_aXvec_s_dout = fifo_aXvec_23__dout;
  assign PEG_Yvec_23_fifo_aXvec_s_empty_n = fifo_aXvec_23__empty_n;
  assign fifo_aXvec_23__read = PEG_Yvec_23_fifo_aXvec_s_read;
  assign PEG_Yvec_23_fifo_inst_in_peek_dout = Yvec_inst_23__dout;
  assign PEG_Yvec_23_fifo_inst_in_peek_empty_n = Yvec_inst_23__empty_n;
  assign PEG_Yvec_23_fifo_inst_in_s_dout = Yvec_inst_23__dout;
  assign PEG_Yvec_23_fifo_inst_in_s_empty_n = Yvec_inst_23__empty_n;
  assign Yvec_inst_23__read = PEG_Yvec_23_fifo_inst_in_s_read;
  assign PEG_Yvec_24_ap_clk = ap_clk;
  assign PEG_Yvec_24__ap_done = PEG_Yvec_24_ap_done;
  assign PEG_Yvec_24__ap_idle = PEG_Yvec_24_ap_idle;
  assign PEG_Yvec_24__ap_ready = PEG_Yvec_24_ap_ready;
  assign PEG_Yvec_24_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_24_ap_start = PEG_Yvec_24__ap_start;
  assign fifo_Y_pe_24__din = PEG_Yvec_24_fifo_Y_out_din;
  assign PEG_Yvec_24_fifo_Y_out_full_n = fifo_Y_pe_24__full_n;
  assign fifo_Y_pe_24__write = PEG_Yvec_24_fifo_Y_out_write;
  assign PEG_Yvec_24_fifo_aXvec_peek_dout = fifo_aXvec_24__dout;
  assign PEG_Yvec_24_fifo_aXvec_peek_empty_n = fifo_aXvec_24__empty_n;
  assign PEG_Yvec_24_fifo_aXvec_s_dout = fifo_aXvec_24__dout;
  assign PEG_Yvec_24_fifo_aXvec_s_empty_n = fifo_aXvec_24__empty_n;
  assign fifo_aXvec_24__read = PEG_Yvec_24_fifo_aXvec_s_read;
  assign PEG_Yvec_24_fifo_inst_in_peek_dout = Yvec_inst_24__dout;
  assign PEG_Yvec_24_fifo_inst_in_peek_empty_n = Yvec_inst_24__empty_n;
  assign PEG_Yvec_24_fifo_inst_in_s_dout = Yvec_inst_24__dout;
  assign PEG_Yvec_24_fifo_inst_in_s_empty_n = Yvec_inst_24__empty_n;
  assign Yvec_inst_24__read = PEG_Yvec_24_fifo_inst_in_s_read;
  assign PEG_Yvec_25_ap_clk = ap_clk;
  assign PEG_Yvec_25__ap_done = PEG_Yvec_25_ap_done;
  assign PEG_Yvec_25__ap_idle = PEG_Yvec_25_ap_idle;
  assign PEG_Yvec_25__ap_ready = PEG_Yvec_25_ap_ready;
  assign PEG_Yvec_25_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_25_ap_start = PEG_Yvec_25__ap_start;
  assign fifo_Y_pe_25__din = PEG_Yvec_25_fifo_Y_out_din;
  assign PEG_Yvec_25_fifo_Y_out_full_n = fifo_Y_pe_25__full_n;
  assign fifo_Y_pe_25__write = PEG_Yvec_25_fifo_Y_out_write;
  assign PEG_Yvec_25_fifo_aXvec_peek_dout = fifo_aXvec_25__dout;
  assign PEG_Yvec_25_fifo_aXvec_peek_empty_n = fifo_aXvec_25__empty_n;
  assign PEG_Yvec_25_fifo_aXvec_s_dout = fifo_aXvec_25__dout;
  assign PEG_Yvec_25_fifo_aXvec_s_empty_n = fifo_aXvec_25__empty_n;
  assign fifo_aXvec_25__read = PEG_Yvec_25_fifo_aXvec_s_read;
  assign PEG_Yvec_25_fifo_inst_in_peek_dout = Yvec_inst_25__dout;
  assign PEG_Yvec_25_fifo_inst_in_peek_empty_n = Yvec_inst_25__empty_n;
  assign PEG_Yvec_25_fifo_inst_in_s_dout = Yvec_inst_25__dout;
  assign PEG_Yvec_25_fifo_inst_in_s_empty_n = Yvec_inst_25__empty_n;
  assign Yvec_inst_25__read = PEG_Yvec_25_fifo_inst_in_s_read;
  assign PEG_Yvec_26_ap_clk = ap_clk;
  assign PEG_Yvec_26__ap_done = PEG_Yvec_26_ap_done;
  assign PEG_Yvec_26__ap_idle = PEG_Yvec_26_ap_idle;
  assign PEG_Yvec_26__ap_ready = PEG_Yvec_26_ap_ready;
  assign PEG_Yvec_26_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_26_ap_start = PEG_Yvec_26__ap_start;
  assign fifo_Y_pe_26__din = PEG_Yvec_26_fifo_Y_out_din;
  assign PEG_Yvec_26_fifo_Y_out_full_n = fifo_Y_pe_26__full_n;
  assign fifo_Y_pe_26__write = PEG_Yvec_26_fifo_Y_out_write;
  assign PEG_Yvec_26_fifo_aXvec_peek_dout = fifo_aXvec_26__dout;
  assign PEG_Yvec_26_fifo_aXvec_peek_empty_n = fifo_aXvec_26__empty_n;
  assign PEG_Yvec_26_fifo_aXvec_s_dout = fifo_aXvec_26__dout;
  assign PEG_Yvec_26_fifo_aXvec_s_empty_n = fifo_aXvec_26__empty_n;
  assign fifo_aXvec_26__read = PEG_Yvec_26_fifo_aXvec_s_read;
  assign PEG_Yvec_26_fifo_inst_in_peek_dout = Yvec_inst_26__dout;
  assign PEG_Yvec_26_fifo_inst_in_peek_empty_n = Yvec_inst_26__empty_n;
  assign PEG_Yvec_26_fifo_inst_in_s_dout = Yvec_inst_26__dout;
  assign PEG_Yvec_26_fifo_inst_in_s_empty_n = Yvec_inst_26__empty_n;
  assign Yvec_inst_26__read = PEG_Yvec_26_fifo_inst_in_s_read;
  assign PEG_Yvec_27_ap_clk = ap_clk;
  assign PEG_Yvec_27__ap_done = PEG_Yvec_27_ap_done;
  assign PEG_Yvec_27__ap_idle = PEG_Yvec_27_ap_idle;
  assign PEG_Yvec_27__ap_ready = PEG_Yvec_27_ap_ready;
  assign PEG_Yvec_27_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_27_ap_start = PEG_Yvec_27__ap_start;
  assign fifo_Y_pe_27__din = PEG_Yvec_27_fifo_Y_out_din;
  assign PEG_Yvec_27_fifo_Y_out_full_n = fifo_Y_pe_27__full_n;
  assign fifo_Y_pe_27__write = PEG_Yvec_27_fifo_Y_out_write;
  assign PEG_Yvec_27_fifo_aXvec_peek_dout = fifo_aXvec_27__dout;
  assign PEG_Yvec_27_fifo_aXvec_peek_empty_n = fifo_aXvec_27__empty_n;
  assign PEG_Yvec_27_fifo_aXvec_s_dout = fifo_aXvec_27__dout;
  assign PEG_Yvec_27_fifo_aXvec_s_empty_n = fifo_aXvec_27__empty_n;
  assign fifo_aXvec_27__read = PEG_Yvec_27_fifo_aXvec_s_read;
  assign PEG_Yvec_27_fifo_inst_in_peek_dout = Yvec_inst_27__dout;
  assign PEG_Yvec_27_fifo_inst_in_peek_empty_n = Yvec_inst_27__empty_n;
  assign PEG_Yvec_27_fifo_inst_in_s_dout = Yvec_inst_27__dout;
  assign PEG_Yvec_27_fifo_inst_in_s_empty_n = Yvec_inst_27__empty_n;
  assign Yvec_inst_27__read = PEG_Yvec_27_fifo_inst_in_s_read;
  assign PEG_Yvec_28_ap_clk = ap_clk;
  assign PEG_Yvec_28__ap_done = PEG_Yvec_28_ap_done;
  assign PEG_Yvec_28__ap_idle = PEG_Yvec_28_ap_idle;
  assign PEG_Yvec_28__ap_ready = PEG_Yvec_28_ap_ready;
  assign PEG_Yvec_28_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_28_ap_start = PEG_Yvec_28__ap_start;
  assign fifo_Y_pe_28__din = PEG_Yvec_28_fifo_Y_out_din;
  assign PEG_Yvec_28_fifo_Y_out_full_n = fifo_Y_pe_28__full_n;
  assign fifo_Y_pe_28__write = PEG_Yvec_28_fifo_Y_out_write;
  assign PEG_Yvec_28_fifo_aXvec_peek_dout = fifo_aXvec_28__dout;
  assign PEG_Yvec_28_fifo_aXvec_peek_empty_n = fifo_aXvec_28__empty_n;
  assign PEG_Yvec_28_fifo_aXvec_s_dout = fifo_aXvec_28__dout;
  assign PEG_Yvec_28_fifo_aXvec_s_empty_n = fifo_aXvec_28__empty_n;
  assign fifo_aXvec_28__read = PEG_Yvec_28_fifo_aXvec_s_read;
  assign PEG_Yvec_28_fifo_inst_in_peek_dout = Yvec_inst_28__dout;
  assign PEG_Yvec_28_fifo_inst_in_peek_empty_n = Yvec_inst_28__empty_n;
  assign PEG_Yvec_28_fifo_inst_in_s_dout = Yvec_inst_28__dout;
  assign PEG_Yvec_28_fifo_inst_in_s_empty_n = Yvec_inst_28__empty_n;
  assign Yvec_inst_28__read = PEG_Yvec_28_fifo_inst_in_s_read;
  assign PEG_Yvec_29_ap_clk = ap_clk;
  assign PEG_Yvec_29__ap_done = PEG_Yvec_29_ap_done;
  assign PEG_Yvec_29__ap_idle = PEG_Yvec_29_ap_idle;
  assign PEG_Yvec_29__ap_ready = PEG_Yvec_29_ap_ready;
  assign PEG_Yvec_29_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_29_ap_start = PEG_Yvec_29__ap_start;
  assign fifo_Y_pe_29__din = PEG_Yvec_29_fifo_Y_out_din;
  assign PEG_Yvec_29_fifo_Y_out_full_n = fifo_Y_pe_29__full_n;
  assign fifo_Y_pe_29__write = PEG_Yvec_29_fifo_Y_out_write;
  assign PEG_Yvec_29_fifo_aXvec_peek_dout = fifo_aXvec_29__dout;
  assign PEG_Yvec_29_fifo_aXvec_peek_empty_n = fifo_aXvec_29__empty_n;
  assign PEG_Yvec_29_fifo_aXvec_s_dout = fifo_aXvec_29__dout;
  assign PEG_Yvec_29_fifo_aXvec_s_empty_n = fifo_aXvec_29__empty_n;
  assign fifo_aXvec_29__read = PEG_Yvec_29_fifo_aXvec_s_read;
  assign PEG_Yvec_29_fifo_inst_in_peek_dout = Yvec_inst_29__dout;
  assign PEG_Yvec_29_fifo_inst_in_peek_empty_n = Yvec_inst_29__empty_n;
  assign PEG_Yvec_29_fifo_inst_in_s_dout = Yvec_inst_29__dout;
  assign PEG_Yvec_29_fifo_inst_in_s_empty_n = Yvec_inst_29__empty_n;
  assign Yvec_inst_29__read = PEG_Yvec_29_fifo_inst_in_s_read;
  assign PEG_Yvec_30_ap_clk = ap_clk;
  assign PEG_Yvec_30__ap_done = PEG_Yvec_30_ap_done;
  assign PEG_Yvec_30__ap_idle = PEG_Yvec_30_ap_idle;
  assign PEG_Yvec_30__ap_ready = PEG_Yvec_30_ap_ready;
  assign PEG_Yvec_30_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_30_ap_start = PEG_Yvec_30__ap_start;
  assign fifo_Y_pe_30__din = PEG_Yvec_30_fifo_Y_out_din;
  assign PEG_Yvec_30_fifo_Y_out_full_n = fifo_Y_pe_30__full_n;
  assign fifo_Y_pe_30__write = PEG_Yvec_30_fifo_Y_out_write;
  assign PEG_Yvec_30_fifo_aXvec_peek_dout = fifo_aXvec_30__dout;
  assign PEG_Yvec_30_fifo_aXvec_peek_empty_n = fifo_aXvec_30__empty_n;
  assign PEG_Yvec_30_fifo_aXvec_s_dout = fifo_aXvec_30__dout;
  assign PEG_Yvec_30_fifo_aXvec_s_empty_n = fifo_aXvec_30__empty_n;
  assign fifo_aXvec_30__read = PEG_Yvec_30_fifo_aXvec_s_read;
  assign PEG_Yvec_30_fifo_inst_in_peek_dout = Yvec_inst_30__dout;
  assign PEG_Yvec_30_fifo_inst_in_peek_empty_n = Yvec_inst_30__empty_n;
  assign PEG_Yvec_30_fifo_inst_in_s_dout = Yvec_inst_30__dout;
  assign PEG_Yvec_30_fifo_inst_in_s_empty_n = Yvec_inst_30__empty_n;
  assign Yvec_inst_30__read = PEG_Yvec_30_fifo_inst_in_s_read;
  assign PEG_Yvec_31_ap_clk = ap_clk;
  assign PEG_Yvec_31__ap_done = PEG_Yvec_31_ap_done;
  assign PEG_Yvec_31__ap_idle = PEG_Yvec_31_ap_idle;
  assign PEG_Yvec_31__ap_ready = PEG_Yvec_31_ap_ready;
  assign PEG_Yvec_31_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_31_ap_start = PEG_Yvec_31__ap_start;
  assign fifo_Y_pe_31__din = PEG_Yvec_31_fifo_Y_out_din;
  assign PEG_Yvec_31_fifo_Y_out_full_n = fifo_Y_pe_31__full_n;
  assign fifo_Y_pe_31__write = PEG_Yvec_31_fifo_Y_out_write;
  assign PEG_Yvec_31_fifo_aXvec_peek_dout = fifo_aXvec_31__dout;
  assign PEG_Yvec_31_fifo_aXvec_peek_empty_n = fifo_aXvec_31__empty_n;
  assign PEG_Yvec_31_fifo_aXvec_s_dout = fifo_aXvec_31__dout;
  assign PEG_Yvec_31_fifo_aXvec_s_empty_n = fifo_aXvec_31__empty_n;
  assign fifo_aXvec_31__read = PEG_Yvec_31_fifo_aXvec_s_read;
  assign PEG_Yvec_31_fifo_inst_in_peek_dout = Yvec_inst_31__dout;
  assign PEG_Yvec_31_fifo_inst_in_peek_empty_n = Yvec_inst_31__empty_n;
  assign PEG_Yvec_31_fifo_inst_in_s_dout = Yvec_inst_31__dout;
  assign PEG_Yvec_31_fifo_inst_in_s_empty_n = Yvec_inst_31__empty_n;
  assign Yvec_inst_31__read = PEG_Yvec_31_fifo_inst_in_s_read;
  assign PEG_Yvec_32_ap_clk = ap_clk;
  assign PEG_Yvec_32__ap_done = PEG_Yvec_32_ap_done;
  assign PEG_Yvec_32__ap_idle = PEG_Yvec_32_ap_idle;
  assign PEG_Yvec_32__ap_ready = PEG_Yvec_32_ap_ready;
  assign PEG_Yvec_32_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_32_ap_start = PEG_Yvec_32__ap_start;
  assign fifo_Y_pe_32__din = PEG_Yvec_32_fifo_Y_out_din;
  assign PEG_Yvec_32_fifo_Y_out_full_n = fifo_Y_pe_32__full_n;
  assign fifo_Y_pe_32__write = PEG_Yvec_32_fifo_Y_out_write;
  assign PEG_Yvec_32_fifo_aXvec_peek_dout = fifo_aXvec_32__dout;
  assign PEG_Yvec_32_fifo_aXvec_peek_empty_n = fifo_aXvec_32__empty_n;
  assign PEG_Yvec_32_fifo_aXvec_s_dout = fifo_aXvec_32__dout;
  assign PEG_Yvec_32_fifo_aXvec_s_empty_n = fifo_aXvec_32__empty_n;
  assign fifo_aXvec_32__read = PEG_Yvec_32_fifo_aXvec_s_read;
  assign PEG_Yvec_32_fifo_inst_in_peek_dout = Yvec_inst_32__dout;
  assign PEG_Yvec_32_fifo_inst_in_peek_empty_n = Yvec_inst_32__empty_n;
  assign PEG_Yvec_32_fifo_inst_in_s_dout = Yvec_inst_32__dout;
  assign PEG_Yvec_32_fifo_inst_in_s_empty_n = Yvec_inst_32__empty_n;
  assign Yvec_inst_32__read = PEG_Yvec_32_fifo_inst_in_s_read;
  assign PEG_Yvec_33_ap_clk = ap_clk;
  assign PEG_Yvec_33__ap_done = PEG_Yvec_33_ap_done;
  assign PEG_Yvec_33__ap_idle = PEG_Yvec_33_ap_idle;
  assign PEG_Yvec_33__ap_ready = PEG_Yvec_33_ap_ready;
  assign PEG_Yvec_33_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_33_ap_start = PEG_Yvec_33__ap_start;
  assign fifo_Y_pe_33__din = PEG_Yvec_33_fifo_Y_out_din;
  assign PEG_Yvec_33_fifo_Y_out_full_n = fifo_Y_pe_33__full_n;
  assign fifo_Y_pe_33__write = PEG_Yvec_33_fifo_Y_out_write;
  assign PEG_Yvec_33_fifo_aXvec_peek_dout = fifo_aXvec_33__dout;
  assign PEG_Yvec_33_fifo_aXvec_peek_empty_n = fifo_aXvec_33__empty_n;
  assign PEG_Yvec_33_fifo_aXvec_s_dout = fifo_aXvec_33__dout;
  assign PEG_Yvec_33_fifo_aXvec_s_empty_n = fifo_aXvec_33__empty_n;
  assign fifo_aXvec_33__read = PEG_Yvec_33_fifo_aXvec_s_read;
  assign PEG_Yvec_33_fifo_inst_in_peek_dout = Yvec_inst_33__dout;
  assign PEG_Yvec_33_fifo_inst_in_peek_empty_n = Yvec_inst_33__empty_n;
  assign PEG_Yvec_33_fifo_inst_in_s_dout = Yvec_inst_33__dout;
  assign PEG_Yvec_33_fifo_inst_in_s_empty_n = Yvec_inst_33__empty_n;
  assign Yvec_inst_33__read = PEG_Yvec_33_fifo_inst_in_s_read;
  assign PEG_Yvec_34_ap_clk = ap_clk;
  assign PEG_Yvec_34__ap_done = PEG_Yvec_34_ap_done;
  assign PEG_Yvec_34__ap_idle = PEG_Yvec_34_ap_idle;
  assign PEG_Yvec_34__ap_ready = PEG_Yvec_34_ap_ready;
  assign PEG_Yvec_34_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_34_ap_start = PEG_Yvec_34__ap_start;
  assign fifo_Y_pe_34__din = PEG_Yvec_34_fifo_Y_out_din;
  assign PEG_Yvec_34_fifo_Y_out_full_n = fifo_Y_pe_34__full_n;
  assign fifo_Y_pe_34__write = PEG_Yvec_34_fifo_Y_out_write;
  assign PEG_Yvec_34_fifo_aXvec_peek_dout = fifo_aXvec_34__dout;
  assign PEG_Yvec_34_fifo_aXvec_peek_empty_n = fifo_aXvec_34__empty_n;
  assign PEG_Yvec_34_fifo_aXvec_s_dout = fifo_aXvec_34__dout;
  assign PEG_Yvec_34_fifo_aXvec_s_empty_n = fifo_aXvec_34__empty_n;
  assign fifo_aXvec_34__read = PEG_Yvec_34_fifo_aXvec_s_read;
  assign PEG_Yvec_34_fifo_inst_in_peek_dout = Yvec_inst_34__dout;
  assign PEG_Yvec_34_fifo_inst_in_peek_empty_n = Yvec_inst_34__empty_n;
  assign PEG_Yvec_34_fifo_inst_in_s_dout = Yvec_inst_34__dout;
  assign PEG_Yvec_34_fifo_inst_in_s_empty_n = Yvec_inst_34__empty_n;
  assign Yvec_inst_34__read = PEG_Yvec_34_fifo_inst_in_s_read;
  assign PEG_Yvec_35_ap_clk = ap_clk;
  assign PEG_Yvec_35__ap_done = PEG_Yvec_35_ap_done;
  assign PEG_Yvec_35__ap_idle = PEG_Yvec_35_ap_idle;
  assign PEG_Yvec_35__ap_ready = PEG_Yvec_35_ap_ready;
  assign PEG_Yvec_35_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_35_ap_start = PEG_Yvec_35__ap_start;
  assign fifo_Y_pe_35__din = PEG_Yvec_35_fifo_Y_out_din;
  assign PEG_Yvec_35_fifo_Y_out_full_n = fifo_Y_pe_35__full_n;
  assign fifo_Y_pe_35__write = PEG_Yvec_35_fifo_Y_out_write;
  assign PEG_Yvec_35_fifo_aXvec_peek_dout = fifo_aXvec_35__dout;
  assign PEG_Yvec_35_fifo_aXvec_peek_empty_n = fifo_aXvec_35__empty_n;
  assign PEG_Yvec_35_fifo_aXvec_s_dout = fifo_aXvec_35__dout;
  assign PEG_Yvec_35_fifo_aXvec_s_empty_n = fifo_aXvec_35__empty_n;
  assign fifo_aXvec_35__read = PEG_Yvec_35_fifo_aXvec_s_read;
  assign PEG_Yvec_35_fifo_inst_in_peek_dout = Yvec_inst_35__dout;
  assign PEG_Yvec_35_fifo_inst_in_peek_empty_n = Yvec_inst_35__empty_n;
  assign PEG_Yvec_35_fifo_inst_in_s_dout = Yvec_inst_35__dout;
  assign PEG_Yvec_35_fifo_inst_in_s_empty_n = Yvec_inst_35__empty_n;
  assign Yvec_inst_35__read = PEG_Yvec_35_fifo_inst_in_s_read;
  assign PEG_Yvec_36_ap_clk = ap_clk;
  assign PEG_Yvec_36__ap_done = PEG_Yvec_36_ap_done;
  assign PEG_Yvec_36__ap_idle = PEG_Yvec_36_ap_idle;
  assign PEG_Yvec_36__ap_ready = PEG_Yvec_36_ap_ready;
  assign PEG_Yvec_36_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_36_ap_start = PEG_Yvec_36__ap_start;
  assign fifo_Y_pe_36__din = PEG_Yvec_36_fifo_Y_out_din;
  assign PEG_Yvec_36_fifo_Y_out_full_n = fifo_Y_pe_36__full_n;
  assign fifo_Y_pe_36__write = PEG_Yvec_36_fifo_Y_out_write;
  assign PEG_Yvec_36_fifo_aXvec_peek_dout = fifo_aXvec_36__dout;
  assign PEG_Yvec_36_fifo_aXvec_peek_empty_n = fifo_aXvec_36__empty_n;
  assign PEG_Yvec_36_fifo_aXvec_s_dout = fifo_aXvec_36__dout;
  assign PEG_Yvec_36_fifo_aXvec_s_empty_n = fifo_aXvec_36__empty_n;
  assign fifo_aXvec_36__read = PEG_Yvec_36_fifo_aXvec_s_read;
  assign PEG_Yvec_36_fifo_inst_in_peek_dout = Yvec_inst_36__dout;
  assign PEG_Yvec_36_fifo_inst_in_peek_empty_n = Yvec_inst_36__empty_n;
  assign PEG_Yvec_36_fifo_inst_in_s_dout = Yvec_inst_36__dout;
  assign PEG_Yvec_36_fifo_inst_in_s_empty_n = Yvec_inst_36__empty_n;
  assign Yvec_inst_36__read = PEG_Yvec_36_fifo_inst_in_s_read;
  assign PEG_Yvec_37_ap_clk = ap_clk;
  assign PEG_Yvec_37__ap_done = PEG_Yvec_37_ap_done;
  assign PEG_Yvec_37__ap_idle = PEG_Yvec_37_ap_idle;
  assign PEG_Yvec_37__ap_ready = PEG_Yvec_37_ap_ready;
  assign PEG_Yvec_37_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_37_ap_start = PEG_Yvec_37__ap_start;
  assign fifo_Y_pe_37__din = PEG_Yvec_37_fifo_Y_out_din;
  assign PEG_Yvec_37_fifo_Y_out_full_n = fifo_Y_pe_37__full_n;
  assign fifo_Y_pe_37__write = PEG_Yvec_37_fifo_Y_out_write;
  assign PEG_Yvec_37_fifo_aXvec_peek_dout = fifo_aXvec_37__dout;
  assign PEG_Yvec_37_fifo_aXvec_peek_empty_n = fifo_aXvec_37__empty_n;
  assign PEG_Yvec_37_fifo_aXvec_s_dout = fifo_aXvec_37__dout;
  assign PEG_Yvec_37_fifo_aXvec_s_empty_n = fifo_aXvec_37__empty_n;
  assign fifo_aXvec_37__read = PEG_Yvec_37_fifo_aXvec_s_read;
  assign PEG_Yvec_37_fifo_inst_in_peek_dout = Yvec_inst_37__dout;
  assign PEG_Yvec_37_fifo_inst_in_peek_empty_n = Yvec_inst_37__empty_n;
  assign PEG_Yvec_37_fifo_inst_in_s_dout = Yvec_inst_37__dout;
  assign PEG_Yvec_37_fifo_inst_in_s_empty_n = Yvec_inst_37__empty_n;
  assign Yvec_inst_37__read = PEG_Yvec_37_fifo_inst_in_s_read;
  assign PEG_Yvec_38_ap_clk = ap_clk;
  assign PEG_Yvec_38__ap_done = PEG_Yvec_38_ap_done;
  assign PEG_Yvec_38__ap_idle = PEG_Yvec_38_ap_idle;
  assign PEG_Yvec_38__ap_ready = PEG_Yvec_38_ap_ready;
  assign PEG_Yvec_38_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_38_ap_start = PEG_Yvec_38__ap_start;
  assign fifo_Y_pe_38__din = PEG_Yvec_38_fifo_Y_out_din;
  assign PEG_Yvec_38_fifo_Y_out_full_n = fifo_Y_pe_38__full_n;
  assign fifo_Y_pe_38__write = PEG_Yvec_38_fifo_Y_out_write;
  assign PEG_Yvec_38_fifo_aXvec_peek_dout = fifo_aXvec_38__dout;
  assign PEG_Yvec_38_fifo_aXvec_peek_empty_n = fifo_aXvec_38__empty_n;
  assign PEG_Yvec_38_fifo_aXvec_s_dout = fifo_aXvec_38__dout;
  assign PEG_Yvec_38_fifo_aXvec_s_empty_n = fifo_aXvec_38__empty_n;
  assign fifo_aXvec_38__read = PEG_Yvec_38_fifo_aXvec_s_read;
  assign PEG_Yvec_38_fifo_inst_in_peek_dout = Yvec_inst_38__dout;
  assign PEG_Yvec_38_fifo_inst_in_peek_empty_n = Yvec_inst_38__empty_n;
  assign PEG_Yvec_38_fifo_inst_in_s_dout = Yvec_inst_38__dout;
  assign PEG_Yvec_38_fifo_inst_in_s_empty_n = Yvec_inst_38__empty_n;
  assign Yvec_inst_38__read = PEG_Yvec_38_fifo_inst_in_s_read;
  assign PEG_Yvec_39_ap_clk = ap_clk;
  assign PEG_Yvec_39__ap_done = PEG_Yvec_39_ap_done;
  assign PEG_Yvec_39__ap_idle = PEG_Yvec_39_ap_idle;
  assign PEG_Yvec_39__ap_ready = PEG_Yvec_39_ap_ready;
  assign PEG_Yvec_39_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_39_ap_start = PEG_Yvec_39__ap_start;
  assign fifo_Y_pe_39__din = PEG_Yvec_39_fifo_Y_out_din;
  assign PEG_Yvec_39_fifo_Y_out_full_n = fifo_Y_pe_39__full_n;
  assign fifo_Y_pe_39__write = PEG_Yvec_39_fifo_Y_out_write;
  assign PEG_Yvec_39_fifo_aXvec_peek_dout = fifo_aXvec_39__dout;
  assign PEG_Yvec_39_fifo_aXvec_peek_empty_n = fifo_aXvec_39__empty_n;
  assign PEG_Yvec_39_fifo_aXvec_s_dout = fifo_aXvec_39__dout;
  assign PEG_Yvec_39_fifo_aXvec_s_empty_n = fifo_aXvec_39__empty_n;
  assign fifo_aXvec_39__read = PEG_Yvec_39_fifo_aXvec_s_read;
  assign PEG_Yvec_39_fifo_inst_in_peek_dout = Yvec_inst_39__dout;
  assign PEG_Yvec_39_fifo_inst_in_peek_empty_n = Yvec_inst_39__empty_n;
  assign PEG_Yvec_39_fifo_inst_in_s_dout = Yvec_inst_39__dout;
  assign PEG_Yvec_39_fifo_inst_in_s_empty_n = Yvec_inst_39__empty_n;
  assign Yvec_inst_39__read = PEG_Yvec_39_fifo_inst_in_s_read;
  assign PEG_Yvec_40_ap_clk = ap_clk;
  assign PEG_Yvec_40__ap_done = PEG_Yvec_40_ap_done;
  assign PEG_Yvec_40__ap_idle = PEG_Yvec_40_ap_idle;
  assign PEG_Yvec_40__ap_ready = PEG_Yvec_40_ap_ready;
  assign PEG_Yvec_40_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_40_ap_start = PEG_Yvec_40__ap_start;
  assign fifo_Y_pe_40__din = PEG_Yvec_40_fifo_Y_out_din;
  assign PEG_Yvec_40_fifo_Y_out_full_n = fifo_Y_pe_40__full_n;
  assign fifo_Y_pe_40__write = PEG_Yvec_40_fifo_Y_out_write;
  assign PEG_Yvec_40_fifo_aXvec_peek_dout = fifo_aXvec_40__dout;
  assign PEG_Yvec_40_fifo_aXvec_peek_empty_n = fifo_aXvec_40__empty_n;
  assign PEG_Yvec_40_fifo_aXvec_s_dout = fifo_aXvec_40__dout;
  assign PEG_Yvec_40_fifo_aXvec_s_empty_n = fifo_aXvec_40__empty_n;
  assign fifo_aXvec_40__read = PEG_Yvec_40_fifo_aXvec_s_read;
  assign PEG_Yvec_40_fifo_inst_in_peek_dout = Yvec_inst_40__dout;
  assign PEG_Yvec_40_fifo_inst_in_peek_empty_n = Yvec_inst_40__empty_n;
  assign PEG_Yvec_40_fifo_inst_in_s_dout = Yvec_inst_40__dout;
  assign PEG_Yvec_40_fifo_inst_in_s_empty_n = Yvec_inst_40__empty_n;
  assign Yvec_inst_40__read = PEG_Yvec_40_fifo_inst_in_s_read;
  assign PEG_Yvec_41_ap_clk = ap_clk;
  assign PEG_Yvec_41__ap_done = PEG_Yvec_41_ap_done;
  assign PEG_Yvec_41__ap_idle = PEG_Yvec_41_ap_idle;
  assign PEG_Yvec_41__ap_ready = PEG_Yvec_41_ap_ready;
  assign PEG_Yvec_41_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_41_ap_start = PEG_Yvec_41__ap_start;
  assign fifo_Y_pe_41__din = PEG_Yvec_41_fifo_Y_out_din;
  assign PEG_Yvec_41_fifo_Y_out_full_n = fifo_Y_pe_41__full_n;
  assign fifo_Y_pe_41__write = PEG_Yvec_41_fifo_Y_out_write;
  assign PEG_Yvec_41_fifo_aXvec_peek_dout = fifo_aXvec_41__dout;
  assign PEG_Yvec_41_fifo_aXvec_peek_empty_n = fifo_aXvec_41__empty_n;
  assign PEG_Yvec_41_fifo_aXvec_s_dout = fifo_aXvec_41__dout;
  assign PEG_Yvec_41_fifo_aXvec_s_empty_n = fifo_aXvec_41__empty_n;
  assign fifo_aXvec_41__read = PEG_Yvec_41_fifo_aXvec_s_read;
  assign PEG_Yvec_41_fifo_inst_in_peek_dout = Yvec_inst_41__dout;
  assign PEG_Yvec_41_fifo_inst_in_peek_empty_n = Yvec_inst_41__empty_n;
  assign PEG_Yvec_41_fifo_inst_in_s_dout = Yvec_inst_41__dout;
  assign PEG_Yvec_41_fifo_inst_in_s_empty_n = Yvec_inst_41__empty_n;
  assign Yvec_inst_41__read = PEG_Yvec_41_fifo_inst_in_s_read;
  assign PEG_Yvec_42_ap_clk = ap_clk;
  assign PEG_Yvec_42__ap_done = PEG_Yvec_42_ap_done;
  assign PEG_Yvec_42__ap_idle = PEG_Yvec_42_ap_idle;
  assign PEG_Yvec_42__ap_ready = PEG_Yvec_42_ap_ready;
  assign PEG_Yvec_42_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_42_ap_start = PEG_Yvec_42__ap_start;
  assign fifo_Y_pe_42__din = PEG_Yvec_42_fifo_Y_out_din;
  assign PEG_Yvec_42_fifo_Y_out_full_n = fifo_Y_pe_42__full_n;
  assign fifo_Y_pe_42__write = PEG_Yvec_42_fifo_Y_out_write;
  assign PEG_Yvec_42_fifo_aXvec_peek_dout = fifo_aXvec_42__dout;
  assign PEG_Yvec_42_fifo_aXvec_peek_empty_n = fifo_aXvec_42__empty_n;
  assign PEG_Yvec_42_fifo_aXvec_s_dout = fifo_aXvec_42__dout;
  assign PEG_Yvec_42_fifo_aXvec_s_empty_n = fifo_aXvec_42__empty_n;
  assign fifo_aXvec_42__read = PEG_Yvec_42_fifo_aXvec_s_read;
  assign PEG_Yvec_42_fifo_inst_in_peek_dout = Yvec_inst_42__dout;
  assign PEG_Yvec_42_fifo_inst_in_peek_empty_n = Yvec_inst_42__empty_n;
  assign PEG_Yvec_42_fifo_inst_in_s_dout = Yvec_inst_42__dout;
  assign PEG_Yvec_42_fifo_inst_in_s_empty_n = Yvec_inst_42__empty_n;
  assign Yvec_inst_42__read = PEG_Yvec_42_fifo_inst_in_s_read;
  assign PEG_Yvec_43_ap_clk = ap_clk;
  assign PEG_Yvec_43__ap_done = PEG_Yvec_43_ap_done;
  assign PEG_Yvec_43__ap_idle = PEG_Yvec_43_ap_idle;
  assign PEG_Yvec_43__ap_ready = PEG_Yvec_43_ap_ready;
  assign PEG_Yvec_43_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_43_ap_start = PEG_Yvec_43__ap_start;
  assign fifo_Y_pe_43__din = PEG_Yvec_43_fifo_Y_out_din;
  assign PEG_Yvec_43_fifo_Y_out_full_n = fifo_Y_pe_43__full_n;
  assign fifo_Y_pe_43__write = PEG_Yvec_43_fifo_Y_out_write;
  assign PEG_Yvec_43_fifo_aXvec_peek_dout = fifo_aXvec_43__dout;
  assign PEG_Yvec_43_fifo_aXvec_peek_empty_n = fifo_aXvec_43__empty_n;
  assign PEG_Yvec_43_fifo_aXvec_s_dout = fifo_aXvec_43__dout;
  assign PEG_Yvec_43_fifo_aXvec_s_empty_n = fifo_aXvec_43__empty_n;
  assign fifo_aXvec_43__read = PEG_Yvec_43_fifo_aXvec_s_read;
  assign PEG_Yvec_43_fifo_inst_in_peek_dout = Yvec_inst_43__dout;
  assign PEG_Yvec_43_fifo_inst_in_peek_empty_n = Yvec_inst_43__empty_n;
  assign PEG_Yvec_43_fifo_inst_in_s_dout = Yvec_inst_43__dout;
  assign PEG_Yvec_43_fifo_inst_in_s_empty_n = Yvec_inst_43__empty_n;
  assign Yvec_inst_43__read = PEG_Yvec_43_fifo_inst_in_s_read;
  assign PEG_Yvec_44_ap_clk = ap_clk;
  assign PEG_Yvec_44__ap_done = PEG_Yvec_44_ap_done;
  assign PEG_Yvec_44__ap_idle = PEG_Yvec_44_ap_idle;
  assign PEG_Yvec_44__ap_ready = PEG_Yvec_44_ap_ready;
  assign PEG_Yvec_44_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_44_ap_start = PEG_Yvec_44__ap_start;
  assign fifo_Y_pe_44__din = PEG_Yvec_44_fifo_Y_out_din;
  assign PEG_Yvec_44_fifo_Y_out_full_n = fifo_Y_pe_44__full_n;
  assign fifo_Y_pe_44__write = PEG_Yvec_44_fifo_Y_out_write;
  assign PEG_Yvec_44_fifo_aXvec_peek_dout = fifo_aXvec_44__dout;
  assign PEG_Yvec_44_fifo_aXvec_peek_empty_n = fifo_aXvec_44__empty_n;
  assign PEG_Yvec_44_fifo_aXvec_s_dout = fifo_aXvec_44__dout;
  assign PEG_Yvec_44_fifo_aXvec_s_empty_n = fifo_aXvec_44__empty_n;
  assign fifo_aXvec_44__read = PEG_Yvec_44_fifo_aXvec_s_read;
  assign PEG_Yvec_44_fifo_inst_in_peek_dout = Yvec_inst_44__dout;
  assign PEG_Yvec_44_fifo_inst_in_peek_empty_n = Yvec_inst_44__empty_n;
  assign PEG_Yvec_44_fifo_inst_in_s_dout = Yvec_inst_44__dout;
  assign PEG_Yvec_44_fifo_inst_in_s_empty_n = Yvec_inst_44__empty_n;
  assign Yvec_inst_44__read = PEG_Yvec_44_fifo_inst_in_s_read;
  assign PEG_Yvec_45_ap_clk = ap_clk;
  assign PEG_Yvec_45__ap_done = PEG_Yvec_45_ap_done;
  assign PEG_Yvec_45__ap_idle = PEG_Yvec_45_ap_idle;
  assign PEG_Yvec_45__ap_ready = PEG_Yvec_45_ap_ready;
  assign PEG_Yvec_45_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_45_ap_start = PEG_Yvec_45__ap_start;
  assign fifo_Y_pe_45__din = PEG_Yvec_45_fifo_Y_out_din;
  assign PEG_Yvec_45_fifo_Y_out_full_n = fifo_Y_pe_45__full_n;
  assign fifo_Y_pe_45__write = PEG_Yvec_45_fifo_Y_out_write;
  assign PEG_Yvec_45_fifo_aXvec_peek_dout = fifo_aXvec_45__dout;
  assign PEG_Yvec_45_fifo_aXvec_peek_empty_n = fifo_aXvec_45__empty_n;
  assign PEG_Yvec_45_fifo_aXvec_s_dout = fifo_aXvec_45__dout;
  assign PEG_Yvec_45_fifo_aXvec_s_empty_n = fifo_aXvec_45__empty_n;
  assign fifo_aXvec_45__read = PEG_Yvec_45_fifo_aXvec_s_read;
  assign PEG_Yvec_45_fifo_inst_in_peek_dout = Yvec_inst_45__dout;
  assign PEG_Yvec_45_fifo_inst_in_peek_empty_n = Yvec_inst_45__empty_n;
  assign PEG_Yvec_45_fifo_inst_in_s_dout = Yvec_inst_45__dout;
  assign PEG_Yvec_45_fifo_inst_in_s_empty_n = Yvec_inst_45__empty_n;
  assign Yvec_inst_45__read = PEG_Yvec_45_fifo_inst_in_s_read;
  assign PEG_Yvec_46_ap_clk = ap_clk;
  assign PEG_Yvec_46__ap_done = PEG_Yvec_46_ap_done;
  assign PEG_Yvec_46__ap_idle = PEG_Yvec_46_ap_idle;
  assign PEG_Yvec_46__ap_ready = PEG_Yvec_46_ap_ready;
  assign PEG_Yvec_46_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_46_ap_start = PEG_Yvec_46__ap_start;
  assign fifo_Y_pe_46__din = PEG_Yvec_46_fifo_Y_out_din;
  assign PEG_Yvec_46_fifo_Y_out_full_n = fifo_Y_pe_46__full_n;
  assign fifo_Y_pe_46__write = PEG_Yvec_46_fifo_Y_out_write;
  assign PEG_Yvec_46_fifo_aXvec_peek_dout = fifo_aXvec_46__dout;
  assign PEG_Yvec_46_fifo_aXvec_peek_empty_n = fifo_aXvec_46__empty_n;
  assign PEG_Yvec_46_fifo_aXvec_s_dout = fifo_aXvec_46__dout;
  assign PEG_Yvec_46_fifo_aXvec_s_empty_n = fifo_aXvec_46__empty_n;
  assign fifo_aXvec_46__read = PEG_Yvec_46_fifo_aXvec_s_read;
  assign PEG_Yvec_46_fifo_inst_in_peek_dout = Yvec_inst_46__dout;
  assign PEG_Yvec_46_fifo_inst_in_peek_empty_n = Yvec_inst_46__empty_n;
  assign PEG_Yvec_46_fifo_inst_in_s_dout = Yvec_inst_46__dout;
  assign PEG_Yvec_46_fifo_inst_in_s_empty_n = Yvec_inst_46__empty_n;
  assign Yvec_inst_46__read = PEG_Yvec_46_fifo_inst_in_s_read;
  assign PEG_Yvec_47_ap_clk = ap_clk;
  assign PEG_Yvec_47__ap_done = PEG_Yvec_47_ap_done;
  assign PEG_Yvec_47__ap_idle = PEG_Yvec_47_ap_idle;
  assign PEG_Yvec_47__ap_ready = PEG_Yvec_47_ap_ready;
  assign PEG_Yvec_47_ap_rst_n = ap_rst_n;
  assign PEG_Yvec_47_ap_start = PEG_Yvec_47__ap_start;
  assign fifo_Y_pe_47__din = PEG_Yvec_47_fifo_Y_out_din;
  assign PEG_Yvec_47_fifo_Y_out_full_n = fifo_Y_pe_47__full_n;
  assign fifo_Y_pe_47__write = PEG_Yvec_47_fifo_Y_out_write;
  assign PEG_Yvec_47_fifo_aXvec_peek_dout = fifo_aXvec_47__dout;
  assign PEG_Yvec_47_fifo_aXvec_peek_empty_n = fifo_aXvec_47__empty_n;
  assign PEG_Yvec_47_fifo_aXvec_s_dout = fifo_aXvec_47__dout;
  assign PEG_Yvec_47_fifo_aXvec_s_empty_n = fifo_aXvec_47__empty_n;
  assign fifo_aXvec_47__read = PEG_Yvec_47_fifo_aXvec_s_read;
  assign PEG_Yvec_47_fifo_inst_in_peek_dout = Yvec_inst_47__dout;
  assign PEG_Yvec_47_fifo_inst_in_peek_empty_n = Yvec_inst_47__empty_n;
  assign PEG_Yvec_47_fifo_inst_in_s_dout = Yvec_inst_47__dout;
  assign PEG_Yvec_47_fifo_inst_in_s_empty_n = Yvec_inst_47__empty_n;
  assign Yvec_inst_47__read = PEG_Yvec_47_fifo_inst_in_s_read;
  assign black_hole_float_v16_0_ap_clk = ap_clk;
  assign black_hole_float_v16_0_ap_rst_n = ap_rst_n;
  assign black_hole_float_v16_0_ap_start = black_hole_float_v16_0__ap_start;
  assign black_hole_float_v16_0_fifo_in_peek_dout = fifo_X_pe_48__dout;
  assign black_hole_float_v16_0_fifo_in_peek_empty_n = fifo_X_pe_48__empty_n;
  assign black_hole_float_v16_0_fifo_in_s_dout = fifo_X_pe_48__dout;
  assign black_hole_float_v16_0_fifo_in_s_empty_n = fifo_X_pe_48__empty_n;
  assign fifo_X_pe_48__read = black_hole_float_v16_0_fifo_in_s_read;
  assign black_hole_int_0_ap_clk = ap_clk;
  assign black_hole_int_0_ap_rst_n = ap_rst_n;
  assign black_hole_int_0_ap_start = black_hole_int_0__ap_start;
  assign black_hole_int_0_fifo_in_peek_dout = PE_inst_48__dout;
  assign black_hole_int_0_fifo_in_peek_empty_n = PE_inst_48__empty_n;
  assign black_hole_int_0_fifo_in_s_dout = PE_inst_48__dout;
  assign black_hole_int_0_fifo_in_s_empty_n = PE_inst_48__empty_n;
  assign PE_inst_48__read = black_hole_int_0_fifo_in_s_read;
  assign read_A_0_A_len = read_A_0___NUM_A_LEN__q0;
  assign read_A_0_A_read_addr_offset = read_A_0___edge_list_ch_0__q0;
  assign edge_list_ch_0_read_addr__din = read_A_0_A_read_addr_s_din;
  assign read_A_0_A_read_addr_s_full_n = edge_list_ch_0_read_addr__full_n;
  assign edge_list_ch_0_read_addr__write = read_A_0_A_read_addr_s_write;
  assign read_A_0_A_read_data_peek_dout = { 1'b0 , edge_list_ch_0_read_data__dout };
  assign read_A_0_A_read_data_peek_empty_n = edge_list_ch_0_read_data__empty_n;
  assign read_A_0_A_read_data_s_dout = { 1'b0 , edge_list_ch_0_read_data__dout };
  assign read_A_0_A_read_data_s_empty_n = edge_list_ch_0_read_data__empty_n;
  assign edge_list_ch_0_read_data__read = read_A_0_A_read_data_s_read;
  assign read_A_0_A_write_addr_offset = read_A_0___edge_list_ch_0__q0;
  assign edge_list_ch_0_write_addr__din = read_A_0_A_write_addr_s_din;
  assign read_A_0_A_write_addr_s_full_n = edge_list_ch_0_write_addr__full_n;
  assign edge_list_ch_0_write_addr__write = read_A_0_A_write_addr_s_write;
  assign edge_list_ch_0_write_data__din = read_A_0_A_write_data_din;
  assign read_A_0_A_write_data_full_n = edge_list_ch_0_write_data__full_n;
  assign edge_list_ch_0_write_data__write = read_A_0_A_write_data_write;
  assign read_A_0_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_0_write_resp__dout };
  assign read_A_0_A_write_resp_peek_empty_n = edge_list_ch_0_write_resp__empty_n;
  assign read_A_0_A_write_resp_s_dout = { 1'b0 , edge_list_ch_0_write_resp__dout };
  assign read_A_0_A_write_resp_s_empty_n = edge_list_ch_0_write_resp__empty_n;
  assign edge_list_ch_0_write_resp__read = read_A_0_A_write_resp_s_read;
  assign read_A_0_P_N = read_A_0___P_N__q0;
  assign read_A_0_ap_clk = ap_clk;
  assign read_A_0__ap_done = read_A_0_ap_done;
  assign read_A_0__ap_idle = read_A_0_ap_idle;
  assign read_A_0__ap_ready = read_A_0_ap_ready;
  assign read_A_0_ap_rst_n = ap_rst_n;
  assign read_A_0_ap_start = read_A_0__ap_start;
  assign fifo_A_0__din = read_A_0_fifo_A_din;
  assign read_A_0_fifo_A_full_n = fifo_A_0__full_n;
  assign fifo_A_0__write = read_A_0_fifo_A_write;
  assign read_A_1_A_len = read_A_1___NUM_A_LEN__q0;
  assign read_A_1_A_read_addr_offset = read_A_1___edge_list_ch_1__q0;
  assign edge_list_ch_1_read_addr__din = read_A_1_A_read_addr_s_din;
  assign read_A_1_A_read_addr_s_full_n = edge_list_ch_1_read_addr__full_n;
  assign edge_list_ch_1_read_addr__write = read_A_1_A_read_addr_s_write;
  assign read_A_1_A_read_data_peek_dout = { 1'b0 , edge_list_ch_1_read_data__dout };
  assign read_A_1_A_read_data_peek_empty_n = edge_list_ch_1_read_data__empty_n;
  assign read_A_1_A_read_data_s_dout = { 1'b0 , edge_list_ch_1_read_data__dout };
  assign read_A_1_A_read_data_s_empty_n = edge_list_ch_1_read_data__empty_n;
  assign edge_list_ch_1_read_data__read = read_A_1_A_read_data_s_read;
  assign read_A_1_A_write_addr_offset = read_A_1___edge_list_ch_1__q0;
  assign edge_list_ch_1_write_addr__din = read_A_1_A_write_addr_s_din;
  assign read_A_1_A_write_addr_s_full_n = edge_list_ch_1_write_addr__full_n;
  assign edge_list_ch_1_write_addr__write = read_A_1_A_write_addr_s_write;
  assign edge_list_ch_1_write_data__din = read_A_1_A_write_data_din;
  assign read_A_1_A_write_data_full_n = edge_list_ch_1_write_data__full_n;
  assign edge_list_ch_1_write_data__write = read_A_1_A_write_data_write;
  assign read_A_1_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_1_write_resp__dout };
  assign read_A_1_A_write_resp_peek_empty_n = edge_list_ch_1_write_resp__empty_n;
  assign read_A_1_A_write_resp_s_dout = { 1'b0 , edge_list_ch_1_write_resp__dout };
  assign read_A_1_A_write_resp_s_empty_n = edge_list_ch_1_write_resp__empty_n;
  assign edge_list_ch_1_write_resp__read = read_A_1_A_write_resp_s_read;
  assign read_A_1_P_N = read_A_1___P_N__q0;
  assign read_A_1_ap_clk = ap_clk;
  assign read_A_1__ap_done = read_A_1_ap_done;
  assign read_A_1__ap_idle = read_A_1_ap_idle;
  assign read_A_1__ap_ready = read_A_1_ap_ready;
  assign read_A_1_ap_rst_n = ap_rst_n;
  assign read_A_1_ap_start = read_A_1__ap_start;
  assign fifo_A_1__din = read_A_1_fifo_A_din;
  assign read_A_1_fifo_A_full_n = fifo_A_1__full_n;
  assign fifo_A_1__write = read_A_1_fifo_A_write;
  assign read_A_2_A_len = read_A_2___NUM_A_LEN__q0;
  assign read_A_2_A_read_addr_offset = read_A_2___edge_list_ch_2__q0;
  assign edge_list_ch_2_read_addr__din = read_A_2_A_read_addr_s_din;
  assign read_A_2_A_read_addr_s_full_n = edge_list_ch_2_read_addr__full_n;
  assign edge_list_ch_2_read_addr__write = read_A_2_A_read_addr_s_write;
  assign read_A_2_A_read_data_peek_dout = { 1'b0 , edge_list_ch_2_read_data__dout };
  assign read_A_2_A_read_data_peek_empty_n = edge_list_ch_2_read_data__empty_n;
  assign read_A_2_A_read_data_s_dout = { 1'b0 , edge_list_ch_2_read_data__dout };
  assign read_A_2_A_read_data_s_empty_n = edge_list_ch_2_read_data__empty_n;
  assign edge_list_ch_2_read_data__read = read_A_2_A_read_data_s_read;
  assign read_A_2_A_write_addr_offset = read_A_2___edge_list_ch_2__q0;
  assign edge_list_ch_2_write_addr__din = read_A_2_A_write_addr_s_din;
  assign read_A_2_A_write_addr_s_full_n = edge_list_ch_2_write_addr__full_n;
  assign edge_list_ch_2_write_addr__write = read_A_2_A_write_addr_s_write;
  assign edge_list_ch_2_write_data__din = read_A_2_A_write_data_din;
  assign read_A_2_A_write_data_full_n = edge_list_ch_2_write_data__full_n;
  assign edge_list_ch_2_write_data__write = read_A_2_A_write_data_write;
  assign read_A_2_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_2_write_resp__dout };
  assign read_A_2_A_write_resp_peek_empty_n = edge_list_ch_2_write_resp__empty_n;
  assign read_A_2_A_write_resp_s_dout = { 1'b0 , edge_list_ch_2_write_resp__dout };
  assign read_A_2_A_write_resp_s_empty_n = edge_list_ch_2_write_resp__empty_n;
  assign edge_list_ch_2_write_resp__read = read_A_2_A_write_resp_s_read;
  assign read_A_2_P_N = read_A_2___P_N__q0;
  assign read_A_2_ap_clk = ap_clk;
  assign read_A_2__ap_done = read_A_2_ap_done;
  assign read_A_2__ap_idle = read_A_2_ap_idle;
  assign read_A_2__ap_ready = read_A_2_ap_ready;
  assign read_A_2_ap_rst_n = ap_rst_n;
  assign read_A_2_ap_start = read_A_2__ap_start;
  assign fifo_A_2__din = read_A_2_fifo_A_din;
  assign read_A_2_fifo_A_full_n = fifo_A_2__full_n;
  assign fifo_A_2__write = read_A_2_fifo_A_write;
  assign read_A_3_A_len = read_A_3___NUM_A_LEN__q0;
  assign read_A_3_A_read_addr_offset = read_A_3___edge_list_ch_3__q0;
  assign edge_list_ch_3_read_addr__din = read_A_3_A_read_addr_s_din;
  assign read_A_3_A_read_addr_s_full_n = edge_list_ch_3_read_addr__full_n;
  assign edge_list_ch_3_read_addr__write = read_A_3_A_read_addr_s_write;
  assign read_A_3_A_read_data_peek_dout = { 1'b0 , edge_list_ch_3_read_data__dout };
  assign read_A_3_A_read_data_peek_empty_n = edge_list_ch_3_read_data__empty_n;
  assign read_A_3_A_read_data_s_dout = { 1'b0 , edge_list_ch_3_read_data__dout };
  assign read_A_3_A_read_data_s_empty_n = edge_list_ch_3_read_data__empty_n;
  assign edge_list_ch_3_read_data__read = read_A_3_A_read_data_s_read;
  assign read_A_3_A_write_addr_offset = read_A_3___edge_list_ch_3__q0;
  assign edge_list_ch_3_write_addr__din = read_A_3_A_write_addr_s_din;
  assign read_A_3_A_write_addr_s_full_n = edge_list_ch_3_write_addr__full_n;
  assign edge_list_ch_3_write_addr__write = read_A_3_A_write_addr_s_write;
  assign edge_list_ch_3_write_data__din = read_A_3_A_write_data_din;
  assign read_A_3_A_write_data_full_n = edge_list_ch_3_write_data__full_n;
  assign edge_list_ch_3_write_data__write = read_A_3_A_write_data_write;
  assign read_A_3_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_3_write_resp__dout };
  assign read_A_3_A_write_resp_peek_empty_n = edge_list_ch_3_write_resp__empty_n;
  assign read_A_3_A_write_resp_s_dout = { 1'b0 , edge_list_ch_3_write_resp__dout };
  assign read_A_3_A_write_resp_s_empty_n = edge_list_ch_3_write_resp__empty_n;
  assign edge_list_ch_3_write_resp__read = read_A_3_A_write_resp_s_read;
  assign read_A_3_P_N = read_A_3___P_N__q0;
  assign read_A_3_ap_clk = ap_clk;
  assign read_A_3__ap_done = read_A_3_ap_done;
  assign read_A_3__ap_idle = read_A_3_ap_idle;
  assign read_A_3__ap_ready = read_A_3_ap_ready;
  assign read_A_3_ap_rst_n = ap_rst_n;
  assign read_A_3_ap_start = read_A_3__ap_start;
  assign fifo_A_3__din = read_A_3_fifo_A_din;
  assign read_A_3_fifo_A_full_n = fifo_A_3__full_n;
  assign fifo_A_3__write = read_A_3_fifo_A_write;
  assign read_A_4_A_len = read_A_4___NUM_A_LEN__q0;
  assign read_A_4_A_read_addr_offset = read_A_4___edge_list_ch_4__q0;
  assign edge_list_ch_4_read_addr__din = read_A_4_A_read_addr_s_din;
  assign read_A_4_A_read_addr_s_full_n = edge_list_ch_4_read_addr__full_n;
  assign edge_list_ch_4_read_addr__write = read_A_4_A_read_addr_s_write;
  assign read_A_4_A_read_data_peek_dout = { 1'b0 , edge_list_ch_4_read_data__dout };
  assign read_A_4_A_read_data_peek_empty_n = edge_list_ch_4_read_data__empty_n;
  assign read_A_4_A_read_data_s_dout = { 1'b0 , edge_list_ch_4_read_data__dout };
  assign read_A_4_A_read_data_s_empty_n = edge_list_ch_4_read_data__empty_n;
  assign edge_list_ch_4_read_data__read = read_A_4_A_read_data_s_read;
  assign read_A_4_A_write_addr_offset = read_A_4___edge_list_ch_4__q0;
  assign edge_list_ch_4_write_addr__din = read_A_4_A_write_addr_s_din;
  assign read_A_4_A_write_addr_s_full_n = edge_list_ch_4_write_addr__full_n;
  assign edge_list_ch_4_write_addr__write = read_A_4_A_write_addr_s_write;
  assign edge_list_ch_4_write_data__din = read_A_4_A_write_data_din;
  assign read_A_4_A_write_data_full_n = edge_list_ch_4_write_data__full_n;
  assign edge_list_ch_4_write_data__write = read_A_4_A_write_data_write;
  assign read_A_4_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_4_write_resp__dout };
  assign read_A_4_A_write_resp_peek_empty_n = edge_list_ch_4_write_resp__empty_n;
  assign read_A_4_A_write_resp_s_dout = { 1'b0 , edge_list_ch_4_write_resp__dout };
  assign read_A_4_A_write_resp_s_empty_n = edge_list_ch_4_write_resp__empty_n;
  assign edge_list_ch_4_write_resp__read = read_A_4_A_write_resp_s_read;
  assign read_A_4_P_N = read_A_4___P_N__q0;
  assign read_A_4_ap_clk = ap_clk;
  assign read_A_4__ap_done = read_A_4_ap_done;
  assign read_A_4__ap_idle = read_A_4_ap_idle;
  assign read_A_4__ap_ready = read_A_4_ap_ready;
  assign read_A_4_ap_rst_n = ap_rst_n;
  assign read_A_4_ap_start = read_A_4__ap_start;
  assign fifo_A_4__din = read_A_4_fifo_A_din;
  assign read_A_4_fifo_A_full_n = fifo_A_4__full_n;
  assign fifo_A_4__write = read_A_4_fifo_A_write;
  assign read_A_5_A_len = read_A_5___NUM_A_LEN__q0;
  assign read_A_5_A_read_addr_offset = read_A_5___edge_list_ch_5__q0;
  assign edge_list_ch_5_read_addr__din = read_A_5_A_read_addr_s_din;
  assign read_A_5_A_read_addr_s_full_n = edge_list_ch_5_read_addr__full_n;
  assign edge_list_ch_5_read_addr__write = read_A_5_A_read_addr_s_write;
  assign read_A_5_A_read_data_peek_dout = { 1'b0 , edge_list_ch_5_read_data__dout };
  assign read_A_5_A_read_data_peek_empty_n = edge_list_ch_5_read_data__empty_n;
  assign read_A_5_A_read_data_s_dout = { 1'b0 , edge_list_ch_5_read_data__dout };
  assign read_A_5_A_read_data_s_empty_n = edge_list_ch_5_read_data__empty_n;
  assign edge_list_ch_5_read_data__read = read_A_5_A_read_data_s_read;
  assign read_A_5_A_write_addr_offset = read_A_5___edge_list_ch_5__q0;
  assign edge_list_ch_5_write_addr__din = read_A_5_A_write_addr_s_din;
  assign read_A_5_A_write_addr_s_full_n = edge_list_ch_5_write_addr__full_n;
  assign edge_list_ch_5_write_addr__write = read_A_5_A_write_addr_s_write;
  assign edge_list_ch_5_write_data__din = read_A_5_A_write_data_din;
  assign read_A_5_A_write_data_full_n = edge_list_ch_5_write_data__full_n;
  assign edge_list_ch_5_write_data__write = read_A_5_A_write_data_write;
  assign read_A_5_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_5_write_resp__dout };
  assign read_A_5_A_write_resp_peek_empty_n = edge_list_ch_5_write_resp__empty_n;
  assign read_A_5_A_write_resp_s_dout = { 1'b0 , edge_list_ch_5_write_resp__dout };
  assign read_A_5_A_write_resp_s_empty_n = edge_list_ch_5_write_resp__empty_n;
  assign edge_list_ch_5_write_resp__read = read_A_5_A_write_resp_s_read;
  assign read_A_5_P_N = read_A_5___P_N__q0;
  assign read_A_5_ap_clk = ap_clk;
  assign read_A_5__ap_done = read_A_5_ap_done;
  assign read_A_5__ap_idle = read_A_5_ap_idle;
  assign read_A_5__ap_ready = read_A_5_ap_ready;
  assign read_A_5_ap_rst_n = ap_rst_n;
  assign read_A_5_ap_start = read_A_5__ap_start;
  assign fifo_A_5__din = read_A_5_fifo_A_din;
  assign read_A_5_fifo_A_full_n = fifo_A_5__full_n;
  assign fifo_A_5__write = read_A_5_fifo_A_write;
  assign read_A_6_A_len = read_A_6___NUM_A_LEN__q0;
  assign read_A_6_A_read_addr_offset = read_A_6___edge_list_ch_6__q0;
  assign edge_list_ch_6_read_addr__din = read_A_6_A_read_addr_s_din;
  assign read_A_6_A_read_addr_s_full_n = edge_list_ch_6_read_addr__full_n;
  assign edge_list_ch_6_read_addr__write = read_A_6_A_read_addr_s_write;
  assign read_A_6_A_read_data_peek_dout = { 1'b0 , edge_list_ch_6_read_data__dout };
  assign read_A_6_A_read_data_peek_empty_n = edge_list_ch_6_read_data__empty_n;
  assign read_A_6_A_read_data_s_dout = { 1'b0 , edge_list_ch_6_read_data__dout };
  assign read_A_6_A_read_data_s_empty_n = edge_list_ch_6_read_data__empty_n;
  assign edge_list_ch_6_read_data__read = read_A_6_A_read_data_s_read;
  assign read_A_6_A_write_addr_offset = read_A_6___edge_list_ch_6__q0;
  assign edge_list_ch_6_write_addr__din = read_A_6_A_write_addr_s_din;
  assign read_A_6_A_write_addr_s_full_n = edge_list_ch_6_write_addr__full_n;
  assign edge_list_ch_6_write_addr__write = read_A_6_A_write_addr_s_write;
  assign edge_list_ch_6_write_data__din = read_A_6_A_write_data_din;
  assign read_A_6_A_write_data_full_n = edge_list_ch_6_write_data__full_n;
  assign edge_list_ch_6_write_data__write = read_A_6_A_write_data_write;
  assign read_A_6_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_6_write_resp__dout };
  assign read_A_6_A_write_resp_peek_empty_n = edge_list_ch_6_write_resp__empty_n;
  assign read_A_6_A_write_resp_s_dout = { 1'b0 , edge_list_ch_6_write_resp__dout };
  assign read_A_6_A_write_resp_s_empty_n = edge_list_ch_6_write_resp__empty_n;
  assign edge_list_ch_6_write_resp__read = read_A_6_A_write_resp_s_read;
  assign read_A_6_P_N = read_A_6___P_N__q0;
  assign read_A_6_ap_clk = ap_clk;
  assign read_A_6__ap_done = read_A_6_ap_done;
  assign read_A_6__ap_idle = read_A_6_ap_idle;
  assign read_A_6__ap_ready = read_A_6_ap_ready;
  assign read_A_6_ap_rst_n = ap_rst_n;
  assign read_A_6_ap_start = read_A_6__ap_start;
  assign fifo_A_6__din = read_A_6_fifo_A_din;
  assign read_A_6_fifo_A_full_n = fifo_A_6__full_n;
  assign fifo_A_6__write = read_A_6_fifo_A_write;
  assign read_A_7_A_len = read_A_7___NUM_A_LEN__q0;
  assign read_A_7_A_read_addr_offset = read_A_7___edge_list_ch_7__q0;
  assign edge_list_ch_7_read_addr__din = read_A_7_A_read_addr_s_din;
  assign read_A_7_A_read_addr_s_full_n = edge_list_ch_7_read_addr__full_n;
  assign edge_list_ch_7_read_addr__write = read_A_7_A_read_addr_s_write;
  assign read_A_7_A_read_data_peek_dout = { 1'b0 , edge_list_ch_7_read_data__dout };
  assign read_A_7_A_read_data_peek_empty_n = edge_list_ch_7_read_data__empty_n;
  assign read_A_7_A_read_data_s_dout = { 1'b0 , edge_list_ch_7_read_data__dout };
  assign read_A_7_A_read_data_s_empty_n = edge_list_ch_7_read_data__empty_n;
  assign edge_list_ch_7_read_data__read = read_A_7_A_read_data_s_read;
  assign read_A_7_A_write_addr_offset = read_A_7___edge_list_ch_7__q0;
  assign edge_list_ch_7_write_addr__din = read_A_7_A_write_addr_s_din;
  assign read_A_7_A_write_addr_s_full_n = edge_list_ch_7_write_addr__full_n;
  assign edge_list_ch_7_write_addr__write = read_A_7_A_write_addr_s_write;
  assign edge_list_ch_7_write_data__din = read_A_7_A_write_data_din;
  assign read_A_7_A_write_data_full_n = edge_list_ch_7_write_data__full_n;
  assign edge_list_ch_7_write_data__write = read_A_7_A_write_data_write;
  assign read_A_7_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_7_write_resp__dout };
  assign read_A_7_A_write_resp_peek_empty_n = edge_list_ch_7_write_resp__empty_n;
  assign read_A_7_A_write_resp_s_dout = { 1'b0 , edge_list_ch_7_write_resp__dout };
  assign read_A_7_A_write_resp_s_empty_n = edge_list_ch_7_write_resp__empty_n;
  assign edge_list_ch_7_write_resp__read = read_A_7_A_write_resp_s_read;
  assign read_A_7_P_N = read_A_7___P_N__q0;
  assign read_A_7_ap_clk = ap_clk;
  assign read_A_7__ap_done = read_A_7_ap_done;
  assign read_A_7__ap_idle = read_A_7_ap_idle;
  assign read_A_7__ap_ready = read_A_7_ap_ready;
  assign read_A_7_ap_rst_n = ap_rst_n;
  assign read_A_7_ap_start = read_A_7__ap_start;
  assign fifo_A_7__din = read_A_7_fifo_A_din;
  assign read_A_7_fifo_A_full_n = fifo_A_7__full_n;
  assign fifo_A_7__write = read_A_7_fifo_A_write;
  assign read_A_8_A_len = read_A_8___NUM_A_LEN__q0;
  assign read_A_8_A_read_addr_offset = read_A_8___edge_list_ch_8__q0;
  assign edge_list_ch_8_read_addr__din = read_A_8_A_read_addr_s_din;
  assign read_A_8_A_read_addr_s_full_n = edge_list_ch_8_read_addr__full_n;
  assign edge_list_ch_8_read_addr__write = read_A_8_A_read_addr_s_write;
  assign read_A_8_A_read_data_peek_dout = { 1'b0 , edge_list_ch_8_read_data__dout };
  assign read_A_8_A_read_data_peek_empty_n = edge_list_ch_8_read_data__empty_n;
  assign read_A_8_A_read_data_s_dout = { 1'b0 , edge_list_ch_8_read_data__dout };
  assign read_A_8_A_read_data_s_empty_n = edge_list_ch_8_read_data__empty_n;
  assign edge_list_ch_8_read_data__read = read_A_8_A_read_data_s_read;
  assign read_A_8_A_write_addr_offset = read_A_8___edge_list_ch_8__q0;
  assign edge_list_ch_8_write_addr__din = read_A_8_A_write_addr_s_din;
  assign read_A_8_A_write_addr_s_full_n = edge_list_ch_8_write_addr__full_n;
  assign edge_list_ch_8_write_addr__write = read_A_8_A_write_addr_s_write;
  assign edge_list_ch_8_write_data__din = read_A_8_A_write_data_din;
  assign read_A_8_A_write_data_full_n = edge_list_ch_8_write_data__full_n;
  assign edge_list_ch_8_write_data__write = read_A_8_A_write_data_write;
  assign read_A_8_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_8_write_resp__dout };
  assign read_A_8_A_write_resp_peek_empty_n = edge_list_ch_8_write_resp__empty_n;
  assign read_A_8_A_write_resp_s_dout = { 1'b0 , edge_list_ch_8_write_resp__dout };
  assign read_A_8_A_write_resp_s_empty_n = edge_list_ch_8_write_resp__empty_n;
  assign edge_list_ch_8_write_resp__read = read_A_8_A_write_resp_s_read;
  assign read_A_8_P_N = read_A_8___P_N__q0;
  assign read_A_8_ap_clk = ap_clk;
  assign read_A_8__ap_done = read_A_8_ap_done;
  assign read_A_8__ap_idle = read_A_8_ap_idle;
  assign read_A_8__ap_ready = read_A_8_ap_ready;
  assign read_A_8_ap_rst_n = ap_rst_n;
  assign read_A_8_ap_start = read_A_8__ap_start;
  assign fifo_A_8__din = read_A_8_fifo_A_din;
  assign read_A_8_fifo_A_full_n = fifo_A_8__full_n;
  assign fifo_A_8__write = read_A_8_fifo_A_write;
  assign read_A_9_A_len = read_A_9___NUM_A_LEN__q0;
  assign read_A_9_A_read_addr_offset = read_A_9___edge_list_ch_9__q0;
  assign edge_list_ch_9_read_addr__din = read_A_9_A_read_addr_s_din;
  assign read_A_9_A_read_addr_s_full_n = edge_list_ch_9_read_addr__full_n;
  assign edge_list_ch_9_read_addr__write = read_A_9_A_read_addr_s_write;
  assign read_A_9_A_read_data_peek_dout = { 1'b0 , edge_list_ch_9_read_data__dout };
  assign read_A_9_A_read_data_peek_empty_n = edge_list_ch_9_read_data__empty_n;
  assign read_A_9_A_read_data_s_dout = { 1'b0 , edge_list_ch_9_read_data__dout };
  assign read_A_9_A_read_data_s_empty_n = edge_list_ch_9_read_data__empty_n;
  assign edge_list_ch_9_read_data__read = read_A_9_A_read_data_s_read;
  assign read_A_9_A_write_addr_offset = read_A_9___edge_list_ch_9__q0;
  assign edge_list_ch_9_write_addr__din = read_A_9_A_write_addr_s_din;
  assign read_A_9_A_write_addr_s_full_n = edge_list_ch_9_write_addr__full_n;
  assign edge_list_ch_9_write_addr__write = read_A_9_A_write_addr_s_write;
  assign edge_list_ch_9_write_data__din = read_A_9_A_write_data_din;
  assign read_A_9_A_write_data_full_n = edge_list_ch_9_write_data__full_n;
  assign edge_list_ch_9_write_data__write = read_A_9_A_write_data_write;
  assign read_A_9_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_9_write_resp__dout };
  assign read_A_9_A_write_resp_peek_empty_n = edge_list_ch_9_write_resp__empty_n;
  assign read_A_9_A_write_resp_s_dout = { 1'b0 , edge_list_ch_9_write_resp__dout };
  assign read_A_9_A_write_resp_s_empty_n = edge_list_ch_9_write_resp__empty_n;
  assign edge_list_ch_9_write_resp__read = read_A_9_A_write_resp_s_read;
  assign read_A_9_P_N = read_A_9___P_N__q0;
  assign read_A_9_ap_clk = ap_clk;
  assign read_A_9__ap_done = read_A_9_ap_done;
  assign read_A_9__ap_idle = read_A_9_ap_idle;
  assign read_A_9__ap_ready = read_A_9_ap_ready;
  assign read_A_9_ap_rst_n = ap_rst_n;
  assign read_A_9_ap_start = read_A_9__ap_start;
  assign fifo_A_9__din = read_A_9_fifo_A_din;
  assign read_A_9_fifo_A_full_n = fifo_A_9__full_n;
  assign fifo_A_9__write = read_A_9_fifo_A_write;
  assign read_A_10_A_len = read_A_10___NUM_A_LEN__q0;
  assign read_A_10_A_read_addr_offset = read_A_10___edge_list_ch_10__q0;
  assign edge_list_ch_10_read_addr__din = read_A_10_A_read_addr_s_din;
  assign read_A_10_A_read_addr_s_full_n = edge_list_ch_10_read_addr__full_n;
  assign edge_list_ch_10_read_addr__write = read_A_10_A_read_addr_s_write;
  assign read_A_10_A_read_data_peek_dout = { 1'b0 , edge_list_ch_10_read_data__dout };
  assign read_A_10_A_read_data_peek_empty_n = edge_list_ch_10_read_data__empty_n;
  assign read_A_10_A_read_data_s_dout = { 1'b0 , edge_list_ch_10_read_data__dout };
  assign read_A_10_A_read_data_s_empty_n = edge_list_ch_10_read_data__empty_n;
  assign edge_list_ch_10_read_data__read = read_A_10_A_read_data_s_read;
  assign read_A_10_A_write_addr_offset = read_A_10___edge_list_ch_10__q0;
  assign edge_list_ch_10_write_addr__din = read_A_10_A_write_addr_s_din;
  assign read_A_10_A_write_addr_s_full_n = edge_list_ch_10_write_addr__full_n;
  assign edge_list_ch_10_write_addr__write = read_A_10_A_write_addr_s_write;
  assign edge_list_ch_10_write_data__din = read_A_10_A_write_data_din;
  assign read_A_10_A_write_data_full_n = edge_list_ch_10_write_data__full_n;
  assign edge_list_ch_10_write_data__write = read_A_10_A_write_data_write;
  assign read_A_10_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_10_write_resp__dout };
  assign read_A_10_A_write_resp_peek_empty_n = edge_list_ch_10_write_resp__empty_n;
  assign read_A_10_A_write_resp_s_dout = { 1'b0 , edge_list_ch_10_write_resp__dout };
  assign read_A_10_A_write_resp_s_empty_n = edge_list_ch_10_write_resp__empty_n;
  assign edge_list_ch_10_write_resp__read = read_A_10_A_write_resp_s_read;
  assign read_A_10_P_N = read_A_10___P_N__q0;
  assign read_A_10_ap_clk = ap_clk;
  assign read_A_10__ap_done = read_A_10_ap_done;
  assign read_A_10__ap_idle = read_A_10_ap_idle;
  assign read_A_10__ap_ready = read_A_10_ap_ready;
  assign read_A_10_ap_rst_n = ap_rst_n;
  assign read_A_10_ap_start = read_A_10__ap_start;
  assign fifo_A_10__din = read_A_10_fifo_A_din;
  assign read_A_10_fifo_A_full_n = fifo_A_10__full_n;
  assign fifo_A_10__write = read_A_10_fifo_A_write;
  assign read_A_11_A_len = read_A_11___NUM_A_LEN__q0;
  assign read_A_11_A_read_addr_offset = read_A_11___edge_list_ch_11__q0;
  assign edge_list_ch_11_read_addr__din = read_A_11_A_read_addr_s_din;
  assign read_A_11_A_read_addr_s_full_n = edge_list_ch_11_read_addr__full_n;
  assign edge_list_ch_11_read_addr__write = read_A_11_A_read_addr_s_write;
  assign read_A_11_A_read_data_peek_dout = { 1'b0 , edge_list_ch_11_read_data__dout };
  assign read_A_11_A_read_data_peek_empty_n = edge_list_ch_11_read_data__empty_n;
  assign read_A_11_A_read_data_s_dout = { 1'b0 , edge_list_ch_11_read_data__dout };
  assign read_A_11_A_read_data_s_empty_n = edge_list_ch_11_read_data__empty_n;
  assign edge_list_ch_11_read_data__read = read_A_11_A_read_data_s_read;
  assign read_A_11_A_write_addr_offset = read_A_11___edge_list_ch_11__q0;
  assign edge_list_ch_11_write_addr__din = read_A_11_A_write_addr_s_din;
  assign read_A_11_A_write_addr_s_full_n = edge_list_ch_11_write_addr__full_n;
  assign edge_list_ch_11_write_addr__write = read_A_11_A_write_addr_s_write;
  assign edge_list_ch_11_write_data__din = read_A_11_A_write_data_din;
  assign read_A_11_A_write_data_full_n = edge_list_ch_11_write_data__full_n;
  assign edge_list_ch_11_write_data__write = read_A_11_A_write_data_write;
  assign read_A_11_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_11_write_resp__dout };
  assign read_A_11_A_write_resp_peek_empty_n = edge_list_ch_11_write_resp__empty_n;
  assign read_A_11_A_write_resp_s_dout = { 1'b0 , edge_list_ch_11_write_resp__dout };
  assign read_A_11_A_write_resp_s_empty_n = edge_list_ch_11_write_resp__empty_n;
  assign edge_list_ch_11_write_resp__read = read_A_11_A_write_resp_s_read;
  assign read_A_11_P_N = read_A_11___P_N__q0;
  assign read_A_11_ap_clk = ap_clk;
  assign read_A_11__ap_done = read_A_11_ap_done;
  assign read_A_11__ap_idle = read_A_11_ap_idle;
  assign read_A_11__ap_ready = read_A_11_ap_ready;
  assign read_A_11_ap_rst_n = ap_rst_n;
  assign read_A_11_ap_start = read_A_11__ap_start;
  assign fifo_A_11__din = read_A_11_fifo_A_din;
  assign read_A_11_fifo_A_full_n = fifo_A_11__full_n;
  assign fifo_A_11__write = read_A_11_fifo_A_write;
  assign read_A_12_A_len = read_A_12___NUM_A_LEN__q0;
  assign read_A_12_A_read_addr_offset = read_A_12___edge_list_ch_12__q0;
  assign edge_list_ch_12_read_addr__din = read_A_12_A_read_addr_s_din;
  assign read_A_12_A_read_addr_s_full_n = edge_list_ch_12_read_addr__full_n;
  assign edge_list_ch_12_read_addr__write = read_A_12_A_read_addr_s_write;
  assign read_A_12_A_read_data_peek_dout = { 1'b0 , edge_list_ch_12_read_data__dout };
  assign read_A_12_A_read_data_peek_empty_n = edge_list_ch_12_read_data__empty_n;
  assign read_A_12_A_read_data_s_dout = { 1'b0 , edge_list_ch_12_read_data__dout };
  assign read_A_12_A_read_data_s_empty_n = edge_list_ch_12_read_data__empty_n;
  assign edge_list_ch_12_read_data__read = read_A_12_A_read_data_s_read;
  assign read_A_12_A_write_addr_offset = read_A_12___edge_list_ch_12__q0;
  assign edge_list_ch_12_write_addr__din = read_A_12_A_write_addr_s_din;
  assign read_A_12_A_write_addr_s_full_n = edge_list_ch_12_write_addr__full_n;
  assign edge_list_ch_12_write_addr__write = read_A_12_A_write_addr_s_write;
  assign edge_list_ch_12_write_data__din = read_A_12_A_write_data_din;
  assign read_A_12_A_write_data_full_n = edge_list_ch_12_write_data__full_n;
  assign edge_list_ch_12_write_data__write = read_A_12_A_write_data_write;
  assign read_A_12_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_12_write_resp__dout };
  assign read_A_12_A_write_resp_peek_empty_n = edge_list_ch_12_write_resp__empty_n;
  assign read_A_12_A_write_resp_s_dout = { 1'b0 , edge_list_ch_12_write_resp__dout };
  assign read_A_12_A_write_resp_s_empty_n = edge_list_ch_12_write_resp__empty_n;
  assign edge_list_ch_12_write_resp__read = read_A_12_A_write_resp_s_read;
  assign read_A_12_P_N = read_A_12___P_N__q0;
  assign read_A_12_ap_clk = ap_clk;
  assign read_A_12__ap_done = read_A_12_ap_done;
  assign read_A_12__ap_idle = read_A_12_ap_idle;
  assign read_A_12__ap_ready = read_A_12_ap_ready;
  assign read_A_12_ap_rst_n = ap_rst_n;
  assign read_A_12_ap_start = read_A_12__ap_start;
  assign fifo_A_12__din = read_A_12_fifo_A_din;
  assign read_A_12_fifo_A_full_n = fifo_A_12__full_n;
  assign fifo_A_12__write = read_A_12_fifo_A_write;
  assign read_A_13_A_len = read_A_13___NUM_A_LEN__q0;
  assign read_A_13_A_read_addr_offset = read_A_13___edge_list_ch_13__q0;
  assign edge_list_ch_13_read_addr__din = read_A_13_A_read_addr_s_din;
  assign read_A_13_A_read_addr_s_full_n = edge_list_ch_13_read_addr__full_n;
  assign edge_list_ch_13_read_addr__write = read_A_13_A_read_addr_s_write;
  assign read_A_13_A_read_data_peek_dout = { 1'b0 , edge_list_ch_13_read_data__dout };
  assign read_A_13_A_read_data_peek_empty_n = edge_list_ch_13_read_data__empty_n;
  assign read_A_13_A_read_data_s_dout = { 1'b0 , edge_list_ch_13_read_data__dout };
  assign read_A_13_A_read_data_s_empty_n = edge_list_ch_13_read_data__empty_n;
  assign edge_list_ch_13_read_data__read = read_A_13_A_read_data_s_read;
  assign read_A_13_A_write_addr_offset = read_A_13___edge_list_ch_13__q0;
  assign edge_list_ch_13_write_addr__din = read_A_13_A_write_addr_s_din;
  assign read_A_13_A_write_addr_s_full_n = edge_list_ch_13_write_addr__full_n;
  assign edge_list_ch_13_write_addr__write = read_A_13_A_write_addr_s_write;
  assign edge_list_ch_13_write_data__din = read_A_13_A_write_data_din;
  assign read_A_13_A_write_data_full_n = edge_list_ch_13_write_data__full_n;
  assign edge_list_ch_13_write_data__write = read_A_13_A_write_data_write;
  assign read_A_13_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_13_write_resp__dout };
  assign read_A_13_A_write_resp_peek_empty_n = edge_list_ch_13_write_resp__empty_n;
  assign read_A_13_A_write_resp_s_dout = { 1'b0 , edge_list_ch_13_write_resp__dout };
  assign read_A_13_A_write_resp_s_empty_n = edge_list_ch_13_write_resp__empty_n;
  assign edge_list_ch_13_write_resp__read = read_A_13_A_write_resp_s_read;
  assign read_A_13_P_N = read_A_13___P_N__q0;
  assign read_A_13_ap_clk = ap_clk;
  assign read_A_13__ap_done = read_A_13_ap_done;
  assign read_A_13__ap_idle = read_A_13_ap_idle;
  assign read_A_13__ap_ready = read_A_13_ap_ready;
  assign read_A_13_ap_rst_n = ap_rst_n;
  assign read_A_13_ap_start = read_A_13__ap_start;
  assign fifo_A_13__din = read_A_13_fifo_A_din;
  assign read_A_13_fifo_A_full_n = fifo_A_13__full_n;
  assign fifo_A_13__write = read_A_13_fifo_A_write;
  assign read_A_14_A_len = read_A_14___NUM_A_LEN__q0;
  assign read_A_14_A_read_addr_offset = read_A_14___edge_list_ch_14__q0;
  assign edge_list_ch_14_read_addr__din = read_A_14_A_read_addr_s_din;
  assign read_A_14_A_read_addr_s_full_n = edge_list_ch_14_read_addr__full_n;
  assign edge_list_ch_14_read_addr__write = read_A_14_A_read_addr_s_write;
  assign read_A_14_A_read_data_peek_dout = { 1'b0 , edge_list_ch_14_read_data__dout };
  assign read_A_14_A_read_data_peek_empty_n = edge_list_ch_14_read_data__empty_n;
  assign read_A_14_A_read_data_s_dout = { 1'b0 , edge_list_ch_14_read_data__dout };
  assign read_A_14_A_read_data_s_empty_n = edge_list_ch_14_read_data__empty_n;
  assign edge_list_ch_14_read_data__read = read_A_14_A_read_data_s_read;
  assign read_A_14_A_write_addr_offset = read_A_14___edge_list_ch_14__q0;
  assign edge_list_ch_14_write_addr__din = read_A_14_A_write_addr_s_din;
  assign read_A_14_A_write_addr_s_full_n = edge_list_ch_14_write_addr__full_n;
  assign edge_list_ch_14_write_addr__write = read_A_14_A_write_addr_s_write;
  assign edge_list_ch_14_write_data__din = read_A_14_A_write_data_din;
  assign read_A_14_A_write_data_full_n = edge_list_ch_14_write_data__full_n;
  assign edge_list_ch_14_write_data__write = read_A_14_A_write_data_write;
  assign read_A_14_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_14_write_resp__dout };
  assign read_A_14_A_write_resp_peek_empty_n = edge_list_ch_14_write_resp__empty_n;
  assign read_A_14_A_write_resp_s_dout = { 1'b0 , edge_list_ch_14_write_resp__dout };
  assign read_A_14_A_write_resp_s_empty_n = edge_list_ch_14_write_resp__empty_n;
  assign edge_list_ch_14_write_resp__read = read_A_14_A_write_resp_s_read;
  assign read_A_14_P_N = read_A_14___P_N__q0;
  assign read_A_14_ap_clk = ap_clk;
  assign read_A_14__ap_done = read_A_14_ap_done;
  assign read_A_14__ap_idle = read_A_14_ap_idle;
  assign read_A_14__ap_ready = read_A_14_ap_ready;
  assign read_A_14_ap_rst_n = ap_rst_n;
  assign read_A_14_ap_start = read_A_14__ap_start;
  assign fifo_A_14__din = read_A_14_fifo_A_din;
  assign read_A_14_fifo_A_full_n = fifo_A_14__full_n;
  assign fifo_A_14__write = read_A_14_fifo_A_write;
  assign read_A_15_A_len = read_A_15___NUM_A_LEN__q0;
  assign read_A_15_A_read_addr_offset = read_A_15___edge_list_ch_15__q0;
  assign edge_list_ch_15_read_addr__din = read_A_15_A_read_addr_s_din;
  assign read_A_15_A_read_addr_s_full_n = edge_list_ch_15_read_addr__full_n;
  assign edge_list_ch_15_read_addr__write = read_A_15_A_read_addr_s_write;
  assign read_A_15_A_read_data_peek_dout = { 1'b0 , edge_list_ch_15_read_data__dout };
  assign read_A_15_A_read_data_peek_empty_n = edge_list_ch_15_read_data__empty_n;
  assign read_A_15_A_read_data_s_dout = { 1'b0 , edge_list_ch_15_read_data__dout };
  assign read_A_15_A_read_data_s_empty_n = edge_list_ch_15_read_data__empty_n;
  assign edge_list_ch_15_read_data__read = read_A_15_A_read_data_s_read;
  assign read_A_15_A_write_addr_offset = read_A_15___edge_list_ch_15__q0;
  assign edge_list_ch_15_write_addr__din = read_A_15_A_write_addr_s_din;
  assign read_A_15_A_write_addr_s_full_n = edge_list_ch_15_write_addr__full_n;
  assign edge_list_ch_15_write_addr__write = read_A_15_A_write_addr_s_write;
  assign edge_list_ch_15_write_data__din = read_A_15_A_write_data_din;
  assign read_A_15_A_write_data_full_n = edge_list_ch_15_write_data__full_n;
  assign edge_list_ch_15_write_data__write = read_A_15_A_write_data_write;
  assign read_A_15_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_15_write_resp__dout };
  assign read_A_15_A_write_resp_peek_empty_n = edge_list_ch_15_write_resp__empty_n;
  assign read_A_15_A_write_resp_s_dout = { 1'b0 , edge_list_ch_15_write_resp__dout };
  assign read_A_15_A_write_resp_s_empty_n = edge_list_ch_15_write_resp__empty_n;
  assign edge_list_ch_15_write_resp__read = read_A_15_A_write_resp_s_read;
  assign read_A_15_P_N = read_A_15___P_N__q0;
  assign read_A_15_ap_clk = ap_clk;
  assign read_A_15__ap_done = read_A_15_ap_done;
  assign read_A_15__ap_idle = read_A_15_ap_idle;
  assign read_A_15__ap_ready = read_A_15_ap_ready;
  assign read_A_15_ap_rst_n = ap_rst_n;
  assign read_A_15_ap_start = read_A_15__ap_start;
  assign fifo_A_15__din = read_A_15_fifo_A_din;
  assign read_A_15_fifo_A_full_n = fifo_A_15__full_n;
  assign fifo_A_15__write = read_A_15_fifo_A_write;
  assign read_A_16_A_len = read_A_16___NUM_A_LEN__q0;
  assign read_A_16_A_read_addr_offset = read_A_16___edge_list_ch_16__q0;
  assign edge_list_ch_16_read_addr__din = read_A_16_A_read_addr_s_din;
  assign read_A_16_A_read_addr_s_full_n = edge_list_ch_16_read_addr__full_n;
  assign edge_list_ch_16_read_addr__write = read_A_16_A_read_addr_s_write;
  assign read_A_16_A_read_data_peek_dout = { 1'b0 , edge_list_ch_16_read_data__dout };
  assign read_A_16_A_read_data_peek_empty_n = edge_list_ch_16_read_data__empty_n;
  assign read_A_16_A_read_data_s_dout = { 1'b0 , edge_list_ch_16_read_data__dout };
  assign read_A_16_A_read_data_s_empty_n = edge_list_ch_16_read_data__empty_n;
  assign edge_list_ch_16_read_data__read = read_A_16_A_read_data_s_read;
  assign read_A_16_A_write_addr_offset = read_A_16___edge_list_ch_16__q0;
  assign edge_list_ch_16_write_addr__din = read_A_16_A_write_addr_s_din;
  assign read_A_16_A_write_addr_s_full_n = edge_list_ch_16_write_addr__full_n;
  assign edge_list_ch_16_write_addr__write = read_A_16_A_write_addr_s_write;
  assign edge_list_ch_16_write_data__din = read_A_16_A_write_data_din;
  assign read_A_16_A_write_data_full_n = edge_list_ch_16_write_data__full_n;
  assign edge_list_ch_16_write_data__write = read_A_16_A_write_data_write;
  assign read_A_16_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_16_write_resp__dout };
  assign read_A_16_A_write_resp_peek_empty_n = edge_list_ch_16_write_resp__empty_n;
  assign read_A_16_A_write_resp_s_dout = { 1'b0 , edge_list_ch_16_write_resp__dout };
  assign read_A_16_A_write_resp_s_empty_n = edge_list_ch_16_write_resp__empty_n;
  assign edge_list_ch_16_write_resp__read = read_A_16_A_write_resp_s_read;
  assign read_A_16_P_N = read_A_16___P_N__q0;
  assign read_A_16_ap_clk = ap_clk;
  assign read_A_16__ap_done = read_A_16_ap_done;
  assign read_A_16__ap_idle = read_A_16_ap_idle;
  assign read_A_16__ap_ready = read_A_16_ap_ready;
  assign read_A_16_ap_rst_n = ap_rst_n;
  assign read_A_16_ap_start = read_A_16__ap_start;
  assign fifo_A_16__din = read_A_16_fifo_A_din;
  assign read_A_16_fifo_A_full_n = fifo_A_16__full_n;
  assign fifo_A_16__write = read_A_16_fifo_A_write;
  assign read_A_17_A_len = read_A_17___NUM_A_LEN__q0;
  assign read_A_17_A_read_addr_offset = read_A_17___edge_list_ch_17__q0;
  assign edge_list_ch_17_read_addr__din = read_A_17_A_read_addr_s_din;
  assign read_A_17_A_read_addr_s_full_n = edge_list_ch_17_read_addr__full_n;
  assign edge_list_ch_17_read_addr__write = read_A_17_A_read_addr_s_write;
  assign read_A_17_A_read_data_peek_dout = { 1'b0 , edge_list_ch_17_read_data__dout };
  assign read_A_17_A_read_data_peek_empty_n = edge_list_ch_17_read_data__empty_n;
  assign read_A_17_A_read_data_s_dout = { 1'b0 , edge_list_ch_17_read_data__dout };
  assign read_A_17_A_read_data_s_empty_n = edge_list_ch_17_read_data__empty_n;
  assign edge_list_ch_17_read_data__read = read_A_17_A_read_data_s_read;
  assign read_A_17_A_write_addr_offset = read_A_17___edge_list_ch_17__q0;
  assign edge_list_ch_17_write_addr__din = read_A_17_A_write_addr_s_din;
  assign read_A_17_A_write_addr_s_full_n = edge_list_ch_17_write_addr__full_n;
  assign edge_list_ch_17_write_addr__write = read_A_17_A_write_addr_s_write;
  assign edge_list_ch_17_write_data__din = read_A_17_A_write_data_din;
  assign read_A_17_A_write_data_full_n = edge_list_ch_17_write_data__full_n;
  assign edge_list_ch_17_write_data__write = read_A_17_A_write_data_write;
  assign read_A_17_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_17_write_resp__dout };
  assign read_A_17_A_write_resp_peek_empty_n = edge_list_ch_17_write_resp__empty_n;
  assign read_A_17_A_write_resp_s_dout = { 1'b0 , edge_list_ch_17_write_resp__dout };
  assign read_A_17_A_write_resp_s_empty_n = edge_list_ch_17_write_resp__empty_n;
  assign edge_list_ch_17_write_resp__read = read_A_17_A_write_resp_s_read;
  assign read_A_17_P_N = read_A_17___P_N__q0;
  assign read_A_17_ap_clk = ap_clk;
  assign read_A_17__ap_done = read_A_17_ap_done;
  assign read_A_17__ap_idle = read_A_17_ap_idle;
  assign read_A_17__ap_ready = read_A_17_ap_ready;
  assign read_A_17_ap_rst_n = ap_rst_n;
  assign read_A_17_ap_start = read_A_17__ap_start;
  assign fifo_A_17__din = read_A_17_fifo_A_din;
  assign read_A_17_fifo_A_full_n = fifo_A_17__full_n;
  assign fifo_A_17__write = read_A_17_fifo_A_write;
  assign read_A_18_A_len = read_A_18___NUM_A_LEN__q0;
  assign read_A_18_A_read_addr_offset = read_A_18___edge_list_ch_18__q0;
  assign edge_list_ch_18_read_addr__din = read_A_18_A_read_addr_s_din;
  assign read_A_18_A_read_addr_s_full_n = edge_list_ch_18_read_addr__full_n;
  assign edge_list_ch_18_read_addr__write = read_A_18_A_read_addr_s_write;
  assign read_A_18_A_read_data_peek_dout = { 1'b0 , edge_list_ch_18_read_data__dout };
  assign read_A_18_A_read_data_peek_empty_n = edge_list_ch_18_read_data__empty_n;
  assign read_A_18_A_read_data_s_dout = { 1'b0 , edge_list_ch_18_read_data__dout };
  assign read_A_18_A_read_data_s_empty_n = edge_list_ch_18_read_data__empty_n;
  assign edge_list_ch_18_read_data__read = read_A_18_A_read_data_s_read;
  assign read_A_18_A_write_addr_offset = read_A_18___edge_list_ch_18__q0;
  assign edge_list_ch_18_write_addr__din = read_A_18_A_write_addr_s_din;
  assign read_A_18_A_write_addr_s_full_n = edge_list_ch_18_write_addr__full_n;
  assign edge_list_ch_18_write_addr__write = read_A_18_A_write_addr_s_write;
  assign edge_list_ch_18_write_data__din = read_A_18_A_write_data_din;
  assign read_A_18_A_write_data_full_n = edge_list_ch_18_write_data__full_n;
  assign edge_list_ch_18_write_data__write = read_A_18_A_write_data_write;
  assign read_A_18_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_18_write_resp__dout };
  assign read_A_18_A_write_resp_peek_empty_n = edge_list_ch_18_write_resp__empty_n;
  assign read_A_18_A_write_resp_s_dout = { 1'b0 , edge_list_ch_18_write_resp__dout };
  assign read_A_18_A_write_resp_s_empty_n = edge_list_ch_18_write_resp__empty_n;
  assign edge_list_ch_18_write_resp__read = read_A_18_A_write_resp_s_read;
  assign read_A_18_P_N = read_A_18___P_N__q0;
  assign read_A_18_ap_clk = ap_clk;
  assign read_A_18__ap_done = read_A_18_ap_done;
  assign read_A_18__ap_idle = read_A_18_ap_idle;
  assign read_A_18__ap_ready = read_A_18_ap_ready;
  assign read_A_18_ap_rst_n = ap_rst_n;
  assign read_A_18_ap_start = read_A_18__ap_start;
  assign fifo_A_18__din = read_A_18_fifo_A_din;
  assign read_A_18_fifo_A_full_n = fifo_A_18__full_n;
  assign fifo_A_18__write = read_A_18_fifo_A_write;
  assign read_A_19_A_len = read_A_19___NUM_A_LEN__q0;
  assign read_A_19_A_read_addr_offset = read_A_19___edge_list_ch_19__q0;
  assign edge_list_ch_19_read_addr__din = read_A_19_A_read_addr_s_din;
  assign read_A_19_A_read_addr_s_full_n = edge_list_ch_19_read_addr__full_n;
  assign edge_list_ch_19_read_addr__write = read_A_19_A_read_addr_s_write;
  assign read_A_19_A_read_data_peek_dout = { 1'b0 , edge_list_ch_19_read_data__dout };
  assign read_A_19_A_read_data_peek_empty_n = edge_list_ch_19_read_data__empty_n;
  assign read_A_19_A_read_data_s_dout = { 1'b0 , edge_list_ch_19_read_data__dout };
  assign read_A_19_A_read_data_s_empty_n = edge_list_ch_19_read_data__empty_n;
  assign edge_list_ch_19_read_data__read = read_A_19_A_read_data_s_read;
  assign read_A_19_A_write_addr_offset = read_A_19___edge_list_ch_19__q0;
  assign edge_list_ch_19_write_addr__din = read_A_19_A_write_addr_s_din;
  assign read_A_19_A_write_addr_s_full_n = edge_list_ch_19_write_addr__full_n;
  assign edge_list_ch_19_write_addr__write = read_A_19_A_write_addr_s_write;
  assign edge_list_ch_19_write_data__din = read_A_19_A_write_data_din;
  assign read_A_19_A_write_data_full_n = edge_list_ch_19_write_data__full_n;
  assign edge_list_ch_19_write_data__write = read_A_19_A_write_data_write;
  assign read_A_19_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_19_write_resp__dout };
  assign read_A_19_A_write_resp_peek_empty_n = edge_list_ch_19_write_resp__empty_n;
  assign read_A_19_A_write_resp_s_dout = { 1'b0 , edge_list_ch_19_write_resp__dout };
  assign read_A_19_A_write_resp_s_empty_n = edge_list_ch_19_write_resp__empty_n;
  assign edge_list_ch_19_write_resp__read = read_A_19_A_write_resp_s_read;
  assign read_A_19_P_N = read_A_19___P_N__q0;
  assign read_A_19_ap_clk = ap_clk;
  assign read_A_19__ap_done = read_A_19_ap_done;
  assign read_A_19__ap_idle = read_A_19_ap_idle;
  assign read_A_19__ap_ready = read_A_19_ap_ready;
  assign read_A_19_ap_rst_n = ap_rst_n;
  assign read_A_19_ap_start = read_A_19__ap_start;
  assign fifo_A_19__din = read_A_19_fifo_A_din;
  assign read_A_19_fifo_A_full_n = fifo_A_19__full_n;
  assign fifo_A_19__write = read_A_19_fifo_A_write;
  assign read_A_20_A_len = read_A_20___NUM_A_LEN__q0;
  assign read_A_20_A_read_addr_offset = read_A_20___edge_list_ch_20__q0;
  assign edge_list_ch_20_read_addr__din = read_A_20_A_read_addr_s_din;
  assign read_A_20_A_read_addr_s_full_n = edge_list_ch_20_read_addr__full_n;
  assign edge_list_ch_20_read_addr__write = read_A_20_A_read_addr_s_write;
  assign read_A_20_A_read_data_peek_dout = { 1'b0 , edge_list_ch_20_read_data__dout };
  assign read_A_20_A_read_data_peek_empty_n = edge_list_ch_20_read_data__empty_n;
  assign read_A_20_A_read_data_s_dout = { 1'b0 , edge_list_ch_20_read_data__dout };
  assign read_A_20_A_read_data_s_empty_n = edge_list_ch_20_read_data__empty_n;
  assign edge_list_ch_20_read_data__read = read_A_20_A_read_data_s_read;
  assign read_A_20_A_write_addr_offset = read_A_20___edge_list_ch_20__q0;
  assign edge_list_ch_20_write_addr__din = read_A_20_A_write_addr_s_din;
  assign read_A_20_A_write_addr_s_full_n = edge_list_ch_20_write_addr__full_n;
  assign edge_list_ch_20_write_addr__write = read_A_20_A_write_addr_s_write;
  assign edge_list_ch_20_write_data__din = read_A_20_A_write_data_din;
  assign read_A_20_A_write_data_full_n = edge_list_ch_20_write_data__full_n;
  assign edge_list_ch_20_write_data__write = read_A_20_A_write_data_write;
  assign read_A_20_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_20_write_resp__dout };
  assign read_A_20_A_write_resp_peek_empty_n = edge_list_ch_20_write_resp__empty_n;
  assign read_A_20_A_write_resp_s_dout = { 1'b0 , edge_list_ch_20_write_resp__dout };
  assign read_A_20_A_write_resp_s_empty_n = edge_list_ch_20_write_resp__empty_n;
  assign edge_list_ch_20_write_resp__read = read_A_20_A_write_resp_s_read;
  assign read_A_20_P_N = read_A_20___P_N__q0;
  assign read_A_20_ap_clk = ap_clk;
  assign read_A_20__ap_done = read_A_20_ap_done;
  assign read_A_20__ap_idle = read_A_20_ap_idle;
  assign read_A_20__ap_ready = read_A_20_ap_ready;
  assign read_A_20_ap_rst_n = ap_rst_n;
  assign read_A_20_ap_start = read_A_20__ap_start;
  assign fifo_A_20__din = read_A_20_fifo_A_din;
  assign read_A_20_fifo_A_full_n = fifo_A_20__full_n;
  assign fifo_A_20__write = read_A_20_fifo_A_write;
  assign read_A_21_A_len = read_A_21___NUM_A_LEN__q0;
  assign read_A_21_A_read_addr_offset = read_A_21___edge_list_ch_21__q0;
  assign edge_list_ch_21_read_addr__din = read_A_21_A_read_addr_s_din;
  assign read_A_21_A_read_addr_s_full_n = edge_list_ch_21_read_addr__full_n;
  assign edge_list_ch_21_read_addr__write = read_A_21_A_read_addr_s_write;
  assign read_A_21_A_read_data_peek_dout = { 1'b0 , edge_list_ch_21_read_data__dout };
  assign read_A_21_A_read_data_peek_empty_n = edge_list_ch_21_read_data__empty_n;
  assign read_A_21_A_read_data_s_dout = { 1'b0 , edge_list_ch_21_read_data__dout };
  assign read_A_21_A_read_data_s_empty_n = edge_list_ch_21_read_data__empty_n;
  assign edge_list_ch_21_read_data__read = read_A_21_A_read_data_s_read;
  assign read_A_21_A_write_addr_offset = read_A_21___edge_list_ch_21__q0;
  assign edge_list_ch_21_write_addr__din = read_A_21_A_write_addr_s_din;
  assign read_A_21_A_write_addr_s_full_n = edge_list_ch_21_write_addr__full_n;
  assign edge_list_ch_21_write_addr__write = read_A_21_A_write_addr_s_write;
  assign edge_list_ch_21_write_data__din = read_A_21_A_write_data_din;
  assign read_A_21_A_write_data_full_n = edge_list_ch_21_write_data__full_n;
  assign edge_list_ch_21_write_data__write = read_A_21_A_write_data_write;
  assign read_A_21_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_21_write_resp__dout };
  assign read_A_21_A_write_resp_peek_empty_n = edge_list_ch_21_write_resp__empty_n;
  assign read_A_21_A_write_resp_s_dout = { 1'b0 , edge_list_ch_21_write_resp__dout };
  assign read_A_21_A_write_resp_s_empty_n = edge_list_ch_21_write_resp__empty_n;
  assign edge_list_ch_21_write_resp__read = read_A_21_A_write_resp_s_read;
  assign read_A_21_P_N = read_A_21___P_N__q0;
  assign read_A_21_ap_clk = ap_clk;
  assign read_A_21__ap_done = read_A_21_ap_done;
  assign read_A_21__ap_idle = read_A_21_ap_idle;
  assign read_A_21__ap_ready = read_A_21_ap_ready;
  assign read_A_21_ap_rst_n = ap_rst_n;
  assign read_A_21_ap_start = read_A_21__ap_start;
  assign fifo_A_21__din = read_A_21_fifo_A_din;
  assign read_A_21_fifo_A_full_n = fifo_A_21__full_n;
  assign fifo_A_21__write = read_A_21_fifo_A_write;
  assign read_A_22_A_len = read_A_22___NUM_A_LEN__q0;
  assign read_A_22_A_read_addr_offset = read_A_22___edge_list_ch_22__q0;
  assign edge_list_ch_22_read_addr__din = read_A_22_A_read_addr_s_din;
  assign read_A_22_A_read_addr_s_full_n = edge_list_ch_22_read_addr__full_n;
  assign edge_list_ch_22_read_addr__write = read_A_22_A_read_addr_s_write;
  assign read_A_22_A_read_data_peek_dout = { 1'b0 , edge_list_ch_22_read_data__dout };
  assign read_A_22_A_read_data_peek_empty_n = edge_list_ch_22_read_data__empty_n;
  assign read_A_22_A_read_data_s_dout = { 1'b0 , edge_list_ch_22_read_data__dout };
  assign read_A_22_A_read_data_s_empty_n = edge_list_ch_22_read_data__empty_n;
  assign edge_list_ch_22_read_data__read = read_A_22_A_read_data_s_read;
  assign read_A_22_A_write_addr_offset = read_A_22___edge_list_ch_22__q0;
  assign edge_list_ch_22_write_addr__din = read_A_22_A_write_addr_s_din;
  assign read_A_22_A_write_addr_s_full_n = edge_list_ch_22_write_addr__full_n;
  assign edge_list_ch_22_write_addr__write = read_A_22_A_write_addr_s_write;
  assign edge_list_ch_22_write_data__din = read_A_22_A_write_data_din;
  assign read_A_22_A_write_data_full_n = edge_list_ch_22_write_data__full_n;
  assign edge_list_ch_22_write_data__write = read_A_22_A_write_data_write;
  assign read_A_22_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_22_write_resp__dout };
  assign read_A_22_A_write_resp_peek_empty_n = edge_list_ch_22_write_resp__empty_n;
  assign read_A_22_A_write_resp_s_dout = { 1'b0 , edge_list_ch_22_write_resp__dout };
  assign read_A_22_A_write_resp_s_empty_n = edge_list_ch_22_write_resp__empty_n;
  assign edge_list_ch_22_write_resp__read = read_A_22_A_write_resp_s_read;
  assign read_A_22_P_N = read_A_22___P_N__q0;
  assign read_A_22_ap_clk = ap_clk;
  assign read_A_22__ap_done = read_A_22_ap_done;
  assign read_A_22__ap_idle = read_A_22_ap_idle;
  assign read_A_22__ap_ready = read_A_22_ap_ready;
  assign read_A_22_ap_rst_n = ap_rst_n;
  assign read_A_22_ap_start = read_A_22__ap_start;
  assign fifo_A_22__din = read_A_22_fifo_A_din;
  assign read_A_22_fifo_A_full_n = fifo_A_22__full_n;
  assign fifo_A_22__write = read_A_22_fifo_A_write;
  assign read_A_23_A_len = read_A_23___NUM_A_LEN__q0;
  assign read_A_23_A_read_addr_offset = read_A_23___edge_list_ch_23__q0;
  assign edge_list_ch_23_read_addr__din = read_A_23_A_read_addr_s_din;
  assign read_A_23_A_read_addr_s_full_n = edge_list_ch_23_read_addr__full_n;
  assign edge_list_ch_23_read_addr__write = read_A_23_A_read_addr_s_write;
  assign read_A_23_A_read_data_peek_dout = { 1'b0 , edge_list_ch_23_read_data__dout };
  assign read_A_23_A_read_data_peek_empty_n = edge_list_ch_23_read_data__empty_n;
  assign read_A_23_A_read_data_s_dout = { 1'b0 , edge_list_ch_23_read_data__dout };
  assign read_A_23_A_read_data_s_empty_n = edge_list_ch_23_read_data__empty_n;
  assign edge_list_ch_23_read_data__read = read_A_23_A_read_data_s_read;
  assign read_A_23_A_write_addr_offset = read_A_23___edge_list_ch_23__q0;
  assign edge_list_ch_23_write_addr__din = read_A_23_A_write_addr_s_din;
  assign read_A_23_A_write_addr_s_full_n = edge_list_ch_23_write_addr__full_n;
  assign edge_list_ch_23_write_addr__write = read_A_23_A_write_addr_s_write;
  assign edge_list_ch_23_write_data__din = read_A_23_A_write_data_din;
  assign read_A_23_A_write_data_full_n = edge_list_ch_23_write_data__full_n;
  assign edge_list_ch_23_write_data__write = read_A_23_A_write_data_write;
  assign read_A_23_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_23_write_resp__dout };
  assign read_A_23_A_write_resp_peek_empty_n = edge_list_ch_23_write_resp__empty_n;
  assign read_A_23_A_write_resp_s_dout = { 1'b0 , edge_list_ch_23_write_resp__dout };
  assign read_A_23_A_write_resp_s_empty_n = edge_list_ch_23_write_resp__empty_n;
  assign edge_list_ch_23_write_resp__read = read_A_23_A_write_resp_s_read;
  assign read_A_23_P_N = read_A_23___P_N__q0;
  assign read_A_23_ap_clk = ap_clk;
  assign read_A_23__ap_done = read_A_23_ap_done;
  assign read_A_23__ap_idle = read_A_23_ap_idle;
  assign read_A_23__ap_ready = read_A_23_ap_ready;
  assign read_A_23_ap_rst_n = ap_rst_n;
  assign read_A_23_ap_start = read_A_23__ap_start;
  assign fifo_A_23__din = read_A_23_fifo_A_din;
  assign read_A_23_fifo_A_full_n = fifo_A_23__full_n;
  assign fifo_A_23__write = read_A_23_fifo_A_write;
  assign read_A_24_A_len = read_A_24___NUM_A_LEN__q0;
  assign read_A_24_A_read_addr_offset = read_A_24___edge_list_ch_24__q0;
  assign edge_list_ch_24_read_addr__din = read_A_24_A_read_addr_s_din;
  assign read_A_24_A_read_addr_s_full_n = edge_list_ch_24_read_addr__full_n;
  assign edge_list_ch_24_read_addr__write = read_A_24_A_read_addr_s_write;
  assign read_A_24_A_read_data_peek_dout = { 1'b0 , edge_list_ch_24_read_data__dout };
  assign read_A_24_A_read_data_peek_empty_n = edge_list_ch_24_read_data__empty_n;
  assign read_A_24_A_read_data_s_dout = { 1'b0 , edge_list_ch_24_read_data__dout };
  assign read_A_24_A_read_data_s_empty_n = edge_list_ch_24_read_data__empty_n;
  assign edge_list_ch_24_read_data__read = read_A_24_A_read_data_s_read;
  assign read_A_24_A_write_addr_offset = read_A_24___edge_list_ch_24__q0;
  assign edge_list_ch_24_write_addr__din = read_A_24_A_write_addr_s_din;
  assign read_A_24_A_write_addr_s_full_n = edge_list_ch_24_write_addr__full_n;
  assign edge_list_ch_24_write_addr__write = read_A_24_A_write_addr_s_write;
  assign edge_list_ch_24_write_data__din = read_A_24_A_write_data_din;
  assign read_A_24_A_write_data_full_n = edge_list_ch_24_write_data__full_n;
  assign edge_list_ch_24_write_data__write = read_A_24_A_write_data_write;
  assign read_A_24_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_24_write_resp__dout };
  assign read_A_24_A_write_resp_peek_empty_n = edge_list_ch_24_write_resp__empty_n;
  assign read_A_24_A_write_resp_s_dout = { 1'b0 , edge_list_ch_24_write_resp__dout };
  assign read_A_24_A_write_resp_s_empty_n = edge_list_ch_24_write_resp__empty_n;
  assign edge_list_ch_24_write_resp__read = read_A_24_A_write_resp_s_read;
  assign read_A_24_P_N = read_A_24___P_N__q0;
  assign read_A_24_ap_clk = ap_clk;
  assign read_A_24__ap_done = read_A_24_ap_done;
  assign read_A_24__ap_idle = read_A_24_ap_idle;
  assign read_A_24__ap_ready = read_A_24_ap_ready;
  assign read_A_24_ap_rst_n = ap_rst_n;
  assign read_A_24_ap_start = read_A_24__ap_start;
  assign fifo_A_24__din = read_A_24_fifo_A_din;
  assign read_A_24_fifo_A_full_n = fifo_A_24__full_n;
  assign fifo_A_24__write = read_A_24_fifo_A_write;
  assign read_A_25_A_len = read_A_25___NUM_A_LEN__q0;
  assign read_A_25_A_read_addr_offset = read_A_25___edge_list_ch_25__q0;
  assign edge_list_ch_25_read_addr__din = read_A_25_A_read_addr_s_din;
  assign read_A_25_A_read_addr_s_full_n = edge_list_ch_25_read_addr__full_n;
  assign edge_list_ch_25_read_addr__write = read_A_25_A_read_addr_s_write;
  assign read_A_25_A_read_data_peek_dout = { 1'b0 , edge_list_ch_25_read_data__dout };
  assign read_A_25_A_read_data_peek_empty_n = edge_list_ch_25_read_data__empty_n;
  assign read_A_25_A_read_data_s_dout = { 1'b0 , edge_list_ch_25_read_data__dout };
  assign read_A_25_A_read_data_s_empty_n = edge_list_ch_25_read_data__empty_n;
  assign edge_list_ch_25_read_data__read = read_A_25_A_read_data_s_read;
  assign read_A_25_A_write_addr_offset = read_A_25___edge_list_ch_25__q0;
  assign edge_list_ch_25_write_addr__din = read_A_25_A_write_addr_s_din;
  assign read_A_25_A_write_addr_s_full_n = edge_list_ch_25_write_addr__full_n;
  assign edge_list_ch_25_write_addr__write = read_A_25_A_write_addr_s_write;
  assign edge_list_ch_25_write_data__din = read_A_25_A_write_data_din;
  assign read_A_25_A_write_data_full_n = edge_list_ch_25_write_data__full_n;
  assign edge_list_ch_25_write_data__write = read_A_25_A_write_data_write;
  assign read_A_25_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_25_write_resp__dout };
  assign read_A_25_A_write_resp_peek_empty_n = edge_list_ch_25_write_resp__empty_n;
  assign read_A_25_A_write_resp_s_dout = { 1'b0 , edge_list_ch_25_write_resp__dout };
  assign read_A_25_A_write_resp_s_empty_n = edge_list_ch_25_write_resp__empty_n;
  assign edge_list_ch_25_write_resp__read = read_A_25_A_write_resp_s_read;
  assign read_A_25_P_N = read_A_25___P_N__q0;
  assign read_A_25_ap_clk = ap_clk;
  assign read_A_25__ap_done = read_A_25_ap_done;
  assign read_A_25__ap_idle = read_A_25_ap_idle;
  assign read_A_25__ap_ready = read_A_25_ap_ready;
  assign read_A_25_ap_rst_n = ap_rst_n;
  assign read_A_25_ap_start = read_A_25__ap_start;
  assign fifo_A_25__din = read_A_25_fifo_A_din;
  assign read_A_25_fifo_A_full_n = fifo_A_25__full_n;
  assign fifo_A_25__write = read_A_25_fifo_A_write;
  assign read_A_26_A_len = read_A_26___NUM_A_LEN__q0;
  assign read_A_26_A_read_addr_offset = read_A_26___edge_list_ch_26__q0;
  assign edge_list_ch_26_read_addr__din = read_A_26_A_read_addr_s_din;
  assign read_A_26_A_read_addr_s_full_n = edge_list_ch_26_read_addr__full_n;
  assign edge_list_ch_26_read_addr__write = read_A_26_A_read_addr_s_write;
  assign read_A_26_A_read_data_peek_dout = { 1'b0 , edge_list_ch_26_read_data__dout };
  assign read_A_26_A_read_data_peek_empty_n = edge_list_ch_26_read_data__empty_n;
  assign read_A_26_A_read_data_s_dout = { 1'b0 , edge_list_ch_26_read_data__dout };
  assign read_A_26_A_read_data_s_empty_n = edge_list_ch_26_read_data__empty_n;
  assign edge_list_ch_26_read_data__read = read_A_26_A_read_data_s_read;
  assign read_A_26_A_write_addr_offset = read_A_26___edge_list_ch_26__q0;
  assign edge_list_ch_26_write_addr__din = read_A_26_A_write_addr_s_din;
  assign read_A_26_A_write_addr_s_full_n = edge_list_ch_26_write_addr__full_n;
  assign edge_list_ch_26_write_addr__write = read_A_26_A_write_addr_s_write;
  assign edge_list_ch_26_write_data__din = read_A_26_A_write_data_din;
  assign read_A_26_A_write_data_full_n = edge_list_ch_26_write_data__full_n;
  assign edge_list_ch_26_write_data__write = read_A_26_A_write_data_write;
  assign read_A_26_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_26_write_resp__dout };
  assign read_A_26_A_write_resp_peek_empty_n = edge_list_ch_26_write_resp__empty_n;
  assign read_A_26_A_write_resp_s_dout = { 1'b0 , edge_list_ch_26_write_resp__dout };
  assign read_A_26_A_write_resp_s_empty_n = edge_list_ch_26_write_resp__empty_n;
  assign edge_list_ch_26_write_resp__read = read_A_26_A_write_resp_s_read;
  assign read_A_26_P_N = read_A_26___P_N__q0;
  assign read_A_26_ap_clk = ap_clk;
  assign read_A_26__ap_done = read_A_26_ap_done;
  assign read_A_26__ap_idle = read_A_26_ap_idle;
  assign read_A_26__ap_ready = read_A_26_ap_ready;
  assign read_A_26_ap_rst_n = ap_rst_n;
  assign read_A_26_ap_start = read_A_26__ap_start;
  assign fifo_A_26__din = read_A_26_fifo_A_din;
  assign read_A_26_fifo_A_full_n = fifo_A_26__full_n;
  assign fifo_A_26__write = read_A_26_fifo_A_write;
  assign read_A_27_A_len = read_A_27___NUM_A_LEN__q0;
  assign read_A_27_A_read_addr_offset = read_A_27___edge_list_ch_27__q0;
  assign edge_list_ch_27_read_addr__din = read_A_27_A_read_addr_s_din;
  assign read_A_27_A_read_addr_s_full_n = edge_list_ch_27_read_addr__full_n;
  assign edge_list_ch_27_read_addr__write = read_A_27_A_read_addr_s_write;
  assign read_A_27_A_read_data_peek_dout = { 1'b0 , edge_list_ch_27_read_data__dout };
  assign read_A_27_A_read_data_peek_empty_n = edge_list_ch_27_read_data__empty_n;
  assign read_A_27_A_read_data_s_dout = { 1'b0 , edge_list_ch_27_read_data__dout };
  assign read_A_27_A_read_data_s_empty_n = edge_list_ch_27_read_data__empty_n;
  assign edge_list_ch_27_read_data__read = read_A_27_A_read_data_s_read;
  assign read_A_27_A_write_addr_offset = read_A_27___edge_list_ch_27__q0;
  assign edge_list_ch_27_write_addr__din = read_A_27_A_write_addr_s_din;
  assign read_A_27_A_write_addr_s_full_n = edge_list_ch_27_write_addr__full_n;
  assign edge_list_ch_27_write_addr__write = read_A_27_A_write_addr_s_write;
  assign edge_list_ch_27_write_data__din = read_A_27_A_write_data_din;
  assign read_A_27_A_write_data_full_n = edge_list_ch_27_write_data__full_n;
  assign edge_list_ch_27_write_data__write = read_A_27_A_write_data_write;
  assign read_A_27_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_27_write_resp__dout };
  assign read_A_27_A_write_resp_peek_empty_n = edge_list_ch_27_write_resp__empty_n;
  assign read_A_27_A_write_resp_s_dout = { 1'b0 , edge_list_ch_27_write_resp__dout };
  assign read_A_27_A_write_resp_s_empty_n = edge_list_ch_27_write_resp__empty_n;
  assign edge_list_ch_27_write_resp__read = read_A_27_A_write_resp_s_read;
  assign read_A_27_P_N = read_A_27___P_N__q0;
  assign read_A_27_ap_clk = ap_clk;
  assign read_A_27__ap_done = read_A_27_ap_done;
  assign read_A_27__ap_idle = read_A_27_ap_idle;
  assign read_A_27__ap_ready = read_A_27_ap_ready;
  assign read_A_27_ap_rst_n = ap_rst_n;
  assign read_A_27_ap_start = read_A_27__ap_start;
  assign fifo_A_27__din = read_A_27_fifo_A_din;
  assign read_A_27_fifo_A_full_n = fifo_A_27__full_n;
  assign fifo_A_27__write = read_A_27_fifo_A_write;
  assign read_A_28_A_len = read_A_28___NUM_A_LEN__q0;
  assign read_A_28_A_read_addr_offset = read_A_28___edge_list_ch_28__q0;
  assign edge_list_ch_28_read_addr__din = read_A_28_A_read_addr_s_din;
  assign read_A_28_A_read_addr_s_full_n = edge_list_ch_28_read_addr__full_n;
  assign edge_list_ch_28_read_addr__write = read_A_28_A_read_addr_s_write;
  assign read_A_28_A_read_data_peek_dout = { 1'b0 , edge_list_ch_28_read_data__dout };
  assign read_A_28_A_read_data_peek_empty_n = edge_list_ch_28_read_data__empty_n;
  assign read_A_28_A_read_data_s_dout = { 1'b0 , edge_list_ch_28_read_data__dout };
  assign read_A_28_A_read_data_s_empty_n = edge_list_ch_28_read_data__empty_n;
  assign edge_list_ch_28_read_data__read = read_A_28_A_read_data_s_read;
  assign read_A_28_A_write_addr_offset = read_A_28___edge_list_ch_28__q0;
  assign edge_list_ch_28_write_addr__din = read_A_28_A_write_addr_s_din;
  assign read_A_28_A_write_addr_s_full_n = edge_list_ch_28_write_addr__full_n;
  assign edge_list_ch_28_write_addr__write = read_A_28_A_write_addr_s_write;
  assign edge_list_ch_28_write_data__din = read_A_28_A_write_data_din;
  assign read_A_28_A_write_data_full_n = edge_list_ch_28_write_data__full_n;
  assign edge_list_ch_28_write_data__write = read_A_28_A_write_data_write;
  assign read_A_28_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_28_write_resp__dout };
  assign read_A_28_A_write_resp_peek_empty_n = edge_list_ch_28_write_resp__empty_n;
  assign read_A_28_A_write_resp_s_dout = { 1'b0 , edge_list_ch_28_write_resp__dout };
  assign read_A_28_A_write_resp_s_empty_n = edge_list_ch_28_write_resp__empty_n;
  assign edge_list_ch_28_write_resp__read = read_A_28_A_write_resp_s_read;
  assign read_A_28_P_N = read_A_28___P_N__q0;
  assign read_A_28_ap_clk = ap_clk;
  assign read_A_28__ap_done = read_A_28_ap_done;
  assign read_A_28__ap_idle = read_A_28_ap_idle;
  assign read_A_28__ap_ready = read_A_28_ap_ready;
  assign read_A_28_ap_rst_n = ap_rst_n;
  assign read_A_28_ap_start = read_A_28__ap_start;
  assign fifo_A_28__din = read_A_28_fifo_A_din;
  assign read_A_28_fifo_A_full_n = fifo_A_28__full_n;
  assign fifo_A_28__write = read_A_28_fifo_A_write;
  assign read_A_29_A_len = read_A_29___NUM_A_LEN__q0;
  assign read_A_29_A_read_addr_offset = read_A_29___edge_list_ch_29__q0;
  assign edge_list_ch_29_read_addr__din = read_A_29_A_read_addr_s_din;
  assign read_A_29_A_read_addr_s_full_n = edge_list_ch_29_read_addr__full_n;
  assign edge_list_ch_29_read_addr__write = read_A_29_A_read_addr_s_write;
  assign read_A_29_A_read_data_peek_dout = { 1'b0 , edge_list_ch_29_read_data__dout };
  assign read_A_29_A_read_data_peek_empty_n = edge_list_ch_29_read_data__empty_n;
  assign read_A_29_A_read_data_s_dout = { 1'b0 , edge_list_ch_29_read_data__dout };
  assign read_A_29_A_read_data_s_empty_n = edge_list_ch_29_read_data__empty_n;
  assign edge_list_ch_29_read_data__read = read_A_29_A_read_data_s_read;
  assign read_A_29_A_write_addr_offset = read_A_29___edge_list_ch_29__q0;
  assign edge_list_ch_29_write_addr__din = read_A_29_A_write_addr_s_din;
  assign read_A_29_A_write_addr_s_full_n = edge_list_ch_29_write_addr__full_n;
  assign edge_list_ch_29_write_addr__write = read_A_29_A_write_addr_s_write;
  assign edge_list_ch_29_write_data__din = read_A_29_A_write_data_din;
  assign read_A_29_A_write_data_full_n = edge_list_ch_29_write_data__full_n;
  assign edge_list_ch_29_write_data__write = read_A_29_A_write_data_write;
  assign read_A_29_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_29_write_resp__dout };
  assign read_A_29_A_write_resp_peek_empty_n = edge_list_ch_29_write_resp__empty_n;
  assign read_A_29_A_write_resp_s_dout = { 1'b0 , edge_list_ch_29_write_resp__dout };
  assign read_A_29_A_write_resp_s_empty_n = edge_list_ch_29_write_resp__empty_n;
  assign edge_list_ch_29_write_resp__read = read_A_29_A_write_resp_s_read;
  assign read_A_29_P_N = read_A_29___P_N__q0;
  assign read_A_29_ap_clk = ap_clk;
  assign read_A_29__ap_done = read_A_29_ap_done;
  assign read_A_29__ap_idle = read_A_29_ap_idle;
  assign read_A_29__ap_ready = read_A_29_ap_ready;
  assign read_A_29_ap_rst_n = ap_rst_n;
  assign read_A_29_ap_start = read_A_29__ap_start;
  assign fifo_A_29__din = read_A_29_fifo_A_din;
  assign read_A_29_fifo_A_full_n = fifo_A_29__full_n;
  assign fifo_A_29__write = read_A_29_fifo_A_write;
  assign read_A_30_A_len = read_A_30___NUM_A_LEN__q0;
  assign read_A_30_A_read_addr_offset = read_A_30___edge_list_ch_30__q0;
  assign edge_list_ch_30_read_addr__din = read_A_30_A_read_addr_s_din;
  assign read_A_30_A_read_addr_s_full_n = edge_list_ch_30_read_addr__full_n;
  assign edge_list_ch_30_read_addr__write = read_A_30_A_read_addr_s_write;
  assign read_A_30_A_read_data_peek_dout = { 1'b0 , edge_list_ch_30_read_data__dout };
  assign read_A_30_A_read_data_peek_empty_n = edge_list_ch_30_read_data__empty_n;
  assign read_A_30_A_read_data_s_dout = { 1'b0 , edge_list_ch_30_read_data__dout };
  assign read_A_30_A_read_data_s_empty_n = edge_list_ch_30_read_data__empty_n;
  assign edge_list_ch_30_read_data__read = read_A_30_A_read_data_s_read;
  assign read_A_30_A_write_addr_offset = read_A_30___edge_list_ch_30__q0;
  assign edge_list_ch_30_write_addr__din = read_A_30_A_write_addr_s_din;
  assign read_A_30_A_write_addr_s_full_n = edge_list_ch_30_write_addr__full_n;
  assign edge_list_ch_30_write_addr__write = read_A_30_A_write_addr_s_write;
  assign edge_list_ch_30_write_data__din = read_A_30_A_write_data_din;
  assign read_A_30_A_write_data_full_n = edge_list_ch_30_write_data__full_n;
  assign edge_list_ch_30_write_data__write = read_A_30_A_write_data_write;
  assign read_A_30_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_30_write_resp__dout };
  assign read_A_30_A_write_resp_peek_empty_n = edge_list_ch_30_write_resp__empty_n;
  assign read_A_30_A_write_resp_s_dout = { 1'b0 , edge_list_ch_30_write_resp__dout };
  assign read_A_30_A_write_resp_s_empty_n = edge_list_ch_30_write_resp__empty_n;
  assign edge_list_ch_30_write_resp__read = read_A_30_A_write_resp_s_read;
  assign read_A_30_P_N = read_A_30___P_N__q0;
  assign read_A_30_ap_clk = ap_clk;
  assign read_A_30__ap_done = read_A_30_ap_done;
  assign read_A_30__ap_idle = read_A_30_ap_idle;
  assign read_A_30__ap_ready = read_A_30_ap_ready;
  assign read_A_30_ap_rst_n = ap_rst_n;
  assign read_A_30_ap_start = read_A_30__ap_start;
  assign fifo_A_30__din = read_A_30_fifo_A_din;
  assign read_A_30_fifo_A_full_n = fifo_A_30__full_n;
  assign fifo_A_30__write = read_A_30_fifo_A_write;
  assign read_A_31_A_len = read_A_31___NUM_A_LEN__q0;
  assign read_A_31_A_read_addr_offset = read_A_31___edge_list_ch_31__q0;
  assign edge_list_ch_31_read_addr__din = read_A_31_A_read_addr_s_din;
  assign read_A_31_A_read_addr_s_full_n = edge_list_ch_31_read_addr__full_n;
  assign edge_list_ch_31_read_addr__write = read_A_31_A_read_addr_s_write;
  assign read_A_31_A_read_data_peek_dout = { 1'b0 , edge_list_ch_31_read_data__dout };
  assign read_A_31_A_read_data_peek_empty_n = edge_list_ch_31_read_data__empty_n;
  assign read_A_31_A_read_data_s_dout = { 1'b0 , edge_list_ch_31_read_data__dout };
  assign read_A_31_A_read_data_s_empty_n = edge_list_ch_31_read_data__empty_n;
  assign edge_list_ch_31_read_data__read = read_A_31_A_read_data_s_read;
  assign read_A_31_A_write_addr_offset = read_A_31___edge_list_ch_31__q0;
  assign edge_list_ch_31_write_addr__din = read_A_31_A_write_addr_s_din;
  assign read_A_31_A_write_addr_s_full_n = edge_list_ch_31_write_addr__full_n;
  assign edge_list_ch_31_write_addr__write = read_A_31_A_write_addr_s_write;
  assign edge_list_ch_31_write_data__din = read_A_31_A_write_data_din;
  assign read_A_31_A_write_data_full_n = edge_list_ch_31_write_data__full_n;
  assign edge_list_ch_31_write_data__write = read_A_31_A_write_data_write;
  assign read_A_31_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_31_write_resp__dout };
  assign read_A_31_A_write_resp_peek_empty_n = edge_list_ch_31_write_resp__empty_n;
  assign read_A_31_A_write_resp_s_dout = { 1'b0 , edge_list_ch_31_write_resp__dout };
  assign read_A_31_A_write_resp_s_empty_n = edge_list_ch_31_write_resp__empty_n;
  assign edge_list_ch_31_write_resp__read = read_A_31_A_write_resp_s_read;
  assign read_A_31_P_N = read_A_31___P_N__q0;
  assign read_A_31_ap_clk = ap_clk;
  assign read_A_31__ap_done = read_A_31_ap_done;
  assign read_A_31__ap_idle = read_A_31_ap_idle;
  assign read_A_31__ap_ready = read_A_31_ap_ready;
  assign read_A_31_ap_rst_n = ap_rst_n;
  assign read_A_31_ap_start = read_A_31__ap_start;
  assign fifo_A_31__din = read_A_31_fifo_A_din;
  assign read_A_31_fifo_A_full_n = fifo_A_31__full_n;
  assign fifo_A_31__write = read_A_31_fifo_A_write;
  assign read_A_32_A_len = read_A_32___NUM_A_LEN__q0;
  assign read_A_32_A_read_addr_offset = read_A_32___edge_list_ch_32__q0;
  assign edge_list_ch_32_read_addr__din = read_A_32_A_read_addr_s_din;
  assign read_A_32_A_read_addr_s_full_n = edge_list_ch_32_read_addr__full_n;
  assign edge_list_ch_32_read_addr__write = read_A_32_A_read_addr_s_write;
  assign read_A_32_A_read_data_peek_dout = { 1'b0 , edge_list_ch_32_read_data__dout };
  assign read_A_32_A_read_data_peek_empty_n = edge_list_ch_32_read_data__empty_n;
  assign read_A_32_A_read_data_s_dout = { 1'b0 , edge_list_ch_32_read_data__dout };
  assign read_A_32_A_read_data_s_empty_n = edge_list_ch_32_read_data__empty_n;
  assign edge_list_ch_32_read_data__read = read_A_32_A_read_data_s_read;
  assign read_A_32_A_write_addr_offset = read_A_32___edge_list_ch_32__q0;
  assign edge_list_ch_32_write_addr__din = read_A_32_A_write_addr_s_din;
  assign read_A_32_A_write_addr_s_full_n = edge_list_ch_32_write_addr__full_n;
  assign edge_list_ch_32_write_addr__write = read_A_32_A_write_addr_s_write;
  assign edge_list_ch_32_write_data__din = read_A_32_A_write_data_din;
  assign read_A_32_A_write_data_full_n = edge_list_ch_32_write_data__full_n;
  assign edge_list_ch_32_write_data__write = read_A_32_A_write_data_write;
  assign read_A_32_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_32_write_resp__dout };
  assign read_A_32_A_write_resp_peek_empty_n = edge_list_ch_32_write_resp__empty_n;
  assign read_A_32_A_write_resp_s_dout = { 1'b0 , edge_list_ch_32_write_resp__dout };
  assign read_A_32_A_write_resp_s_empty_n = edge_list_ch_32_write_resp__empty_n;
  assign edge_list_ch_32_write_resp__read = read_A_32_A_write_resp_s_read;
  assign read_A_32_P_N = read_A_32___P_N__q0;
  assign read_A_32_ap_clk = ap_clk;
  assign read_A_32__ap_done = read_A_32_ap_done;
  assign read_A_32__ap_idle = read_A_32_ap_idle;
  assign read_A_32__ap_ready = read_A_32_ap_ready;
  assign read_A_32_ap_rst_n = ap_rst_n;
  assign read_A_32_ap_start = read_A_32__ap_start;
  assign fifo_A_32__din = read_A_32_fifo_A_din;
  assign read_A_32_fifo_A_full_n = fifo_A_32__full_n;
  assign fifo_A_32__write = read_A_32_fifo_A_write;
  assign read_A_33_A_len = read_A_33___NUM_A_LEN__q0;
  assign read_A_33_A_read_addr_offset = read_A_33___edge_list_ch_33__q0;
  assign edge_list_ch_33_read_addr__din = read_A_33_A_read_addr_s_din;
  assign read_A_33_A_read_addr_s_full_n = edge_list_ch_33_read_addr__full_n;
  assign edge_list_ch_33_read_addr__write = read_A_33_A_read_addr_s_write;
  assign read_A_33_A_read_data_peek_dout = { 1'b0 , edge_list_ch_33_read_data__dout };
  assign read_A_33_A_read_data_peek_empty_n = edge_list_ch_33_read_data__empty_n;
  assign read_A_33_A_read_data_s_dout = { 1'b0 , edge_list_ch_33_read_data__dout };
  assign read_A_33_A_read_data_s_empty_n = edge_list_ch_33_read_data__empty_n;
  assign edge_list_ch_33_read_data__read = read_A_33_A_read_data_s_read;
  assign read_A_33_A_write_addr_offset = read_A_33___edge_list_ch_33__q0;
  assign edge_list_ch_33_write_addr__din = read_A_33_A_write_addr_s_din;
  assign read_A_33_A_write_addr_s_full_n = edge_list_ch_33_write_addr__full_n;
  assign edge_list_ch_33_write_addr__write = read_A_33_A_write_addr_s_write;
  assign edge_list_ch_33_write_data__din = read_A_33_A_write_data_din;
  assign read_A_33_A_write_data_full_n = edge_list_ch_33_write_data__full_n;
  assign edge_list_ch_33_write_data__write = read_A_33_A_write_data_write;
  assign read_A_33_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_33_write_resp__dout };
  assign read_A_33_A_write_resp_peek_empty_n = edge_list_ch_33_write_resp__empty_n;
  assign read_A_33_A_write_resp_s_dout = { 1'b0 , edge_list_ch_33_write_resp__dout };
  assign read_A_33_A_write_resp_s_empty_n = edge_list_ch_33_write_resp__empty_n;
  assign edge_list_ch_33_write_resp__read = read_A_33_A_write_resp_s_read;
  assign read_A_33_P_N = read_A_33___P_N__q0;
  assign read_A_33_ap_clk = ap_clk;
  assign read_A_33__ap_done = read_A_33_ap_done;
  assign read_A_33__ap_idle = read_A_33_ap_idle;
  assign read_A_33__ap_ready = read_A_33_ap_ready;
  assign read_A_33_ap_rst_n = ap_rst_n;
  assign read_A_33_ap_start = read_A_33__ap_start;
  assign fifo_A_33__din = read_A_33_fifo_A_din;
  assign read_A_33_fifo_A_full_n = fifo_A_33__full_n;
  assign fifo_A_33__write = read_A_33_fifo_A_write;
  assign read_A_34_A_len = read_A_34___NUM_A_LEN__q0;
  assign read_A_34_A_read_addr_offset = read_A_34___edge_list_ch_34__q0;
  assign edge_list_ch_34_read_addr__din = read_A_34_A_read_addr_s_din;
  assign read_A_34_A_read_addr_s_full_n = edge_list_ch_34_read_addr__full_n;
  assign edge_list_ch_34_read_addr__write = read_A_34_A_read_addr_s_write;
  assign read_A_34_A_read_data_peek_dout = { 1'b0 , edge_list_ch_34_read_data__dout };
  assign read_A_34_A_read_data_peek_empty_n = edge_list_ch_34_read_data__empty_n;
  assign read_A_34_A_read_data_s_dout = { 1'b0 , edge_list_ch_34_read_data__dout };
  assign read_A_34_A_read_data_s_empty_n = edge_list_ch_34_read_data__empty_n;
  assign edge_list_ch_34_read_data__read = read_A_34_A_read_data_s_read;
  assign read_A_34_A_write_addr_offset = read_A_34___edge_list_ch_34__q0;
  assign edge_list_ch_34_write_addr__din = read_A_34_A_write_addr_s_din;
  assign read_A_34_A_write_addr_s_full_n = edge_list_ch_34_write_addr__full_n;
  assign edge_list_ch_34_write_addr__write = read_A_34_A_write_addr_s_write;
  assign edge_list_ch_34_write_data__din = read_A_34_A_write_data_din;
  assign read_A_34_A_write_data_full_n = edge_list_ch_34_write_data__full_n;
  assign edge_list_ch_34_write_data__write = read_A_34_A_write_data_write;
  assign read_A_34_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_34_write_resp__dout };
  assign read_A_34_A_write_resp_peek_empty_n = edge_list_ch_34_write_resp__empty_n;
  assign read_A_34_A_write_resp_s_dout = { 1'b0 , edge_list_ch_34_write_resp__dout };
  assign read_A_34_A_write_resp_s_empty_n = edge_list_ch_34_write_resp__empty_n;
  assign edge_list_ch_34_write_resp__read = read_A_34_A_write_resp_s_read;
  assign read_A_34_P_N = read_A_34___P_N__q0;
  assign read_A_34_ap_clk = ap_clk;
  assign read_A_34__ap_done = read_A_34_ap_done;
  assign read_A_34__ap_idle = read_A_34_ap_idle;
  assign read_A_34__ap_ready = read_A_34_ap_ready;
  assign read_A_34_ap_rst_n = ap_rst_n;
  assign read_A_34_ap_start = read_A_34__ap_start;
  assign fifo_A_34__din = read_A_34_fifo_A_din;
  assign read_A_34_fifo_A_full_n = fifo_A_34__full_n;
  assign fifo_A_34__write = read_A_34_fifo_A_write;
  assign read_A_35_A_len = read_A_35___NUM_A_LEN__q0;
  assign read_A_35_A_read_addr_offset = read_A_35___edge_list_ch_35__q0;
  assign edge_list_ch_35_read_addr__din = read_A_35_A_read_addr_s_din;
  assign read_A_35_A_read_addr_s_full_n = edge_list_ch_35_read_addr__full_n;
  assign edge_list_ch_35_read_addr__write = read_A_35_A_read_addr_s_write;
  assign read_A_35_A_read_data_peek_dout = { 1'b0 , edge_list_ch_35_read_data__dout };
  assign read_A_35_A_read_data_peek_empty_n = edge_list_ch_35_read_data__empty_n;
  assign read_A_35_A_read_data_s_dout = { 1'b0 , edge_list_ch_35_read_data__dout };
  assign read_A_35_A_read_data_s_empty_n = edge_list_ch_35_read_data__empty_n;
  assign edge_list_ch_35_read_data__read = read_A_35_A_read_data_s_read;
  assign read_A_35_A_write_addr_offset = read_A_35___edge_list_ch_35__q0;
  assign edge_list_ch_35_write_addr__din = read_A_35_A_write_addr_s_din;
  assign read_A_35_A_write_addr_s_full_n = edge_list_ch_35_write_addr__full_n;
  assign edge_list_ch_35_write_addr__write = read_A_35_A_write_addr_s_write;
  assign edge_list_ch_35_write_data__din = read_A_35_A_write_data_din;
  assign read_A_35_A_write_data_full_n = edge_list_ch_35_write_data__full_n;
  assign edge_list_ch_35_write_data__write = read_A_35_A_write_data_write;
  assign read_A_35_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_35_write_resp__dout };
  assign read_A_35_A_write_resp_peek_empty_n = edge_list_ch_35_write_resp__empty_n;
  assign read_A_35_A_write_resp_s_dout = { 1'b0 , edge_list_ch_35_write_resp__dout };
  assign read_A_35_A_write_resp_s_empty_n = edge_list_ch_35_write_resp__empty_n;
  assign edge_list_ch_35_write_resp__read = read_A_35_A_write_resp_s_read;
  assign read_A_35_P_N = read_A_35___P_N__q0;
  assign read_A_35_ap_clk = ap_clk;
  assign read_A_35__ap_done = read_A_35_ap_done;
  assign read_A_35__ap_idle = read_A_35_ap_idle;
  assign read_A_35__ap_ready = read_A_35_ap_ready;
  assign read_A_35_ap_rst_n = ap_rst_n;
  assign read_A_35_ap_start = read_A_35__ap_start;
  assign fifo_A_35__din = read_A_35_fifo_A_din;
  assign read_A_35_fifo_A_full_n = fifo_A_35__full_n;
  assign fifo_A_35__write = read_A_35_fifo_A_write;
  assign read_A_36_A_len = read_A_36___NUM_A_LEN__q0;
  assign read_A_36_A_read_addr_offset = read_A_36___edge_list_ch_36__q0;
  assign edge_list_ch_36_read_addr__din = read_A_36_A_read_addr_s_din;
  assign read_A_36_A_read_addr_s_full_n = edge_list_ch_36_read_addr__full_n;
  assign edge_list_ch_36_read_addr__write = read_A_36_A_read_addr_s_write;
  assign read_A_36_A_read_data_peek_dout = { 1'b0 , edge_list_ch_36_read_data__dout };
  assign read_A_36_A_read_data_peek_empty_n = edge_list_ch_36_read_data__empty_n;
  assign read_A_36_A_read_data_s_dout = { 1'b0 , edge_list_ch_36_read_data__dout };
  assign read_A_36_A_read_data_s_empty_n = edge_list_ch_36_read_data__empty_n;
  assign edge_list_ch_36_read_data__read = read_A_36_A_read_data_s_read;
  assign read_A_36_A_write_addr_offset = read_A_36___edge_list_ch_36__q0;
  assign edge_list_ch_36_write_addr__din = read_A_36_A_write_addr_s_din;
  assign read_A_36_A_write_addr_s_full_n = edge_list_ch_36_write_addr__full_n;
  assign edge_list_ch_36_write_addr__write = read_A_36_A_write_addr_s_write;
  assign edge_list_ch_36_write_data__din = read_A_36_A_write_data_din;
  assign read_A_36_A_write_data_full_n = edge_list_ch_36_write_data__full_n;
  assign edge_list_ch_36_write_data__write = read_A_36_A_write_data_write;
  assign read_A_36_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_36_write_resp__dout };
  assign read_A_36_A_write_resp_peek_empty_n = edge_list_ch_36_write_resp__empty_n;
  assign read_A_36_A_write_resp_s_dout = { 1'b0 , edge_list_ch_36_write_resp__dout };
  assign read_A_36_A_write_resp_s_empty_n = edge_list_ch_36_write_resp__empty_n;
  assign edge_list_ch_36_write_resp__read = read_A_36_A_write_resp_s_read;
  assign read_A_36_P_N = read_A_36___P_N__q0;
  assign read_A_36_ap_clk = ap_clk;
  assign read_A_36__ap_done = read_A_36_ap_done;
  assign read_A_36__ap_idle = read_A_36_ap_idle;
  assign read_A_36__ap_ready = read_A_36_ap_ready;
  assign read_A_36_ap_rst_n = ap_rst_n;
  assign read_A_36_ap_start = read_A_36__ap_start;
  assign fifo_A_36__din = read_A_36_fifo_A_din;
  assign read_A_36_fifo_A_full_n = fifo_A_36__full_n;
  assign fifo_A_36__write = read_A_36_fifo_A_write;
  assign read_A_37_A_len = read_A_37___NUM_A_LEN__q0;
  assign read_A_37_A_read_addr_offset = read_A_37___edge_list_ch_37__q0;
  assign edge_list_ch_37_read_addr__din = read_A_37_A_read_addr_s_din;
  assign read_A_37_A_read_addr_s_full_n = edge_list_ch_37_read_addr__full_n;
  assign edge_list_ch_37_read_addr__write = read_A_37_A_read_addr_s_write;
  assign read_A_37_A_read_data_peek_dout = { 1'b0 , edge_list_ch_37_read_data__dout };
  assign read_A_37_A_read_data_peek_empty_n = edge_list_ch_37_read_data__empty_n;
  assign read_A_37_A_read_data_s_dout = { 1'b0 , edge_list_ch_37_read_data__dout };
  assign read_A_37_A_read_data_s_empty_n = edge_list_ch_37_read_data__empty_n;
  assign edge_list_ch_37_read_data__read = read_A_37_A_read_data_s_read;
  assign read_A_37_A_write_addr_offset = read_A_37___edge_list_ch_37__q0;
  assign edge_list_ch_37_write_addr__din = read_A_37_A_write_addr_s_din;
  assign read_A_37_A_write_addr_s_full_n = edge_list_ch_37_write_addr__full_n;
  assign edge_list_ch_37_write_addr__write = read_A_37_A_write_addr_s_write;
  assign edge_list_ch_37_write_data__din = read_A_37_A_write_data_din;
  assign read_A_37_A_write_data_full_n = edge_list_ch_37_write_data__full_n;
  assign edge_list_ch_37_write_data__write = read_A_37_A_write_data_write;
  assign read_A_37_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_37_write_resp__dout };
  assign read_A_37_A_write_resp_peek_empty_n = edge_list_ch_37_write_resp__empty_n;
  assign read_A_37_A_write_resp_s_dout = { 1'b0 , edge_list_ch_37_write_resp__dout };
  assign read_A_37_A_write_resp_s_empty_n = edge_list_ch_37_write_resp__empty_n;
  assign edge_list_ch_37_write_resp__read = read_A_37_A_write_resp_s_read;
  assign read_A_37_P_N = read_A_37___P_N__q0;
  assign read_A_37_ap_clk = ap_clk;
  assign read_A_37__ap_done = read_A_37_ap_done;
  assign read_A_37__ap_idle = read_A_37_ap_idle;
  assign read_A_37__ap_ready = read_A_37_ap_ready;
  assign read_A_37_ap_rst_n = ap_rst_n;
  assign read_A_37_ap_start = read_A_37__ap_start;
  assign fifo_A_37__din = read_A_37_fifo_A_din;
  assign read_A_37_fifo_A_full_n = fifo_A_37__full_n;
  assign fifo_A_37__write = read_A_37_fifo_A_write;
  assign read_A_38_A_len = read_A_38___NUM_A_LEN__q0;
  assign read_A_38_A_read_addr_offset = read_A_38___edge_list_ch_38__q0;
  assign edge_list_ch_38_read_addr__din = read_A_38_A_read_addr_s_din;
  assign read_A_38_A_read_addr_s_full_n = edge_list_ch_38_read_addr__full_n;
  assign edge_list_ch_38_read_addr__write = read_A_38_A_read_addr_s_write;
  assign read_A_38_A_read_data_peek_dout = { 1'b0 , edge_list_ch_38_read_data__dout };
  assign read_A_38_A_read_data_peek_empty_n = edge_list_ch_38_read_data__empty_n;
  assign read_A_38_A_read_data_s_dout = { 1'b0 , edge_list_ch_38_read_data__dout };
  assign read_A_38_A_read_data_s_empty_n = edge_list_ch_38_read_data__empty_n;
  assign edge_list_ch_38_read_data__read = read_A_38_A_read_data_s_read;
  assign read_A_38_A_write_addr_offset = read_A_38___edge_list_ch_38__q0;
  assign edge_list_ch_38_write_addr__din = read_A_38_A_write_addr_s_din;
  assign read_A_38_A_write_addr_s_full_n = edge_list_ch_38_write_addr__full_n;
  assign edge_list_ch_38_write_addr__write = read_A_38_A_write_addr_s_write;
  assign edge_list_ch_38_write_data__din = read_A_38_A_write_data_din;
  assign read_A_38_A_write_data_full_n = edge_list_ch_38_write_data__full_n;
  assign edge_list_ch_38_write_data__write = read_A_38_A_write_data_write;
  assign read_A_38_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_38_write_resp__dout };
  assign read_A_38_A_write_resp_peek_empty_n = edge_list_ch_38_write_resp__empty_n;
  assign read_A_38_A_write_resp_s_dout = { 1'b0 , edge_list_ch_38_write_resp__dout };
  assign read_A_38_A_write_resp_s_empty_n = edge_list_ch_38_write_resp__empty_n;
  assign edge_list_ch_38_write_resp__read = read_A_38_A_write_resp_s_read;
  assign read_A_38_P_N = read_A_38___P_N__q0;
  assign read_A_38_ap_clk = ap_clk;
  assign read_A_38__ap_done = read_A_38_ap_done;
  assign read_A_38__ap_idle = read_A_38_ap_idle;
  assign read_A_38__ap_ready = read_A_38_ap_ready;
  assign read_A_38_ap_rst_n = ap_rst_n;
  assign read_A_38_ap_start = read_A_38__ap_start;
  assign fifo_A_38__din = read_A_38_fifo_A_din;
  assign read_A_38_fifo_A_full_n = fifo_A_38__full_n;
  assign fifo_A_38__write = read_A_38_fifo_A_write;
  assign read_A_39_A_len = read_A_39___NUM_A_LEN__q0;
  assign read_A_39_A_read_addr_offset = read_A_39___edge_list_ch_39__q0;
  assign edge_list_ch_39_read_addr__din = read_A_39_A_read_addr_s_din;
  assign read_A_39_A_read_addr_s_full_n = edge_list_ch_39_read_addr__full_n;
  assign edge_list_ch_39_read_addr__write = read_A_39_A_read_addr_s_write;
  assign read_A_39_A_read_data_peek_dout = { 1'b0 , edge_list_ch_39_read_data__dout };
  assign read_A_39_A_read_data_peek_empty_n = edge_list_ch_39_read_data__empty_n;
  assign read_A_39_A_read_data_s_dout = { 1'b0 , edge_list_ch_39_read_data__dout };
  assign read_A_39_A_read_data_s_empty_n = edge_list_ch_39_read_data__empty_n;
  assign edge_list_ch_39_read_data__read = read_A_39_A_read_data_s_read;
  assign read_A_39_A_write_addr_offset = read_A_39___edge_list_ch_39__q0;
  assign edge_list_ch_39_write_addr__din = read_A_39_A_write_addr_s_din;
  assign read_A_39_A_write_addr_s_full_n = edge_list_ch_39_write_addr__full_n;
  assign edge_list_ch_39_write_addr__write = read_A_39_A_write_addr_s_write;
  assign edge_list_ch_39_write_data__din = read_A_39_A_write_data_din;
  assign read_A_39_A_write_data_full_n = edge_list_ch_39_write_data__full_n;
  assign edge_list_ch_39_write_data__write = read_A_39_A_write_data_write;
  assign read_A_39_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_39_write_resp__dout };
  assign read_A_39_A_write_resp_peek_empty_n = edge_list_ch_39_write_resp__empty_n;
  assign read_A_39_A_write_resp_s_dout = { 1'b0 , edge_list_ch_39_write_resp__dout };
  assign read_A_39_A_write_resp_s_empty_n = edge_list_ch_39_write_resp__empty_n;
  assign edge_list_ch_39_write_resp__read = read_A_39_A_write_resp_s_read;
  assign read_A_39_P_N = read_A_39___P_N__q0;
  assign read_A_39_ap_clk = ap_clk;
  assign read_A_39__ap_done = read_A_39_ap_done;
  assign read_A_39__ap_idle = read_A_39_ap_idle;
  assign read_A_39__ap_ready = read_A_39_ap_ready;
  assign read_A_39_ap_rst_n = ap_rst_n;
  assign read_A_39_ap_start = read_A_39__ap_start;
  assign fifo_A_39__din = read_A_39_fifo_A_din;
  assign read_A_39_fifo_A_full_n = fifo_A_39__full_n;
  assign fifo_A_39__write = read_A_39_fifo_A_write;
  assign read_A_40_A_len = read_A_40___NUM_A_LEN__q0;
  assign read_A_40_A_read_addr_offset = read_A_40___edge_list_ch_40__q0;
  assign edge_list_ch_40_read_addr__din = read_A_40_A_read_addr_s_din;
  assign read_A_40_A_read_addr_s_full_n = edge_list_ch_40_read_addr__full_n;
  assign edge_list_ch_40_read_addr__write = read_A_40_A_read_addr_s_write;
  assign read_A_40_A_read_data_peek_dout = { 1'b0 , edge_list_ch_40_read_data__dout };
  assign read_A_40_A_read_data_peek_empty_n = edge_list_ch_40_read_data__empty_n;
  assign read_A_40_A_read_data_s_dout = { 1'b0 , edge_list_ch_40_read_data__dout };
  assign read_A_40_A_read_data_s_empty_n = edge_list_ch_40_read_data__empty_n;
  assign edge_list_ch_40_read_data__read = read_A_40_A_read_data_s_read;
  assign read_A_40_A_write_addr_offset = read_A_40___edge_list_ch_40__q0;
  assign edge_list_ch_40_write_addr__din = read_A_40_A_write_addr_s_din;
  assign read_A_40_A_write_addr_s_full_n = edge_list_ch_40_write_addr__full_n;
  assign edge_list_ch_40_write_addr__write = read_A_40_A_write_addr_s_write;
  assign edge_list_ch_40_write_data__din = read_A_40_A_write_data_din;
  assign read_A_40_A_write_data_full_n = edge_list_ch_40_write_data__full_n;
  assign edge_list_ch_40_write_data__write = read_A_40_A_write_data_write;
  assign read_A_40_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_40_write_resp__dout };
  assign read_A_40_A_write_resp_peek_empty_n = edge_list_ch_40_write_resp__empty_n;
  assign read_A_40_A_write_resp_s_dout = { 1'b0 , edge_list_ch_40_write_resp__dout };
  assign read_A_40_A_write_resp_s_empty_n = edge_list_ch_40_write_resp__empty_n;
  assign edge_list_ch_40_write_resp__read = read_A_40_A_write_resp_s_read;
  assign read_A_40_P_N = read_A_40___P_N__q0;
  assign read_A_40_ap_clk = ap_clk;
  assign read_A_40__ap_done = read_A_40_ap_done;
  assign read_A_40__ap_idle = read_A_40_ap_idle;
  assign read_A_40__ap_ready = read_A_40_ap_ready;
  assign read_A_40_ap_rst_n = ap_rst_n;
  assign read_A_40_ap_start = read_A_40__ap_start;
  assign fifo_A_40__din = read_A_40_fifo_A_din;
  assign read_A_40_fifo_A_full_n = fifo_A_40__full_n;
  assign fifo_A_40__write = read_A_40_fifo_A_write;
  assign read_A_41_A_len = read_A_41___NUM_A_LEN__q0;
  assign read_A_41_A_read_addr_offset = read_A_41___edge_list_ch_41__q0;
  assign edge_list_ch_41_read_addr__din = read_A_41_A_read_addr_s_din;
  assign read_A_41_A_read_addr_s_full_n = edge_list_ch_41_read_addr__full_n;
  assign edge_list_ch_41_read_addr__write = read_A_41_A_read_addr_s_write;
  assign read_A_41_A_read_data_peek_dout = { 1'b0 , edge_list_ch_41_read_data__dout };
  assign read_A_41_A_read_data_peek_empty_n = edge_list_ch_41_read_data__empty_n;
  assign read_A_41_A_read_data_s_dout = { 1'b0 , edge_list_ch_41_read_data__dout };
  assign read_A_41_A_read_data_s_empty_n = edge_list_ch_41_read_data__empty_n;
  assign edge_list_ch_41_read_data__read = read_A_41_A_read_data_s_read;
  assign read_A_41_A_write_addr_offset = read_A_41___edge_list_ch_41__q0;
  assign edge_list_ch_41_write_addr__din = read_A_41_A_write_addr_s_din;
  assign read_A_41_A_write_addr_s_full_n = edge_list_ch_41_write_addr__full_n;
  assign edge_list_ch_41_write_addr__write = read_A_41_A_write_addr_s_write;
  assign edge_list_ch_41_write_data__din = read_A_41_A_write_data_din;
  assign read_A_41_A_write_data_full_n = edge_list_ch_41_write_data__full_n;
  assign edge_list_ch_41_write_data__write = read_A_41_A_write_data_write;
  assign read_A_41_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_41_write_resp__dout };
  assign read_A_41_A_write_resp_peek_empty_n = edge_list_ch_41_write_resp__empty_n;
  assign read_A_41_A_write_resp_s_dout = { 1'b0 , edge_list_ch_41_write_resp__dout };
  assign read_A_41_A_write_resp_s_empty_n = edge_list_ch_41_write_resp__empty_n;
  assign edge_list_ch_41_write_resp__read = read_A_41_A_write_resp_s_read;
  assign read_A_41_P_N = read_A_41___P_N__q0;
  assign read_A_41_ap_clk = ap_clk;
  assign read_A_41__ap_done = read_A_41_ap_done;
  assign read_A_41__ap_idle = read_A_41_ap_idle;
  assign read_A_41__ap_ready = read_A_41_ap_ready;
  assign read_A_41_ap_rst_n = ap_rst_n;
  assign read_A_41_ap_start = read_A_41__ap_start;
  assign fifo_A_41__din = read_A_41_fifo_A_din;
  assign read_A_41_fifo_A_full_n = fifo_A_41__full_n;
  assign fifo_A_41__write = read_A_41_fifo_A_write;
  assign read_A_42_A_len = read_A_42___NUM_A_LEN__q0;
  assign read_A_42_A_read_addr_offset = read_A_42___edge_list_ch_42__q0;
  assign edge_list_ch_42_read_addr__din = read_A_42_A_read_addr_s_din;
  assign read_A_42_A_read_addr_s_full_n = edge_list_ch_42_read_addr__full_n;
  assign edge_list_ch_42_read_addr__write = read_A_42_A_read_addr_s_write;
  assign read_A_42_A_read_data_peek_dout = { 1'b0 , edge_list_ch_42_read_data__dout };
  assign read_A_42_A_read_data_peek_empty_n = edge_list_ch_42_read_data__empty_n;
  assign read_A_42_A_read_data_s_dout = { 1'b0 , edge_list_ch_42_read_data__dout };
  assign read_A_42_A_read_data_s_empty_n = edge_list_ch_42_read_data__empty_n;
  assign edge_list_ch_42_read_data__read = read_A_42_A_read_data_s_read;
  assign read_A_42_A_write_addr_offset = read_A_42___edge_list_ch_42__q0;
  assign edge_list_ch_42_write_addr__din = read_A_42_A_write_addr_s_din;
  assign read_A_42_A_write_addr_s_full_n = edge_list_ch_42_write_addr__full_n;
  assign edge_list_ch_42_write_addr__write = read_A_42_A_write_addr_s_write;
  assign edge_list_ch_42_write_data__din = read_A_42_A_write_data_din;
  assign read_A_42_A_write_data_full_n = edge_list_ch_42_write_data__full_n;
  assign edge_list_ch_42_write_data__write = read_A_42_A_write_data_write;
  assign read_A_42_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_42_write_resp__dout };
  assign read_A_42_A_write_resp_peek_empty_n = edge_list_ch_42_write_resp__empty_n;
  assign read_A_42_A_write_resp_s_dout = { 1'b0 , edge_list_ch_42_write_resp__dout };
  assign read_A_42_A_write_resp_s_empty_n = edge_list_ch_42_write_resp__empty_n;
  assign edge_list_ch_42_write_resp__read = read_A_42_A_write_resp_s_read;
  assign read_A_42_P_N = read_A_42___P_N__q0;
  assign read_A_42_ap_clk = ap_clk;
  assign read_A_42__ap_done = read_A_42_ap_done;
  assign read_A_42__ap_idle = read_A_42_ap_idle;
  assign read_A_42__ap_ready = read_A_42_ap_ready;
  assign read_A_42_ap_rst_n = ap_rst_n;
  assign read_A_42_ap_start = read_A_42__ap_start;
  assign fifo_A_42__din = read_A_42_fifo_A_din;
  assign read_A_42_fifo_A_full_n = fifo_A_42__full_n;
  assign fifo_A_42__write = read_A_42_fifo_A_write;
  assign read_A_43_A_len = read_A_43___NUM_A_LEN__q0;
  assign read_A_43_A_read_addr_offset = read_A_43___edge_list_ch_43__q0;
  assign edge_list_ch_43_read_addr__din = read_A_43_A_read_addr_s_din;
  assign read_A_43_A_read_addr_s_full_n = edge_list_ch_43_read_addr__full_n;
  assign edge_list_ch_43_read_addr__write = read_A_43_A_read_addr_s_write;
  assign read_A_43_A_read_data_peek_dout = { 1'b0 , edge_list_ch_43_read_data__dout };
  assign read_A_43_A_read_data_peek_empty_n = edge_list_ch_43_read_data__empty_n;
  assign read_A_43_A_read_data_s_dout = { 1'b0 , edge_list_ch_43_read_data__dout };
  assign read_A_43_A_read_data_s_empty_n = edge_list_ch_43_read_data__empty_n;
  assign edge_list_ch_43_read_data__read = read_A_43_A_read_data_s_read;
  assign read_A_43_A_write_addr_offset = read_A_43___edge_list_ch_43__q0;
  assign edge_list_ch_43_write_addr__din = read_A_43_A_write_addr_s_din;
  assign read_A_43_A_write_addr_s_full_n = edge_list_ch_43_write_addr__full_n;
  assign edge_list_ch_43_write_addr__write = read_A_43_A_write_addr_s_write;
  assign edge_list_ch_43_write_data__din = read_A_43_A_write_data_din;
  assign read_A_43_A_write_data_full_n = edge_list_ch_43_write_data__full_n;
  assign edge_list_ch_43_write_data__write = read_A_43_A_write_data_write;
  assign read_A_43_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_43_write_resp__dout };
  assign read_A_43_A_write_resp_peek_empty_n = edge_list_ch_43_write_resp__empty_n;
  assign read_A_43_A_write_resp_s_dout = { 1'b0 , edge_list_ch_43_write_resp__dout };
  assign read_A_43_A_write_resp_s_empty_n = edge_list_ch_43_write_resp__empty_n;
  assign edge_list_ch_43_write_resp__read = read_A_43_A_write_resp_s_read;
  assign read_A_43_P_N = read_A_43___P_N__q0;
  assign read_A_43_ap_clk = ap_clk;
  assign read_A_43__ap_done = read_A_43_ap_done;
  assign read_A_43__ap_idle = read_A_43_ap_idle;
  assign read_A_43__ap_ready = read_A_43_ap_ready;
  assign read_A_43_ap_rst_n = ap_rst_n;
  assign read_A_43_ap_start = read_A_43__ap_start;
  assign fifo_A_43__din = read_A_43_fifo_A_din;
  assign read_A_43_fifo_A_full_n = fifo_A_43__full_n;
  assign fifo_A_43__write = read_A_43_fifo_A_write;
  assign read_A_44_A_len = read_A_44___NUM_A_LEN__q0;
  assign read_A_44_A_read_addr_offset = read_A_44___edge_list_ch_44__q0;
  assign edge_list_ch_44_read_addr__din = read_A_44_A_read_addr_s_din;
  assign read_A_44_A_read_addr_s_full_n = edge_list_ch_44_read_addr__full_n;
  assign edge_list_ch_44_read_addr__write = read_A_44_A_read_addr_s_write;
  assign read_A_44_A_read_data_peek_dout = { 1'b0 , edge_list_ch_44_read_data__dout };
  assign read_A_44_A_read_data_peek_empty_n = edge_list_ch_44_read_data__empty_n;
  assign read_A_44_A_read_data_s_dout = { 1'b0 , edge_list_ch_44_read_data__dout };
  assign read_A_44_A_read_data_s_empty_n = edge_list_ch_44_read_data__empty_n;
  assign edge_list_ch_44_read_data__read = read_A_44_A_read_data_s_read;
  assign read_A_44_A_write_addr_offset = read_A_44___edge_list_ch_44__q0;
  assign edge_list_ch_44_write_addr__din = read_A_44_A_write_addr_s_din;
  assign read_A_44_A_write_addr_s_full_n = edge_list_ch_44_write_addr__full_n;
  assign edge_list_ch_44_write_addr__write = read_A_44_A_write_addr_s_write;
  assign edge_list_ch_44_write_data__din = read_A_44_A_write_data_din;
  assign read_A_44_A_write_data_full_n = edge_list_ch_44_write_data__full_n;
  assign edge_list_ch_44_write_data__write = read_A_44_A_write_data_write;
  assign read_A_44_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_44_write_resp__dout };
  assign read_A_44_A_write_resp_peek_empty_n = edge_list_ch_44_write_resp__empty_n;
  assign read_A_44_A_write_resp_s_dout = { 1'b0 , edge_list_ch_44_write_resp__dout };
  assign read_A_44_A_write_resp_s_empty_n = edge_list_ch_44_write_resp__empty_n;
  assign edge_list_ch_44_write_resp__read = read_A_44_A_write_resp_s_read;
  assign read_A_44_P_N = read_A_44___P_N__q0;
  assign read_A_44_ap_clk = ap_clk;
  assign read_A_44__ap_done = read_A_44_ap_done;
  assign read_A_44__ap_idle = read_A_44_ap_idle;
  assign read_A_44__ap_ready = read_A_44_ap_ready;
  assign read_A_44_ap_rst_n = ap_rst_n;
  assign read_A_44_ap_start = read_A_44__ap_start;
  assign fifo_A_44__din = read_A_44_fifo_A_din;
  assign read_A_44_fifo_A_full_n = fifo_A_44__full_n;
  assign fifo_A_44__write = read_A_44_fifo_A_write;
  assign read_A_45_A_len = read_A_45___NUM_A_LEN__q0;
  assign read_A_45_A_read_addr_offset = read_A_45___edge_list_ch_45__q0;
  assign edge_list_ch_45_read_addr__din = read_A_45_A_read_addr_s_din;
  assign read_A_45_A_read_addr_s_full_n = edge_list_ch_45_read_addr__full_n;
  assign edge_list_ch_45_read_addr__write = read_A_45_A_read_addr_s_write;
  assign read_A_45_A_read_data_peek_dout = { 1'b0 , edge_list_ch_45_read_data__dout };
  assign read_A_45_A_read_data_peek_empty_n = edge_list_ch_45_read_data__empty_n;
  assign read_A_45_A_read_data_s_dout = { 1'b0 , edge_list_ch_45_read_data__dout };
  assign read_A_45_A_read_data_s_empty_n = edge_list_ch_45_read_data__empty_n;
  assign edge_list_ch_45_read_data__read = read_A_45_A_read_data_s_read;
  assign read_A_45_A_write_addr_offset = read_A_45___edge_list_ch_45__q0;
  assign edge_list_ch_45_write_addr__din = read_A_45_A_write_addr_s_din;
  assign read_A_45_A_write_addr_s_full_n = edge_list_ch_45_write_addr__full_n;
  assign edge_list_ch_45_write_addr__write = read_A_45_A_write_addr_s_write;
  assign edge_list_ch_45_write_data__din = read_A_45_A_write_data_din;
  assign read_A_45_A_write_data_full_n = edge_list_ch_45_write_data__full_n;
  assign edge_list_ch_45_write_data__write = read_A_45_A_write_data_write;
  assign read_A_45_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_45_write_resp__dout };
  assign read_A_45_A_write_resp_peek_empty_n = edge_list_ch_45_write_resp__empty_n;
  assign read_A_45_A_write_resp_s_dout = { 1'b0 , edge_list_ch_45_write_resp__dout };
  assign read_A_45_A_write_resp_s_empty_n = edge_list_ch_45_write_resp__empty_n;
  assign edge_list_ch_45_write_resp__read = read_A_45_A_write_resp_s_read;
  assign read_A_45_P_N = read_A_45___P_N__q0;
  assign read_A_45_ap_clk = ap_clk;
  assign read_A_45__ap_done = read_A_45_ap_done;
  assign read_A_45__ap_idle = read_A_45_ap_idle;
  assign read_A_45__ap_ready = read_A_45_ap_ready;
  assign read_A_45_ap_rst_n = ap_rst_n;
  assign read_A_45_ap_start = read_A_45__ap_start;
  assign fifo_A_45__din = read_A_45_fifo_A_din;
  assign read_A_45_fifo_A_full_n = fifo_A_45__full_n;
  assign fifo_A_45__write = read_A_45_fifo_A_write;
  assign read_A_46_A_len = read_A_46___NUM_A_LEN__q0;
  assign read_A_46_A_read_addr_offset = read_A_46___edge_list_ch_46__q0;
  assign edge_list_ch_46_read_addr__din = read_A_46_A_read_addr_s_din;
  assign read_A_46_A_read_addr_s_full_n = edge_list_ch_46_read_addr__full_n;
  assign edge_list_ch_46_read_addr__write = read_A_46_A_read_addr_s_write;
  assign read_A_46_A_read_data_peek_dout = { 1'b0 , edge_list_ch_46_read_data__dout };
  assign read_A_46_A_read_data_peek_empty_n = edge_list_ch_46_read_data__empty_n;
  assign read_A_46_A_read_data_s_dout = { 1'b0 , edge_list_ch_46_read_data__dout };
  assign read_A_46_A_read_data_s_empty_n = edge_list_ch_46_read_data__empty_n;
  assign edge_list_ch_46_read_data__read = read_A_46_A_read_data_s_read;
  assign read_A_46_A_write_addr_offset = read_A_46___edge_list_ch_46__q0;
  assign edge_list_ch_46_write_addr__din = read_A_46_A_write_addr_s_din;
  assign read_A_46_A_write_addr_s_full_n = edge_list_ch_46_write_addr__full_n;
  assign edge_list_ch_46_write_addr__write = read_A_46_A_write_addr_s_write;
  assign edge_list_ch_46_write_data__din = read_A_46_A_write_data_din;
  assign read_A_46_A_write_data_full_n = edge_list_ch_46_write_data__full_n;
  assign edge_list_ch_46_write_data__write = read_A_46_A_write_data_write;
  assign read_A_46_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_46_write_resp__dout };
  assign read_A_46_A_write_resp_peek_empty_n = edge_list_ch_46_write_resp__empty_n;
  assign read_A_46_A_write_resp_s_dout = { 1'b0 , edge_list_ch_46_write_resp__dout };
  assign read_A_46_A_write_resp_s_empty_n = edge_list_ch_46_write_resp__empty_n;
  assign edge_list_ch_46_write_resp__read = read_A_46_A_write_resp_s_read;
  assign read_A_46_P_N = read_A_46___P_N__q0;
  assign read_A_46_ap_clk = ap_clk;
  assign read_A_46__ap_done = read_A_46_ap_done;
  assign read_A_46__ap_idle = read_A_46_ap_idle;
  assign read_A_46__ap_ready = read_A_46_ap_ready;
  assign read_A_46_ap_rst_n = ap_rst_n;
  assign read_A_46_ap_start = read_A_46__ap_start;
  assign fifo_A_46__din = read_A_46_fifo_A_din;
  assign read_A_46_fifo_A_full_n = fifo_A_46__full_n;
  assign fifo_A_46__write = read_A_46_fifo_A_write;
  assign read_A_47_A_len = read_A_47___NUM_A_LEN__q0;
  assign read_A_47_A_read_addr_offset = read_A_47___edge_list_ch_47__q0;
  assign edge_list_ch_47_read_addr__din = read_A_47_A_read_addr_s_din;
  assign read_A_47_A_read_addr_s_full_n = edge_list_ch_47_read_addr__full_n;
  assign edge_list_ch_47_read_addr__write = read_A_47_A_read_addr_s_write;
  assign read_A_47_A_read_data_peek_dout = { 1'b0 , edge_list_ch_47_read_data__dout };
  assign read_A_47_A_read_data_peek_empty_n = edge_list_ch_47_read_data__empty_n;
  assign read_A_47_A_read_data_s_dout = { 1'b0 , edge_list_ch_47_read_data__dout };
  assign read_A_47_A_read_data_s_empty_n = edge_list_ch_47_read_data__empty_n;
  assign edge_list_ch_47_read_data__read = read_A_47_A_read_data_s_read;
  assign read_A_47_A_write_addr_offset = read_A_47___edge_list_ch_47__q0;
  assign edge_list_ch_47_write_addr__din = read_A_47_A_write_addr_s_din;
  assign read_A_47_A_write_addr_s_full_n = edge_list_ch_47_write_addr__full_n;
  assign edge_list_ch_47_write_addr__write = read_A_47_A_write_addr_s_write;
  assign edge_list_ch_47_write_data__din = read_A_47_A_write_data_din;
  assign read_A_47_A_write_data_full_n = edge_list_ch_47_write_data__full_n;
  assign edge_list_ch_47_write_data__write = read_A_47_A_write_data_write;
  assign read_A_47_A_write_resp_peek_dout = { 1'b0 , edge_list_ch_47_write_resp__dout };
  assign read_A_47_A_write_resp_peek_empty_n = edge_list_ch_47_write_resp__empty_n;
  assign read_A_47_A_write_resp_s_dout = { 1'b0 , edge_list_ch_47_write_resp__dout };
  assign read_A_47_A_write_resp_s_empty_n = edge_list_ch_47_write_resp__empty_n;
  assign edge_list_ch_47_write_resp__read = read_A_47_A_write_resp_s_read;
  assign read_A_47_P_N = read_A_47___P_N__q0;
  assign read_A_47_ap_clk = ap_clk;
  assign read_A_47__ap_done = read_A_47_ap_done;
  assign read_A_47__ap_idle = read_A_47_ap_idle;
  assign read_A_47__ap_ready = read_A_47_ap_ready;
  assign read_A_47_ap_rst_n = ap_rst_n;
  assign read_A_47_ap_start = read_A_47__ap_start;
  assign fifo_A_47__din = read_A_47_fifo_A_din;
  assign read_A_47_fifo_A_full_n = fifo_A_47__full_n;
  assign fifo_A_47__write = read_A_47_fifo_A_write;
  assign read_X_0_K = read_X_0___K__q0;
  assign read_X_0_P_N = read_X_0___P_N__q0;
  assign read_X_0_ap_clk = ap_clk;
  assign read_X_0__ap_done = read_X_0_ap_done;
  assign read_X_0__ap_idle = read_X_0_ap_idle;
  assign read_X_0__ap_ready = read_X_0_ap_ready;
  assign read_X_0_ap_rst_n = ap_rst_n;
  assign read_X_0_ap_start = read_X_0__ap_start;
  assign fifo_X_pe_0__din = read_X_0_fifo_X_din;
  assign read_X_0_fifo_X_full_n = fifo_X_pe_0__full_n;
  assign fifo_X_pe_0__write = read_X_0_fifo_X_write;
  assign read_X_0_vec_X_read_addr_offset = read_X_0___vec_X__q0;
  assign vec_X_read_addr__din = read_X_0_vec_X_read_addr_s_din;
  assign read_X_0_vec_X_read_addr_s_full_n = vec_X_read_addr__full_n;
  assign vec_X_read_addr__write = read_X_0_vec_X_read_addr_s_write;
  assign read_X_0_vec_X_read_data_peek_dout = { 1'b0 , vec_X_read_data__dout };
  assign read_X_0_vec_X_read_data_peek_empty_n = vec_X_read_data__empty_n;
  assign read_X_0_vec_X_read_data_s_dout = { 1'b0 , vec_X_read_data__dout };
  assign read_X_0_vec_X_read_data_s_empty_n = vec_X_read_data__empty_n;
  assign vec_X_read_data__read = read_X_0_vec_X_read_data_s_read;
  assign read_X_0_vec_X_write_addr_offset = read_X_0___vec_X__q0;
  assign vec_X_write_addr__din = read_X_0_vec_X_write_addr_s_din;
  assign read_X_0_vec_X_write_addr_s_full_n = vec_X_write_addr__full_n;
  assign vec_X_write_addr__write = read_X_0_vec_X_write_addr_s_write;
  assign vec_X_write_data__din = read_X_0_vec_X_write_data_din;
  assign read_X_0_vec_X_write_data_full_n = vec_X_write_data__full_n;
  assign vec_X_write_data__write = read_X_0_vec_X_write_data_write;
  assign read_X_0_vec_X_write_resp_peek_dout = { 1'b0 , vec_X_write_resp__dout };
  assign read_X_0_vec_X_write_resp_peek_empty_n = vec_X_write_resp__empty_n;
  assign read_X_0_vec_X_write_resp_s_dout = { 1'b0 , vec_X_write_resp__dout };
  assign read_X_0_vec_X_write_resp_s_empty_n = vec_X_write_resp__empty_n;
  assign vec_X_write_resp__read = read_X_0_vec_X_write_resp_s_read;
  assign read_Y_0_M = read_Y_0___M__q0;
  assign read_Y_0_P_N = read_Y_0___P_N__q0;
  assign read_Y_0_Y_read_addr_offset = read_Y_0___vec_Y__q0;
  assign vec_Y_read_addr__din = read_Y_0_Y_read_addr_s_din;
  assign read_Y_0_Y_read_addr_s_full_n = vec_Y_read_addr__full_n;
  assign vec_Y_read_addr__write = read_Y_0_Y_read_addr_s_write;
  assign read_Y_0_Y_read_data_peek_dout = { 1'b0 , vec_Y_read_data__dout };
  assign read_Y_0_Y_read_data_peek_empty_n = vec_Y_read_data__empty_n;
  assign read_Y_0_Y_read_data_s_dout = { 1'b0 , vec_Y_read_data__dout };
  assign read_Y_0_Y_read_data_s_empty_n = vec_Y_read_data__empty_n;
  assign vec_Y_read_data__read = read_Y_0_Y_read_data_s_read;
  assign read_Y_0_Y_write_addr_offset = read_Y_0___vec_Y__q0;
  assign vec_Y_write_addr__din = read_Y_0_Y_write_addr_s_din;
  assign read_Y_0_Y_write_addr_s_full_n = vec_Y_write_addr__full_n;
  assign vec_Y_write_addr__write = read_Y_0_Y_write_addr_s_write;
  assign vec_Y_write_data__din = read_Y_0_Y_write_data_din;
  assign read_Y_0_Y_write_data_full_n = vec_Y_write_data__full_n;
  assign vec_Y_write_data__write = read_Y_0_Y_write_data_write;
  assign read_Y_0_Y_write_resp_peek_dout = { 1'b0 , vec_Y_write_resp__dout };
  assign read_Y_0_Y_write_resp_peek_empty_n = vec_Y_write_resp__empty_n;
  assign read_Y_0_Y_write_resp_s_dout = { 1'b0 , vec_Y_write_resp__dout };
  assign read_Y_0_Y_write_resp_s_empty_n = vec_Y_write_resp__empty_n;
  assign vec_Y_write_resp__read = read_Y_0_Y_write_resp_s_read;
  assign read_Y_0_ap_clk = ap_clk;
  assign read_Y_0__ap_done = read_Y_0_ap_done;
  assign read_Y_0__ap_idle = read_Y_0_ap_idle;
  assign read_Y_0__ap_ready = read_Y_0_ap_ready;
  assign read_Y_0_ap_rst_n = ap_rst_n;
  assign read_Y_0_ap_start = read_Y_0__ap_start;
  assign fifo_Y_in__din = read_Y_0_fifo_Y_din;
  assign read_Y_0_fifo_Y_full_n = fifo_Y_in__full_n;
  assign fifo_Y_in__write = read_Y_0_fifo_Y_write;
  assign read_edge_list_ptr_0_K = read_edge_list_ptr_0___K__q0;
  assign read_edge_list_ptr_0_M = read_edge_list_ptr_0___M__q0;
  assign PE_inst_0__din = read_edge_list_ptr_0_PE_inst_din;
  assign read_edge_list_ptr_0_PE_inst_full_n = PE_inst_0__full_n;
  assign PE_inst_0__write = read_edge_list_ptr_0_PE_inst_write;
  assign read_edge_list_ptr_0_P_N = read_edge_list_ptr_0___P_N__q0;
  assign read_edge_list_ptr_0_ap_clk = ap_clk;
  assign read_edge_list_ptr_0__ap_done = read_edge_list_ptr_0_ap_done;
  assign read_edge_list_ptr_0__ap_idle = read_edge_list_ptr_0_ap_idle;
  assign read_edge_list_ptr_0__ap_ready = read_edge_list_ptr_0_ap_ready;
  assign read_edge_list_ptr_0_ap_rst_n = ap_rst_n;
  assign read_edge_list_ptr_0_ap_start = read_edge_list_ptr_0__ap_start;
  assign read_edge_list_ptr_0_edge_list_ptr_read_addr_offset = read_edge_list_ptr_0___edge_list_ptr__q0;
  assign edge_list_ptr_read_addr__din = read_edge_list_ptr_0_edge_list_ptr_read_addr_s_din;
  assign read_edge_list_ptr_0_edge_list_ptr_read_addr_s_full_n = edge_list_ptr_read_addr__full_n;
  assign edge_list_ptr_read_addr__write = read_edge_list_ptr_0_edge_list_ptr_read_addr_s_write;
  assign read_edge_list_ptr_0_edge_list_ptr_read_data_peek_dout = { 1'b0 , edge_list_ptr_read_data__dout };
  assign read_edge_list_ptr_0_edge_list_ptr_read_data_peek_empty_n = edge_list_ptr_read_data__empty_n;
  assign read_edge_list_ptr_0_edge_list_ptr_read_data_s_dout = { 1'b0 , edge_list_ptr_read_data__dout };
  assign read_edge_list_ptr_0_edge_list_ptr_read_data_s_empty_n = edge_list_ptr_read_data__empty_n;
  assign edge_list_ptr_read_data__read = read_edge_list_ptr_0_edge_list_ptr_read_data_s_read;
  assign read_edge_list_ptr_0_edge_list_ptr_write_addr_offset = read_edge_list_ptr_0___edge_list_ptr__q0;
  assign edge_list_ptr_write_addr__din = read_edge_list_ptr_0_edge_list_ptr_write_addr_s_din;
  assign read_edge_list_ptr_0_edge_list_ptr_write_addr_s_full_n = edge_list_ptr_write_addr__full_n;
  assign edge_list_ptr_write_addr__write = read_edge_list_ptr_0_edge_list_ptr_write_addr_s_write;
  assign edge_list_ptr_write_data__din = read_edge_list_ptr_0_edge_list_ptr_write_data_din;
  assign read_edge_list_ptr_0_edge_list_ptr_write_data_full_n = edge_list_ptr_write_data__full_n;
  assign edge_list_ptr_write_data__write = read_edge_list_ptr_0_edge_list_ptr_write_data_write;
  assign read_edge_list_ptr_0_edge_list_ptr_write_resp_peek_dout = { 1'b0 , edge_list_ptr_write_resp__dout };
  assign read_edge_list_ptr_0_edge_list_ptr_write_resp_peek_empty_n = edge_list_ptr_write_resp__empty_n;
  assign read_edge_list_ptr_0_edge_list_ptr_write_resp_s_dout = { 1'b0 , edge_list_ptr_write_resp__dout };
  assign read_edge_list_ptr_0_edge_list_ptr_write_resp_s_empty_n = edge_list_ptr_write_resp__empty_n;
  assign edge_list_ptr_write_resp__read = read_edge_list_ptr_0_edge_list_ptr_write_resp_s_read;
  assign read_edge_list_ptr_0_num_ite = read_edge_list_ptr_0___NUM_ITE__q0;
  assign write_Y_0_M = write_Y_0___M__q0;
  assign write_Y_0_P_N = write_Y_0___P_N__q0;
  assign write_Y_0_Y_out_read_addr_offset = write_Y_0___vec_Y_out__q0;
  assign vec_Y_out_read_addr__din = write_Y_0_Y_out_read_addr_s_din;
  assign write_Y_0_Y_out_read_addr_s_full_n = vec_Y_out_read_addr__full_n;
  assign vec_Y_out_read_addr__write = write_Y_0_Y_out_read_addr_s_write;
  assign write_Y_0_Y_out_read_data_peek_dout = { 1'b0 , vec_Y_out_read_data__dout };
  assign write_Y_0_Y_out_read_data_peek_empty_n = vec_Y_out_read_data__empty_n;
  assign write_Y_0_Y_out_read_data_s_dout = { 1'b0 , vec_Y_out_read_data__dout };
  assign write_Y_0_Y_out_read_data_s_empty_n = vec_Y_out_read_data__empty_n;
  assign vec_Y_out_read_data__read = write_Y_0_Y_out_read_data_s_read;
  assign write_Y_0_Y_out_write_addr_offset = write_Y_0___vec_Y_out__q0;
  assign vec_Y_out_write_addr__din = write_Y_0_Y_out_write_addr_s_din;
  assign write_Y_0_Y_out_write_addr_s_full_n = vec_Y_out_write_addr__full_n;
  assign vec_Y_out_write_addr__write = write_Y_0_Y_out_write_addr_s_write;
  assign vec_Y_out_write_data__din = write_Y_0_Y_out_write_data_din;
  assign write_Y_0_Y_out_write_data_full_n = vec_Y_out_write_data__full_n;
  assign vec_Y_out_write_data__write = write_Y_0_Y_out_write_data_write;
  assign write_Y_0_Y_out_write_resp_peek_dout = { 1'b0 , vec_Y_out_write_resp__dout };
  assign write_Y_0_Y_out_write_resp_peek_empty_n = vec_Y_out_write_resp__empty_n;
  assign write_Y_0_Y_out_write_resp_s_dout = { 1'b0 , vec_Y_out_write_resp__dout };
  assign write_Y_0_Y_out_write_resp_s_empty_n = vec_Y_out_write_resp__empty_n;
  assign vec_Y_out_write_resp__read = write_Y_0_Y_out_write_resp_s_read;
  assign write_Y_0_ap_clk = ap_clk;
  assign write_Y_0__ap_done = write_Y_0_ap_done;
  assign write_Y_0__ap_idle = write_Y_0_ap_idle;
  assign write_Y_0__ap_ready = write_Y_0_ap_ready;
  assign write_Y_0_ap_rst_n = ap_rst_n;
  assign write_Y_0_ap_start = write_Y_0__ap_start;
  assign write_Y_0_fifo_Y_peek_dout = fifo_Y_out__dout;
  assign write_Y_0_fifo_Y_peek_empty_n = fifo_Y_out__empty_n;
  assign write_Y_0_fifo_Y_s_dout = fifo_Y_out__dout;
  assign write_Y_0_fifo_Y_s_empty_n = fifo_Y_out__empty_n;
  assign fifo_Y_out__read = write_Y_0_fifo_Y_s_read;
  assign edge_list_ch_0__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_0_ARADDR = edge_list_ch_0__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_0_ARBURST = edge_list_ch_0__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_0_ARCACHE = edge_list_ch_0__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_0_ARID = edge_list_ch_0__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_0_ARLEN = edge_list_ch_0__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_0_ARLOCK = edge_list_ch_0__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_0_ARPROT = edge_list_ch_0__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_0_ARQOS = edge_list_ch_0__m_axi_m_axi_ARQOS;
  assign edge_list_ch_0__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_0_ARREADY;
  assign m_axi_edge_list_ch_0_ARSIZE = edge_list_ch_0__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_0_ARVALID = edge_list_ch_0__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_0_AWADDR = edge_list_ch_0__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_0_AWBURST = edge_list_ch_0__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_0_AWCACHE = edge_list_ch_0__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_0_AWID = edge_list_ch_0__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_0_AWLEN = edge_list_ch_0__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_0_AWLOCK = edge_list_ch_0__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_0_AWPROT = edge_list_ch_0__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_0_AWQOS = edge_list_ch_0__m_axi_m_axi_AWQOS;
  assign edge_list_ch_0__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_0_AWREADY;
  assign m_axi_edge_list_ch_0_AWSIZE = edge_list_ch_0__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_0_AWVALID = edge_list_ch_0__m_axi_m_axi_AWVALID;
  assign edge_list_ch_0__m_axi_m_axi_BID = m_axi_edge_list_ch_0_BID;
  assign m_axi_edge_list_ch_0_BREADY = edge_list_ch_0__m_axi_m_axi_BREADY;
  assign edge_list_ch_0__m_axi_m_axi_BRESP = m_axi_edge_list_ch_0_BRESP;
  assign edge_list_ch_0__m_axi_m_axi_BVALID = m_axi_edge_list_ch_0_BVALID;
  assign edge_list_ch_0__m_axi_m_axi_RDATA = m_axi_edge_list_ch_0_RDATA;
  assign edge_list_ch_0__m_axi_m_axi_RID = m_axi_edge_list_ch_0_RID;
  assign edge_list_ch_0__m_axi_m_axi_RLAST = m_axi_edge_list_ch_0_RLAST;
  assign m_axi_edge_list_ch_0_RREADY = edge_list_ch_0__m_axi_m_axi_RREADY;
  assign edge_list_ch_0__m_axi_m_axi_RRESP = m_axi_edge_list_ch_0_RRESP;
  assign edge_list_ch_0__m_axi_m_axi_RVALID = m_axi_edge_list_ch_0_RVALID;
  assign m_axi_edge_list_ch_0_WDATA = edge_list_ch_0__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_0_WLAST = edge_list_ch_0__m_axi_m_axi_WLAST;
  assign edge_list_ch_0__m_axi_m_axi_WREADY = m_axi_edge_list_ch_0_WREADY;
  assign m_axi_edge_list_ch_0_WSTRB = edge_list_ch_0__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_0_WVALID = edge_list_ch_0__m_axi_m_axi_WVALID;
  assign edge_list_ch_0__m_axi_read_addr_din = edge_list_ch_0_read_addr__din;
  assign edge_list_ch_0_read_addr__full_n = edge_list_ch_0__m_axi_read_addr_full_n;
  assign edge_list_ch_0__m_axi_read_addr_write = edge_list_ch_0_read_addr__write;
  assign edge_list_ch_0_read_data__dout = edge_list_ch_0__m_axi_read_data_dout;
  assign edge_list_ch_0_read_data__empty_n = edge_list_ch_0__m_axi_read_data_empty_n;
  assign edge_list_ch_0__m_axi_read_data_read = edge_list_ch_0_read_data__read;
  assign edge_list_ch_0__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_0__m_axi_write_addr_din = edge_list_ch_0_write_addr__din;
  assign edge_list_ch_0_write_addr__full_n = edge_list_ch_0__m_axi_write_addr_full_n;
  assign edge_list_ch_0__m_axi_write_addr_write = edge_list_ch_0_write_addr__write;
  assign edge_list_ch_0__m_axi_write_data_din = edge_list_ch_0_write_data__din;
  assign edge_list_ch_0_write_data__full_n = edge_list_ch_0__m_axi_write_data_full_n;
  assign edge_list_ch_0__m_axi_write_data_write = edge_list_ch_0_write_data__write;
  assign edge_list_ch_0_write_resp__dout = edge_list_ch_0__m_axi_write_resp_dout;
  assign edge_list_ch_0_write_resp__empty_n = edge_list_ch_0__m_axi_write_resp_empty_n;
  assign edge_list_ch_0__m_axi_write_resp_read = edge_list_ch_0_write_resp__read;
  assign edge_list_ch_1__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_1_ARADDR = edge_list_ch_1__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_1_ARBURST = edge_list_ch_1__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_1_ARCACHE = edge_list_ch_1__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_1_ARID = edge_list_ch_1__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_1_ARLEN = edge_list_ch_1__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_1_ARLOCK = edge_list_ch_1__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_1_ARPROT = edge_list_ch_1__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_1_ARQOS = edge_list_ch_1__m_axi_m_axi_ARQOS;
  assign edge_list_ch_1__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_1_ARREADY;
  assign m_axi_edge_list_ch_1_ARSIZE = edge_list_ch_1__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_1_ARVALID = edge_list_ch_1__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_1_AWADDR = edge_list_ch_1__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_1_AWBURST = edge_list_ch_1__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_1_AWCACHE = edge_list_ch_1__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_1_AWID = edge_list_ch_1__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_1_AWLEN = edge_list_ch_1__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_1_AWLOCK = edge_list_ch_1__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_1_AWPROT = edge_list_ch_1__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_1_AWQOS = edge_list_ch_1__m_axi_m_axi_AWQOS;
  assign edge_list_ch_1__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_1_AWREADY;
  assign m_axi_edge_list_ch_1_AWSIZE = edge_list_ch_1__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_1_AWVALID = edge_list_ch_1__m_axi_m_axi_AWVALID;
  assign edge_list_ch_1__m_axi_m_axi_BID = m_axi_edge_list_ch_1_BID;
  assign m_axi_edge_list_ch_1_BREADY = edge_list_ch_1__m_axi_m_axi_BREADY;
  assign edge_list_ch_1__m_axi_m_axi_BRESP = m_axi_edge_list_ch_1_BRESP;
  assign edge_list_ch_1__m_axi_m_axi_BVALID = m_axi_edge_list_ch_1_BVALID;
  assign edge_list_ch_1__m_axi_m_axi_RDATA = m_axi_edge_list_ch_1_RDATA;
  assign edge_list_ch_1__m_axi_m_axi_RID = m_axi_edge_list_ch_1_RID;
  assign edge_list_ch_1__m_axi_m_axi_RLAST = m_axi_edge_list_ch_1_RLAST;
  assign m_axi_edge_list_ch_1_RREADY = edge_list_ch_1__m_axi_m_axi_RREADY;
  assign edge_list_ch_1__m_axi_m_axi_RRESP = m_axi_edge_list_ch_1_RRESP;
  assign edge_list_ch_1__m_axi_m_axi_RVALID = m_axi_edge_list_ch_1_RVALID;
  assign m_axi_edge_list_ch_1_WDATA = edge_list_ch_1__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_1_WLAST = edge_list_ch_1__m_axi_m_axi_WLAST;
  assign edge_list_ch_1__m_axi_m_axi_WREADY = m_axi_edge_list_ch_1_WREADY;
  assign m_axi_edge_list_ch_1_WSTRB = edge_list_ch_1__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_1_WVALID = edge_list_ch_1__m_axi_m_axi_WVALID;
  assign edge_list_ch_1__m_axi_read_addr_din = edge_list_ch_1_read_addr__din;
  assign edge_list_ch_1_read_addr__full_n = edge_list_ch_1__m_axi_read_addr_full_n;
  assign edge_list_ch_1__m_axi_read_addr_write = edge_list_ch_1_read_addr__write;
  assign edge_list_ch_1_read_data__dout = edge_list_ch_1__m_axi_read_data_dout;
  assign edge_list_ch_1_read_data__empty_n = edge_list_ch_1__m_axi_read_data_empty_n;
  assign edge_list_ch_1__m_axi_read_data_read = edge_list_ch_1_read_data__read;
  assign edge_list_ch_1__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_1__m_axi_write_addr_din = edge_list_ch_1_write_addr__din;
  assign edge_list_ch_1_write_addr__full_n = edge_list_ch_1__m_axi_write_addr_full_n;
  assign edge_list_ch_1__m_axi_write_addr_write = edge_list_ch_1_write_addr__write;
  assign edge_list_ch_1__m_axi_write_data_din = edge_list_ch_1_write_data__din;
  assign edge_list_ch_1_write_data__full_n = edge_list_ch_1__m_axi_write_data_full_n;
  assign edge_list_ch_1__m_axi_write_data_write = edge_list_ch_1_write_data__write;
  assign edge_list_ch_1_write_resp__dout = edge_list_ch_1__m_axi_write_resp_dout;
  assign edge_list_ch_1_write_resp__empty_n = edge_list_ch_1__m_axi_write_resp_empty_n;
  assign edge_list_ch_1__m_axi_write_resp_read = edge_list_ch_1_write_resp__read;
  assign edge_list_ch_2__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_2_ARADDR = edge_list_ch_2__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_2_ARBURST = edge_list_ch_2__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_2_ARCACHE = edge_list_ch_2__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_2_ARID = edge_list_ch_2__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_2_ARLEN = edge_list_ch_2__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_2_ARLOCK = edge_list_ch_2__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_2_ARPROT = edge_list_ch_2__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_2_ARQOS = edge_list_ch_2__m_axi_m_axi_ARQOS;
  assign edge_list_ch_2__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_2_ARREADY;
  assign m_axi_edge_list_ch_2_ARSIZE = edge_list_ch_2__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_2_ARVALID = edge_list_ch_2__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_2_AWADDR = edge_list_ch_2__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_2_AWBURST = edge_list_ch_2__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_2_AWCACHE = edge_list_ch_2__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_2_AWID = edge_list_ch_2__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_2_AWLEN = edge_list_ch_2__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_2_AWLOCK = edge_list_ch_2__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_2_AWPROT = edge_list_ch_2__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_2_AWQOS = edge_list_ch_2__m_axi_m_axi_AWQOS;
  assign edge_list_ch_2__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_2_AWREADY;
  assign m_axi_edge_list_ch_2_AWSIZE = edge_list_ch_2__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_2_AWVALID = edge_list_ch_2__m_axi_m_axi_AWVALID;
  assign edge_list_ch_2__m_axi_m_axi_BID = m_axi_edge_list_ch_2_BID;
  assign m_axi_edge_list_ch_2_BREADY = edge_list_ch_2__m_axi_m_axi_BREADY;
  assign edge_list_ch_2__m_axi_m_axi_BRESP = m_axi_edge_list_ch_2_BRESP;
  assign edge_list_ch_2__m_axi_m_axi_BVALID = m_axi_edge_list_ch_2_BVALID;
  assign edge_list_ch_2__m_axi_m_axi_RDATA = m_axi_edge_list_ch_2_RDATA;
  assign edge_list_ch_2__m_axi_m_axi_RID = m_axi_edge_list_ch_2_RID;
  assign edge_list_ch_2__m_axi_m_axi_RLAST = m_axi_edge_list_ch_2_RLAST;
  assign m_axi_edge_list_ch_2_RREADY = edge_list_ch_2__m_axi_m_axi_RREADY;
  assign edge_list_ch_2__m_axi_m_axi_RRESP = m_axi_edge_list_ch_2_RRESP;
  assign edge_list_ch_2__m_axi_m_axi_RVALID = m_axi_edge_list_ch_2_RVALID;
  assign m_axi_edge_list_ch_2_WDATA = edge_list_ch_2__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_2_WLAST = edge_list_ch_2__m_axi_m_axi_WLAST;
  assign edge_list_ch_2__m_axi_m_axi_WREADY = m_axi_edge_list_ch_2_WREADY;
  assign m_axi_edge_list_ch_2_WSTRB = edge_list_ch_2__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_2_WVALID = edge_list_ch_2__m_axi_m_axi_WVALID;
  assign edge_list_ch_2__m_axi_read_addr_din = edge_list_ch_2_read_addr__din;
  assign edge_list_ch_2_read_addr__full_n = edge_list_ch_2__m_axi_read_addr_full_n;
  assign edge_list_ch_2__m_axi_read_addr_write = edge_list_ch_2_read_addr__write;
  assign edge_list_ch_2_read_data__dout = edge_list_ch_2__m_axi_read_data_dout;
  assign edge_list_ch_2_read_data__empty_n = edge_list_ch_2__m_axi_read_data_empty_n;
  assign edge_list_ch_2__m_axi_read_data_read = edge_list_ch_2_read_data__read;
  assign edge_list_ch_2__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_2__m_axi_write_addr_din = edge_list_ch_2_write_addr__din;
  assign edge_list_ch_2_write_addr__full_n = edge_list_ch_2__m_axi_write_addr_full_n;
  assign edge_list_ch_2__m_axi_write_addr_write = edge_list_ch_2_write_addr__write;
  assign edge_list_ch_2__m_axi_write_data_din = edge_list_ch_2_write_data__din;
  assign edge_list_ch_2_write_data__full_n = edge_list_ch_2__m_axi_write_data_full_n;
  assign edge_list_ch_2__m_axi_write_data_write = edge_list_ch_2_write_data__write;
  assign edge_list_ch_2_write_resp__dout = edge_list_ch_2__m_axi_write_resp_dout;
  assign edge_list_ch_2_write_resp__empty_n = edge_list_ch_2__m_axi_write_resp_empty_n;
  assign edge_list_ch_2__m_axi_write_resp_read = edge_list_ch_2_write_resp__read;
  assign edge_list_ch_3__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_3_ARADDR = edge_list_ch_3__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_3_ARBURST = edge_list_ch_3__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_3_ARCACHE = edge_list_ch_3__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_3_ARID = edge_list_ch_3__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_3_ARLEN = edge_list_ch_3__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_3_ARLOCK = edge_list_ch_3__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_3_ARPROT = edge_list_ch_3__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_3_ARQOS = edge_list_ch_3__m_axi_m_axi_ARQOS;
  assign edge_list_ch_3__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_3_ARREADY;
  assign m_axi_edge_list_ch_3_ARSIZE = edge_list_ch_3__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_3_ARVALID = edge_list_ch_3__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_3_AWADDR = edge_list_ch_3__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_3_AWBURST = edge_list_ch_3__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_3_AWCACHE = edge_list_ch_3__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_3_AWID = edge_list_ch_3__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_3_AWLEN = edge_list_ch_3__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_3_AWLOCK = edge_list_ch_3__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_3_AWPROT = edge_list_ch_3__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_3_AWQOS = edge_list_ch_3__m_axi_m_axi_AWQOS;
  assign edge_list_ch_3__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_3_AWREADY;
  assign m_axi_edge_list_ch_3_AWSIZE = edge_list_ch_3__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_3_AWVALID = edge_list_ch_3__m_axi_m_axi_AWVALID;
  assign edge_list_ch_3__m_axi_m_axi_BID = m_axi_edge_list_ch_3_BID;
  assign m_axi_edge_list_ch_3_BREADY = edge_list_ch_3__m_axi_m_axi_BREADY;
  assign edge_list_ch_3__m_axi_m_axi_BRESP = m_axi_edge_list_ch_3_BRESP;
  assign edge_list_ch_3__m_axi_m_axi_BVALID = m_axi_edge_list_ch_3_BVALID;
  assign edge_list_ch_3__m_axi_m_axi_RDATA = m_axi_edge_list_ch_3_RDATA;
  assign edge_list_ch_3__m_axi_m_axi_RID = m_axi_edge_list_ch_3_RID;
  assign edge_list_ch_3__m_axi_m_axi_RLAST = m_axi_edge_list_ch_3_RLAST;
  assign m_axi_edge_list_ch_3_RREADY = edge_list_ch_3__m_axi_m_axi_RREADY;
  assign edge_list_ch_3__m_axi_m_axi_RRESP = m_axi_edge_list_ch_3_RRESP;
  assign edge_list_ch_3__m_axi_m_axi_RVALID = m_axi_edge_list_ch_3_RVALID;
  assign m_axi_edge_list_ch_3_WDATA = edge_list_ch_3__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_3_WLAST = edge_list_ch_3__m_axi_m_axi_WLAST;
  assign edge_list_ch_3__m_axi_m_axi_WREADY = m_axi_edge_list_ch_3_WREADY;
  assign m_axi_edge_list_ch_3_WSTRB = edge_list_ch_3__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_3_WVALID = edge_list_ch_3__m_axi_m_axi_WVALID;
  assign edge_list_ch_3__m_axi_read_addr_din = edge_list_ch_3_read_addr__din;
  assign edge_list_ch_3_read_addr__full_n = edge_list_ch_3__m_axi_read_addr_full_n;
  assign edge_list_ch_3__m_axi_read_addr_write = edge_list_ch_3_read_addr__write;
  assign edge_list_ch_3_read_data__dout = edge_list_ch_3__m_axi_read_data_dout;
  assign edge_list_ch_3_read_data__empty_n = edge_list_ch_3__m_axi_read_data_empty_n;
  assign edge_list_ch_3__m_axi_read_data_read = edge_list_ch_3_read_data__read;
  assign edge_list_ch_3__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_3__m_axi_write_addr_din = edge_list_ch_3_write_addr__din;
  assign edge_list_ch_3_write_addr__full_n = edge_list_ch_3__m_axi_write_addr_full_n;
  assign edge_list_ch_3__m_axi_write_addr_write = edge_list_ch_3_write_addr__write;
  assign edge_list_ch_3__m_axi_write_data_din = edge_list_ch_3_write_data__din;
  assign edge_list_ch_3_write_data__full_n = edge_list_ch_3__m_axi_write_data_full_n;
  assign edge_list_ch_3__m_axi_write_data_write = edge_list_ch_3_write_data__write;
  assign edge_list_ch_3_write_resp__dout = edge_list_ch_3__m_axi_write_resp_dout;
  assign edge_list_ch_3_write_resp__empty_n = edge_list_ch_3__m_axi_write_resp_empty_n;
  assign edge_list_ch_3__m_axi_write_resp_read = edge_list_ch_3_write_resp__read;
  assign edge_list_ch_4__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_4_ARADDR = edge_list_ch_4__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_4_ARBURST = edge_list_ch_4__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_4_ARCACHE = edge_list_ch_4__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_4_ARID = edge_list_ch_4__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_4_ARLEN = edge_list_ch_4__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_4_ARLOCK = edge_list_ch_4__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_4_ARPROT = edge_list_ch_4__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_4_ARQOS = edge_list_ch_4__m_axi_m_axi_ARQOS;
  assign edge_list_ch_4__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_4_ARREADY;
  assign m_axi_edge_list_ch_4_ARSIZE = edge_list_ch_4__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_4_ARVALID = edge_list_ch_4__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_4_AWADDR = edge_list_ch_4__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_4_AWBURST = edge_list_ch_4__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_4_AWCACHE = edge_list_ch_4__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_4_AWID = edge_list_ch_4__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_4_AWLEN = edge_list_ch_4__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_4_AWLOCK = edge_list_ch_4__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_4_AWPROT = edge_list_ch_4__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_4_AWQOS = edge_list_ch_4__m_axi_m_axi_AWQOS;
  assign edge_list_ch_4__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_4_AWREADY;
  assign m_axi_edge_list_ch_4_AWSIZE = edge_list_ch_4__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_4_AWVALID = edge_list_ch_4__m_axi_m_axi_AWVALID;
  assign edge_list_ch_4__m_axi_m_axi_BID = m_axi_edge_list_ch_4_BID;
  assign m_axi_edge_list_ch_4_BREADY = edge_list_ch_4__m_axi_m_axi_BREADY;
  assign edge_list_ch_4__m_axi_m_axi_BRESP = m_axi_edge_list_ch_4_BRESP;
  assign edge_list_ch_4__m_axi_m_axi_BVALID = m_axi_edge_list_ch_4_BVALID;
  assign edge_list_ch_4__m_axi_m_axi_RDATA = m_axi_edge_list_ch_4_RDATA;
  assign edge_list_ch_4__m_axi_m_axi_RID = m_axi_edge_list_ch_4_RID;
  assign edge_list_ch_4__m_axi_m_axi_RLAST = m_axi_edge_list_ch_4_RLAST;
  assign m_axi_edge_list_ch_4_RREADY = edge_list_ch_4__m_axi_m_axi_RREADY;
  assign edge_list_ch_4__m_axi_m_axi_RRESP = m_axi_edge_list_ch_4_RRESP;
  assign edge_list_ch_4__m_axi_m_axi_RVALID = m_axi_edge_list_ch_4_RVALID;
  assign m_axi_edge_list_ch_4_WDATA = edge_list_ch_4__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_4_WLAST = edge_list_ch_4__m_axi_m_axi_WLAST;
  assign edge_list_ch_4__m_axi_m_axi_WREADY = m_axi_edge_list_ch_4_WREADY;
  assign m_axi_edge_list_ch_4_WSTRB = edge_list_ch_4__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_4_WVALID = edge_list_ch_4__m_axi_m_axi_WVALID;
  assign edge_list_ch_4__m_axi_read_addr_din = edge_list_ch_4_read_addr__din;
  assign edge_list_ch_4_read_addr__full_n = edge_list_ch_4__m_axi_read_addr_full_n;
  assign edge_list_ch_4__m_axi_read_addr_write = edge_list_ch_4_read_addr__write;
  assign edge_list_ch_4_read_data__dout = edge_list_ch_4__m_axi_read_data_dout;
  assign edge_list_ch_4_read_data__empty_n = edge_list_ch_4__m_axi_read_data_empty_n;
  assign edge_list_ch_4__m_axi_read_data_read = edge_list_ch_4_read_data__read;
  assign edge_list_ch_4__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_4__m_axi_write_addr_din = edge_list_ch_4_write_addr__din;
  assign edge_list_ch_4_write_addr__full_n = edge_list_ch_4__m_axi_write_addr_full_n;
  assign edge_list_ch_4__m_axi_write_addr_write = edge_list_ch_4_write_addr__write;
  assign edge_list_ch_4__m_axi_write_data_din = edge_list_ch_4_write_data__din;
  assign edge_list_ch_4_write_data__full_n = edge_list_ch_4__m_axi_write_data_full_n;
  assign edge_list_ch_4__m_axi_write_data_write = edge_list_ch_4_write_data__write;
  assign edge_list_ch_4_write_resp__dout = edge_list_ch_4__m_axi_write_resp_dout;
  assign edge_list_ch_4_write_resp__empty_n = edge_list_ch_4__m_axi_write_resp_empty_n;
  assign edge_list_ch_4__m_axi_write_resp_read = edge_list_ch_4_write_resp__read;
  assign edge_list_ch_5__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_5_ARADDR = edge_list_ch_5__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_5_ARBURST = edge_list_ch_5__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_5_ARCACHE = edge_list_ch_5__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_5_ARID = edge_list_ch_5__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_5_ARLEN = edge_list_ch_5__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_5_ARLOCK = edge_list_ch_5__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_5_ARPROT = edge_list_ch_5__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_5_ARQOS = edge_list_ch_5__m_axi_m_axi_ARQOS;
  assign edge_list_ch_5__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_5_ARREADY;
  assign m_axi_edge_list_ch_5_ARSIZE = edge_list_ch_5__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_5_ARVALID = edge_list_ch_5__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_5_AWADDR = edge_list_ch_5__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_5_AWBURST = edge_list_ch_5__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_5_AWCACHE = edge_list_ch_5__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_5_AWID = edge_list_ch_5__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_5_AWLEN = edge_list_ch_5__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_5_AWLOCK = edge_list_ch_5__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_5_AWPROT = edge_list_ch_5__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_5_AWQOS = edge_list_ch_5__m_axi_m_axi_AWQOS;
  assign edge_list_ch_5__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_5_AWREADY;
  assign m_axi_edge_list_ch_5_AWSIZE = edge_list_ch_5__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_5_AWVALID = edge_list_ch_5__m_axi_m_axi_AWVALID;
  assign edge_list_ch_5__m_axi_m_axi_BID = m_axi_edge_list_ch_5_BID;
  assign m_axi_edge_list_ch_5_BREADY = edge_list_ch_5__m_axi_m_axi_BREADY;
  assign edge_list_ch_5__m_axi_m_axi_BRESP = m_axi_edge_list_ch_5_BRESP;
  assign edge_list_ch_5__m_axi_m_axi_BVALID = m_axi_edge_list_ch_5_BVALID;
  assign edge_list_ch_5__m_axi_m_axi_RDATA = m_axi_edge_list_ch_5_RDATA;
  assign edge_list_ch_5__m_axi_m_axi_RID = m_axi_edge_list_ch_5_RID;
  assign edge_list_ch_5__m_axi_m_axi_RLAST = m_axi_edge_list_ch_5_RLAST;
  assign m_axi_edge_list_ch_5_RREADY = edge_list_ch_5__m_axi_m_axi_RREADY;
  assign edge_list_ch_5__m_axi_m_axi_RRESP = m_axi_edge_list_ch_5_RRESP;
  assign edge_list_ch_5__m_axi_m_axi_RVALID = m_axi_edge_list_ch_5_RVALID;
  assign m_axi_edge_list_ch_5_WDATA = edge_list_ch_5__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_5_WLAST = edge_list_ch_5__m_axi_m_axi_WLAST;
  assign edge_list_ch_5__m_axi_m_axi_WREADY = m_axi_edge_list_ch_5_WREADY;
  assign m_axi_edge_list_ch_5_WSTRB = edge_list_ch_5__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_5_WVALID = edge_list_ch_5__m_axi_m_axi_WVALID;
  assign edge_list_ch_5__m_axi_read_addr_din = edge_list_ch_5_read_addr__din;
  assign edge_list_ch_5_read_addr__full_n = edge_list_ch_5__m_axi_read_addr_full_n;
  assign edge_list_ch_5__m_axi_read_addr_write = edge_list_ch_5_read_addr__write;
  assign edge_list_ch_5_read_data__dout = edge_list_ch_5__m_axi_read_data_dout;
  assign edge_list_ch_5_read_data__empty_n = edge_list_ch_5__m_axi_read_data_empty_n;
  assign edge_list_ch_5__m_axi_read_data_read = edge_list_ch_5_read_data__read;
  assign edge_list_ch_5__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_5__m_axi_write_addr_din = edge_list_ch_5_write_addr__din;
  assign edge_list_ch_5_write_addr__full_n = edge_list_ch_5__m_axi_write_addr_full_n;
  assign edge_list_ch_5__m_axi_write_addr_write = edge_list_ch_5_write_addr__write;
  assign edge_list_ch_5__m_axi_write_data_din = edge_list_ch_5_write_data__din;
  assign edge_list_ch_5_write_data__full_n = edge_list_ch_5__m_axi_write_data_full_n;
  assign edge_list_ch_5__m_axi_write_data_write = edge_list_ch_5_write_data__write;
  assign edge_list_ch_5_write_resp__dout = edge_list_ch_5__m_axi_write_resp_dout;
  assign edge_list_ch_5_write_resp__empty_n = edge_list_ch_5__m_axi_write_resp_empty_n;
  assign edge_list_ch_5__m_axi_write_resp_read = edge_list_ch_5_write_resp__read;
  assign edge_list_ch_6__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_6_ARADDR = edge_list_ch_6__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_6_ARBURST = edge_list_ch_6__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_6_ARCACHE = edge_list_ch_6__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_6_ARID = edge_list_ch_6__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_6_ARLEN = edge_list_ch_6__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_6_ARLOCK = edge_list_ch_6__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_6_ARPROT = edge_list_ch_6__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_6_ARQOS = edge_list_ch_6__m_axi_m_axi_ARQOS;
  assign edge_list_ch_6__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_6_ARREADY;
  assign m_axi_edge_list_ch_6_ARSIZE = edge_list_ch_6__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_6_ARVALID = edge_list_ch_6__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_6_AWADDR = edge_list_ch_6__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_6_AWBURST = edge_list_ch_6__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_6_AWCACHE = edge_list_ch_6__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_6_AWID = edge_list_ch_6__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_6_AWLEN = edge_list_ch_6__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_6_AWLOCK = edge_list_ch_6__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_6_AWPROT = edge_list_ch_6__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_6_AWQOS = edge_list_ch_6__m_axi_m_axi_AWQOS;
  assign edge_list_ch_6__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_6_AWREADY;
  assign m_axi_edge_list_ch_6_AWSIZE = edge_list_ch_6__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_6_AWVALID = edge_list_ch_6__m_axi_m_axi_AWVALID;
  assign edge_list_ch_6__m_axi_m_axi_BID = m_axi_edge_list_ch_6_BID;
  assign m_axi_edge_list_ch_6_BREADY = edge_list_ch_6__m_axi_m_axi_BREADY;
  assign edge_list_ch_6__m_axi_m_axi_BRESP = m_axi_edge_list_ch_6_BRESP;
  assign edge_list_ch_6__m_axi_m_axi_BVALID = m_axi_edge_list_ch_6_BVALID;
  assign edge_list_ch_6__m_axi_m_axi_RDATA = m_axi_edge_list_ch_6_RDATA;
  assign edge_list_ch_6__m_axi_m_axi_RID = m_axi_edge_list_ch_6_RID;
  assign edge_list_ch_6__m_axi_m_axi_RLAST = m_axi_edge_list_ch_6_RLAST;
  assign m_axi_edge_list_ch_6_RREADY = edge_list_ch_6__m_axi_m_axi_RREADY;
  assign edge_list_ch_6__m_axi_m_axi_RRESP = m_axi_edge_list_ch_6_RRESP;
  assign edge_list_ch_6__m_axi_m_axi_RVALID = m_axi_edge_list_ch_6_RVALID;
  assign m_axi_edge_list_ch_6_WDATA = edge_list_ch_6__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_6_WLAST = edge_list_ch_6__m_axi_m_axi_WLAST;
  assign edge_list_ch_6__m_axi_m_axi_WREADY = m_axi_edge_list_ch_6_WREADY;
  assign m_axi_edge_list_ch_6_WSTRB = edge_list_ch_6__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_6_WVALID = edge_list_ch_6__m_axi_m_axi_WVALID;
  assign edge_list_ch_6__m_axi_read_addr_din = edge_list_ch_6_read_addr__din;
  assign edge_list_ch_6_read_addr__full_n = edge_list_ch_6__m_axi_read_addr_full_n;
  assign edge_list_ch_6__m_axi_read_addr_write = edge_list_ch_6_read_addr__write;
  assign edge_list_ch_6_read_data__dout = edge_list_ch_6__m_axi_read_data_dout;
  assign edge_list_ch_6_read_data__empty_n = edge_list_ch_6__m_axi_read_data_empty_n;
  assign edge_list_ch_6__m_axi_read_data_read = edge_list_ch_6_read_data__read;
  assign edge_list_ch_6__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_6__m_axi_write_addr_din = edge_list_ch_6_write_addr__din;
  assign edge_list_ch_6_write_addr__full_n = edge_list_ch_6__m_axi_write_addr_full_n;
  assign edge_list_ch_6__m_axi_write_addr_write = edge_list_ch_6_write_addr__write;
  assign edge_list_ch_6__m_axi_write_data_din = edge_list_ch_6_write_data__din;
  assign edge_list_ch_6_write_data__full_n = edge_list_ch_6__m_axi_write_data_full_n;
  assign edge_list_ch_6__m_axi_write_data_write = edge_list_ch_6_write_data__write;
  assign edge_list_ch_6_write_resp__dout = edge_list_ch_6__m_axi_write_resp_dout;
  assign edge_list_ch_6_write_resp__empty_n = edge_list_ch_6__m_axi_write_resp_empty_n;
  assign edge_list_ch_6__m_axi_write_resp_read = edge_list_ch_6_write_resp__read;
  assign edge_list_ch_7__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_7_ARADDR = edge_list_ch_7__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_7_ARBURST = edge_list_ch_7__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_7_ARCACHE = edge_list_ch_7__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_7_ARID = edge_list_ch_7__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_7_ARLEN = edge_list_ch_7__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_7_ARLOCK = edge_list_ch_7__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_7_ARPROT = edge_list_ch_7__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_7_ARQOS = edge_list_ch_7__m_axi_m_axi_ARQOS;
  assign edge_list_ch_7__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_7_ARREADY;
  assign m_axi_edge_list_ch_7_ARSIZE = edge_list_ch_7__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_7_ARVALID = edge_list_ch_7__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_7_AWADDR = edge_list_ch_7__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_7_AWBURST = edge_list_ch_7__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_7_AWCACHE = edge_list_ch_7__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_7_AWID = edge_list_ch_7__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_7_AWLEN = edge_list_ch_7__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_7_AWLOCK = edge_list_ch_7__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_7_AWPROT = edge_list_ch_7__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_7_AWQOS = edge_list_ch_7__m_axi_m_axi_AWQOS;
  assign edge_list_ch_7__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_7_AWREADY;
  assign m_axi_edge_list_ch_7_AWSIZE = edge_list_ch_7__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_7_AWVALID = edge_list_ch_7__m_axi_m_axi_AWVALID;
  assign edge_list_ch_7__m_axi_m_axi_BID = m_axi_edge_list_ch_7_BID;
  assign m_axi_edge_list_ch_7_BREADY = edge_list_ch_7__m_axi_m_axi_BREADY;
  assign edge_list_ch_7__m_axi_m_axi_BRESP = m_axi_edge_list_ch_7_BRESP;
  assign edge_list_ch_7__m_axi_m_axi_BVALID = m_axi_edge_list_ch_7_BVALID;
  assign edge_list_ch_7__m_axi_m_axi_RDATA = m_axi_edge_list_ch_7_RDATA;
  assign edge_list_ch_7__m_axi_m_axi_RID = m_axi_edge_list_ch_7_RID;
  assign edge_list_ch_7__m_axi_m_axi_RLAST = m_axi_edge_list_ch_7_RLAST;
  assign m_axi_edge_list_ch_7_RREADY = edge_list_ch_7__m_axi_m_axi_RREADY;
  assign edge_list_ch_7__m_axi_m_axi_RRESP = m_axi_edge_list_ch_7_RRESP;
  assign edge_list_ch_7__m_axi_m_axi_RVALID = m_axi_edge_list_ch_7_RVALID;
  assign m_axi_edge_list_ch_7_WDATA = edge_list_ch_7__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_7_WLAST = edge_list_ch_7__m_axi_m_axi_WLAST;
  assign edge_list_ch_7__m_axi_m_axi_WREADY = m_axi_edge_list_ch_7_WREADY;
  assign m_axi_edge_list_ch_7_WSTRB = edge_list_ch_7__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_7_WVALID = edge_list_ch_7__m_axi_m_axi_WVALID;
  assign edge_list_ch_7__m_axi_read_addr_din = edge_list_ch_7_read_addr__din;
  assign edge_list_ch_7_read_addr__full_n = edge_list_ch_7__m_axi_read_addr_full_n;
  assign edge_list_ch_7__m_axi_read_addr_write = edge_list_ch_7_read_addr__write;
  assign edge_list_ch_7_read_data__dout = edge_list_ch_7__m_axi_read_data_dout;
  assign edge_list_ch_7_read_data__empty_n = edge_list_ch_7__m_axi_read_data_empty_n;
  assign edge_list_ch_7__m_axi_read_data_read = edge_list_ch_7_read_data__read;
  assign edge_list_ch_7__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_7__m_axi_write_addr_din = edge_list_ch_7_write_addr__din;
  assign edge_list_ch_7_write_addr__full_n = edge_list_ch_7__m_axi_write_addr_full_n;
  assign edge_list_ch_7__m_axi_write_addr_write = edge_list_ch_7_write_addr__write;
  assign edge_list_ch_7__m_axi_write_data_din = edge_list_ch_7_write_data__din;
  assign edge_list_ch_7_write_data__full_n = edge_list_ch_7__m_axi_write_data_full_n;
  assign edge_list_ch_7__m_axi_write_data_write = edge_list_ch_7_write_data__write;
  assign edge_list_ch_7_write_resp__dout = edge_list_ch_7__m_axi_write_resp_dout;
  assign edge_list_ch_7_write_resp__empty_n = edge_list_ch_7__m_axi_write_resp_empty_n;
  assign edge_list_ch_7__m_axi_write_resp_read = edge_list_ch_7_write_resp__read;
  assign edge_list_ch_8__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_8_ARADDR = edge_list_ch_8__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_8_ARBURST = edge_list_ch_8__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_8_ARCACHE = edge_list_ch_8__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_8_ARID = edge_list_ch_8__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_8_ARLEN = edge_list_ch_8__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_8_ARLOCK = edge_list_ch_8__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_8_ARPROT = edge_list_ch_8__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_8_ARQOS = edge_list_ch_8__m_axi_m_axi_ARQOS;
  assign edge_list_ch_8__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_8_ARREADY;
  assign m_axi_edge_list_ch_8_ARSIZE = edge_list_ch_8__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_8_ARVALID = edge_list_ch_8__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_8_AWADDR = edge_list_ch_8__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_8_AWBURST = edge_list_ch_8__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_8_AWCACHE = edge_list_ch_8__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_8_AWID = edge_list_ch_8__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_8_AWLEN = edge_list_ch_8__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_8_AWLOCK = edge_list_ch_8__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_8_AWPROT = edge_list_ch_8__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_8_AWQOS = edge_list_ch_8__m_axi_m_axi_AWQOS;
  assign edge_list_ch_8__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_8_AWREADY;
  assign m_axi_edge_list_ch_8_AWSIZE = edge_list_ch_8__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_8_AWVALID = edge_list_ch_8__m_axi_m_axi_AWVALID;
  assign edge_list_ch_8__m_axi_m_axi_BID = m_axi_edge_list_ch_8_BID;
  assign m_axi_edge_list_ch_8_BREADY = edge_list_ch_8__m_axi_m_axi_BREADY;
  assign edge_list_ch_8__m_axi_m_axi_BRESP = m_axi_edge_list_ch_8_BRESP;
  assign edge_list_ch_8__m_axi_m_axi_BVALID = m_axi_edge_list_ch_8_BVALID;
  assign edge_list_ch_8__m_axi_m_axi_RDATA = m_axi_edge_list_ch_8_RDATA;
  assign edge_list_ch_8__m_axi_m_axi_RID = m_axi_edge_list_ch_8_RID;
  assign edge_list_ch_8__m_axi_m_axi_RLAST = m_axi_edge_list_ch_8_RLAST;
  assign m_axi_edge_list_ch_8_RREADY = edge_list_ch_8__m_axi_m_axi_RREADY;
  assign edge_list_ch_8__m_axi_m_axi_RRESP = m_axi_edge_list_ch_8_RRESP;
  assign edge_list_ch_8__m_axi_m_axi_RVALID = m_axi_edge_list_ch_8_RVALID;
  assign m_axi_edge_list_ch_8_WDATA = edge_list_ch_8__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_8_WLAST = edge_list_ch_8__m_axi_m_axi_WLAST;
  assign edge_list_ch_8__m_axi_m_axi_WREADY = m_axi_edge_list_ch_8_WREADY;
  assign m_axi_edge_list_ch_8_WSTRB = edge_list_ch_8__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_8_WVALID = edge_list_ch_8__m_axi_m_axi_WVALID;
  assign edge_list_ch_8__m_axi_read_addr_din = edge_list_ch_8_read_addr__din;
  assign edge_list_ch_8_read_addr__full_n = edge_list_ch_8__m_axi_read_addr_full_n;
  assign edge_list_ch_8__m_axi_read_addr_write = edge_list_ch_8_read_addr__write;
  assign edge_list_ch_8_read_data__dout = edge_list_ch_8__m_axi_read_data_dout;
  assign edge_list_ch_8_read_data__empty_n = edge_list_ch_8__m_axi_read_data_empty_n;
  assign edge_list_ch_8__m_axi_read_data_read = edge_list_ch_8_read_data__read;
  assign edge_list_ch_8__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_8__m_axi_write_addr_din = edge_list_ch_8_write_addr__din;
  assign edge_list_ch_8_write_addr__full_n = edge_list_ch_8__m_axi_write_addr_full_n;
  assign edge_list_ch_8__m_axi_write_addr_write = edge_list_ch_8_write_addr__write;
  assign edge_list_ch_8__m_axi_write_data_din = edge_list_ch_8_write_data__din;
  assign edge_list_ch_8_write_data__full_n = edge_list_ch_8__m_axi_write_data_full_n;
  assign edge_list_ch_8__m_axi_write_data_write = edge_list_ch_8_write_data__write;
  assign edge_list_ch_8_write_resp__dout = edge_list_ch_8__m_axi_write_resp_dout;
  assign edge_list_ch_8_write_resp__empty_n = edge_list_ch_8__m_axi_write_resp_empty_n;
  assign edge_list_ch_8__m_axi_write_resp_read = edge_list_ch_8_write_resp__read;
  assign edge_list_ch_9__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_9_ARADDR = edge_list_ch_9__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_9_ARBURST = edge_list_ch_9__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_9_ARCACHE = edge_list_ch_9__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_9_ARID = edge_list_ch_9__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_9_ARLEN = edge_list_ch_9__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_9_ARLOCK = edge_list_ch_9__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_9_ARPROT = edge_list_ch_9__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_9_ARQOS = edge_list_ch_9__m_axi_m_axi_ARQOS;
  assign edge_list_ch_9__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_9_ARREADY;
  assign m_axi_edge_list_ch_9_ARSIZE = edge_list_ch_9__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_9_ARVALID = edge_list_ch_9__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_9_AWADDR = edge_list_ch_9__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_9_AWBURST = edge_list_ch_9__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_9_AWCACHE = edge_list_ch_9__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_9_AWID = edge_list_ch_9__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_9_AWLEN = edge_list_ch_9__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_9_AWLOCK = edge_list_ch_9__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_9_AWPROT = edge_list_ch_9__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_9_AWQOS = edge_list_ch_9__m_axi_m_axi_AWQOS;
  assign edge_list_ch_9__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_9_AWREADY;
  assign m_axi_edge_list_ch_9_AWSIZE = edge_list_ch_9__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_9_AWVALID = edge_list_ch_9__m_axi_m_axi_AWVALID;
  assign edge_list_ch_9__m_axi_m_axi_BID = m_axi_edge_list_ch_9_BID;
  assign m_axi_edge_list_ch_9_BREADY = edge_list_ch_9__m_axi_m_axi_BREADY;
  assign edge_list_ch_9__m_axi_m_axi_BRESP = m_axi_edge_list_ch_9_BRESP;
  assign edge_list_ch_9__m_axi_m_axi_BVALID = m_axi_edge_list_ch_9_BVALID;
  assign edge_list_ch_9__m_axi_m_axi_RDATA = m_axi_edge_list_ch_9_RDATA;
  assign edge_list_ch_9__m_axi_m_axi_RID = m_axi_edge_list_ch_9_RID;
  assign edge_list_ch_9__m_axi_m_axi_RLAST = m_axi_edge_list_ch_9_RLAST;
  assign m_axi_edge_list_ch_9_RREADY = edge_list_ch_9__m_axi_m_axi_RREADY;
  assign edge_list_ch_9__m_axi_m_axi_RRESP = m_axi_edge_list_ch_9_RRESP;
  assign edge_list_ch_9__m_axi_m_axi_RVALID = m_axi_edge_list_ch_9_RVALID;
  assign m_axi_edge_list_ch_9_WDATA = edge_list_ch_9__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_9_WLAST = edge_list_ch_9__m_axi_m_axi_WLAST;
  assign edge_list_ch_9__m_axi_m_axi_WREADY = m_axi_edge_list_ch_9_WREADY;
  assign m_axi_edge_list_ch_9_WSTRB = edge_list_ch_9__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_9_WVALID = edge_list_ch_9__m_axi_m_axi_WVALID;
  assign edge_list_ch_9__m_axi_read_addr_din = edge_list_ch_9_read_addr__din;
  assign edge_list_ch_9_read_addr__full_n = edge_list_ch_9__m_axi_read_addr_full_n;
  assign edge_list_ch_9__m_axi_read_addr_write = edge_list_ch_9_read_addr__write;
  assign edge_list_ch_9_read_data__dout = edge_list_ch_9__m_axi_read_data_dout;
  assign edge_list_ch_9_read_data__empty_n = edge_list_ch_9__m_axi_read_data_empty_n;
  assign edge_list_ch_9__m_axi_read_data_read = edge_list_ch_9_read_data__read;
  assign edge_list_ch_9__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_9__m_axi_write_addr_din = edge_list_ch_9_write_addr__din;
  assign edge_list_ch_9_write_addr__full_n = edge_list_ch_9__m_axi_write_addr_full_n;
  assign edge_list_ch_9__m_axi_write_addr_write = edge_list_ch_9_write_addr__write;
  assign edge_list_ch_9__m_axi_write_data_din = edge_list_ch_9_write_data__din;
  assign edge_list_ch_9_write_data__full_n = edge_list_ch_9__m_axi_write_data_full_n;
  assign edge_list_ch_9__m_axi_write_data_write = edge_list_ch_9_write_data__write;
  assign edge_list_ch_9_write_resp__dout = edge_list_ch_9__m_axi_write_resp_dout;
  assign edge_list_ch_9_write_resp__empty_n = edge_list_ch_9__m_axi_write_resp_empty_n;
  assign edge_list_ch_9__m_axi_write_resp_read = edge_list_ch_9_write_resp__read;
  assign edge_list_ch_10__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_10_ARADDR = edge_list_ch_10__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_10_ARBURST = edge_list_ch_10__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_10_ARCACHE = edge_list_ch_10__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_10_ARID = edge_list_ch_10__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_10_ARLEN = edge_list_ch_10__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_10_ARLOCK = edge_list_ch_10__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_10_ARPROT = edge_list_ch_10__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_10_ARQOS = edge_list_ch_10__m_axi_m_axi_ARQOS;
  assign edge_list_ch_10__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_10_ARREADY;
  assign m_axi_edge_list_ch_10_ARSIZE = edge_list_ch_10__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_10_ARVALID = edge_list_ch_10__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_10_AWADDR = edge_list_ch_10__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_10_AWBURST = edge_list_ch_10__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_10_AWCACHE = edge_list_ch_10__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_10_AWID = edge_list_ch_10__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_10_AWLEN = edge_list_ch_10__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_10_AWLOCK = edge_list_ch_10__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_10_AWPROT = edge_list_ch_10__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_10_AWQOS = edge_list_ch_10__m_axi_m_axi_AWQOS;
  assign edge_list_ch_10__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_10_AWREADY;
  assign m_axi_edge_list_ch_10_AWSIZE = edge_list_ch_10__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_10_AWVALID = edge_list_ch_10__m_axi_m_axi_AWVALID;
  assign edge_list_ch_10__m_axi_m_axi_BID = m_axi_edge_list_ch_10_BID;
  assign m_axi_edge_list_ch_10_BREADY = edge_list_ch_10__m_axi_m_axi_BREADY;
  assign edge_list_ch_10__m_axi_m_axi_BRESP = m_axi_edge_list_ch_10_BRESP;
  assign edge_list_ch_10__m_axi_m_axi_BVALID = m_axi_edge_list_ch_10_BVALID;
  assign edge_list_ch_10__m_axi_m_axi_RDATA = m_axi_edge_list_ch_10_RDATA;
  assign edge_list_ch_10__m_axi_m_axi_RID = m_axi_edge_list_ch_10_RID;
  assign edge_list_ch_10__m_axi_m_axi_RLAST = m_axi_edge_list_ch_10_RLAST;
  assign m_axi_edge_list_ch_10_RREADY = edge_list_ch_10__m_axi_m_axi_RREADY;
  assign edge_list_ch_10__m_axi_m_axi_RRESP = m_axi_edge_list_ch_10_RRESP;
  assign edge_list_ch_10__m_axi_m_axi_RVALID = m_axi_edge_list_ch_10_RVALID;
  assign m_axi_edge_list_ch_10_WDATA = edge_list_ch_10__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_10_WLAST = edge_list_ch_10__m_axi_m_axi_WLAST;
  assign edge_list_ch_10__m_axi_m_axi_WREADY = m_axi_edge_list_ch_10_WREADY;
  assign m_axi_edge_list_ch_10_WSTRB = edge_list_ch_10__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_10_WVALID = edge_list_ch_10__m_axi_m_axi_WVALID;
  assign edge_list_ch_10__m_axi_read_addr_din = edge_list_ch_10_read_addr__din;
  assign edge_list_ch_10_read_addr__full_n = edge_list_ch_10__m_axi_read_addr_full_n;
  assign edge_list_ch_10__m_axi_read_addr_write = edge_list_ch_10_read_addr__write;
  assign edge_list_ch_10_read_data__dout = edge_list_ch_10__m_axi_read_data_dout;
  assign edge_list_ch_10_read_data__empty_n = edge_list_ch_10__m_axi_read_data_empty_n;
  assign edge_list_ch_10__m_axi_read_data_read = edge_list_ch_10_read_data__read;
  assign edge_list_ch_10__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_10__m_axi_write_addr_din = edge_list_ch_10_write_addr__din;
  assign edge_list_ch_10_write_addr__full_n = edge_list_ch_10__m_axi_write_addr_full_n;
  assign edge_list_ch_10__m_axi_write_addr_write = edge_list_ch_10_write_addr__write;
  assign edge_list_ch_10__m_axi_write_data_din = edge_list_ch_10_write_data__din;
  assign edge_list_ch_10_write_data__full_n = edge_list_ch_10__m_axi_write_data_full_n;
  assign edge_list_ch_10__m_axi_write_data_write = edge_list_ch_10_write_data__write;
  assign edge_list_ch_10_write_resp__dout = edge_list_ch_10__m_axi_write_resp_dout;
  assign edge_list_ch_10_write_resp__empty_n = edge_list_ch_10__m_axi_write_resp_empty_n;
  assign edge_list_ch_10__m_axi_write_resp_read = edge_list_ch_10_write_resp__read;
  assign edge_list_ch_11__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_11_ARADDR = edge_list_ch_11__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_11_ARBURST = edge_list_ch_11__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_11_ARCACHE = edge_list_ch_11__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_11_ARID = edge_list_ch_11__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_11_ARLEN = edge_list_ch_11__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_11_ARLOCK = edge_list_ch_11__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_11_ARPROT = edge_list_ch_11__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_11_ARQOS = edge_list_ch_11__m_axi_m_axi_ARQOS;
  assign edge_list_ch_11__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_11_ARREADY;
  assign m_axi_edge_list_ch_11_ARSIZE = edge_list_ch_11__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_11_ARVALID = edge_list_ch_11__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_11_AWADDR = edge_list_ch_11__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_11_AWBURST = edge_list_ch_11__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_11_AWCACHE = edge_list_ch_11__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_11_AWID = edge_list_ch_11__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_11_AWLEN = edge_list_ch_11__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_11_AWLOCK = edge_list_ch_11__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_11_AWPROT = edge_list_ch_11__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_11_AWQOS = edge_list_ch_11__m_axi_m_axi_AWQOS;
  assign edge_list_ch_11__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_11_AWREADY;
  assign m_axi_edge_list_ch_11_AWSIZE = edge_list_ch_11__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_11_AWVALID = edge_list_ch_11__m_axi_m_axi_AWVALID;
  assign edge_list_ch_11__m_axi_m_axi_BID = m_axi_edge_list_ch_11_BID;
  assign m_axi_edge_list_ch_11_BREADY = edge_list_ch_11__m_axi_m_axi_BREADY;
  assign edge_list_ch_11__m_axi_m_axi_BRESP = m_axi_edge_list_ch_11_BRESP;
  assign edge_list_ch_11__m_axi_m_axi_BVALID = m_axi_edge_list_ch_11_BVALID;
  assign edge_list_ch_11__m_axi_m_axi_RDATA = m_axi_edge_list_ch_11_RDATA;
  assign edge_list_ch_11__m_axi_m_axi_RID = m_axi_edge_list_ch_11_RID;
  assign edge_list_ch_11__m_axi_m_axi_RLAST = m_axi_edge_list_ch_11_RLAST;
  assign m_axi_edge_list_ch_11_RREADY = edge_list_ch_11__m_axi_m_axi_RREADY;
  assign edge_list_ch_11__m_axi_m_axi_RRESP = m_axi_edge_list_ch_11_RRESP;
  assign edge_list_ch_11__m_axi_m_axi_RVALID = m_axi_edge_list_ch_11_RVALID;
  assign m_axi_edge_list_ch_11_WDATA = edge_list_ch_11__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_11_WLAST = edge_list_ch_11__m_axi_m_axi_WLAST;
  assign edge_list_ch_11__m_axi_m_axi_WREADY = m_axi_edge_list_ch_11_WREADY;
  assign m_axi_edge_list_ch_11_WSTRB = edge_list_ch_11__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_11_WVALID = edge_list_ch_11__m_axi_m_axi_WVALID;
  assign edge_list_ch_11__m_axi_read_addr_din = edge_list_ch_11_read_addr__din;
  assign edge_list_ch_11_read_addr__full_n = edge_list_ch_11__m_axi_read_addr_full_n;
  assign edge_list_ch_11__m_axi_read_addr_write = edge_list_ch_11_read_addr__write;
  assign edge_list_ch_11_read_data__dout = edge_list_ch_11__m_axi_read_data_dout;
  assign edge_list_ch_11_read_data__empty_n = edge_list_ch_11__m_axi_read_data_empty_n;
  assign edge_list_ch_11__m_axi_read_data_read = edge_list_ch_11_read_data__read;
  assign edge_list_ch_11__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_11__m_axi_write_addr_din = edge_list_ch_11_write_addr__din;
  assign edge_list_ch_11_write_addr__full_n = edge_list_ch_11__m_axi_write_addr_full_n;
  assign edge_list_ch_11__m_axi_write_addr_write = edge_list_ch_11_write_addr__write;
  assign edge_list_ch_11__m_axi_write_data_din = edge_list_ch_11_write_data__din;
  assign edge_list_ch_11_write_data__full_n = edge_list_ch_11__m_axi_write_data_full_n;
  assign edge_list_ch_11__m_axi_write_data_write = edge_list_ch_11_write_data__write;
  assign edge_list_ch_11_write_resp__dout = edge_list_ch_11__m_axi_write_resp_dout;
  assign edge_list_ch_11_write_resp__empty_n = edge_list_ch_11__m_axi_write_resp_empty_n;
  assign edge_list_ch_11__m_axi_write_resp_read = edge_list_ch_11_write_resp__read;
  assign edge_list_ch_12__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_12_ARADDR = edge_list_ch_12__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_12_ARBURST = edge_list_ch_12__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_12_ARCACHE = edge_list_ch_12__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_12_ARID = edge_list_ch_12__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_12_ARLEN = edge_list_ch_12__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_12_ARLOCK = edge_list_ch_12__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_12_ARPROT = edge_list_ch_12__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_12_ARQOS = edge_list_ch_12__m_axi_m_axi_ARQOS;
  assign edge_list_ch_12__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_12_ARREADY;
  assign m_axi_edge_list_ch_12_ARSIZE = edge_list_ch_12__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_12_ARVALID = edge_list_ch_12__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_12_AWADDR = edge_list_ch_12__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_12_AWBURST = edge_list_ch_12__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_12_AWCACHE = edge_list_ch_12__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_12_AWID = edge_list_ch_12__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_12_AWLEN = edge_list_ch_12__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_12_AWLOCK = edge_list_ch_12__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_12_AWPROT = edge_list_ch_12__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_12_AWQOS = edge_list_ch_12__m_axi_m_axi_AWQOS;
  assign edge_list_ch_12__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_12_AWREADY;
  assign m_axi_edge_list_ch_12_AWSIZE = edge_list_ch_12__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_12_AWVALID = edge_list_ch_12__m_axi_m_axi_AWVALID;
  assign edge_list_ch_12__m_axi_m_axi_BID = m_axi_edge_list_ch_12_BID;
  assign m_axi_edge_list_ch_12_BREADY = edge_list_ch_12__m_axi_m_axi_BREADY;
  assign edge_list_ch_12__m_axi_m_axi_BRESP = m_axi_edge_list_ch_12_BRESP;
  assign edge_list_ch_12__m_axi_m_axi_BVALID = m_axi_edge_list_ch_12_BVALID;
  assign edge_list_ch_12__m_axi_m_axi_RDATA = m_axi_edge_list_ch_12_RDATA;
  assign edge_list_ch_12__m_axi_m_axi_RID = m_axi_edge_list_ch_12_RID;
  assign edge_list_ch_12__m_axi_m_axi_RLAST = m_axi_edge_list_ch_12_RLAST;
  assign m_axi_edge_list_ch_12_RREADY = edge_list_ch_12__m_axi_m_axi_RREADY;
  assign edge_list_ch_12__m_axi_m_axi_RRESP = m_axi_edge_list_ch_12_RRESP;
  assign edge_list_ch_12__m_axi_m_axi_RVALID = m_axi_edge_list_ch_12_RVALID;
  assign m_axi_edge_list_ch_12_WDATA = edge_list_ch_12__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_12_WLAST = edge_list_ch_12__m_axi_m_axi_WLAST;
  assign edge_list_ch_12__m_axi_m_axi_WREADY = m_axi_edge_list_ch_12_WREADY;
  assign m_axi_edge_list_ch_12_WSTRB = edge_list_ch_12__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_12_WVALID = edge_list_ch_12__m_axi_m_axi_WVALID;
  assign edge_list_ch_12__m_axi_read_addr_din = edge_list_ch_12_read_addr__din;
  assign edge_list_ch_12_read_addr__full_n = edge_list_ch_12__m_axi_read_addr_full_n;
  assign edge_list_ch_12__m_axi_read_addr_write = edge_list_ch_12_read_addr__write;
  assign edge_list_ch_12_read_data__dout = edge_list_ch_12__m_axi_read_data_dout;
  assign edge_list_ch_12_read_data__empty_n = edge_list_ch_12__m_axi_read_data_empty_n;
  assign edge_list_ch_12__m_axi_read_data_read = edge_list_ch_12_read_data__read;
  assign edge_list_ch_12__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_12__m_axi_write_addr_din = edge_list_ch_12_write_addr__din;
  assign edge_list_ch_12_write_addr__full_n = edge_list_ch_12__m_axi_write_addr_full_n;
  assign edge_list_ch_12__m_axi_write_addr_write = edge_list_ch_12_write_addr__write;
  assign edge_list_ch_12__m_axi_write_data_din = edge_list_ch_12_write_data__din;
  assign edge_list_ch_12_write_data__full_n = edge_list_ch_12__m_axi_write_data_full_n;
  assign edge_list_ch_12__m_axi_write_data_write = edge_list_ch_12_write_data__write;
  assign edge_list_ch_12_write_resp__dout = edge_list_ch_12__m_axi_write_resp_dout;
  assign edge_list_ch_12_write_resp__empty_n = edge_list_ch_12__m_axi_write_resp_empty_n;
  assign edge_list_ch_12__m_axi_write_resp_read = edge_list_ch_12_write_resp__read;
  assign edge_list_ch_13__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_13_ARADDR = edge_list_ch_13__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_13_ARBURST = edge_list_ch_13__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_13_ARCACHE = edge_list_ch_13__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_13_ARID = edge_list_ch_13__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_13_ARLEN = edge_list_ch_13__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_13_ARLOCK = edge_list_ch_13__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_13_ARPROT = edge_list_ch_13__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_13_ARQOS = edge_list_ch_13__m_axi_m_axi_ARQOS;
  assign edge_list_ch_13__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_13_ARREADY;
  assign m_axi_edge_list_ch_13_ARSIZE = edge_list_ch_13__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_13_ARVALID = edge_list_ch_13__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_13_AWADDR = edge_list_ch_13__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_13_AWBURST = edge_list_ch_13__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_13_AWCACHE = edge_list_ch_13__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_13_AWID = edge_list_ch_13__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_13_AWLEN = edge_list_ch_13__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_13_AWLOCK = edge_list_ch_13__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_13_AWPROT = edge_list_ch_13__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_13_AWQOS = edge_list_ch_13__m_axi_m_axi_AWQOS;
  assign edge_list_ch_13__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_13_AWREADY;
  assign m_axi_edge_list_ch_13_AWSIZE = edge_list_ch_13__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_13_AWVALID = edge_list_ch_13__m_axi_m_axi_AWVALID;
  assign edge_list_ch_13__m_axi_m_axi_BID = m_axi_edge_list_ch_13_BID;
  assign m_axi_edge_list_ch_13_BREADY = edge_list_ch_13__m_axi_m_axi_BREADY;
  assign edge_list_ch_13__m_axi_m_axi_BRESP = m_axi_edge_list_ch_13_BRESP;
  assign edge_list_ch_13__m_axi_m_axi_BVALID = m_axi_edge_list_ch_13_BVALID;
  assign edge_list_ch_13__m_axi_m_axi_RDATA = m_axi_edge_list_ch_13_RDATA;
  assign edge_list_ch_13__m_axi_m_axi_RID = m_axi_edge_list_ch_13_RID;
  assign edge_list_ch_13__m_axi_m_axi_RLAST = m_axi_edge_list_ch_13_RLAST;
  assign m_axi_edge_list_ch_13_RREADY = edge_list_ch_13__m_axi_m_axi_RREADY;
  assign edge_list_ch_13__m_axi_m_axi_RRESP = m_axi_edge_list_ch_13_RRESP;
  assign edge_list_ch_13__m_axi_m_axi_RVALID = m_axi_edge_list_ch_13_RVALID;
  assign m_axi_edge_list_ch_13_WDATA = edge_list_ch_13__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_13_WLAST = edge_list_ch_13__m_axi_m_axi_WLAST;
  assign edge_list_ch_13__m_axi_m_axi_WREADY = m_axi_edge_list_ch_13_WREADY;
  assign m_axi_edge_list_ch_13_WSTRB = edge_list_ch_13__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_13_WVALID = edge_list_ch_13__m_axi_m_axi_WVALID;
  assign edge_list_ch_13__m_axi_read_addr_din = edge_list_ch_13_read_addr__din;
  assign edge_list_ch_13_read_addr__full_n = edge_list_ch_13__m_axi_read_addr_full_n;
  assign edge_list_ch_13__m_axi_read_addr_write = edge_list_ch_13_read_addr__write;
  assign edge_list_ch_13_read_data__dout = edge_list_ch_13__m_axi_read_data_dout;
  assign edge_list_ch_13_read_data__empty_n = edge_list_ch_13__m_axi_read_data_empty_n;
  assign edge_list_ch_13__m_axi_read_data_read = edge_list_ch_13_read_data__read;
  assign edge_list_ch_13__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_13__m_axi_write_addr_din = edge_list_ch_13_write_addr__din;
  assign edge_list_ch_13_write_addr__full_n = edge_list_ch_13__m_axi_write_addr_full_n;
  assign edge_list_ch_13__m_axi_write_addr_write = edge_list_ch_13_write_addr__write;
  assign edge_list_ch_13__m_axi_write_data_din = edge_list_ch_13_write_data__din;
  assign edge_list_ch_13_write_data__full_n = edge_list_ch_13__m_axi_write_data_full_n;
  assign edge_list_ch_13__m_axi_write_data_write = edge_list_ch_13_write_data__write;
  assign edge_list_ch_13_write_resp__dout = edge_list_ch_13__m_axi_write_resp_dout;
  assign edge_list_ch_13_write_resp__empty_n = edge_list_ch_13__m_axi_write_resp_empty_n;
  assign edge_list_ch_13__m_axi_write_resp_read = edge_list_ch_13_write_resp__read;
  assign edge_list_ch_14__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_14_ARADDR = edge_list_ch_14__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_14_ARBURST = edge_list_ch_14__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_14_ARCACHE = edge_list_ch_14__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_14_ARID = edge_list_ch_14__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_14_ARLEN = edge_list_ch_14__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_14_ARLOCK = edge_list_ch_14__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_14_ARPROT = edge_list_ch_14__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_14_ARQOS = edge_list_ch_14__m_axi_m_axi_ARQOS;
  assign edge_list_ch_14__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_14_ARREADY;
  assign m_axi_edge_list_ch_14_ARSIZE = edge_list_ch_14__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_14_ARVALID = edge_list_ch_14__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_14_AWADDR = edge_list_ch_14__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_14_AWBURST = edge_list_ch_14__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_14_AWCACHE = edge_list_ch_14__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_14_AWID = edge_list_ch_14__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_14_AWLEN = edge_list_ch_14__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_14_AWLOCK = edge_list_ch_14__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_14_AWPROT = edge_list_ch_14__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_14_AWQOS = edge_list_ch_14__m_axi_m_axi_AWQOS;
  assign edge_list_ch_14__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_14_AWREADY;
  assign m_axi_edge_list_ch_14_AWSIZE = edge_list_ch_14__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_14_AWVALID = edge_list_ch_14__m_axi_m_axi_AWVALID;
  assign edge_list_ch_14__m_axi_m_axi_BID = m_axi_edge_list_ch_14_BID;
  assign m_axi_edge_list_ch_14_BREADY = edge_list_ch_14__m_axi_m_axi_BREADY;
  assign edge_list_ch_14__m_axi_m_axi_BRESP = m_axi_edge_list_ch_14_BRESP;
  assign edge_list_ch_14__m_axi_m_axi_BVALID = m_axi_edge_list_ch_14_BVALID;
  assign edge_list_ch_14__m_axi_m_axi_RDATA = m_axi_edge_list_ch_14_RDATA;
  assign edge_list_ch_14__m_axi_m_axi_RID = m_axi_edge_list_ch_14_RID;
  assign edge_list_ch_14__m_axi_m_axi_RLAST = m_axi_edge_list_ch_14_RLAST;
  assign m_axi_edge_list_ch_14_RREADY = edge_list_ch_14__m_axi_m_axi_RREADY;
  assign edge_list_ch_14__m_axi_m_axi_RRESP = m_axi_edge_list_ch_14_RRESP;
  assign edge_list_ch_14__m_axi_m_axi_RVALID = m_axi_edge_list_ch_14_RVALID;
  assign m_axi_edge_list_ch_14_WDATA = edge_list_ch_14__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_14_WLAST = edge_list_ch_14__m_axi_m_axi_WLAST;
  assign edge_list_ch_14__m_axi_m_axi_WREADY = m_axi_edge_list_ch_14_WREADY;
  assign m_axi_edge_list_ch_14_WSTRB = edge_list_ch_14__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_14_WVALID = edge_list_ch_14__m_axi_m_axi_WVALID;
  assign edge_list_ch_14__m_axi_read_addr_din = edge_list_ch_14_read_addr__din;
  assign edge_list_ch_14_read_addr__full_n = edge_list_ch_14__m_axi_read_addr_full_n;
  assign edge_list_ch_14__m_axi_read_addr_write = edge_list_ch_14_read_addr__write;
  assign edge_list_ch_14_read_data__dout = edge_list_ch_14__m_axi_read_data_dout;
  assign edge_list_ch_14_read_data__empty_n = edge_list_ch_14__m_axi_read_data_empty_n;
  assign edge_list_ch_14__m_axi_read_data_read = edge_list_ch_14_read_data__read;
  assign edge_list_ch_14__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_14__m_axi_write_addr_din = edge_list_ch_14_write_addr__din;
  assign edge_list_ch_14_write_addr__full_n = edge_list_ch_14__m_axi_write_addr_full_n;
  assign edge_list_ch_14__m_axi_write_addr_write = edge_list_ch_14_write_addr__write;
  assign edge_list_ch_14__m_axi_write_data_din = edge_list_ch_14_write_data__din;
  assign edge_list_ch_14_write_data__full_n = edge_list_ch_14__m_axi_write_data_full_n;
  assign edge_list_ch_14__m_axi_write_data_write = edge_list_ch_14_write_data__write;
  assign edge_list_ch_14_write_resp__dout = edge_list_ch_14__m_axi_write_resp_dout;
  assign edge_list_ch_14_write_resp__empty_n = edge_list_ch_14__m_axi_write_resp_empty_n;
  assign edge_list_ch_14__m_axi_write_resp_read = edge_list_ch_14_write_resp__read;
  assign edge_list_ch_15__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_15_ARADDR = edge_list_ch_15__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_15_ARBURST = edge_list_ch_15__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_15_ARCACHE = edge_list_ch_15__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_15_ARID = edge_list_ch_15__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_15_ARLEN = edge_list_ch_15__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_15_ARLOCK = edge_list_ch_15__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_15_ARPROT = edge_list_ch_15__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_15_ARQOS = edge_list_ch_15__m_axi_m_axi_ARQOS;
  assign edge_list_ch_15__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_15_ARREADY;
  assign m_axi_edge_list_ch_15_ARSIZE = edge_list_ch_15__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_15_ARVALID = edge_list_ch_15__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_15_AWADDR = edge_list_ch_15__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_15_AWBURST = edge_list_ch_15__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_15_AWCACHE = edge_list_ch_15__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_15_AWID = edge_list_ch_15__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_15_AWLEN = edge_list_ch_15__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_15_AWLOCK = edge_list_ch_15__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_15_AWPROT = edge_list_ch_15__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_15_AWQOS = edge_list_ch_15__m_axi_m_axi_AWQOS;
  assign edge_list_ch_15__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_15_AWREADY;
  assign m_axi_edge_list_ch_15_AWSIZE = edge_list_ch_15__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_15_AWVALID = edge_list_ch_15__m_axi_m_axi_AWVALID;
  assign edge_list_ch_15__m_axi_m_axi_BID = m_axi_edge_list_ch_15_BID;
  assign m_axi_edge_list_ch_15_BREADY = edge_list_ch_15__m_axi_m_axi_BREADY;
  assign edge_list_ch_15__m_axi_m_axi_BRESP = m_axi_edge_list_ch_15_BRESP;
  assign edge_list_ch_15__m_axi_m_axi_BVALID = m_axi_edge_list_ch_15_BVALID;
  assign edge_list_ch_15__m_axi_m_axi_RDATA = m_axi_edge_list_ch_15_RDATA;
  assign edge_list_ch_15__m_axi_m_axi_RID = m_axi_edge_list_ch_15_RID;
  assign edge_list_ch_15__m_axi_m_axi_RLAST = m_axi_edge_list_ch_15_RLAST;
  assign m_axi_edge_list_ch_15_RREADY = edge_list_ch_15__m_axi_m_axi_RREADY;
  assign edge_list_ch_15__m_axi_m_axi_RRESP = m_axi_edge_list_ch_15_RRESP;
  assign edge_list_ch_15__m_axi_m_axi_RVALID = m_axi_edge_list_ch_15_RVALID;
  assign m_axi_edge_list_ch_15_WDATA = edge_list_ch_15__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_15_WLAST = edge_list_ch_15__m_axi_m_axi_WLAST;
  assign edge_list_ch_15__m_axi_m_axi_WREADY = m_axi_edge_list_ch_15_WREADY;
  assign m_axi_edge_list_ch_15_WSTRB = edge_list_ch_15__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_15_WVALID = edge_list_ch_15__m_axi_m_axi_WVALID;
  assign edge_list_ch_15__m_axi_read_addr_din = edge_list_ch_15_read_addr__din;
  assign edge_list_ch_15_read_addr__full_n = edge_list_ch_15__m_axi_read_addr_full_n;
  assign edge_list_ch_15__m_axi_read_addr_write = edge_list_ch_15_read_addr__write;
  assign edge_list_ch_15_read_data__dout = edge_list_ch_15__m_axi_read_data_dout;
  assign edge_list_ch_15_read_data__empty_n = edge_list_ch_15__m_axi_read_data_empty_n;
  assign edge_list_ch_15__m_axi_read_data_read = edge_list_ch_15_read_data__read;
  assign edge_list_ch_15__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_15__m_axi_write_addr_din = edge_list_ch_15_write_addr__din;
  assign edge_list_ch_15_write_addr__full_n = edge_list_ch_15__m_axi_write_addr_full_n;
  assign edge_list_ch_15__m_axi_write_addr_write = edge_list_ch_15_write_addr__write;
  assign edge_list_ch_15__m_axi_write_data_din = edge_list_ch_15_write_data__din;
  assign edge_list_ch_15_write_data__full_n = edge_list_ch_15__m_axi_write_data_full_n;
  assign edge_list_ch_15__m_axi_write_data_write = edge_list_ch_15_write_data__write;
  assign edge_list_ch_15_write_resp__dout = edge_list_ch_15__m_axi_write_resp_dout;
  assign edge_list_ch_15_write_resp__empty_n = edge_list_ch_15__m_axi_write_resp_empty_n;
  assign edge_list_ch_15__m_axi_write_resp_read = edge_list_ch_15_write_resp__read;
  assign edge_list_ch_16__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_16_ARADDR = edge_list_ch_16__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_16_ARBURST = edge_list_ch_16__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_16_ARCACHE = edge_list_ch_16__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_16_ARID = edge_list_ch_16__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_16_ARLEN = edge_list_ch_16__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_16_ARLOCK = edge_list_ch_16__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_16_ARPROT = edge_list_ch_16__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_16_ARQOS = edge_list_ch_16__m_axi_m_axi_ARQOS;
  assign edge_list_ch_16__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_16_ARREADY;
  assign m_axi_edge_list_ch_16_ARSIZE = edge_list_ch_16__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_16_ARVALID = edge_list_ch_16__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_16_AWADDR = edge_list_ch_16__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_16_AWBURST = edge_list_ch_16__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_16_AWCACHE = edge_list_ch_16__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_16_AWID = edge_list_ch_16__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_16_AWLEN = edge_list_ch_16__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_16_AWLOCK = edge_list_ch_16__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_16_AWPROT = edge_list_ch_16__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_16_AWQOS = edge_list_ch_16__m_axi_m_axi_AWQOS;
  assign edge_list_ch_16__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_16_AWREADY;
  assign m_axi_edge_list_ch_16_AWSIZE = edge_list_ch_16__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_16_AWVALID = edge_list_ch_16__m_axi_m_axi_AWVALID;
  assign edge_list_ch_16__m_axi_m_axi_BID = m_axi_edge_list_ch_16_BID;
  assign m_axi_edge_list_ch_16_BREADY = edge_list_ch_16__m_axi_m_axi_BREADY;
  assign edge_list_ch_16__m_axi_m_axi_BRESP = m_axi_edge_list_ch_16_BRESP;
  assign edge_list_ch_16__m_axi_m_axi_BVALID = m_axi_edge_list_ch_16_BVALID;
  assign edge_list_ch_16__m_axi_m_axi_RDATA = m_axi_edge_list_ch_16_RDATA;
  assign edge_list_ch_16__m_axi_m_axi_RID = m_axi_edge_list_ch_16_RID;
  assign edge_list_ch_16__m_axi_m_axi_RLAST = m_axi_edge_list_ch_16_RLAST;
  assign m_axi_edge_list_ch_16_RREADY = edge_list_ch_16__m_axi_m_axi_RREADY;
  assign edge_list_ch_16__m_axi_m_axi_RRESP = m_axi_edge_list_ch_16_RRESP;
  assign edge_list_ch_16__m_axi_m_axi_RVALID = m_axi_edge_list_ch_16_RVALID;
  assign m_axi_edge_list_ch_16_WDATA = edge_list_ch_16__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_16_WLAST = edge_list_ch_16__m_axi_m_axi_WLAST;
  assign edge_list_ch_16__m_axi_m_axi_WREADY = m_axi_edge_list_ch_16_WREADY;
  assign m_axi_edge_list_ch_16_WSTRB = edge_list_ch_16__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_16_WVALID = edge_list_ch_16__m_axi_m_axi_WVALID;
  assign edge_list_ch_16__m_axi_read_addr_din = edge_list_ch_16_read_addr__din;
  assign edge_list_ch_16_read_addr__full_n = edge_list_ch_16__m_axi_read_addr_full_n;
  assign edge_list_ch_16__m_axi_read_addr_write = edge_list_ch_16_read_addr__write;
  assign edge_list_ch_16_read_data__dout = edge_list_ch_16__m_axi_read_data_dout;
  assign edge_list_ch_16_read_data__empty_n = edge_list_ch_16__m_axi_read_data_empty_n;
  assign edge_list_ch_16__m_axi_read_data_read = edge_list_ch_16_read_data__read;
  assign edge_list_ch_16__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_16__m_axi_write_addr_din = edge_list_ch_16_write_addr__din;
  assign edge_list_ch_16_write_addr__full_n = edge_list_ch_16__m_axi_write_addr_full_n;
  assign edge_list_ch_16__m_axi_write_addr_write = edge_list_ch_16_write_addr__write;
  assign edge_list_ch_16__m_axi_write_data_din = edge_list_ch_16_write_data__din;
  assign edge_list_ch_16_write_data__full_n = edge_list_ch_16__m_axi_write_data_full_n;
  assign edge_list_ch_16__m_axi_write_data_write = edge_list_ch_16_write_data__write;
  assign edge_list_ch_16_write_resp__dout = edge_list_ch_16__m_axi_write_resp_dout;
  assign edge_list_ch_16_write_resp__empty_n = edge_list_ch_16__m_axi_write_resp_empty_n;
  assign edge_list_ch_16__m_axi_write_resp_read = edge_list_ch_16_write_resp__read;
  assign edge_list_ch_17__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_17_ARADDR = edge_list_ch_17__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_17_ARBURST = edge_list_ch_17__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_17_ARCACHE = edge_list_ch_17__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_17_ARID = edge_list_ch_17__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_17_ARLEN = edge_list_ch_17__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_17_ARLOCK = edge_list_ch_17__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_17_ARPROT = edge_list_ch_17__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_17_ARQOS = edge_list_ch_17__m_axi_m_axi_ARQOS;
  assign edge_list_ch_17__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_17_ARREADY;
  assign m_axi_edge_list_ch_17_ARSIZE = edge_list_ch_17__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_17_ARVALID = edge_list_ch_17__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_17_AWADDR = edge_list_ch_17__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_17_AWBURST = edge_list_ch_17__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_17_AWCACHE = edge_list_ch_17__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_17_AWID = edge_list_ch_17__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_17_AWLEN = edge_list_ch_17__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_17_AWLOCK = edge_list_ch_17__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_17_AWPROT = edge_list_ch_17__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_17_AWQOS = edge_list_ch_17__m_axi_m_axi_AWQOS;
  assign edge_list_ch_17__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_17_AWREADY;
  assign m_axi_edge_list_ch_17_AWSIZE = edge_list_ch_17__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_17_AWVALID = edge_list_ch_17__m_axi_m_axi_AWVALID;
  assign edge_list_ch_17__m_axi_m_axi_BID = m_axi_edge_list_ch_17_BID;
  assign m_axi_edge_list_ch_17_BREADY = edge_list_ch_17__m_axi_m_axi_BREADY;
  assign edge_list_ch_17__m_axi_m_axi_BRESP = m_axi_edge_list_ch_17_BRESP;
  assign edge_list_ch_17__m_axi_m_axi_BVALID = m_axi_edge_list_ch_17_BVALID;
  assign edge_list_ch_17__m_axi_m_axi_RDATA = m_axi_edge_list_ch_17_RDATA;
  assign edge_list_ch_17__m_axi_m_axi_RID = m_axi_edge_list_ch_17_RID;
  assign edge_list_ch_17__m_axi_m_axi_RLAST = m_axi_edge_list_ch_17_RLAST;
  assign m_axi_edge_list_ch_17_RREADY = edge_list_ch_17__m_axi_m_axi_RREADY;
  assign edge_list_ch_17__m_axi_m_axi_RRESP = m_axi_edge_list_ch_17_RRESP;
  assign edge_list_ch_17__m_axi_m_axi_RVALID = m_axi_edge_list_ch_17_RVALID;
  assign m_axi_edge_list_ch_17_WDATA = edge_list_ch_17__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_17_WLAST = edge_list_ch_17__m_axi_m_axi_WLAST;
  assign edge_list_ch_17__m_axi_m_axi_WREADY = m_axi_edge_list_ch_17_WREADY;
  assign m_axi_edge_list_ch_17_WSTRB = edge_list_ch_17__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_17_WVALID = edge_list_ch_17__m_axi_m_axi_WVALID;
  assign edge_list_ch_17__m_axi_read_addr_din = edge_list_ch_17_read_addr__din;
  assign edge_list_ch_17_read_addr__full_n = edge_list_ch_17__m_axi_read_addr_full_n;
  assign edge_list_ch_17__m_axi_read_addr_write = edge_list_ch_17_read_addr__write;
  assign edge_list_ch_17_read_data__dout = edge_list_ch_17__m_axi_read_data_dout;
  assign edge_list_ch_17_read_data__empty_n = edge_list_ch_17__m_axi_read_data_empty_n;
  assign edge_list_ch_17__m_axi_read_data_read = edge_list_ch_17_read_data__read;
  assign edge_list_ch_17__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_17__m_axi_write_addr_din = edge_list_ch_17_write_addr__din;
  assign edge_list_ch_17_write_addr__full_n = edge_list_ch_17__m_axi_write_addr_full_n;
  assign edge_list_ch_17__m_axi_write_addr_write = edge_list_ch_17_write_addr__write;
  assign edge_list_ch_17__m_axi_write_data_din = edge_list_ch_17_write_data__din;
  assign edge_list_ch_17_write_data__full_n = edge_list_ch_17__m_axi_write_data_full_n;
  assign edge_list_ch_17__m_axi_write_data_write = edge_list_ch_17_write_data__write;
  assign edge_list_ch_17_write_resp__dout = edge_list_ch_17__m_axi_write_resp_dout;
  assign edge_list_ch_17_write_resp__empty_n = edge_list_ch_17__m_axi_write_resp_empty_n;
  assign edge_list_ch_17__m_axi_write_resp_read = edge_list_ch_17_write_resp__read;
  assign edge_list_ch_18__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_18_ARADDR = edge_list_ch_18__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_18_ARBURST = edge_list_ch_18__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_18_ARCACHE = edge_list_ch_18__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_18_ARID = edge_list_ch_18__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_18_ARLEN = edge_list_ch_18__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_18_ARLOCK = edge_list_ch_18__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_18_ARPROT = edge_list_ch_18__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_18_ARQOS = edge_list_ch_18__m_axi_m_axi_ARQOS;
  assign edge_list_ch_18__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_18_ARREADY;
  assign m_axi_edge_list_ch_18_ARSIZE = edge_list_ch_18__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_18_ARVALID = edge_list_ch_18__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_18_AWADDR = edge_list_ch_18__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_18_AWBURST = edge_list_ch_18__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_18_AWCACHE = edge_list_ch_18__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_18_AWID = edge_list_ch_18__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_18_AWLEN = edge_list_ch_18__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_18_AWLOCK = edge_list_ch_18__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_18_AWPROT = edge_list_ch_18__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_18_AWQOS = edge_list_ch_18__m_axi_m_axi_AWQOS;
  assign edge_list_ch_18__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_18_AWREADY;
  assign m_axi_edge_list_ch_18_AWSIZE = edge_list_ch_18__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_18_AWVALID = edge_list_ch_18__m_axi_m_axi_AWVALID;
  assign edge_list_ch_18__m_axi_m_axi_BID = m_axi_edge_list_ch_18_BID;
  assign m_axi_edge_list_ch_18_BREADY = edge_list_ch_18__m_axi_m_axi_BREADY;
  assign edge_list_ch_18__m_axi_m_axi_BRESP = m_axi_edge_list_ch_18_BRESP;
  assign edge_list_ch_18__m_axi_m_axi_BVALID = m_axi_edge_list_ch_18_BVALID;
  assign edge_list_ch_18__m_axi_m_axi_RDATA = m_axi_edge_list_ch_18_RDATA;
  assign edge_list_ch_18__m_axi_m_axi_RID = m_axi_edge_list_ch_18_RID;
  assign edge_list_ch_18__m_axi_m_axi_RLAST = m_axi_edge_list_ch_18_RLAST;
  assign m_axi_edge_list_ch_18_RREADY = edge_list_ch_18__m_axi_m_axi_RREADY;
  assign edge_list_ch_18__m_axi_m_axi_RRESP = m_axi_edge_list_ch_18_RRESP;
  assign edge_list_ch_18__m_axi_m_axi_RVALID = m_axi_edge_list_ch_18_RVALID;
  assign m_axi_edge_list_ch_18_WDATA = edge_list_ch_18__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_18_WLAST = edge_list_ch_18__m_axi_m_axi_WLAST;
  assign edge_list_ch_18__m_axi_m_axi_WREADY = m_axi_edge_list_ch_18_WREADY;
  assign m_axi_edge_list_ch_18_WSTRB = edge_list_ch_18__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_18_WVALID = edge_list_ch_18__m_axi_m_axi_WVALID;
  assign edge_list_ch_18__m_axi_read_addr_din = edge_list_ch_18_read_addr__din;
  assign edge_list_ch_18_read_addr__full_n = edge_list_ch_18__m_axi_read_addr_full_n;
  assign edge_list_ch_18__m_axi_read_addr_write = edge_list_ch_18_read_addr__write;
  assign edge_list_ch_18_read_data__dout = edge_list_ch_18__m_axi_read_data_dout;
  assign edge_list_ch_18_read_data__empty_n = edge_list_ch_18__m_axi_read_data_empty_n;
  assign edge_list_ch_18__m_axi_read_data_read = edge_list_ch_18_read_data__read;
  assign edge_list_ch_18__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_18__m_axi_write_addr_din = edge_list_ch_18_write_addr__din;
  assign edge_list_ch_18_write_addr__full_n = edge_list_ch_18__m_axi_write_addr_full_n;
  assign edge_list_ch_18__m_axi_write_addr_write = edge_list_ch_18_write_addr__write;
  assign edge_list_ch_18__m_axi_write_data_din = edge_list_ch_18_write_data__din;
  assign edge_list_ch_18_write_data__full_n = edge_list_ch_18__m_axi_write_data_full_n;
  assign edge_list_ch_18__m_axi_write_data_write = edge_list_ch_18_write_data__write;
  assign edge_list_ch_18_write_resp__dout = edge_list_ch_18__m_axi_write_resp_dout;
  assign edge_list_ch_18_write_resp__empty_n = edge_list_ch_18__m_axi_write_resp_empty_n;
  assign edge_list_ch_18__m_axi_write_resp_read = edge_list_ch_18_write_resp__read;
  assign edge_list_ch_19__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_19_ARADDR = edge_list_ch_19__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_19_ARBURST = edge_list_ch_19__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_19_ARCACHE = edge_list_ch_19__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_19_ARID = edge_list_ch_19__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_19_ARLEN = edge_list_ch_19__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_19_ARLOCK = edge_list_ch_19__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_19_ARPROT = edge_list_ch_19__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_19_ARQOS = edge_list_ch_19__m_axi_m_axi_ARQOS;
  assign edge_list_ch_19__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_19_ARREADY;
  assign m_axi_edge_list_ch_19_ARSIZE = edge_list_ch_19__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_19_ARVALID = edge_list_ch_19__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_19_AWADDR = edge_list_ch_19__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_19_AWBURST = edge_list_ch_19__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_19_AWCACHE = edge_list_ch_19__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_19_AWID = edge_list_ch_19__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_19_AWLEN = edge_list_ch_19__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_19_AWLOCK = edge_list_ch_19__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_19_AWPROT = edge_list_ch_19__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_19_AWQOS = edge_list_ch_19__m_axi_m_axi_AWQOS;
  assign edge_list_ch_19__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_19_AWREADY;
  assign m_axi_edge_list_ch_19_AWSIZE = edge_list_ch_19__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_19_AWVALID = edge_list_ch_19__m_axi_m_axi_AWVALID;
  assign edge_list_ch_19__m_axi_m_axi_BID = m_axi_edge_list_ch_19_BID;
  assign m_axi_edge_list_ch_19_BREADY = edge_list_ch_19__m_axi_m_axi_BREADY;
  assign edge_list_ch_19__m_axi_m_axi_BRESP = m_axi_edge_list_ch_19_BRESP;
  assign edge_list_ch_19__m_axi_m_axi_BVALID = m_axi_edge_list_ch_19_BVALID;
  assign edge_list_ch_19__m_axi_m_axi_RDATA = m_axi_edge_list_ch_19_RDATA;
  assign edge_list_ch_19__m_axi_m_axi_RID = m_axi_edge_list_ch_19_RID;
  assign edge_list_ch_19__m_axi_m_axi_RLAST = m_axi_edge_list_ch_19_RLAST;
  assign m_axi_edge_list_ch_19_RREADY = edge_list_ch_19__m_axi_m_axi_RREADY;
  assign edge_list_ch_19__m_axi_m_axi_RRESP = m_axi_edge_list_ch_19_RRESP;
  assign edge_list_ch_19__m_axi_m_axi_RVALID = m_axi_edge_list_ch_19_RVALID;
  assign m_axi_edge_list_ch_19_WDATA = edge_list_ch_19__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_19_WLAST = edge_list_ch_19__m_axi_m_axi_WLAST;
  assign edge_list_ch_19__m_axi_m_axi_WREADY = m_axi_edge_list_ch_19_WREADY;
  assign m_axi_edge_list_ch_19_WSTRB = edge_list_ch_19__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_19_WVALID = edge_list_ch_19__m_axi_m_axi_WVALID;
  assign edge_list_ch_19__m_axi_read_addr_din = edge_list_ch_19_read_addr__din;
  assign edge_list_ch_19_read_addr__full_n = edge_list_ch_19__m_axi_read_addr_full_n;
  assign edge_list_ch_19__m_axi_read_addr_write = edge_list_ch_19_read_addr__write;
  assign edge_list_ch_19_read_data__dout = edge_list_ch_19__m_axi_read_data_dout;
  assign edge_list_ch_19_read_data__empty_n = edge_list_ch_19__m_axi_read_data_empty_n;
  assign edge_list_ch_19__m_axi_read_data_read = edge_list_ch_19_read_data__read;
  assign edge_list_ch_19__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_19__m_axi_write_addr_din = edge_list_ch_19_write_addr__din;
  assign edge_list_ch_19_write_addr__full_n = edge_list_ch_19__m_axi_write_addr_full_n;
  assign edge_list_ch_19__m_axi_write_addr_write = edge_list_ch_19_write_addr__write;
  assign edge_list_ch_19__m_axi_write_data_din = edge_list_ch_19_write_data__din;
  assign edge_list_ch_19_write_data__full_n = edge_list_ch_19__m_axi_write_data_full_n;
  assign edge_list_ch_19__m_axi_write_data_write = edge_list_ch_19_write_data__write;
  assign edge_list_ch_19_write_resp__dout = edge_list_ch_19__m_axi_write_resp_dout;
  assign edge_list_ch_19_write_resp__empty_n = edge_list_ch_19__m_axi_write_resp_empty_n;
  assign edge_list_ch_19__m_axi_write_resp_read = edge_list_ch_19_write_resp__read;
  assign edge_list_ch_20__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_20_ARADDR = edge_list_ch_20__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_20_ARBURST = edge_list_ch_20__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_20_ARCACHE = edge_list_ch_20__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_20_ARID = edge_list_ch_20__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_20_ARLEN = edge_list_ch_20__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_20_ARLOCK = edge_list_ch_20__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_20_ARPROT = edge_list_ch_20__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_20_ARQOS = edge_list_ch_20__m_axi_m_axi_ARQOS;
  assign edge_list_ch_20__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_20_ARREADY;
  assign m_axi_edge_list_ch_20_ARSIZE = edge_list_ch_20__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_20_ARVALID = edge_list_ch_20__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_20_AWADDR = edge_list_ch_20__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_20_AWBURST = edge_list_ch_20__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_20_AWCACHE = edge_list_ch_20__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_20_AWID = edge_list_ch_20__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_20_AWLEN = edge_list_ch_20__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_20_AWLOCK = edge_list_ch_20__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_20_AWPROT = edge_list_ch_20__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_20_AWQOS = edge_list_ch_20__m_axi_m_axi_AWQOS;
  assign edge_list_ch_20__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_20_AWREADY;
  assign m_axi_edge_list_ch_20_AWSIZE = edge_list_ch_20__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_20_AWVALID = edge_list_ch_20__m_axi_m_axi_AWVALID;
  assign edge_list_ch_20__m_axi_m_axi_BID = m_axi_edge_list_ch_20_BID;
  assign m_axi_edge_list_ch_20_BREADY = edge_list_ch_20__m_axi_m_axi_BREADY;
  assign edge_list_ch_20__m_axi_m_axi_BRESP = m_axi_edge_list_ch_20_BRESP;
  assign edge_list_ch_20__m_axi_m_axi_BVALID = m_axi_edge_list_ch_20_BVALID;
  assign edge_list_ch_20__m_axi_m_axi_RDATA = m_axi_edge_list_ch_20_RDATA;
  assign edge_list_ch_20__m_axi_m_axi_RID = m_axi_edge_list_ch_20_RID;
  assign edge_list_ch_20__m_axi_m_axi_RLAST = m_axi_edge_list_ch_20_RLAST;
  assign m_axi_edge_list_ch_20_RREADY = edge_list_ch_20__m_axi_m_axi_RREADY;
  assign edge_list_ch_20__m_axi_m_axi_RRESP = m_axi_edge_list_ch_20_RRESP;
  assign edge_list_ch_20__m_axi_m_axi_RVALID = m_axi_edge_list_ch_20_RVALID;
  assign m_axi_edge_list_ch_20_WDATA = edge_list_ch_20__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_20_WLAST = edge_list_ch_20__m_axi_m_axi_WLAST;
  assign edge_list_ch_20__m_axi_m_axi_WREADY = m_axi_edge_list_ch_20_WREADY;
  assign m_axi_edge_list_ch_20_WSTRB = edge_list_ch_20__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_20_WVALID = edge_list_ch_20__m_axi_m_axi_WVALID;
  assign edge_list_ch_20__m_axi_read_addr_din = edge_list_ch_20_read_addr__din;
  assign edge_list_ch_20_read_addr__full_n = edge_list_ch_20__m_axi_read_addr_full_n;
  assign edge_list_ch_20__m_axi_read_addr_write = edge_list_ch_20_read_addr__write;
  assign edge_list_ch_20_read_data__dout = edge_list_ch_20__m_axi_read_data_dout;
  assign edge_list_ch_20_read_data__empty_n = edge_list_ch_20__m_axi_read_data_empty_n;
  assign edge_list_ch_20__m_axi_read_data_read = edge_list_ch_20_read_data__read;
  assign edge_list_ch_20__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_20__m_axi_write_addr_din = edge_list_ch_20_write_addr__din;
  assign edge_list_ch_20_write_addr__full_n = edge_list_ch_20__m_axi_write_addr_full_n;
  assign edge_list_ch_20__m_axi_write_addr_write = edge_list_ch_20_write_addr__write;
  assign edge_list_ch_20__m_axi_write_data_din = edge_list_ch_20_write_data__din;
  assign edge_list_ch_20_write_data__full_n = edge_list_ch_20__m_axi_write_data_full_n;
  assign edge_list_ch_20__m_axi_write_data_write = edge_list_ch_20_write_data__write;
  assign edge_list_ch_20_write_resp__dout = edge_list_ch_20__m_axi_write_resp_dout;
  assign edge_list_ch_20_write_resp__empty_n = edge_list_ch_20__m_axi_write_resp_empty_n;
  assign edge_list_ch_20__m_axi_write_resp_read = edge_list_ch_20_write_resp__read;
  assign edge_list_ch_21__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_21_ARADDR = edge_list_ch_21__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_21_ARBURST = edge_list_ch_21__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_21_ARCACHE = edge_list_ch_21__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_21_ARID = edge_list_ch_21__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_21_ARLEN = edge_list_ch_21__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_21_ARLOCK = edge_list_ch_21__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_21_ARPROT = edge_list_ch_21__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_21_ARQOS = edge_list_ch_21__m_axi_m_axi_ARQOS;
  assign edge_list_ch_21__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_21_ARREADY;
  assign m_axi_edge_list_ch_21_ARSIZE = edge_list_ch_21__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_21_ARVALID = edge_list_ch_21__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_21_AWADDR = edge_list_ch_21__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_21_AWBURST = edge_list_ch_21__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_21_AWCACHE = edge_list_ch_21__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_21_AWID = edge_list_ch_21__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_21_AWLEN = edge_list_ch_21__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_21_AWLOCK = edge_list_ch_21__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_21_AWPROT = edge_list_ch_21__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_21_AWQOS = edge_list_ch_21__m_axi_m_axi_AWQOS;
  assign edge_list_ch_21__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_21_AWREADY;
  assign m_axi_edge_list_ch_21_AWSIZE = edge_list_ch_21__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_21_AWVALID = edge_list_ch_21__m_axi_m_axi_AWVALID;
  assign edge_list_ch_21__m_axi_m_axi_BID = m_axi_edge_list_ch_21_BID;
  assign m_axi_edge_list_ch_21_BREADY = edge_list_ch_21__m_axi_m_axi_BREADY;
  assign edge_list_ch_21__m_axi_m_axi_BRESP = m_axi_edge_list_ch_21_BRESP;
  assign edge_list_ch_21__m_axi_m_axi_BVALID = m_axi_edge_list_ch_21_BVALID;
  assign edge_list_ch_21__m_axi_m_axi_RDATA = m_axi_edge_list_ch_21_RDATA;
  assign edge_list_ch_21__m_axi_m_axi_RID = m_axi_edge_list_ch_21_RID;
  assign edge_list_ch_21__m_axi_m_axi_RLAST = m_axi_edge_list_ch_21_RLAST;
  assign m_axi_edge_list_ch_21_RREADY = edge_list_ch_21__m_axi_m_axi_RREADY;
  assign edge_list_ch_21__m_axi_m_axi_RRESP = m_axi_edge_list_ch_21_RRESP;
  assign edge_list_ch_21__m_axi_m_axi_RVALID = m_axi_edge_list_ch_21_RVALID;
  assign m_axi_edge_list_ch_21_WDATA = edge_list_ch_21__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_21_WLAST = edge_list_ch_21__m_axi_m_axi_WLAST;
  assign edge_list_ch_21__m_axi_m_axi_WREADY = m_axi_edge_list_ch_21_WREADY;
  assign m_axi_edge_list_ch_21_WSTRB = edge_list_ch_21__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_21_WVALID = edge_list_ch_21__m_axi_m_axi_WVALID;
  assign edge_list_ch_21__m_axi_read_addr_din = edge_list_ch_21_read_addr__din;
  assign edge_list_ch_21_read_addr__full_n = edge_list_ch_21__m_axi_read_addr_full_n;
  assign edge_list_ch_21__m_axi_read_addr_write = edge_list_ch_21_read_addr__write;
  assign edge_list_ch_21_read_data__dout = edge_list_ch_21__m_axi_read_data_dout;
  assign edge_list_ch_21_read_data__empty_n = edge_list_ch_21__m_axi_read_data_empty_n;
  assign edge_list_ch_21__m_axi_read_data_read = edge_list_ch_21_read_data__read;
  assign edge_list_ch_21__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_21__m_axi_write_addr_din = edge_list_ch_21_write_addr__din;
  assign edge_list_ch_21_write_addr__full_n = edge_list_ch_21__m_axi_write_addr_full_n;
  assign edge_list_ch_21__m_axi_write_addr_write = edge_list_ch_21_write_addr__write;
  assign edge_list_ch_21__m_axi_write_data_din = edge_list_ch_21_write_data__din;
  assign edge_list_ch_21_write_data__full_n = edge_list_ch_21__m_axi_write_data_full_n;
  assign edge_list_ch_21__m_axi_write_data_write = edge_list_ch_21_write_data__write;
  assign edge_list_ch_21_write_resp__dout = edge_list_ch_21__m_axi_write_resp_dout;
  assign edge_list_ch_21_write_resp__empty_n = edge_list_ch_21__m_axi_write_resp_empty_n;
  assign edge_list_ch_21__m_axi_write_resp_read = edge_list_ch_21_write_resp__read;
  assign edge_list_ch_22__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_22_ARADDR = edge_list_ch_22__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_22_ARBURST = edge_list_ch_22__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_22_ARCACHE = edge_list_ch_22__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_22_ARID = edge_list_ch_22__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_22_ARLEN = edge_list_ch_22__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_22_ARLOCK = edge_list_ch_22__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_22_ARPROT = edge_list_ch_22__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_22_ARQOS = edge_list_ch_22__m_axi_m_axi_ARQOS;
  assign edge_list_ch_22__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_22_ARREADY;
  assign m_axi_edge_list_ch_22_ARSIZE = edge_list_ch_22__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_22_ARVALID = edge_list_ch_22__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_22_AWADDR = edge_list_ch_22__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_22_AWBURST = edge_list_ch_22__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_22_AWCACHE = edge_list_ch_22__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_22_AWID = edge_list_ch_22__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_22_AWLEN = edge_list_ch_22__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_22_AWLOCK = edge_list_ch_22__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_22_AWPROT = edge_list_ch_22__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_22_AWQOS = edge_list_ch_22__m_axi_m_axi_AWQOS;
  assign edge_list_ch_22__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_22_AWREADY;
  assign m_axi_edge_list_ch_22_AWSIZE = edge_list_ch_22__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_22_AWVALID = edge_list_ch_22__m_axi_m_axi_AWVALID;
  assign edge_list_ch_22__m_axi_m_axi_BID = m_axi_edge_list_ch_22_BID;
  assign m_axi_edge_list_ch_22_BREADY = edge_list_ch_22__m_axi_m_axi_BREADY;
  assign edge_list_ch_22__m_axi_m_axi_BRESP = m_axi_edge_list_ch_22_BRESP;
  assign edge_list_ch_22__m_axi_m_axi_BVALID = m_axi_edge_list_ch_22_BVALID;
  assign edge_list_ch_22__m_axi_m_axi_RDATA = m_axi_edge_list_ch_22_RDATA;
  assign edge_list_ch_22__m_axi_m_axi_RID = m_axi_edge_list_ch_22_RID;
  assign edge_list_ch_22__m_axi_m_axi_RLAST = m_axi_edge_list_ch_22_RLAST;
  assign m_axi_edge_list_ch_22_RREADY = edge_list_ch_22__m_axi_m_axi_RREADY;
  assign edge_list_ch_22__m_axi_m_axi_RRESP = m_axi_edge_list_ch_22_RRESP;
  assign edge_list_ch_22__m_axi_m_axi_RVALID = m_axi_edge_list_ch_22_RVALID;
  assign m_axi_edge_list_ch_22_WDATA = edge_list_ch_22__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_22_WLAST = edge_list_ch_22__m_axi_m_axi_WLAST;
  assign edge_list_ch_22__m_axi_m_axi_WREADY = m_axi_edge_list_ch_22_WREADY;
  assign m_axi_edge_list_ch_22_WSTRB = edge_list_ch_22__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_22_WVALID = edge_list_ch_22__m_axi_m_axi_WVALID;
  assign edge_list_ch_22__m_axi_read_addr_din = edge_list_ch_22_read_addr__din;
  assign edge_list_ch_22_read_addr__full_n = edge_list_ch_22__m_axi_read_addr_full_n;
  assign edge_list_ch_22__m_axi_read_addr_write = edge_list_ch_22_read_addr__write;
  assign edge_list_ch_22_read_data__dout = edge_list_ch_22__m_axi_read_data_dout;
  assign edge_list_ch_22_read_data__empty_n = edge_list_ch_22__m_axi_read_data_empty_n;
  assign edge_list_ch_22__m_axi_read_data_read = edge_list_ch_22_read_data__read;
  assign edge_list_ch_22__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_22__m_axi_write_addr_din = edge_list_ch_22_write_addr__din;
  assign edge_list_ch_22_write_addr__full_n = edge_list_ch_22__m_axi_write_addr_full_n;
  assign edge_list_ch_22__m_axi_write_addr_write = edge_list_ch_22_write_addr__write;
  assign edge_list_ch_22__m_axi_write_data_din = edge_list_ch_22_write_data__din;
  assign edge_list_ch_22_write_data__full_n = edge_list_ch_22__m_axi_write_data_full_n;
  assign edge_list_ch_22__m_axi_write_data_write = edge_list_ch_22_write_data__write;
  assign edge_list_ch_22_write_resp__dout = edge_list_ch_22__m_axi_write_resp_dout;
  assign edge_list_ch_22_write_resp__empty_n = edge_list_ch_22__m_axi_write_resp_empty_n;
  assign edge_list_ch_22__m_axi_write_resp_read = edge_list_ch_22_write_resp__read;
  assign edge_list_ch_23__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_23_ARADDR = edge_list_ch_23__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_23_ARBURST = edge_list_ch_23__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_23_ARCACHE = edge_list_ch_23__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_23_ARID = edge_list_ch_23__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_23_ARLEN = edge_list_ch_23__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_23_ARLOCK = edge_list_ch_23__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_23_ARPROT = edge_list_ch_23__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_23_ARQOS = edge_list_ch_23__m_axi_m_axi_ARQOS;
  assign edge_list_ch_23__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_23_ARREADY;
  assign m_axi_edge_list_ch_23_ARSIZE = edge_list_ch_23__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_23_ARVALID = edge_list_ch_23__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_23_AWADDR = edge_list_ch_23__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_23_AWBURST = edge_list_ch_23__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_23_AWCACHE = edge_list_ch_23__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_23_AWID = edge_list_ch_23__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_23_AWLEN = edge_list_ch_23__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_23_AWLOCK = edge_list_ch_23__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_23_AWPROT = edge_list_ch_23__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_23_AWQOS = edge_list_ch_23__m_axi_m_axi_AWQOS;
  assign edge_list_ch_23__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_23_AWREADY;
  assign m_axi_edge_list_ch_23_AWSIZE = edge_list_ch_23__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_23_AWVALID = edge_list_ch_23__m_axi_m_axi_AWVALID;
  assign edge_list_ch_23__m_axi_m_axi_BID = m_axi_edge_list_ch_23_BID;
  assign m_axi_edge_list_ch_23_BREADY = edge_list_ch_23__m_axi_m_axi_BREADY;
  assign edge_list_ch_23__m_axi_m_axi_BRESP = m_axi_edge_list_ch_23_BRESP;
  assign edge_list_ch_23__m_axi_m_axi_BVALID = m_axi_edge_list_ch_23_BVALID;
  assign edge_list_ch_23__m_axi_m_axi_RDATA = m_axi_edge_list_ch_23_RDATA;
  assign edge_list_ch_23__m_axi_m_axi_RID = m_axi_edge_list_ch_23_RID;
  assign edge_list_ch_23__m_axi_m_axi_RLAST = m_axi_edge_list_ch_23_RLAST;
  assign m_axi_edge_list_ch_23_RREADY = edge_list_ch_23__m_axi_m_axi_RREADY;
  assign edge_list_ch_23__m_axi_m_axi_RRESP = m_axi_edge_list_ch_23_RRESP;
  assign edge_list_ch_23__m_axi_m_axi_RVALID = m_axi_edge_list_ch_23_RVALID;
  assign m_axi_edge_list_ch_23_WDATA = edge_list_ch_23__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_23_WLAST = edge_list_ch_23__m_axi_m_axi_WLAST;
  assign edge_list_ch_23__m_axi_m_axi_WREADY = m_axi_edge_list_ch_23_WREADY;
  assign m_axi_edge_list_ch_23_WSTRB = edge_list_ch_23__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_23_WVALID = edge_list_ch_23__m_axi_m_axi_WVALID;
  assign edge_list_ch_23__m_axi_read_addr_din = edge_list_ch_23_read_addr__din;
  assign edge_list_ch_23_read_addr__full_n = edge_list_ch_23__m_axi_read_addr_full_n;
  assign edge_list_ch_23__m_axi_read_addr_write = edge_list_ch_23_read_addr__write;
  assign edge_list_ch_23_read_data__dout = edge_list_ch_23__m_axi_read_data_dout;
  assign edge_list_ch_23_read_data__empty_n = edge_list_ch_23__m_axi_read_data_empty_n;
  assign edge_list_ch_23__m_axi_read_data_read = edge_list_ch_23_read_data__read;
  assign edge_list_ch_23__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_23__m_axi_write_addr_din = edge_list_ch_23_write_addr__din;
  assign edge_list_ch_23_write_addr__full_n = edge_list_ch_23__m_axi_write_addr_full_n;
  assign edge_list_ch_23__m_axi_write_addr_write = edge_list_ch_23_write_addr__write;
  assign edge_list_ch_23__m_axi_write_data_din = edge_list_ch_23_write_data__din;
  assign edge_list_ch_23_write_data__full_n = edge_list_ch_23__m_axi_write_data_full_n;
  assign edge_list_ch_23__m_axi_write_data_write = edge_list_ch_23_write_data__write;
  assign edge_list_ch_23_write_resp__dout = edge_list_ch_23__m_axi_write_resp_dout;
  assign edge_list_ch_23_write_resp__empty_n = edge_list_ch_23__m_axi_write_resp_empty_n;
  assign edge_list_ch_23__m_axi_write_resp_read = edge_list_ch_23_write_resp__read;
  assign edge_list_ch_24__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_24_ARADDR = edge_list_ch_24__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_24_ARBURST = edge_list_ch_24__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_24_ARCACHE = edge_list_ch_24__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_24_ARID = edge_list_ch_24__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_24_ARLEN = edge_list_ch_24__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_24_ARLOCK = edge_list_ch_24__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_24_ARPROT = edge_list_ch_24__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_24_ARQOS = edge_list_ch_24__m_axi_m_axi_ARQOS;
  assign edge_list_ch_24__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_24_ARREADY;
  assign m_axi_edge_list_ch_24_ARSIZE = edge_list_ch_24__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_24_ARVALID = edge_list_ch_24__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_24_AWADDR = edge_list_ch_24__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_24_AWBURST = edge_list_ch_24__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_24_AWCACHE = edge_list_ch_24__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_24_AWID = edge_list_ch_24__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_24_AWLEN = edge_list_ch_24__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_24_AWLOCK = edge_list_ch_24__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_24_AWPROT = edge_list_ch_24__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_24_AWQOS = edge_list_ch_24__m_axi_m_axi_AWQOS;
  assign edge_list_ch_24__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_24_AWREADY;
  assign m_axi_edge_list_ch_24_AWSIZE = edge_list_ch_24__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_24_AWVALID = edge_list_ch_24__m_axi_m_axi_AWVALID;
  assign edge_list_ch_24__m_axi_m_axi_BID = m_axi_edge_list_ch_24_BID;
  assign m_axi_edge_list_ch_24_BREADY = edge_list_ch_24__m_axi_m_axi_BREADY;
  assign edge_list_ch_24__m_axi_m_axi_BRESP = m_axi_edge_list_ch_24_BRESP;
  assign edge_list_ch_24__m_axi_m_axi_BVALID = m_axi_edge_list_ch_24_BVALID;
  assign edge_list_ch_24__m_axi_m_axi_RDATA = m_axi_edge_list_ch_24_RDATA;
  assign edge_list_ch_24__m_axi_m_axi_RID = m_axi_edge_list_ch_24_RID;
  assign edge_list_ch_24__m_axi_m_axi_RLAST = m_axi_edge_list_ch_24_RLAST;
  assign m_axi_edge_list_ch_24_RREADY = edge_list_ch_24__m_axi_m_axi_RREADY;
  assign edge_list_ch_24__m_axi_m_axi_RRESP = m_axi_edge_list_ch_24_RRESP;
  assign edge_list_ch_24__m_axi_m_axi_RVALID = m_axi_edge_list_ch_24_RVALID;
  assign m_axi_edge_list_ch_24_WDATA = edge_list_ch_24__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_24_WLAST = edge_list_ch_24__m_axi_m_axi_WLAST;
  assign edge_list_ch_24__m_axi_m_axi_WREADY = m_axi_edge_list_ch_24_WREADY;
  assign m_axi_edge_list_ch_24_WSTRB = edge_list_ch_24__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_24_WVALID = edge_list_ch_24__m_axi_m_axi_WVALID;
  assign edge_list_ch_24__m_axi_read_addr_din = edge_list_ch_24_read_addr__din;
  assign edge_list_ch_24_read_addr__full_n = edge_list_ch_24__m_axi_read_addr_full_n;
  assign edge_list_ch_24__m_axi_read_addr_write = edge_list_ch_24_read_addr__write;
  assign edge_list_ch_24_read_data__dout = edge_list_ch_24__m_axi_read_data_dout;
  assign edge_list_ch_24_read_data__empty_n = edge_list_ch_24__m_axi_read_data_empty_n;
  assign edge_list_ch_24__m_axi_read_data_read = edge_list_ch_24_read_data__read;
  assign edge_list_ch_24__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_24__m_axi_write_addr_din = edge_list_ch_24_write_addr__din;
  assign edge_list_ch_24_write_addr__full_n = edge_list_ch_24__m_axi_write_addr_full_n;
  assign edge_list_ch_24__m_axi_write_addr_write = edge_list_ch_24_write_addr__write;
  assign edge_list_ch_24__m_axi_write_data_din = edge_list_ch_24_write_data__din;
  assign edge_list_ch_24_write_data__full_n = edge_list_ch_24__m_axi_write_data_full_n;
  assign edge_list_ch_24__m_axi_write_data_write = edge_list_ch_24_write_data__write;
  assign edge_list_ch_24_write_resp__dout = edge_list_ch_24__m_axi_write_resp_dout;
  assign edge_list_ch_24_write_resp__empty_n = edge_list_ch_24__m_axi_write_resp_empty_n;
  assign edge_list_ch_24__m_axi_write_resp_read = edge_list_ch_24_write_resp__read;
  assign edge_list_ch_25__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_25_ARADDR = edge_list_ch_25__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_25_ARBURST = edge_list_ch_25__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_25_ARCACHE = edge_list_ch_25__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_25_ARID = edge_list_ch_25__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_25_ARLEN = edge_list_ch_25__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_25_ARLOCK = edge_list_ch_25__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_25_ARPROT = edge_list_ch_25__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_25_ARQOS = edge_list_ch_25__m_axi_m_axi_ARQOS;
  assign edge_list_ch_25__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_25_ARREADY;
  assign m_axi_edge_list_ch_25_ARSIZE = edge_list_ch_25__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_25_ARVALID = edge_list_ch_25__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_25_AWADDR = edge_list_ch_25__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_25_AWBURST = edge_list_ch_25__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_25_AWCACHE = edge_list_ch_25__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_25_AWID = edge_list_ch_25__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_25_AWLEN = edge_list_ch_25__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_25_AWLOCK = edge_list_ch_25__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_25_AWPROT = edge_list_ch_25__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_25_AWQOS = edge_list_ch_25__m_axi_m_axi_AWQOS;
  assign edge_list_ch_25__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_25_AWREADY;
  assign m_axi_edge_list_ch_25_AWSIZE = edge_list_ch_25__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_25_AWVALID = edge_list_ch_25__m_axi_m_axi_AWVALID;
  assign edge_list_ch_25__m_axi_m_axi_BID = m_axi_edge_list_ch_25_BID;
  assign m_axi_edge_list_ch_25_BREADY = edge_list_ch_25__m_axi_m_axi_BREADY;
  assign edge_list_ch_25__m_axi_m_axi_BRESP = m_axi_edge_list_ch_25_BRESP;
  assign edge_list_ch_25__m_axi_m_axi_BVALID = m_axi_edge_list_ch_25_BVALID;
  assign edge_list_ch_25__m_axi_m_axi_RDATA = m_axi_edge_list_ch_25_RDATA;
  assign edge_list_ch_25__m_axi_m_axi_RID = m_axi_edge_list_ch_25_RID;
  assign edge_list_ch_25__m_axi_m_axi_RLAST = m_axi_edge_list_ch_25_RLAST;
  assign m_axi_edge_list_ch_25_RREADY = edge_list_ch_25__m_axi_m_axi_RREADY;
  assign edge_list_ch_25__m_axi_m_axi_RRESP = m_axi_edge_list_ch_25_RRESP;
  assign edge_list_ch_25__m_axi_m_axi_RVALID = m_axi_edge_list_ch_25_RVALID;
  assign m_axi_edge_list_ch_25_WDATA = edge_list_ch_25__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_25_WLAST = edge_list_ch_25__m_axi_m_axi_WLAST;
  assign edge_list_ch_25__m_axi_m_axi_WREADY = m_axi_edge_list_ch_25_WREADY;
  assign m_axi_edge_list_ch_25_WSTRB = edge_list_ch_25__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_25_WVALID = edge_list_ch_25__m_axi_m_axi_WVALID;
  assign edge_list_ch_25__m_axi_read_addr_din = edge_list_ch_25_read_addr__din;
  assign edge_list_ch_25_read_addr__full_n = edge_list_ch_25__m_axi_read_addr_full_n;
  assign edge_list_ch_25__m_axi_read_addr_write = edge_list_ch_25_read_addr__write;
  assign edge_list_ch_25_read_data__dout = edge_list_ch_25__m_axi_read_data_dout;
  assign edge_list_ch_25_read_data__empty_n = edge_list_ch_25__m_axi_read_data_empty_n;
  assign edge_list_ch_25__m_axi_read_data_read = edge_list_ch_25_read_data__read;
  assign edge_list_ch_25__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_25__m_axi_write_addr_din = edge_list_ch_25_write_addr__din;
  assign edge_list_ch_25_write_addr__full_n = edge_list_ch_25__m_axi_write_addr_full_n;
  assign edge_list_ch_25__m_axi_write_addr_write = edge_list_ch_25_write_addr__write;
  assign edge_list_ch_25__m_axi_write_data_din = edge_list_ch_25_write_data__din;
  assign edge_list_ch_25_write_data__full_n = edge_list_ch_25__m_axi_write_data_full_n;
  assign edge_list_ch_25__m_axi_write_data_write = edge_list_ch_25_write_data__write;
  assign edge_list_ch_25_write_resp__dout = edge_list_ch_25__m_axi_write_resp_dout;
  assign edge_list_ch_25_write_resp__empty_n = edge_list_ch_25__m_axi_write_resp_empty_n;
  assign edge_list_ch_25__m_axi_write_resp_read = edge_list_ch_25_write_resp__read;
  assign edge_list_ch_26__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_26_ARADDR = edge_list_ch_26__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_26_ARBURST = edge_list_ch_26__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_26_ARCACHE = edge_list_ch_26__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_26_ARID = edge_list_ch_26__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_26_ARLEN = edge_list_ch_26__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_26_ARLOCK = edge_list_ch_26__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_26_ARPROT = edge_list_ch_26__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_26_ARQOS = edge_list_ch_26__m_axi_m_axi_ARQOS;
  assign edge_list_ch_26__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_26_ARREADY;
  assign m_axi_edge_list_ch_26_ARSIZE = edge_list_ch_26__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_26_ARVALID = edge_list_ch_26__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_26_AWADDR = edge_list_ch_26__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_26_AWBURST = edge_list_ch_26__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_26_AWCACHE = edge_list_ch_26__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_26_AWID = edge_list_ch_26__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_26_AWLEN = edge_list_ch_26__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_26_AWLOCK = edge_list_ch_26__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_26_AWPROT = edge_list_ch_26__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_26_AWQOS = edge_list_ch_26__m_axi_m_axi_AWQOS;
  assign edge_list_ch_26__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_26_AWREADY;
  assign m_axi_edge_list_ch_26_AWSIZE = edge_list_ch_26__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_26_AWVALID = edge_list_ch_26__m_axi_m_axi_AWVALID;
  assign edge_list_ch_26__m_axi_m_axi_BID = m_axi_edge_list_ch_26_BID;
  assign m_axi_edge_list_ch_26_BREADY = edge_list_ch_26__m_axi_m_axi_BREADY;
  assign edge_list_ch_26__m_axi_m_axi_BRESP = m_axi_edge_list_ch_26_BRESP;
  assign edge_list_ch_26__m_axi_m_axi_BVALID = m_axi_edge_list_ch_26_BVALID;
  assign edge_list_ch_26__m_axi_m_axi_RDATA = m_axi_edge_list_ch_26_RDATA;
  assign edge_list_ch_26__m_axi_m_axi_RID = m_axi_edge_list_ch_26_RID;
  assign edge_list_ch_26__m_axi_m_axi_RLAST = m_axi_edge_list_ch_26_RLAST;
  assign m_axi_edge_list_ch_26_RREADY = edge_list_ch_26__m_axi_m_axi_RREADY;
  assign edge_list_ch_26__m_axi_m_axi_RRESP = m_axi_edge_list_ch_26_RRESP;
  assign edge_list_ch_26__m_axi_m_axi_RVALID = m_axi_edge_list_ch_26_RVALID;
  assign m_axi_edge_list_ch_26_WDATA = edge_list_ch_26__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_26_WLAST = edge_list_ch_26__m_axi_m_axi_WLAST;
  assign edge_list_ch_26__m_axi_m_axi_WREADY = m_axi_edge_list_ch_26_WREADY;
  assign m_axi_edge_list_ch_26_WSTRB = edge_list_ch_26__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_26_WVALID = edge_list_ch_26__m_axi_m_axi_WVALID;
  assign edge_list_ch_26__m_axi_read_addr_din = edge_list_ch_26_read_addr__din;
  assign edge_list_ch_26_read_addr__full_n = edge_list_ch_26__m_axi_read_addr_full_n;
  assign edge_list_ch_26__m_axi_read_addr_write = edge_list_ch_26_read_addr__write;
  assign edge_list_ch_26_read_data__dout = edge_list_ch_26__m_axi_read_data_dout;
  assign edge_list_ch_26_read_data__empty_n = edge_list_ch_26__m_axi_read_data_empty_n;
  assign edge_list_ch_26__m_axi_read_data_read = edge_list_ch_26_read_data__read;
  assign edge_list_ch_26__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_26__m_axi_write_addr_din = edge_list_ch_26_write_addr__din;
  assign edge_list_ch_26_write_addr__full_n = edge_list_ch_26__m_axi_write_addr_full_n;
  assign edge_list_ch_26__m_axi_write_addr_write = edge_list_ch_26_write_addr__write;
  assign edge_list_ch_26__m_axi_write_data_din = edge_list_ch_26_write_data__din;
  assign edge_list_ch_26_write_data__full_n = edge_list_ch_26__m_axi_write_data_full_n;
  assign edge_list_ch_26__m_axi_write_data_write = edge_list_ch_26_write_data__write;
  assign edge_list_ch_26_write_resp__dout = edge_list_ch_26__m_axi_write_resp_dout;
  assign edge_list_ch_26_write_resp__empty_n = edge_list_ch_26__m_axi_write_resp_empty_n;
  assign edge_list_ch_26__m_axi_write_resp_read = edge_list_ch_26_write_resp__read;
  assign edge_list_ch_27__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_27_ARADDR = edge_list_ch_27__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_27_ARBURST = edge_list_ch_27__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_27_ARCACHE = edge_list_ch_27__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_27_ARID = edge_list_ch_27__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_27_ARLEN = edge_list_ch_27__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_27_ARLOCK = edge_list_ch_27__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_27_ARPROT = edge_list_ch_27__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_27_ARQOS = edge_list_ch_27__m_axi_m_axi_ARQOS;
  assign edge_list_ch_27__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_27_ARREADY;
  assign m_axi_edge_list_ch_27_ARSIZE = edge_list_ch_27__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_27_ARVALID = edge_list_ch_27__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_27_AWADDR = edge_list_ch_27__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_27_AWBURST = edge_list_ch_27__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_27_AWCACHE = edge_list_ch_27__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_27_AWID = edge_list_ch_27__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_27_AWLEN = edge_list_ch_27__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_27_AWLOCK = edge_list_ch_27__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_27_AWPROT = edge_list_ch_27__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_27_AWQOS = edge_list_ch_27__m_axi_m_axi_AWQOS;
  assign edge_list_ch_27__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_27_AWREADY;
  assign m_axi_edge_list_ch_27_AWSIZE = edge_list_ch_27__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_27_AWVALID = edge_list_ch_27__m_axi_m_axi_AWVALID;
  assign edge_list_ch_27__m_axi_m_axi_BID = m_axi_edge_list_ch_27_BID;
  assign m_axi_edge_list_ch_27_BREADY = edge_list_ch_27__m_axi_m_axi_BREADY;
  assign edge_list_ch_27__m_axi_m_axi_BRESP = m_axi_edge_list_ch_27_BRESP;
  assign edge_list_ch_27__m_axi_m_axi_BVALID = m_axi_edge_list_ch_27_BVALID;
  assign edge_list_ch_27__m_axi_m_axi_RDATA = m_axi_edge_list_ch_27_RDATA;
  assign edge_list_ch_27__m_axi_m_axi_RID = m_axi_edge_list_ch_27_RID;
  assign edge_list_ch_27__m_axi_m_axi_RLAST = m_axi_edge_list_ch_27_RLAST;
  assign m_axi_edge_list_ch_27_RREADY = edge_list_ch_27__m_axi_m_axi_RREADY;
  assign edge_list_ch_27__m_axi_m_axi_RRESP = m_axi_edge_list_ch_27_RRESP;
  assign edge_list_ch_27__m_axi_m_axi_RVALID = m_axi_edge_list_ch_27_RVALID;
  assign m_axi_edge_list_ch_27_WDATA = edge_list_ch_27__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_27_WLAST = edge_list_ch_27__m_axi_m_axi_WLAST;
  assign edge_list_ch_27__m_axi_m_axi_WREADY = m_axi_edge_list_ch_27_WREADY;
  assign m_axi_edge_list_ch_27_WSTRB = edge_list_ch_27__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_27_WVALID = edge_list_ch_27__m_axi_m_axi_WVALID;
  assign edge_list_ch_27__m_axi_read_addr_din = edge_list_ch_27_read_addr__din;
  assign edge_list_ch_27_read_addr__full_n = edge_list_ch_27__m_axi_read_addr_full_n;
  assign edge_list_ch_27__m_axi_read_addr_write = edge_list_ch_27_read_addr__write;
  assign edge_list_ch_27_read_data__dout = edge_list_ch_27__m_axi_read_data_dout;
  assign edge_list_ch_27_read_data__empty_n = edge_list_ch_27__m_axi_read_data_empty_n;
  assign edge_list_ch_27__m_axi_read_data_read = edge_list_ch_27_read_data__read;
  assign edge_list_ch_27__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_27__m_axi_write_addr_din = edge_list_ch_27_write_addr__din;
  assign edge_list_ch_27_write_addr__full_n = edge_list_ch_27__m_axi_write_addr_full_n;
  assign edge_list_ch_27__m_axi_write_addr_write = edge_list_ch_27_write_addr__write;
  assign edge_list_ch_27__m_axi_write_data_din = edge_list_ch_27_write_data__din;
  assign edge_list_ch_27_write_data__full_n = edge_list_ch_27__m_axi_write_data_full_n;
  assign edge_list_ch_27__m_axi_write_data_write = edge_list_ch_27_write_data__write;
  assign edge_list_ch_27_write_resp__dout = edge_list_ch_27__m_axi_write_resp_dout;
  assign edge_list_ch_27_write_resp__empty_n = edge_list_ch_27__m_axi_write_resp_empty_n;
  assign edge_list_ch_27__m_axi_write_resp_read = edge_list_ch_27_write_resp__read;
  assign edge_list_ch_28__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_28_ARADDR = edge_list_ch_28__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_28_ARBURST = edge_list_ch_28__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_28_ARCACHE = edge_list_ch_28__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_28_ARID = edge_list_ch_28__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_28_ARLEN = edge_list_ch_28__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_28_ARLOCK = edge_list_ch_28__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_28_ARPROT = edge_list_ch_28__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_28_ARQOS = edge_list_ch_28__m_axi_m_axi_ARQOS;
  assign edge_list_ch_28__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_28_ARREADY;
  assign m_axi_edge_list_ch_28_ARSIZE = edge_list_ch_28__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_28_ARVALID = edge_list_ch_28__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_28_AWADDR = edge_list_ch_28__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_28_AWBURST = edge_list_ch_28__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_28_AWCACHE = edge_list_ch_28__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_28_AWID = edge_list_ch_28__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_28_AWLEN = edge_list_ch_28__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_28_AWLOCK = edge_list_ch_28__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_28_AWPROT = edge_list_ch_28__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_28_AWQOS = edge_list_ch_28__m_axi_m_axi_AWQOS;
  assign edge_list_ch_28__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_28_AWREADY;
  assign m_axi_edge_list_ch_28_AWSIZE = edge_list_ch_28__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_28_AWVALID = edge_list_ch_28__m_axi_m_axi_AWVALID;
  assign edge_list_ch_28__m_axi_m_axi_BID = m_axi_edge_list_ch_28_BID;
  assign m_axi_edge_list_ch_28_BREADY = edge_list_ch_28__m_axi_m_axi_BREADY;
  assign edge_list_ch_28__m_axi_m_axi_BRESP = m_axi_edge_list_ch_28_BRESP;
  assign edge_list_ch_28__m_axi_m_axi_BVALID = m_axi_edge_list_ch_28_BVALID;
  assign edge_list_ch_28__m_axi_m_axi_RDATA = m_axi_edge_list_ch_28_RDATA;
  assign edge_list_ch_28__m_axi_m_axi_RID = m_axi_edge_list_ch_28_RID;
  assign edge_list_ch_28__m_axi_m_axi_RLAST = m_axi_edge_list_ch_28_RLAST;
  assign m_axi_edge_list_ch_28_RREADY = edge_list_ch_28__m_axi_m_axi_RREADY;
  assign edge_list_ch_28__m_axi_m_axi_RRESP = m_axi_edge_list_ch_28_RRESP;
  assign edge_list_ch_28__m_axi_m_axi_RVALID = m_axi_edge_list_ch_28_RVALID;
  assign m_axi_edge_list_ch_28_WDATA = edge_list_ch_28__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_28_WLAST = edge_list_ch_28__m_axi_m_axi_WLAST;
  assign edge_list_ch_28__m_axi_m_axi_WREADY = m_axi_edge_list_ch_28_WREADY;
  assign m_axi_edge_list_ch_28_WSTRB = edge_list_ch_28__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_28_WVALID = edge_list_ch_28__m_axi_m_axi_WVALID;
  assign edge_list_ch_28__m_axi_read_addr_din = edge_list_ch_28_read_addr__din;
  assign edge_list_ch_28_read_addr__full_n = edge_list_ch_28__m_axi_read_addr_full_n;
  assign edge_list_ch_28__m_axi_read_addr_write = edge_list_ch_28_read_addr__write;
  assign edge_list_ch_28_read_data__dout = edge_list_ch_28__m_axi_read_data_dout;
  assign edge_list_ch_28_read_data__empty_n = edge_list_ch_28__m_axi_read_data_empty_n;
  assign edge_list_ch_28__m_axi_read_data_read = edge_list_ch_28_read_data__read;
  assign edge_list_ch_28__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_28__m_axi_write_addr_din = edge_list_ch_28_write_addr__din;
  assign edge_list_ch_28_write_addr__full_n = edge_list_ch_28__m_axi_write_addr_full_n;
  assign edge_list_ch_28__m_axi_write_addr_write = edge_list_ch_28_write_addr__write;
  assign edge_list_ch_28__m_axi_write_data_din = edge_list_ch_28_write_data__din;
  assign edge_list_ch_28_write_data__full_n = edge_list_ch_28__m_axi_write_data_full_n;
  assign edge_list_ch_28__m_axi_write_data_write = edge_list_ch_28_write_data__write;
  assign edge_list_ch_28_write_resp__dout = edge_list_ch_28__m_axi_write_resp_dout;
  assign edge_list_ch_28_write_resp__empty_n = edge_list_ch_28__m_axi_write_resp_empty_n;
  assign edge_list_ch_28__m_axi_write_resp_read = edge_list_ch_28_write_resp__read;
  assign edge_list_ch_29__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_29_ARADDR = edge_list_ch_29__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_29_ARBURST = edge_list_ch_29__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_29_ARCACHE = edge_list_ch_29__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_29_ARID = edge_list_ch_29__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_29_ARLEN = edge_list_ch_29__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_29_ARLOCK = edge_list_ch_29__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_29_ARPROT = edge_list_ch_29__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_29_ARQOS = edge_list_ch_29__m_axi_m_axi_ARQOS;
  assign edge_list_ch_29__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_29_ARREADY;
  assign m_axi_edge_list_ch_29_ARSIZE = edge_list_ch_29__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_29_ARVALID = edge_list_ch_29__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_29_AWADDR = edge_list_ch_29__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_29_AWBURST = edge_list_ch_29__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_29_AWCACHE = edge_list_ch_29__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_29_AWID = edge_list_ch_29__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_29_AWLEN = edge_list_ch_29__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_29_AWLOCK = edge_list_ch_29__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_29_AWPROT = edge_list_ch_29__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_29_AWQOS = edge_list_ch_29__m_axi_m_axi_AWQOS;
  assign edge_list_ch_29__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_29_AWREADY;
  assign m_axi_edge_list_ch_29_AWSIZE = edge_list_ch_29__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_29_AWVALID = edge_list_ch_29__m_axi_m_axi_AWVALID;
  assign edge_list_ch_29__m_axi_m_axi_BID = m_axi_edge_list_ch_29_BID;
  assign m_axi_edge_list_ch_29_BREADY = edge_list_ch_29__m_axi_m_axi_BREADY;
  assign edge_list_ch_29__m_axi_m_axi_BRESP = m_axi_edge_list_ch_29_BRESP;
  assign edge_list_ch_29__m_axi_m_axi_BVALID = m_axi_edge_list_ch_29_BVALID;
  assign edge_list_ch_29__m_axi_m_axi_RDATA = m_axi_edge_list_ch_29_RDATA;
  assign edge_list_ch_29__m_axi_m_axi_RID = m_axi_edge_list_ch_29_RID;
  assign edge_list_ch_29__m_axi_m_axi_RLAST = m_axi_edge_list_ch_29_RLAST;
  assign m_axi_edge_list_ch_29_RREADY = edge_list_ch_29__m_axi_m_axi_RREADY;
  assign edge_list_ch_29__m_axi_m_axi_RRESP = m_axi_edge_list_ch_29_RRESP;
  assign edge_list_ch_29__m_axi_m_axi_RVALID = m_axi_edge_list_ch_29_RVALID;
  assign m_axi_edge_list_ch_29_WDATA = edge_list_ch_29__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_29_WLAST = edge_list_ch_29__m_axi_m_axi_WLAST;
  assign edge_list_ch_29__m_axi_m_axi_WREADY = m_axi_edge_list_ch_29_WREADY;
  assign m_axi_edge_list_ch_29_WSTRB = edge_list_ch_29__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_29_WVALID = edge_list_ch_29__m_axi_m_axi_WVALID;
  assign edge_list_ch_29__m_axi_read_addr_din = edge_list_ch_29_read_addr__din;
  assign edge_list_ch_29_read_addr__full_n = edge_list_ch_29__m_axi_read_addr_full_n;
  assign edge_list_ch_29__m_axi_read_addr_write = edge_list_ch_29_read_addr__write;
  assign edge_list_ch_29_read_data__dout = edge_list_ch_29__m_axi_read_data_dout;
  assign edge_list_ch_29_read_data__empty_n = edge_list_ch_29__m_axi_read_data_empty_n;
  assign edge_list_ch_29__m_axi_read_data_read = edge_list_ch_29_read_data__read;
  assign edge_list_ch_29__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_29__m_axi_write_addr_din = edge_list_ch_29_write_addr__din;
  assign edge_list_ch_29_write_addr__full_n = edge_list_ch_29__m_axi_write_addr_full_n;
  assign edge_list_ch_29__m_axi_write_addr_write = edge_list_ch_29_write_addr__write;
  assign edge_list_ch_29__m_axi_write_data_din = edge_list_ch_29_write_data__din;
  assign edge_list_ch_29_write_data__full_n = edge_list_ch_29__m_axi_write_data_full_n;
  assign edge_list_ch_29__m_axi_write_data_write = edge_list_ch_29_write_data__write;
  assign edge_list_ch_29_write_resp__dout = edge_list_ch_29__m_axi_write_resp_dout;
  assign edge_list_ch_29_write_resp__empty_n = edge_list_ch_29__m_axi_write_resp_empty_n;
  assign edge_list_ch_29__m_axi_write_resp_read = edge_list_ch_29_write_resp__read;
  assign edge_list_ch_30__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_30_ARADDR = edge_list_ch_30__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_30_ARBURST = edge_list_ch_30__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_30_ARCACHE = edge_list_ch_30__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_30_ARID = edge_list_ch_30__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_30_ARLEN = edge_list_ch_30__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_30_ARLOCK = edge_list_ch_30__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_30_ARPROT = edge_list_ch_30__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_30_ARQOS = edge_list_ch_30__m_axi_m_axi_ARQOS;
  assign edge_list_ch_30__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_30_ARREADY;
  assign m_axi_edge_list_ch_30_ARSIZE = edge_list_ch_30__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_30_ARVALID = edge_list_ch_30__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_30_AWADDR = edge_list_ch_30__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_30_AWBURST = edge_list_ch_30__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_30_AWCACHE = edge_list_ch_30__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_30_AWID = edge_list_ch_30__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_30_AWLEN = edge_list_ch_30__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_30_AWLOCK = edge_list_ch_30__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_30_AWPROT = edge_list_ch_30__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_30_AWQOS = edge_list_ch_30__m_axi_m_axi_AWQOS;
  assign edge_list_ch_30__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_30_AWREADY;
  assign m_axi_edge_list_ch_30_AWSIZE = edge_list_ch_30__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_30_AWVALID = edge_list_ch_30__m_axi_m_axi_AWVALID;
  assign edge_list_ch_30__m_axi_m_axi_BID = m_axi_edge_list_ch_30_BID;
  assign m_axi_edge_list_ch_30_BREADY = edge_list_ch_30__m_axi_m_axi_BREADY;
  assign edge_list_ch_30__m_axi_m_axi_BRESP = m_axi_edge_list_ch_30_BRESP;
  assign edge_list_ch_30__m_axi_m_axi_BVALID = m_axi_edge_list_ch_30_BVALID;
  assign edge_list_ch_30__m_axi_m_axi_RDATA = m_axi_edge_list_ch_30_RDATA;
  assign edge_list_ch_30__m_axi_m_axi_RID = m_axi_edge_list_ch_30_RID;
  assign edge_list_ch_30__m_axi_m_axi_RLAST = m_axi_edge_list_ch_30_RLAST;
  assign m_axi_edge_list_ch_30_RREADY = edge_list_ch_30__m_axi_m_axi_RREADY;
  assign edge_list_ch_30__m_axi_m_axi_RRESP = m_axi_edge_list_ch_30_RRESP;
  assign edge_list_ch_30__m_axi_m_axi_RVALID = m_axi_edge_list_ch_30_RVALID;
  assign m_axi_edge_list_ch_30_WDATA = edge_list_ch_30__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_30_WLAST = edge_list_ch_30__m_axi_m_axi_WLAST;
  assign edge_list_ch_30__m_axi_m_axi_WREADY = m_axi_edge_list_ch_30_WREADY;
  assign m_axi_edge_list_ch_30_WSTRB = edge_list_ch_30__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_30_WVALID = edge_list_ch_30__m_axi_m_axi_WVALID;
  assign edge_list_ch_30__m_axi_read_addr_din = edge_list_ch_30_read_addr__din;
  assign edge_list_ch_30_read_addr__full_n = edge_list_ch_30__m_axi_read_addr_full_n;
  assign edge_list_ch_30__m_axi_read_addr_write = edge_list_ch_30_read_addr__write;
  assign edge_list_ch_30_read_data__dout = edge_list_ch_30__m_axi_read_data_dout;
  assign edge_list_ch_30_read_data__empty_n = edge_list_ch_30__m_axi_read_data_empty_n;
  assign edge_list_ch_30__m_axi_read_data_read = edge_list_ch_30_read_data__read;
  assign edge_list_ch_30__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_30__m_axi_write_addr_din = edge_list_ch_30_write_addr__din;
  assign edge_list_ch_30_write_addr__full_n = edge_list_ch_30__m_axi_write_addr_full_n;
  assign edge_list_ch_30__m_axi_write_addr_write = edge_list_ch_30_write_addr__write;
  assign edge_list_ch_30__m_axi_write_data_din = edge_list_ch_30_write_data__din;
  assign edge_list_ch_30_write_data__full_n = edge_list_ch_30__m_axi_write_data_full_n;
  assign edge_list_ch_30__m_axi_write_data_write = edge_list_ch_30_write_data__write;
  assign edge_list_ch_30_write_resp__dout = edge_list_ch_30__m_axi_write_resp_dout;
  assign edge_list_ch_30_write_resp__empty_n = edge_list_ch_30__m_axi_write_resp_empty_n;
  assign edge_list_ch_30__m_axi_write_resp_read = edge_list_ch_30_write_resp__read;
  assign edge_list_ch_31__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_31_ARADDR = edge_list_ch_31__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_31_ARBURST = edge_list_ch_31__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_31_ARCACHE = edge_list_ch_31__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_31_ARID = edge_list_ch_31__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_31_ARLEN = edge_list_ch_31__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_31_ARLOCK = edge_list_ch_31__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_31_ARPROT = edge_list_ch_31__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_31_ARQOS = edge_list_ch_31__m_axi_m_axi_ARQOS;
  assign edge_list_ch_31__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_31_ARREADY;
  assign m_axi_edge_list_ch_31_ARSIZE = edge_list_ch_31__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_31_ARVALID = edge_list_ch_31__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_31_AWADDR = edge_list_ch_31__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_31_AWBURST = edge_list_ch_31__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_31_AWCACHE = edge_list_ch_31__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_31_AWID = edge_list_ch_31__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_31_AWLEN = edge_list_ch_31__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_31_AWLOCK = edge_list_ch_31__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_31_AWPROT = edge_list_ch_31__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_31_AWQOS = edge_list_ch_31__m_axi_m_axi_AWQOS;
  assign edge_list_ch_31__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_31_AWREADY;
  assign m_axi_edge_list_ch_31_AWSIZE = edge_list_ch_31__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_31_AWVALID = edge_list_ch_31__m_axi_m_axi_AWVALID;
  assign edge_list_ch_31__m_axi_m_axi_BID = m_axi_edge_list_ch_31_BID;
  assign m_axi_edge_list_ch_31_BREADY = edge_list_ch_31__m_axi_m_axi_BREADY;
  assign edge_list_ch_31__m_axi_m_axi_BRESP = m_axi_edge_list_ch_31_BRESP;
  assign edge_list_ch_31__m_axi_m_axi_BVALID = m_axi_edge_list_ch_31_BVALID;
  assign edge_list_ch_31__m_axi_m_axi_RDATA = m_axi_edge_list_ch_31_RDATA;
  assign edge_list_ch_31__m_axi_m_axi_RID = m_axi_edge_list_ch_31_RID;
  assign edge_list_ch_31__m_axi_m_axi_RLAST = m_axi_edge_list_ch_31_RLAST;
  assign m_axi_edge_list_ch_31_RREADY = edge_list_ch_31__m_axi_m_axi_RREADY;
  assign edge_list_ch_31__m_axi_m_axi_RRESP = m_axi_edge_list_ch_31_RRESP;
  assign edge_list_ch_31__m_axi_m_axi_RVALID = m_axi_edge_list_ch_31_RVALID;
  assign m_axi_edge_list_ch_31_WDATA = edge_list_ch_31__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_31_WLAST = edge_list_ch_31__m_axi_m_axi_WLAST;
  assign edge_list_ch_31__m_axi_m_axi_WREADY = m_axi_edge_list_ch_31_WREADY;
  assign m_axi_edge_list_ch_31_WSTRB = edge_list_ch_31__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_31_WVALID = edge_list_ch_31__m_axi_m_axi_WVALID;
  assign edge_list_ch_31__m_axi_read_addr_din = edge_list_ch_31_read_addr__din;
  assign edge_list_ch_31_read_addr__full_n = edge_list_ch_31__m_axi_read_addr_full_n;
  assign edge_list_ch_31__m_axi_read_addr_write = edge_list_ch_31_read_addr__write;
  assign edge_list_ch_31_read_data__dout = edge_list_ch_31__m_axi_read_data_dout;
  assign edge_list_ch_31_read_data__empty_n = edge_list_ch_31__m_axi_read_data_empty_n;
  assign edge_list_ch_31__m_axi_read_data_read = edge_list_ch_31_read_data__read;
  assign edge_list_ch_31__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_31__m_axi_write_addr_din = edge_list_ch_31_write_addr__din;
  assign edge_list_ch_31_write_addr__full_n = edge_list_ch_31__m_axi_write_addr_full_n;
  assign edge_list_ch_31__m_axi_write_addr_write = edge_list_ch_31_write_addr__write;
  assign edge_list_ch_31__m_axi_write_data_din = edge_list_ch_31_write_data__din;
  assign edge_list_ch_31_write_data__full_n = edge_list_ch_31__m_axi_write_data_full_n;
  assign edge_list_ch_31__m_axi_write_data_write = edge_list_ch_31_write_data__write;
  assign edge_list_ch_31_write_resp__dout = edge_list_ch_31__m_axi_write_resp_dout;
  assign edge_list_ch_31_write_resp__empty_n = edge_list_ch_31__m_axi_write_resp_empty_n;
  assign edge_list_ch_31__m_axi_write_resp_read = edge_list_ch_31_write_resp__read;
  assign edge_list_ch_32__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_32_ARADDR = edge_list_ch_32__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_32_ARBURST = edge_list_ch_32__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_32_ARCACHE = edge_list_ch_32__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_32_ARID = edge_list_ch_32__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_32_ARLEN = edge_list_ch_32__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_32_ARLOCK = edge_list_ch_32__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_32_ARPROT = edge_list_ch_32__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_32_ARQOS = edge_list_ch_32__m_axi_m_axi_ARQOS;
  assign edge_list_ch_32__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_32_ARREADY;
  assign m_axi_edge_list_ch_32_ARSIZE = edge_list_ch_32__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_32_ARVALID = edge_list_ch_32__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_32_AWADDR = edge_list_ch_32__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_32_AWBURST = edge_list_ch_32__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_32_AWCACHE = edge_list_ch_32__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_32_AWID = edge_list_ch_32__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_32_AWLEN = edge_list_ch_32__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_32_AWLOCK = edge_list_ch_32__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_32_AWPROT = edge_list_ch_32__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_32_AWQOS = edge_list_ch_32__m_axi_m_axi_AWQOS;
  assign edge_list_ch_32__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_32_AWREADY;
  assign m_axi_edge_list_ch_32_AWSIZE = edge_list_ch_32__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_32_AWVALID = edge_list_ch_32__m_axi_m_axi_AWVALID;
  assign edge_list_ch_32__m_axi_m_axi_BID = m_axi_edge_list_ch_32_BID;
  assign m_axi_edge_list_ch_32_BREADY = edge_list_ch_32__m_axi_m_axi_BREADY;
  assign edge_list_ch_32__m_axi_m_axi_BRESP = m_axi_edge_list_ch_32_BRESP;
  assign edge_list_ch_32__m_axi_m_axi_BVALID = m_axi_edge_list_ch_32_BVALID;
  assign edge_list_ch_32__m_axi_m_axi_RDATA = m_axi_edge_list_ch_32_RDATA;
  assign edge_list_ch_32__m_axi_m_axi_RID = m_axi_edge_list_ch_32_RID;
  assign edge_list_ch_32__m_axi_m_axi_RLAST = m_axi_edge_list_ch_32_RLAST;
  assign m_axi_edge_list_ch_32_RREADY = edge_list_ch_32__m_axi_m_axi_RREADY;
  assign edge_list_ch_32__m_axi_m_axi_RRESP = m_axi_edge_list_ch_32_RRESP;
  assign edge_list_ch_32__m_axi_m_axi_RVALID = m_axi_edge_list_ch_32_RVALID;
  assign m_axi_edge_list_ch_32_WDATA = edge_list_ch_32__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_32_WLAST = edge_list_ch_32__m_axi_m_axi_WLAST;
  assign edge_list_ch_32__m_axi_m_axi_WREADY = m_axi_edge_list_ch_32_WREADY;
  assign m_axi_edge_list_ch_32_WSTRB = edge_list_ch_32__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_32_WVALID = edge_list_ch_32__m_axi_m_axi_WVALID;
  assign edge_list_ch_32__m_axi_read_addr_din = edge_list_ch_32_read_addr__din;
  assign edge_list_ch_32_read_addr__full_n = edge_list_ch_32__m_axi_read_addr_full_n;
  assign edge_list_ch_32__m_axi_read_addr_write = edge_list_ch_32_read_addr__write;
  assign edge_list_ch_32_read_data__dout = edge_list_ch_32__m_axi_read_data_dout;
  assign edge_list_ch_32_read_data__empty_n = edge_list_ch_32__m_axi_read_data_empty_n;
  assign edge_list_ch_32__m_axi_read_data_read = edge_list_ch_32_read_data__read;
  assign edge_list_ch_32__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_32__m_axi_write_addr_din = edge_list_ch_32_write_addr__din;
  assign edge_list_ch_32_write_addr__full_n = edge_list_ch_32__m_axi_write_addr_full_n;
  assign edge_list_ch_32__m_axi_write_addr_write = edge_list_ch_32_write_addr__write;
  assign edge_list_ch_32__m_axi_write_data_din = edge_list_ch_32_write_data__din;
  assign edge_list_ch_32_write_data__full_n = edge_list_ch_32__m_axi_write_data_full_n;
  assign edge_list_ch_32__m_axi_write_data_write = edge_list_ch_32_write_data__write;
  assign edge_list_ch_32_write_resp__dout = edge_list_ch_32__m_axi_write_resp_dout;
  assign edge_list_ch_32_write_resp__empty_n = edge_list_ch_32__m_axi_write_resp_empty_n;
  assign edge_list_ch_32__m_axi_write_resp_read = edge_list_ch_32_write_resp__read;
  assign edge_list_ch_33__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_33_ARADDR = edge_list_ch_33__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_33_ARBURST = edge_list_ch_33__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_33_ARCACHE = edge_list_ch_33__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_33_ARID = edge_list_ch_33__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_33_ARLEN = edge_list_ch_33__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_33_ARLOCK = edge_list_ch_33__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_33_ARPROT = edge_list_ch_33__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_33_ARQOS = edge_list_ch_33__m_axi_m_axi_ARQOS;
  assign edge_list_ch_33__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_33_ARREADY;
  assign m_axi_edge_list_ch_33_ARSIZE = edge_list_ch_33__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_33_ARVALID = edge_list_ch_33__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_33_AWADDR = edge_list_ch_33__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_33_AWBURST = edge_list_ch_33__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_33_AWCACHE = edge_list_ch_33__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_33_AWID = edge_list_ch_33__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_33_AWLEN = edge_list_ch_33__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_33_AWLOCK = edge_list_ch_33__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_33_AWPROT = edge_list_ch_33__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_33_AWQOS = edge_list_ch_33__m_axi_m_axi_AWQOS;
  assign edge_list_ch_33__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_33_AWREADY;
  assign m_axi_edge_list_ch_33_AWSIZE = edge_list_ch_33__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_33_AWVALID = edge_list_ch_33__m_axi_m_axi_AWVALID;
  assign edge_list_ch_33__m_axi_m_axi_BID = m_axi_edge_list_ch_33_BID;
  assign m_axi_edge_list_ch_33_BREADY = edge_list_ch_33__m_axi_m_axi_BREADY;
  assign edge_list_ch_33__m_axi_m_axi_BRESP = m_axi_edge_list_ch_33_BRESP;
  assign edge_list_ch_33__m_axi_m_axi_BVALID = m_axi_edge_list_ch_33_BVALID;
  assign edge_list_ch_33__m_axi_m_axi_RDATA = m_axi_edge_list_ch_33_RDATA;
  assign edge_list_ch_33__m_axi_m_axi_RID = m_axi_edge_list_ch_33_RID;
  assign edge_list_ch_33__m_axi_m_axi_RLAST = m_axi_edge_list_ch_33_RLAST;
  assign m_axi_edge_list_ch_33_RREADY = edge_list_ch_33__m_axi_m_axi_RREADY;
  assign edge_list_ch_33__m_axi_m_axi_RRESP = m_axi_edge_list_ch_33_RRESP;
  assign edge_list_ch_33__m_axi_m_axi_RVALID = m_axi_edge_list_ch_33_RVALID;
  assign m_axi_edge_list_ch_33_WDATA = edge_list_ch_33__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_33_WLAST = edge_list_ch_33__m_axi_m_axi_WLAST;
  assign edge_list_ch_33__m_axi_m_axi_WREADY = m_axi_edge_list_ch_33_WREADY;
  assign m_axi_edge_list_ch_33_WSTRB = edge_list_ch_33__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_33_WVALID = edge_list_ch_33__m_axi_m_axi_WVALID;
  assign edge_list_ch_33__m_axi_read_addr_din = edge_list_ch_33_read_addr__din;
  assign edge_list_ch_33_read_addr__full_n = edge_list_ch_33__m_axi_read_addr_full_n;
  assign edge_list_ch_33__m_axi_read_addr_write = edge_list_ch_33_read_addr__write;
  assign edge_list_ch_33_read_data__dout = edge_list_ch_33__m_axi_read_data_dout;
  assign edge_list_ch_33_read_data__empty_n = edge_list_ch_33__m_axi_read_data_empty_n;
  assign edge_list_ch_33__m_axi_read_data_read = edge_list_ch_33_read_data__read;
  assign edge_list_ch_33__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_33__m_axi_write_addr_din = edge_list_ch_33_write_addr__din;
  assign edge_list_ch_33_write_addr__full_n = edge_list_ch_33__m_axi_write_addr_full_n;
  assign edge_list_ch_33__m_axi_write_addr_write = edge_list_ch_33_write_addr__write;
  assign edge_list_ch_33__m_axi_write_data_din = edge_list_ch_33_write_data__din;
  assign edge_list_ch_33_write_data__full_n = edge_list_ch_33__m_axi_write_data_full_n;
  assign edge_list_ch_33__m_axi_write_data_write = edge_list_ch_33_write_data__write;
  assign edge_list_ch_33_write_resp__dout = edge_list_ch_33__m_axi_write_resp_dout;
  assign edge_list_ch_33_write_resp__empty_n = edge_list_ch_33__m_axi_write_resp_empty_n;
  assign edge_list_ch_33__m_axi_write_resp_read = edge_list_ch_33_write_resp__read;
  assign edge_list_ch_34__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_34_ARADDR = edge_list_ch_34__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_34_ARBURST = edge_list_ch_34__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_34_ARCACHE = edge_list_ch_34__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_34_ARID = edge_list_ch_34__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_34_ARLEN = edge_list_ch_34__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_34_ARLOCK = edge_list_ch_34__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_34_ARPROT = edge_list_ch_34__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_34_ARQOS = edge_list_ch_34__m_axi_m_axi_ARQOS;
  assign edge_list_ch_34__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_34_ARREADY;
  assign m_axi_edge_list_ch_34_ARSIZE = edge_list_ch_34__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_34_ARVALID = edge_list_ch_34__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_34_AWADDR = edge_list_ch_34__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_34_AWBURST = edge_list_ch_34__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_34_AWCACHE = edge_list_ch_34__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_34_AWID = edge_list_ch_34__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_34_AWLEN = edge_list_ch_34__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_34_AWLOCK = edge_list_ch_34__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_34_AWPROT = edge_list_ch_34__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_34_AWQOS = edge_list_ch_34__m_axi_m_axi_AWQOS;
  assign edge_list_ch_34__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_34_AWREADY;
  assign m_axi_edge_list_ch_34_AWSIZE = edge_list_ch_34__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_34_AWVALID = edge_list_ch_34__m_axi_m_axi_AWVALID;
  assign edge_list_ch_34__m_axi_m_axi_BID = m_axi_edge_list_ch_34_BID;
  assign m_axi_edge_list_ch_34_BREADY = edge_list_ch_34__m_axi_m_axi_BREADY;
  assign edge_list_ch_34__m_axi_m_axi_BRESP = m_axi_edge_list_ch_34_BRESP;
  assign edge_list_ch_34__m_axi_m_axi_BVALID = m_axi_edge_list_ch_34_BVALID;
  assign edge_list_ch_34__m_axi_m_axi_RDATA = m_axi_edge_list_ch_34_RDATA;
  assign edge_list_ch_34__m_axi_m_axi_RID = m_axi_edge_list_ch_34_RID;
  assign edge_list_ch_34__m_axi_m_axi_RLAST = m_axi_edge_list_ch_34_RLAST;
  assign m_axi_edge_list_ch_34_RREADY = edge_list_ch_34__m_axi_m_axi_RREADY;
  assign edge_list_ch_34__m_axi_m_axi_RRESP = m_axi_edge_list_ch_34_RRESP;
  assign edge_list_ch_34__m_axi_m_axi_RVALID = m_axi_edge_list_ch_34_RVALID;
  assign m_axi_edge_list_ch_34_WDATA = edge_list_ch_34__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_34_WLAST = edge_list_ch_34__m_axi_m_axi_WLAST;
  assign edge_list_ch_34__m_axi_m_axi_WREADY = m_axi_edge_list_ch_34_WREADY;
  assign m_axi_edge_list_ch_34_WSTRB = edge_list_ch_34__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_34_WVALID = edge_list_ch_34__m_axi_m_axi_WVALID;
  assign edge_list_ch_34__m_axi_read_addr_din = edge_list_ch_34_read_addr__din;
  assign edge_list_ch_34_read_addr__full_n = edge_list_ch_34__m_axi_read_addr_full_n;
  assign edge_list_ch_34__m_axi_read_addr_write = edge_list_ch_34_read_addr__write;
  assign edge_list_ch_34_read_data__dout = edge_list_ch_34__m_axi_read_data_dout;
  assign edge_list_ch_34_read_data__empty_n = edge_list_ch_34__m_axi_read_data_empty_n;
  assign edge_list_ch_34__m_axi_read_data_read = edge_list_ch_34_read_data__read;
  assign edge_list_ch_34__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_34__m_axi_write_addr_din = edge_list_ch_34_write_addr__din;
  assign edge_list_ch_34_write_addr__full_n = edge_list_ch_34__m_axi_write_addr_full_n;
  assign edge_list_ch_34__m_axi_write_addr_write = edge_list_ch_34_write_addr__write;
  assign edge_list_ch_34__m_axi_write_data_din = edge_list_ch_34_write_data__din;
  assign edge_list_ch_34_write_data__full_n = edge_list_ch_34__m_axi_write_data_full_n;
  assign edge_list_ch_34__m_axi_write_data_write = edge_list_ch_34_write_data__write;
  assign edge_list_ch_34_write_resp__dout = edge_list_ch_34__m_axi_write_resp_dout;
  assign edge_list_ch_34_write_resp__empty_n = edge_list_ch_34__m_axi_write_resp_empty_n;
  assign edge_list_ch_34__m_axi_write_resp_read = edge_list_ch_34_write_resp__read;
  assign edge_list_ch_35__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_35_ARADDR = edge_list_ch_35__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_35_ARBURST = edge_list_ch_35__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_35_ARCACHE = edge_list_ch_35__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_35_ARID = edge_list_ch_35__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_35_ARLEN = edge_list_ch_35__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_35_ARLOCK = edge_list_ch_35__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_35_ARPROT = edge_list_ch_35__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_35_ARQOS = edge_list_ch_35__m_axi_m_axi_ARQOS;
  assign edge_list_ch_35__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_35_ARREADY;
  assign m_axi_edge_list_ch_35_ARSIZE = edge_list_ch_35__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_35_ARVALID = edge_list_ch_35__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_35_AWADDR = edge_list_ch_35__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_35_AWBURST = edge_list_ch_35__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_35_AWCACHE = edge_list_ch_35__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_35_AWID = edge_list_ch_35__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_35_AWLEN = edge_list_ch_35__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_35_AWLOCK = edge_list_ch_35__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_35_AWPROT = edge_list_ch_35__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_35_AWQOS = edge_list_ch_35__m_axi_m_axi_AWQOS;
  assign edge_list_ch_35__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_35_AWREADY;
  assign m_axi_edge_list_ch_35_AWSIZE = edge_list_ch_35__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_35_AWVALID = edge_list_ch_35__m_axi_m_axi_AWVALID;
  assign edge_list_ch_35__m_axi_m_axi_BID = m_axi_edge_list_ch_35_BID;
  assign m_axi_edge_list_ch_35_BREADY = edge_list_ch_35__m_axi_m_axi_BREADY;
  assign edge_list_ch_35__m_axi_m_axi_BRESP = m_axi_edge_list_ch_35_BRESP;
  assign edge_list_ch_35__m_axi_m_axi_BVALID = m_axi_edge_list_ch_35_BVALID;
  assign edge_list_ch_35__m_axi_m_axi_RDATA = m_axi_edge_list_ch_35_RDATA;
  assign edge_list_ch_35__m_axi_m_axi_RID = m_axi_edge_list_ch_35_RID;
  assign edge_list_ch_35__m_axi_m_axi_RLAST = m_axi_edge_list_ch_35_RLAST;
  assign m_axi_edge_list_ch_35_RREADY = edge_list_ch_35__m_axi_m_axi_RREADY;
  assign edge_list_ch_35__m_axi_m_axi_RRESP = m_axi_edge_list_ch_35_RRESP;
  assign edge_list_ch_35__m_axi_m_axi_RVALID = m_axi_edge_list_ch_35_RVALID;
  assign m_axi_edge_list_ch_35_WDATA = edge_list_ch_35__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_35_WLAST = edge_list_ch_35__m_axi_m_axi_WLAST;
  assign edge_list_ch_35__m_axi_m_axi_WREADY = m_axi_edge_list_ch_35_WREADY;
  assign m_axi_edge_list_ch_35_WSTRB = edge_list_ch_35__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_35_WVALID = edge_list_ch_35__m_axi_m_axi_WVALID;
  assign edge_list_ch_35__m_axi_read_addr_din = edge_list_ch_35_read_addr__din;
  assign edge_list_ch_35_read_addr__full_n = edge_list_ch_35__m_axi_read_addr_full_n;
  assign edge_list_ch_35__m_axi_read_addr_write = edge_list_ch_35_read_addr__write;
  assign edge_list_ch_35_read_data__dout = edge_list_ch_35__m_axi_read_data_dout;
  assign edge_list_ch_35_read_data__empty_n = edge_list_ch_35__m_axi_read_data_empty_n;
  assign edge_list_ch_35__m_axi_read_data_read = edge_list_ch_35_read_data__read;
  assign edge_list_ch_35__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_35__m_axi_write_addr_din = edge_list_ch_35_write_addr__din;
  assign edge_list_ch_35_write_addr__full_n = edge_list_ch_35__m_axi_write_addr_full_n;
  assign edge_list_ch_35__m_axi_write_addr_write = edge_list_ch_35_write_addr__write;
  assign edge_list_ch_35__m_axi_write_data_din = edge_list_ch_35_write_data__din;
  assign edge_list_ch_35_write_data__full_n = edge_list_ch_35__m_axi_write_data_full_n;
  assign edge_list_ch_35__m_axi_write_data_write = edge_list_ch_35_write_data__write;
  assign edge_list_ch_35_write_resp__dout = edge_list_ch_35__m_axi_write_resp_dout;
  assign edge_list_ch_35_write_resp__empty_n = edge_list_ch_35__m_axi_write_resp_empty_n;
  assign edge_list_ch_35__m_axi_write_resp_read = edge_list_ch_35_write_resp__read;
  assign edge_list_ch_36__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_36_ARADDR = edge_list_ch_36__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_36_ARBURST = edge_list_ch_36__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_36_ARCACHE = edge_list_ch_36__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_36_ARID = edge_list_ch_36__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_36_ARLEN = edge_list_ch_36__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_36_ARLOCK = edge_list_ch_36__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_36_ARPROT = edge_list_ch_36__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_36_ARQOS = edge_list_ch_36__m_axi_m_axi_ARQOS;
  assign edge_list_ch_36__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_36_ARREADY;
  assign m_axi_edge_list_ch_36_ARSIZE = edge_list_ch_36__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_36_ARVALID = edge_list_ch_36__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_36_AWADDR = edge_list_ch_36__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_36_AWBURST = edge_list_ch_36__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_36_AWCACHE = edge_list_ch_36__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_36_AWID = edge_list_ch_36__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_36_AWLEN = edge_list_ch_36__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_36_AWLOCK = edge_list_ch_36__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_36_AWPROT = edge_list_ch_36__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_36_AWQOS = edge_list_ch_36__m_axi_m_axi_AWQOS;
  assign edge_list_ch_36__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_36_AWREADY;
  assign m_axi_edge_list_ch_36_AWSIZE = edge_list_ch_36__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_36_AWVALID = edge_list_ch_36__m_axi_m_axi_AWVALID;
  assign edge_list_ch_36__m_axi_m_axi_BID = m_axi_edge_list_ch_36_BID;
  assign m_axi_edge_list_ch_36_BREADY = edge_list_ch_36__m_axi_m_axi_BREADY;
  assign edge_list_ch_36__m_axi_m_axi_BRESP = m_axi_edge_list_ch_36_BRESP;
  assign edge_list_ch_36__m_axi_m_axi_BVALID = m_axi_edge_list_ch_36_BVALID;
  assign edge_list_ch_36__m_axi_m_axi_RDATA = m_axi_edge_list_ch_36_RDATA;
  assign edge_list_ch_36__m_axi_m_axi_RID = m_axi_edge_list_ch_36_RID;
  assign edge_list_ch_36__m_axi_m_axi_RLAST = m_axi_edge_list_ch_36_RLAST;
  assign m_axi_edge_list_ch_36_RREADY = edge_list_ch_36__m_axi_m_axi_RREADY;
  assign edge_list_ch_36__m_axi_m_axi_RRESP = m_axi_edge_list_ch_36_RRESP;
  assign edge_list_ch_36__m_axi_m_axi_RVALID = m_axi_edge_list_ch_36_RVALID;
  assign m_axi_edge_list_ch_36_WDATA = edge_list_ch_36__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_36_WLAST = edge_list_ch_36__m_axi_m_axi_WLAST;
  assign edge_list_ch_36__m_axi_m_axi_WREADY = m_axi_edge_list_ch_36_WREADY;
  assign m_axi_edge_list_ch_36_WSTRB = edge_list_ch_36__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_36_WVALID = edge_list_ch_36__m_axi_m_axi_WVALID;
  assign edge_list_ch_36__m_axi_read_addr_din = edge_list_ch_36_read_addr__din;
  assign edge_list_ch_36_read_addr__full_n = edge_list_ch_36__m_axi_read_addr_full_n;
  assign edge_list_ch_36__m_axi_read_addr_write = edge_list_ch_36_read_addr__write;
  assign edge_list_ch_36_read_data__dout = edge_list_ch_36__m_axi_read_data_dout;
  assign edge_list_ch_36_read_data__empty_n = edge_list_ch_36__m_axi_read_data_empty_n;
  assign edge_list_ch_36__m_axi_read_data_read = edge_list_ch_36_read_data__read;
  assign edge_list_ch_36__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_36__m_axi_write_addr_din = edge_list_ch_36_write_addr__din;
  assign edge_list_ch_36_write_addr__full_n = edge_list_ch_36__m_axi_write_addr_full_n;
  assign edge_list_ch_36__m_axi_write_addr_write = edge_list_ch_36_write_addr__write;
  assign edge_list_ch_36__m_axi_write_data_din = edge_list_ch_36_write_data__din;
  assign edge_list_ch_36_write_data__full_n = edge_list_ch_36__m_axi_write_data_full_n;
  assign edge_list_ch_36__m_axi_write_data_write = edge_list_ch_36_write_data__write;
  assign edge_list_ch_36_write_resp__dout = edge_list_ch_36__m_axi_write_resp_dout;
  assign edge_list_ch_36_write_resp__empty_n = edge_list_ch_36__m_axi_write_resp_empty_n;
  assign edge_list_ch_36__m_axi_write_resp_read = edge_list_ch_36_write_resp__read;
  assign edge_list_ch_37__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_37_ARADDR = edge_list_ch_37__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_37_ARBURST = edge_list_ch_37__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_37_ARCACHE = edge_list_ch_37__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_37_ARID = edge_list_ch_37__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_37_ARLEN = edge_list_ch_37__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_37_ARLOCK = edge_list_ch_37__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_37_ARPROT = edge_list_ch_37__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_37_ARQOS = edge_list_ch_37__m_axi_m_axi_ARQOS;
  assign edge_list_ch_37__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_37_ARREADY;
  assign m_axi_edge_list_ch_37_ARSIZE = edge_list_ch_37__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_37_ARVALID = edge_list_ch_37__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_37_AWADDR = edge_list_ch_37__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_37_AWBURST = edge_list_ch_37__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_37_AWCACHE = edge_list_ch_37__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_37_AWID = edge_list_ch_37__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_37_AWLEN = edge_list_ch_37__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_37_AWLOCK = edge_list_ch_37__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_37_AWPROT = edge_list_ch_37__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_37_AWQOS = edge_list_ch_37__m_axi_m_axi_AWQOS;
  assign edge_list_ch_37__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_37_AWREADY;
  assign m_axi_edge_list_ch_37_AWSIZE = edge_list_ch_37__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_37_AWVALID = edge_list_ch_37__m_axi_m_axi_AWVALID;
  assign edge_list_ch_37__m_axi_m_axi_BID = m_axi_edge_list_ch_37_BID;
  assign m_axi_edge_list_ch_37_BREADY = edge_list_ch_37__m_axi_m_axi_BREADY;
  assign edge_list_ch_37__m_axi_m_axi_BRESP = m_axi_edge_list_ch_37_BRESP;
  assign edge_list_ch_37__m_axi_m_axi_BVALID = m_axi_edge_list_ch_37_BVALID;
  assign edge_list_ch_37__m_axi_m_axi_RDATA = m_axi_edge_list_ch_37_RDATA;
  assign edge_list_ch_37__m_axi_m_axi_RID = m_axi_edge_list_ch_37_RID;
  assign edge_list_ch_37__m_axi_m_axi_RLAST = m_axi_edge_list_ch_37_RLAST;
  assign m_axi_edge_list_ch_37_RREADY = edge_list_ch_37__m_axi_m_axi_RREADY;
  assign edge_list_ch_37__m_axi_m_axi_RRESP = m_axi_edge_list_ch_37_RRESP;
  assign edge_list_ch_37__m_axi_m_axi_RVALID = m_axi_edge_list_ch_37_RVALID;
  assign m_axi_edge_list_ch_37_WDATA = edge_list_ch_37__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_37_WLAST = edge_list_ch_37__m_axi_m_axi_WLAST;
  assign edge_list_ch_37__m_axi_m_axi_WREADY = m_axi_edge_list_ch_37_WREADY;
  assign m_axi_edge_list_ch_37_WSTRB = edge_list_ch_37__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_37_WVALID = edge_list_ch_37__m_axi_m_axi_WVALID;
  assign edge_list_ch_37__m_axi_read_addr_din = edge_list_ch_37_read_addr__din;
  assign edge_list_ch_37_read_addr__full_n = edge_list_ch_37__m_axi_read_addr_full_n;
  assign edge_list_ch_37__m_axi_read_addr_write = edge_list_ch_37_read_addr__write;
  assign edge_list_ch_37_read_data__dout = edge_list_ch_37__m_axi_read_data_dout;
  assign edge_list_ch_37_read_data__empty_n = edge_list_ch_37__m_axi_read_data_empty_n;
  assign edge_list_ch_37__m_axi_read_data_read = edge_list_ch_37_read_data__read;
  assign edge_list_ch_37__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_37__m_axi_write_addr_din = edge_list_ch_37_write_addr__din;
  assign edge_list_ch_37_write_addr__full_n = edge_list_ch_37__m_axi_write_addr_full_n;
  assign edge_list_ch_37__m_axi_write_addr_write = edge_list_ch_37_write_addr__write;
  assign edge_list_ch_37__m_axi_write_data_din = edge_list_ch_37_write_data__din;
  assign edge_list_ch_37_write_data__full_n = edge_list_ch_37__m_axi_write_data_full_n;
  assign edge_list_ch_37__m_axi_write_data_write = edge_list_ch_37_write_data__write;
  assign edge_list_ch_37_write_resp__dout = edge_list_ch_37__m_axi_write_resp_dout;
  assign edge_list_ch_37_write_resp__empty_n = edge_list_ch_37__m_axi_write_resp_empty_n;
  assign edge_list_ch_37__m_axi_write_resp_read = edge_list_ch_37_write_resp__read;
  assign edge_list_ch_38__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_38_ARADDR = edge_list_ch_38__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_38_ARBURST = edge_list_ch_38__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_38_ARCACHE = edge_list_ch_38__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_38_ARID = edge_list_ch_38__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_38_ARLEN = edge_list_ch_38__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_38_ARLOCK = edge_list_ch_38__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_38_ARPROT = edge_list_ch_38__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_38_ARQOS = edge_list_ch_38__m_axi_m_axi_ARQOS;
  assign edge_list_ch_38__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_38_ARREADY;
  assign m_axi_edge_list_ch_38_ARSIZE = edge_list_ch_38__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_38_ARVALID = edge_list_ch_38__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_38_AWADDR = edge_list_ch_38__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_38_AWBURST = edge_list_ch_38__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_38_AWCACHE = edge_list_ch_38__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_38_AWID = edge_list_ch_38__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_38_AWLEN = edge_list_ch_38__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_38_AWLOCK = edge_list_ch_38__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_38_AWPROT = edge_list_ch_38__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_38_AWQOS = edge_list_ch_38__m_axi_m_axi_AWQOS;
  assign edge_list_ch_38__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_38_AWREADY;
  assign m_axi_edge_list_ch_38_AWSIZE = edge_list_ch_38__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_38_AWVALID = edge_list_ch_38__m_axi_m_axi_AWVALID;
  assign edge_list_ch_38__m_axi_m_axi_BID = m_axi_edge_list_ch_38_BID;
  assign m_axi_edge_list_ch_38_BREADY = edge_list_ch_38__m_axi_m_axi_BREADY;
  assign edge_list_ch_38__m_axi_m_axi_BRESP = m_axi_edge_list_ch_38_BRESP;
  assign edge_list_ch_38__m_axi_m_axi_BVALID = m_axi_edge_list_ch_38_BVALID;
  assign edge_list_ch_38__m_axi_m_axi_RDATA = m_axi_edge_list_ch_38_RDATA;
  assign edge_list_ch_38__m_axi_m_axi_RID = m_axi_edge_list_ch_38_RID;
  assign edge_list_ch_38__m_axi_m_axi_RLAST = m_axi_edge_list_ch_38_RLAST;
  assign m_axi_edge_list_ch_38_RREADY = edge_list_ch_38__m_axi_m_axi_RREADY;
  assign edge_list_ch_38__m_axi_m_axi_RRESP = m_axi_edge_list_ch_38_RRESP;
  assign edge_list_ch_38__m_axi_m_axi_RVALID = m_axi_edge_list_ch_38_RVALID;
  assign m_axi_edge_list_ch_38_WDATA = edge_list_ch_38__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_38_WLAST = edge_list_ch_38__m_axi_m_axi_WLAST;
  assign edge_list_ch_38__m_axi_m_axi_WREADY = m_axi_edge_list_ch_38_WREADY;
  assign m_axi_edge_list_ch_38_WSTRB = edge_list_ch_38__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_38_WVALID = edge_list_ch_38__m_axi_m_axi_WVALID;
  assign edge_list_ch_38__m_axi_read_addr_din = edge_list_ch_38_read_addr__din;
  assign edge_list_ch_38_read_addr__full_n = edge_list_ch_38__m_axi_read_addr_full_n;
  assign edge_list_ch_38__m_axi_read_addr_write = edge_list_ch_38_read_addr__write;
  assign edge_list_ch_38_read_data__dout = edge_list_ch_38__m_axi_read_data_dout;
  assign edge_list_ch_38_read_data__empty_n = edge_list_ch_38__m_axi_read_data_empty_n;
  assign edge_list_ch_38__m_axi_read_data_read = edge_list_ch_38_read_data__read;
  assign edge_list_ch_38__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_38__m_axi_write_addr_din = edge_list_ch_38_write_addr__din;
  assign edge_list_ch_38_write_addr__full_n = edge_list_ch_38__m_axi_write_addr_full_n;
  assign edge_list_ch_38__m_axi_write_addr_write = edge_list_ch_38_write_addr__write;
  assign edge_list_ch_38__m_axi_write_data_din = edge_list_ch_38_write_data__din;
  assign edge_list_ch_38_write_data__full_n = edge_list_ch_38__m_axi_write_data_full_n;
  assign edge_list_ch_38__m_axi_write_data_write = edge_list_ch_38_write_data__write;
  assign edge_list_ch_38_write_resp__dout = edge_list_ch_38__m_axi_write_resp_dout;
  assign edge_list_ch_38_write_resp__empty_n = edge_list_ch_38__m_axi_write_resp_empty_n;
  assign edge_list_ch_38__m_axi_write_resp_read = edge_list_ch_38_write_resp__read;
  assign edge_list_ch_39__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_39_ARADDR = edge_list_ch_39__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_39_ARBURST = edge_list_ch_39__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_39_ARCACHE = edge_list_ch_39__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_39_ARID = edge_list_ch_39__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_39_ARLEN = edge_list_ch_39__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_39_ARLOCK = edge_list_ch_39__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_39_ARPROT = edge_list_ch_39__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_39_ARQOS = edge_list_ch_39__m_axi_m_axi_ARQOS;
  assign edge_list_ch_39__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_39_ARREADY;
  assign m_axi_edge_list_ch_39_ARSIZE = edge_list_ch_39__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_39_ARVALID = edge_list_ch_39__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_39_AWADDR = edge_list_ch_39__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_39_AWBURST = edge_list_ch_39__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_39_AWCACHE = edge_list_ch_39__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_39_AWID = edge_list_ch_39__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_39_AWLEN = edge_list_ch_39__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_39_AWLOCK = edge_list_ch_39__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_39_AWPROT = edge_list_ch_39__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_39_AWQOS = edge_list_ch_39__m_axi_m_axi_AWQOS;
  assign edge_list_ch_39__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_39_AWREADY;
  assign m_axi_edge_list_ch_39_AWSIZE = edge_list_ch_39__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_39_AWVALID = edge_list_ch_39__m_axi_m_axi_AWVALID;
  assign edge_list_ch_39__m_axi_m_axi_BID = m_axi_edge_list_ch_39_BID;
  assign m_axi_edge_list_ch_39_BREADY = edge_list_ch_39__m_axi_m_axi_BREADY;
  assign edge_list_ch_39__m_axi_m_axi_BRESP = m_axi_edge_list_ch_39_BRESP;
  assign edge_list_ch_39__m_axi_m_axi_BVALID = m_axi_edge_list_ch_39_BVALID;
  assign edge_list_ch_39__m_axi_m_axi_RDATA = m_axi_edge_list_ch_39_RDATA;
  assign edge_list_ch_39__m_axi_m_axi_RID = m_axi_edge_list_ch_39_RID;
  assign edge_list_ch_39__m_axi_m_axi_RLAST = m_axi_edge_list_ch_39_RLAST;
  assign m_axi_edge_list_ch_39_RREADY = edge_list_ch_39__m_axi_m_axi_RREADY;
  assign edge_list_ch_39__m_axi_m_axi_RRESP = m_axi_edge_list_ch_39_RRESP;
  assign edge_list_ch_39__m_axi_m_axi_RVALID = m_axi_edge_list_ch_39_RVALID;
  assign m_axi_edge_list_ch_39_WDATA = edge_list_ch_39__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_39_WLAST = edge_list_ch_39__m_axi_m_axi_WLAST;
  assign edge_list_ch_39__m_axi_m_axi_WREADY = m_axi_edge_list_ch_39_WREADY;
  assign m_axi_edge_list_ch_39_WSTRB = edge_list_ch_39__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_39_WVALID = edge_list_ch_39__m_axi_m_axi_WVALID;
  assign edge_list_ch_39__m_axi_read_addr_din = edge_list_ch_39_read_addr__din;
  assign edge_list_ch_39_read_addr__full_n = edge_list_ch_39__m_axi_read_addr_full_n;
  assign edge_list_ch_39__m_axi_read_addr_write = edge_list_ch_39_read_addr__write;
  assign edge_list_ch_39_read_data__dout = edge_list_ch_39__m_axi_read_data_dout;
  assign edge_list_ch_39_read_data__empty_n = edge_list_ch_39__m_axi_read_data_empty_n;
  assign edge_list_ch_39__m_axi_read_data_read = edge_list_ch_39_read_data__read;
  assign edge_list_ch_39__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_39__m_axi_write_addr_din = edge_list_ch_39_write_addr__din;
  assign edge_list_ch_39_write_addr__full_n = edge_list_ch_39__m_axi_write_addr_full_n;
  assign edge_list_ch_39__m_axi_write_addr_write = edge_list_ch_39_write_addr__write;
  assign edge_list_ch_39__m_axi_write_data_din = edge_list_ch_39_write_data__din;
  assign edge_list_ch_39_write_data__full_n = edge_list_ch_39__m_axi_write_data_full_n;
  assign edge_list_ch_39__m_axi_write_data_write = edge_list_ch_39_write_data__write;
  assign edge_list_ch_39_write_resp__dout = edge_list_ch_39__m_axi_write_resp_dout;
  assign edge_list_ch_39_write_resp__empty_n = edge_list_ch_39__m_axi_write_resp_empty_n;
  assign edge_list_ch_39__m_axi_write_resp_read = edge_list_ch_39_write_resp__read;
  assign edge_list_ch_40__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_40_ARADDR = edge_list_ch_40__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_40_ARBURST = edge_list_ch_40__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_40_ARCACHE = edge_list_ch_40__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_40_ARID = edge_list_ch_40__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_40_ARLEN = edge_list_ch_40__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_40_ARLOCK = edge_list_ch_40__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_40_ARPROT = edge_list_ch_40__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_40_ARQOS = edge_list_ch_40__m_axi_m_axi_ARQOS;
  assign edge_list_ch_40__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_40_ARREADY;
  assign m_axi_edge_list_ch_40_ARSIZE = edge_list_ch_40__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_40_ARVALID = edge_list_ch_40__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_40_AWADDR = edge_list_ch_40__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_40_AWBURST = edge_list_ch_40__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_40_AWCACHE = edge_list_ch_40__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_40_AWID = edge_list_ch_40__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_40_AWLEN = edge_list_ch_40__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_40_AWLOCK = edge_list_ch_40__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_40_AWPROT = edge_list_ch_40__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_40_AWQOS = edge_list_ch_40__m_axi_m_axi_AWQOS;
  assign edge_list_ch_40__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_40_AWREADY;
  assign m_axi_edge_list_ch_40_AWSIZE = edge_list_ch_40__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_40_AWVALID = edge_list_ch_40__m_axi_m_axi_AWVALID;
  assign edge_list_ch_40__m_axi_m_axi_BID = m_axi_edge_list_ch_40_BID;
  assign m_axi_edge_list_ch_40_BREADY = edge_list_ch_40__m_axi_m_axi_BREADY;
  assign edge_list_ch_40__m_axi_m_axi_BRESP = m_axi_edge_list_ch_40_BRESP;
  assign edge_list_ch_40__m_axi_m_axi_BVALID = m_axi_edge_list_ch_40_BVALID;
  assign edge_list_ch_40__m_axi_m_axi_RDATA = m_axi_edge_list_ch_40_RDATA;
  assign edge_list_ch_40__m_axi_m_axi_RID = m_axi_edge_list_ch_40_RID;
  assign edge_list_ch_40__m_axi_m_axi_RLAST = m_axi_edge_list_ch_40_RLAST;
  assign m_axi_edge_list_ch_40_RREADY = edge_list_ch_40__m_axi_m_axi_RREADY;
  assign edge_list_ch_40__m_axi_m_axi_RRESP = m_axi_edge_list_ch_40_RRESP;
  assign edge_list_ch_40__m_axi_m_axi_RVALID = m_axi_edge_list_ch_40_RVALID;
  assign m_axi_edge_list_ch_40_WDATA = edge_list_ch_40__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_40_WLAST = edge_list_ch_40__m_axi_m_axi_WLAST;
  assign edge_list_ch_40__m_axi_m_axi_WREADY = m_axi_edge_list_ch_40_WREADY;
  assign m_axi_edge_list_ch_40_WSTRB = edge_list_ch_40__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_40_WVALID = edge_list_ch_40__m_axi_m_axi_WVALID;
  assign edge_list_ch_40__m_axi_read_addr_din = edge_list_ch_40_read_addr__din;
  assign edge_list_ch_40_read_addr__full_n = edge_list_ch_40__m_axi_read_addr_full_n;
  assign edge_list_ch_40__m_axi_read_addr_write = edge_list_ch_40_read_addr__write;
  assign edge_list_ch_40_read_data__dout = edge_list_ch_40__m_axi_read_data_dout;
  assign edge_list_ch_40_read_data__empty_n = edge_list_ch_40__m_axi_read_data_empty_n;
  assign edge_list_ch_40__m_axi_read_data_read = edge_list_ch_40_read_data__read;
  assign edge_list_ch_40__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_40__m_axi_write_addr_din = edge_list_ch_40_write_addr__din;
  assign edge_list_ch_40_write_addr__full_n = edge_list_ch_40__m_axi_write_addr_full_n;
  assign edge_list_ch_40__m_axi_write_addr_write = edge_list_ch_40_write_addr__write;
  assign edge_list_ch_40__m_axi_write_data_din = edge_list_ch_40_write_data__din;
  assign edge_list_ch_40_write_data__full_n = edge_list_ch_40__m_axi_write_data_full_n;
  assign edge_list_ch_40__m_axi_write_data_write = edge_list_ch_40_write_data__write;
  assign edge_list_ch_40_write_resp__dout = edge_list_ch_40__m_axi_write_resp_dout;
  assign edge_list_ch_40_write_resp__empty_n = edge_list_ch_40__m_axi_write_resp_empty_n;
  assign edge_list_ch_40__m_axi_write_resp_read = edge_list_ch_40_write_resp__read;
  assign edge_list_ch_41__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_41_ARADDR = edge_list_ch_41__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_41_ARBURST = edge_list_ch_41__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_41_ARCACHE = edge_list_ch_41__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_41_ARID = edge_list_ch_41__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_41_ARLEN = edge_list_ch_41__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_41_ARLOCK = edge_list_ch_41__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_41_ARPROT = edge_list_ch_41__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_41_ARQOS = edge_list_ch_41__m_axi_m_axi_ARQOS;
  assign edge_list_ch_41__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_41_ARREADY;
  assign m_axi_edge_list_ch_41_ARSIZE = edge_list_ch_41__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_41_ARVALID = edge_list_ch_41__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_41_AWADDR = edge_list_ch_41__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_41_AWBURST = edge_list_ch_41__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_41_AWCACHE = edge_list_ch_41__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_41_AWID = edge_list_ch_41__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_41_AWLEN = edge_list_ch_41__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_41_AWLOCK = edge_list_ch_41__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_41_AWPROT = edge_list_ch_41__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_41_AWQOS = edge_list_ch_41__m_axi_m_axi_AWQOS;
  assign edge_list_ch_41__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_41_AWREADY;
  assign m_axi_edge_list_ch_41_AWSIZE = edge_list_ch_41__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_41_AWVALID = edge_list_ch_41__m_axi_m_axi_AWVALID;
  assign edge_list_ch_41__m_axi_m_axi_BID = m_axi_edge_list_ch_41_BID;
  assign m_axi_edge_list_ch_41_BREADY = edge_list_ch_41__m_axi_m_axi_BREADY;
  assign edge_list_ch_41__m_axi_m_axi_BRESP = m_axi_edge_list_ch_41_BRESP;
  assign edge_list_ch_41__m_axi_m_axi_BVALID = m_axi_edge_list_ch_41_BVALID;
  assign edge_list_ch_41__m_axi_m_axi_RDATA = m_axi_edge_list_ch_41_RDATA;
  assign edge_list_ch_41__m_axi_m_axi_RID = m_axi_edge_list_ch_41_RID;
  assign edge_list_ch_41__m_axi_m_axi_RLAST = m_axi_edge_list_ch_41_RLAST;
  assign m_axi_edge_list_ch_41_RREADY = edge_list_ch_41__m_axi_m_axi_RREADY;
  assign edge_list_ch_41__m_axi_m_axi_RRESP = m_axi_edge_list_ch_41_RRESP;
  assign edge_list_ch_41__m_axi_m_axi_RVALID = m_axi_edge_list_ch_41_RVALID;
  assign m_axi_edge_list_ch_41_WDATA = edge_list_ch_41__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_41_WLAST = edge_list_ch_41__m_axi_m_axi_WLAST;
  assign edge_list_ch_41__m_axi_m_axi_WREADY = m_axi_edge_list_ch_41_WREADY;
  assign m_axi_edge_list_ch_41_WSTRB = edge_list_ch_41__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_41_WVALID = edge_list_ch_41__m_axi_m_axi_WVALID;
  assign edge_list_ch_41__m_axi_read_addr_din = edge_list_ch_41_read_addr__din;
  assign edge_list_ch_41_read_addr__full_n = edge_list_ch_41__m_axi_read_addr_full_n;
  assign edge_list_ch_41__m_axi_read_addr_write = edge_list_ch_41_read_addr__write;
  assign edge_list_ch_41_read_data__dout = edge_list_ch_41__m_axi_read_data_dout;
  assign edge_list_ch_41_read_data__empty_n = edge_list_ch_41__m_axi_read_data_empty_n;
  assign edge_list_ch_41__m_axi_read_data_read = edge_list_ch_41_read_data__read;
  assign edge_list_ch_41__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_41__m_axi_write_addr_din = edge_list_ch_41_write_addr__din;
  assign edge_list_ch_41_write_addr__full_n = edge_list_ch_41__m_axi_write_addr_full_n;
  assign edge_list_ch_41__m_axi_write_addr_write = edge_list_ch_41_write_addr__write;
  assign edge_list_ch_41__m_axi_write_data_din = edge_list_ch_41_write_data__din;
  assign edge_list_ch_41_write_data__full_n = edge_list_ch_41__m_axi_write_data_full_n;
  assign edge_list_ch_41__m_axi_write_data_write = edge_list_ch_41_write_data__write;
  assign edge_list_ch_41_write_resp__dout = edge_list_ch_41__m_axi_write_resp_dout;
  assign edge_list_ch_41_write_resp__empty_n = edge_list_ch_41__m_axi_write_resp_empty_n;
  assign edge_list_ch_41__m_axi_write_resp_read = edge_list_ch_41_write_resp__read;
  assign edge_list_ch_42__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_42_ARADDR = edge_list_ch_42__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_42_ARBURST = edge_list_ch_42__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_42_ARCACHE = edge_list_ch_42__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_42_ARID = edge_list_ch_42__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_42_ARLEN = edge_list_ch_42__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_42_ARLOCK = edge_list_ch_42__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_42_ARPROT = edge_list_ch_42__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_42_ARQOS = edge_list_ch_42__m_axi_m_axi_ARQOS;
  assign edge_list_ch_42__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_42_ARREADY;
  assign m_axi_edge_list_ch_42_ARSIZE = edge_list_ch_42__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_42_ARVALID = edge_list_ch_42__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_42_AWADDR = edge_list_ch_42__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_42_AWBURST = edge_list_ch_42__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_42_AWCACHE = edge_list_ch_42__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_42_AWID = edge_list_ch_42__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_42_AWLEN = edge_list_ch_42__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_42_AWLOCK = edge_list_ch_42__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_42_AWPROT = edge_list_ch_42__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_42_AWQOS = edge_list_ch_42__m_axi_m_axi_AWQOS;
  assign edge_list_ch_42__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_42_AWREADY;
  assign m_axi_edge_list_ch_42_AWSIZE = edge_list_ch_42__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_42_AWVALID = edge_list_ch_42__m_axi_m_axi_AWVALID;
  assign edge_list_ch_42__m_axi_m_axi_BID = m_axi_edge_list_ch_42_BID;
  assign m_axi_edge_list_ch_42_BREADY = edge_list_ch_42__m_axi_m_axi_BREADY;
  assign edge_list_ch_42__m_axi_m_axi_BRESP = m_axi_edge_list_ch_42_BRESP;
  assign edge_list_ch_42__m_axi_m_axi_BVALID = m_axi_edge_list_ch_42_BVALID;
  assign edge_list_ch_42__m_axi_m_axi_RDATA = m_axi_edge_list_ch_42_RDATA;
  assign edge_list_ch_42__m_axi_m_axi_RID = m_axi_edge_list_ch_42_RID;
  assign edge_list_ch_42__m_axi_m_axi_RLAST = m_axi_edge_list_ch_42_RLAST;
  assign m_axi_edge_list_ch_42_RREADY = edge_list_ch_42__m_axi_m_axi_RREADY;
  assign edge_list_ch_42__m_axi_m_axi_RRESP = m_axi_edge_list_ch_42_RRESP;
  assign edge_list_ch_42__m_axi_m_axi_RVALID = m_axi_edge_list_ch_42_RVALID;
  assign m_axi_edge_list_ch_42_WDATA = edge_list_ch_42__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_42_WLAST = edge_list_ch_42__m_axi_m_axi_WLAST;
  assign edge_list_ch_42__m_axi_m_axi_WREADY = m_axi_edge_list_ch_42_WREADY;
  assign m_axi_edge_list_ch_42_WSTRB = edge_list_ch_42__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_42_WVALID = edge_list_ch_42__m_axi_m_axi_WVALID;
  assign edge_list_ch_42__m_axi_read_addr_din = edge_list_ch_42_read_addr__din;
  assign edge_list_ch_42_read_addr__full_n = edge_list_ch_42__m_axi_read_addr_full_n;
  assign edge_list_ch_42__m_axi_read_addr_write = edge_list_ch_42_read_addr__write;
  assign edge_list_ch_42_read_data__dout = edge_list_ch_42__m_axi_read_data_dout;
  assign edge_list_ch_42_read_data__empty_n = edge_list_ch_42__m_axi_read_data_empty_n;
  assign edge_list_ch_42__m_axi_read_data_read = edge_list_ch_42_read_data__read;
  assign edge_list_ch_42__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_42__m_axi_write_addr_din = edge_list_ch_42_write_addr__din;
  assign edge_list_ch_42_write_addr__full_n = edge_list_ch_42__m_axi_write_addr_full_n;
  assign edge_list_ch_42__m_axi_write_addr_write = edge_list_ch_42_write_addr__write;
  assign edge_list_ch_42__m_axi_write_data_din = edge_list_ch_42_write_data__din;
  assign edge_list_ch_42_write_data__full_n = edge_list_ch_42__m_axi_write_data_full_n;
  assign edge_list_ch_42__m_axi_write_data_write = edge_list_ch_42_write_data__write;
  assign edge_list_ch_42_write_resp__dout = edge_list_ch_42__m_axi_write_resp_dout;
  assign edge_list_ch_42_write_resp__empty_n = edge_list_ch_42__m_axi_write_resp_empty_n;
  assign edge_list_ch_42__m_axi_write_resp_read = edge_list_ch_42_write_resp__read;
  assign edge_list_ch_43__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_43_ARADDR = edge_list_ch_43__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_43_ARBURST = edge_list_ch_43__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_43_ARCACHE = edge_list_ch_43__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_43_ARID = edge_list_ch_43__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_43_ARLEN = edge_list_ch_43__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_43_ARLOCK = edge_list_ch_43__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_43_ARPROT = edge_list_ch_43__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_43_ARQOS = edge_list_ch_43__m_axi_m_axi_ARQOS;
  assign edge_list_ch_43__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_43_ARREADY;
  assign m_axi_edge_list_ch_43_ARSIZE = edge_list_ch_43__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_43_ARVALID = edge_list_ch_43__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_43_AWADDR = edge_list_ch_43__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_43_AWBURST = edge_list_ch_43__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_43_AWCACHE = edge_list_ch_43__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_43_AWID = edge_list_ch_43__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_43_AWLEN = edge_list_ch_43__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_43_AWLOCK = edge_list_ch_43__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_43_AWPROT = edge_list_ch_43__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_43_AWQOS = edge_list_ch_43__m_axi_m_axi_AWQOS;
  assign edge_list_ch_43__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_43_AWREADY;
  assign m_axi_edge_list_ch_43_AWSIZE = edge_list_ch_43__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_43_AWVALID = edge_list_ch_43__m_axi_m_axi_AWVALID;
  assign edge_list_ch_43__m_axi_m_axi_BID = m_axi_edge_list_ch_43_BID;
  assign m_axi_edge_list_ch_43_BREADY = edge_list_ch_43__m_axi_m_axi_BREADY;
  assign edge_list_ch_43__m_axi_m_axi_BRESP = m_axi_edge_list_ch_43_BRESP;
  assign edge_list_ch_43__m_axi_m_axi_BVALID = m_axi_edge_list_ch_43_BVALID;
  assign edge_list_ch_43__m_axi_m_axi_RDATA = m_axi_edge_list_ch_43_RDATA;
  assign edge_list_ch_43__m_axi_m_axi_RID = m_axi_edge_list_ch_43_RID;
  assign edge_list_ch_43__m_axi_m_axi_RLAST = m_axi_edge_list_ch_43_RLAST;
  assign m_axi_edge_list_ch_43_RREADY = edge_list_ch_43__m_axi_m_axi_RREADY;
  assign edge_list_ch_43__m_axi_m_axi_RRESP = m_axi_edge_list_ch_43_RRESP;
  assign edge_list_ch_43__m_axi_m_axi_RVALID = m_axi_edge_list_ch_43_RVALID;
  assign m_axi_edge_list_ch_43_WDATA = edge_list_ch_43__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_43_WLAST = edge_list_ch_43__m_axi_m_axi_WLAST;
  assign edge_list_ch_43__m_axi_m_axi_WREADY = m_axi_edge_list_ch_43_WREADY;
  assign m_axi_edge_list_ch_43_WSTRB = edge_list_ch_43__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_43_WVALID = edge_list_ch_43__m_axi_m_axi_WVALID;
  assign edge_list_ch_43__m_axi_read_addr_din = edge_list_ch_43_read_addr__din;
  assign edge_list_ch_43_read_addr__full_n = edge_list_ch_43__m_axi_read_addr_full_n;
  assign edge_list_ch_43__m_axi_read_addr_write = edge_list_ch_43_read_addr__write;
  assign edge_list_ch_43_read_data__dout = edge_list_ch_43__m_axi_read_data_dout;
  assign edge_list_ch_43_read_data__empty_n = edge_list_ch_43__m_axi_read_data_empty_n;
  assign edge_list_ch_43__m_axi_read_data_read = edge_list_ch_43_read_data__read;
  assign edge_list_ch_43__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_43__m_axi_write_addr_din = edge_list_ch_43_write_addr__din;
  assign edge_list_ch_43_write_addr__full_n = edge_list_ch_43__m_axi_write_addr_full_n;
  assign edge_list_ch_43__m_axi_write_addr_write = edge_list_ch_43_write_addr__write;
  assign edge_list_ch_43__m_axi_write_data_din = edge_list_ch_43_write_data__din;
  assign edge_list_ch_43_write_data__full_n = edge_list_ch_43__m_axi_write_data_full_n;
  assign edge_list_ch_43__m_axi_write_data_write = edge_list_ch_43_write_data__write;
  assign edge_list_ch_43_write_resp__dout = edge_list_ch_43__m_axi_write_resp_dout;
  assign edge_list_ch_43_write_resp__empty_n = edge_list_ch_43__m_axi_write_resp_empty_n;
  assign edge_list_ch_43__m_axi_write_resp_read = edge_list_ch_43_write_resp__read;
  assign edge_list_ch_44__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_44_ARADDR = edge_list_ch_44__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_44_ARBURST = edge_list_ch_44__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_44_ARCACHE = edge_list_ch_44__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_44_ARID = edge_list_ch_44__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_44_ARLEN = edge_list_ch_44__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_44_ARLOCK = edge_list_ch_44__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_44_ARPROT = edge_list_ch_44__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_44_ARQOS = edge_list_ch_44__m_axi_m_axi_ARQOS;
  assign edge_list_ch_44__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_44_ARREADY;
  assign m_axi_edge_list_ch_44_ARSIZE = edge_list_ch_44__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_44_ARVALID = edge_list_ch_44__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_44_AWADDR = edge_list_ch_44__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_44_AWBURST = edge_list_ch_44__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_44_AWCACHE = edge_list_ch_44__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_44_AWID = edge_list_ch_44__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_44_AWLEN = edge_list_ch_44__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_44_AWLOCK = edge_list_ch_44__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_44_AWPROT = edge_list_ch_44__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_44_AWQOS = edge_list_ch_44__m_axi_m_axi_AWQOS;
  assign edge_list_ch_44__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_44_AWREADY;
  assign m_axi_edge_list_ch_44_AWSIZE = edge_list_ch_44__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_44_AWVALID = edge_list_ch_44__m_axi_m_axi_AWVALID;
  assign edge_list_ch_44__m_axi_m_axi_BID = m_axi_edge_list_ch_44_BID;
  assign m_axi_edge_list_ch_44_BREADY = edge_list_ch_44__m_axi_m_axi_BREADY;
  assign edge_list_ch_44__m_axi_m_axi_BRESP = m_axi_edge_list_ch_44_BRESP;
  assign edge_list_ch_44__m_axi_m_axi_BVALID = m_axi_edge_list_ch_44_BVALID;
  assign edge_list_ch_44__m_axi_m_axi_RDATA = m_axi_edge_list_ch_44_RDATA;
  assign edge_list_ch_44__m_axi_m_axi_RID = m_axi_edge_list_ch_44_RID;
  assign edge_list_ch_44__m_axi_m_axi_RLAST = m_axi_edge_list_ch_44_RLAST;
  assign m_axi_edge_list_ch_44_RREADY = edge_list_ch_44__m_axi_m_axi_RREADY;
  assign edge_list_ch_44__m_axi_m_axi_RRESP = m_axi_edge_list_ch_44_RRESP;
  assign edge_list_ch_44__m_axi_m_axi_RVALID = m_axi_edge_list_ch_44_RVALID;
  assign m_axi_edge_list_ch_44_WDATA = edge_list_ch_44__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_44_WLAST = edge_list_ch_44__m_axi_m_axi_WLAST;
  assign edge_list_ch_44__m_axi_m_axi_WREADY = m_axi_edge_list_ch_44_WREADY;
  assign m_axi_edge_list_ch_44_WSTRB = edge_list_ch_44__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_44_WVALID = edge_list_ch_44__m_axi_m_axi_WVALID;
  assign edge_list_ch_44__m_axi_read_addr_din = edge_list_ch_44_read_addr__din;
  assign edge_list_ch_44_read_addr__full_n = edge_list_ch_44__m_axi_read_addr_full_n;
  assign edge_list_ch_44__m_axi_read_addr_write = edge_list_ch_44_read_addr__write;
  assign edge_list_ch_44_read_data__dout = edge_list_ch_44__m_axi_read_data_dout;
  assign edge_list_ch_44_read_data__empty_n = edge_list_ch_44__m_axi_read_data_empty_n;
  assign edge_list_ch_44__m_axi_read_data_read = edge_list_ch_44_read_data__read;
  assign edge_list_ch_44__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_44__m_axi_write_addr_din = edge_list_ch_44_write_addr__din;
  assign edge_list_ch_44_write_addr__full_n = edge_list_ch_44__m_axi_write_addr_full_n;
  assign edge_list_ch_44__m_axi_write_addr_write = edge_list_ch_44_write_addr__write;
  assign edge_list_ch_44__m_axi_write_data_din = edge_list_ch_44_write_data__din;
  assign edge_list_ch_44_write_data__full_n = edge_list_ch_44__m_axi_write_data_full_n;
  assign edge_list_ch_44__m_axi_write_data_write = edge_list_ch_44_write_data__write;
  assign edge_list_ch_44_write_resp__dout = edge_list_ch_44__m_axi_write_resp_dout;
  assign edge_list_ch_44_write_resp__empty_n = edge_list_ch_44__m_axi_write_resp_empty_n;
  assign edge_list_ch_44__m_axi_write_resp_read = edge_list_ch_44_write_resp__read;
  assign edge_list_ch_45__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_45_ARADDR = edge_list_ch_45__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_45_ARBURST = edge_list_ch_45__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_45_ARCACHE = edge_list_ch_45__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_45_ARID = edge_list_ch_45__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_45_ARLEN = edge_list_ch_45__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_45_ARLOCK = edge_list_ch_45__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_45_ARPROT = edge_list_ch_45__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_45_ARQOS = edge_list_ch_45__m_axi_m_axi_ARQOS;
  assign edge_list_ch_45__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_45_ARREADY;
  assign m_axi_edge_list_ch_45_ARSIZE = edge_list_ch_45__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_45_ARVALID = edge_list_ch_45__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_45_AWADDR = edge_list_ch_45__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_45_AWBURST = edge_list_ch_45__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_45_AWCACHE = edge_list_ch_45__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_45_AWID = edge_list_ch_45__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_45_AWLEN = edge_list_ch_45__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_45_AWLOCK = edge_list_ch_45__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_45_AWPROT = edge_list_ch_45__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_45_AWQOS = edge_list_ch_45__m_axi_m_axi_AWQOS;
  assign edge_list_ch_45__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_45_AWREADY;
  assign m_axi_edge_list_ch_45_AWSIZE = edge_list_ch_45__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_45_AWVALID = edge_list_ch_45__m_axi_m_axi_AWVALID;
  assign edge_list_ch_45__m_axi_m_axi_BID = m_axi_edge_list_ch_45_BID;
  assign m_axi_edge_list_ch_45_BREADY = edge_list_ch_45__m_axi_m_axi_BREADY;
  assign edge_list_ch_45__m_axi_m_axi_BRESP = m_axi_edge_list_ch_45_BRESP;
  assign edge_list_ch_45__m_axi_m_axi_BVALID = m_axi_edge_list_ch_45_BVALID;
  assign edge_list_ch_45__m_axi_m_axi_RDATA = m_axi_edge_list_ch_45_RDATA;
  assign edge_list_ch_45__m_axi_m_axi_RID = m_axi_edge_list_ch_45_RID;
  assign edge_list_ch_45__m_axi_m_axi_RLAST = m_axi_edge_list_ch_45_RLAST;
  assign m_axi_edge_list_ch_45_RREADY = edge_list_ch_45__m_axi_m_axi_RREADY;
  assign edge_list_ch_45__m_axi_m_axi_RRESP = m_axi_edge_list_ch_45_RRESP;
  assign edge_list_ch_45__m_axi_m_axi_RVALID = m_axi_edge_list_ch_45_RVALID;
  assign m_axi_edge_list_ch_45_WDATA = edge_list_ch_45__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_45_WLAST = edge_list_ch_45__m_axi_m_axi_WLAST;
  assign edge_list_ch_45__m_axi_m_axi_WREADY = m_axi_edge_list_ch_45_WREADY;
  assign m_axi_edge_list_ch_45_WSTRB = edge_list_ch_45__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_45_WVALID = edge_list_ch_45__m_axi_m_axi_WVALID;
  assign edge_list_ch_45__m_axi_read_addr_din = edge_list_ch_45_read_addr__din;
  assign edge_list_ch_45_read_addr__full_n = edge_list_ch_45__m_axi_read_addr_full_n;
  assign edge_list_ch_45__m_axi_read_addr_write = edge_list_ch_45_read_addr__write;
  assign edge_list_ch_45_read_data__dout = edge_list_ch_45__m_axi_read_data_dout;
  assign edge_list_ch_45_read_data__empty_n = edge_list_ch_45__m_axi_read_data_empty_n;
  assign edge_list_ch_45__m_axi_read_data_read = edge_list_ch_45_read_data__read;
  assign edge_list_ch_45__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_45__m_axi_write_addr_din = edge_list_ch_45_write_addr__din;
  assign edge_list_ch_45_write_addr__full_n = edge_list_ch_45__m_axi_write_addr_full_n;
  assign edge_list_ch_45__m_axi_write_addr_write = edge_list_ch_45_write_addr__write;
  assign edge_list_ch_45__m_axi_write_data_din = edge_list_ch_45_write_data__din;
  assign edge_list_ch_45_write_data__full_n = edge_list_ch_45__m_axi_write_data_full_n;
  assign edge_list_ch_45__m_axi_write_data_write = edge_list_ch_45_write_data__write;
  assign edge_list_ch_45_write_resp__dout = edge_list_ch_45__m_axi_write_resp_dout;
  assign edge_list_ch_45_write_resp__empty_n = edge_list_ch_45__m_axi_write_resp_empty_n;
  assign edge_list_ch_45__m_axi_write_resp_read = edge_list_ch_45_write_resp__read;
  assign edge_list_ch_46__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_46_ARADDR = edge_list_ch_46__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_46_ARBURST = edge_list_ch_46__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_46_ARCACHE = edge_list_ch_46__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_46_ARID = edge_list_ch_46__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_46_ARLEN = edge_list_ch_46__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_46_ARLOCK = edge_list_ch_46__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_46_ARPROT = edge_list_ch_46__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_46_ARQOS = edge_list_ch_46__m_axi_m_axi_ARQOS;
  assign edge_list_ch_46__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_46_ARREADY;
  assign m_axi_edge_list_ch_46_ARSIZE = edge_list_ch_46__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_46_ARVALID = edge_list_ch_46__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_46_AWADDR = edge_list_ch_46__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_46_AWBURST = edge_list_ch_46__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_46_AWCACHE = edge_list_ch_46__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_46_AWID = edge_list_ch_46__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_46_AWLEN = edge_list_ch_46__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_46_AWLOCK = edge_list_ch_46__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_46_AWPROT = edge_list_ch_46__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_46_AWQOS = edge_list_ch_46__m_axi_m_axi_AWQOS;
  assign edge_list_ch_46__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_46_AWREADY;
  assign m_axi_edge_list_ch_46_AWSIZE = edge_list_ch_46__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_46_AWVALID = edge_list_ch_46__m_axi_m_axi_AWVALID;
  assign edge_list_ch_46__m_axi_m_axi_BID = m_axi_edge_list_ch_46_BID;
  assign m_axi_edge_list_ch_46_BREADY = edge_list_ch_46__m_axi_m_axi_BREADY;
  assign edge_list_ch_46__m_axi_m_axi_BRESP = m_axi_edge_list_ch_46_BRESP;
  assign edge_list_ch_46__m_axi_m_axi_BVALID = m_axi_edge_list_ch_46_BVALID;
  assign edge_list_ch_46__m_axi_m_axi_RDATA = m_axi_edge_list_ch_46_RDATA;
  assign edge_list_ch_46__m_axi_m_axi_RID = m_axi_edge_list_ch_46_RID;
  assign edge_list_ch_46__m_axi_m_axi_RLAST = m_axi_edge_list_ch_46_RLAST;
  assign m_axi_edge_list_ch_46_RREADY = edge_list_ch_46__m_axi_m_axi_RREADY;
  assign edge_list_ch_46__m_axi_m_axi_RRESP = m_axi_edge_list_ch_46_RRESP;
  assign edge_list_ch_46__m_axi_m_axi_RVALID = m_axi_edge_list_ch_46_RVALID;
  assign m_axi_edge_list_ch_46_WDATA = edge_list_ch_46__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_46_WLAST = edge_list_ch_46__m_axi_m_axi_WLAST;
  assign edge_list_ch_46__m_axi_m_axi_WREADY = m_axi_edge_list_ch_46_WREADY;
  assign m_axi_edge_list_ch_46_WSTRB = edge_list_ch_46__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_46_WVALID = edge_list_ch_46__m_axi_m_axi_WVALID;
  assign edge_list_ch_46__m_axi_read_addr_din = edge_list_ch_46_read_addr__din;
  assign edge_list_ch_46_read_addr__full_n = edge_list_ch_46__m_axi_read_addr_full_n;
  assign edge_list_ch_46__m_axi_read_addr_write = edge_list_ch_46_read_addr__write;
  assign edge_list_ch_46_read_data__dout = edge_list_ch_46__m_axi_read_data_dout;
  assign edge_list_ch_46_read_data__empty_n = edge_list_ch_46__m_axi_read_data_empty_n;
  assign edge_list_ch_46__m_axi_read_data_read = edge_list_ch_46_read_data__read;
  assign edge_list_ch_46__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_46__m_axi_write_addr_din = edge_list_ch_46_write_addr__din;
  assign edge_list_ch_46_write_addr__full_n = edge_list_ch_46__m_axi_write_addr_full_n;
  assign edge_list_ch_46__m_axi_write_addr_write = edge_list_ch_46_write_addr__write;
  assign edge_list_ch_46__m_axi_write_data_din = edge_list_ch_46_write_data__din;
  assign edge_list_ch_46_write_data__full_n = edge_list_ch_46__m_axi_write_data_full_n;
  assign edge_list_ch_46__m_axi_write_data_write = edge_list_ch_46_write_data__write;
  assign edge_list_ch_46_write_resp__dout = edge_list_ch_46__m_axi_write_resp_dout;
  assign edge_list_ch_46_write_resp__empty_n = edge_list_ch_46__m_axi_write_resp_empty_n;
  assign edge_list_ch_46__m_axi_write_resp_read = edge_list_ch_46_write_resp__read;
  assign edge_list_ch_47__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ch_47_ARADDR = edge_list_ch_47__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ch_47_ARBURST = edge_list_ch_47__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ch_47_ARCACHE = edge_list_ch_47__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ch_47_ARID = edge_list_ch_47__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ch_47_ARLEN = edge_list_ch_47__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ch_47_ARLOCK = edge_list_ch_47__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ch_47_ARPROT = edge_list_ch_47__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ch_47_ARQOS = edge_list_ch_47__m_axi_m_axi_ARQOS;
  assign edge_list_ch_47__m_axi_m_axi_ARREADY = m_axi_edge_list_ch_47_ARREADY;
  assign m_axi_edge_list_ch_47_ARSIZE = edge_list_ch_47__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ch_47_ARVALID = edge_list_ch_47__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ch_47_AWADDR = edge_list_ch_47__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ch_47_AWBURST = edge_list_ch_47__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ch_47_AWCACHE = edge_list_ch_47__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ch_47_AWID = edge_list_ch_47__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ch_47_AWLEN = edge_list_ch_47__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ch_47_AWLOCK = edge_list_ch_47__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ch_47_AWPROT = edge_list_ch_47__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ch_47_AWQOS = edge_list_ch_47__m_axi_m_axi_AWQOS;
  assign edge_list_ch_47__m_axi_m_axi_AWREADY = m_axi_edge_list_ch_47_AWREADY;
  assign m_axi_edge_list_ch_47_AWSIZE = edge_list_ch_47__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ch_47_AWVALID = edge_list_ch_47__m_axi_m_axi_AWVALID;
  assign edge_list_ch_47__m_axi_m_axi_BID = m_axi_edge_list_ch_47_BID;
  assign m_axi_edge_list_ch_47_BREADY = edge_list_ch_47__m_axi_m_axi_BREADY;
  assign edge_list_ch_47__m_axi_m_axi_BRESP = m_axi_edge_list_ch_47_BRESP;
  assign edge_list_ch_47__m_axi_m_axi_BVALID = m_axi_edge_list_ch_47_BVALID;
  assign edge_list_ch_47__m_axi_m_axi_RDATA = m_axi_edge_list_ch_47_RDATA;
  assign edge_list_ch_47__m_axi_m_axi_RID = m_axi_edge_list_ch_47_RID;
  assign edge_list_ch_47__m_axi_m_axi_RLAST = m_axi_edge_list_ch_47_RLAST;
  assign m_axi_edge_list_ch_47_RREADY = edge_list_ch_47__m_axi_m_axi_RREADY;
  assign edge_list_ch_47__m_axi_m_axi_RRESP = m_axi_edge_list_ch_47_RRESP;
  assign edge_list_ch_47__m_axi_m_axi_RVALID = m_axi_edge_list_ch_47_RVALID;
  assign m_axi_edge_list_ch_47_WDATA = edge_list_ch_47__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ch_47_WLAST = edge_list_ch_47__m_axi_m_axi_WLAST;
  assign edge_list_ch_47__m_axi_m_axi_WREADY = m_axi_edge_list_ch_47_WREADY;
  assign m_axi_edge_list_ch_47_WSTRB = edge_list_ch_47__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ch_47_WVALID = edge_list_ch_47__m_axi_m_axi_WVALID;
  assign edge_list_ch_47__m_axi_read_addr_din = edge_list_ch_47_read_addr__din;
  assign edge_list_ch_47_read_addr__full_n = edge_list_ch_47__m_axi_read_addr_full_n;
  assign edge_list_ch_47__m_axi_read_addr_write = edge_list_ch_47_read_addr__write;
  assign edge_list_ch_47_read_data__dout = edge_list_ch_47__m_axi_read_data_dout;
  assign edge_list_ch_47_read_data__empty_n = edge_list_ch_47__m_axi_read_data_empty_n;
  assign edge_list_ch_47__m_axi_read_data_read = edge_list_ch_47_read_data__read;
  assign edge_list_ch_47__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ch_47__m_axi_write_addr_din = edge_list_ch_47_write_addr__din;
  assign edge_list_ch_47_write_addr__full_n = edge_list_ch_47__m_axi_write_addr_full_n;
  assign edge_list_ch_47__m_axi_write_addr_write = edge_list_ch_47_write_addr__write;
  assign edge_list_ch_47__m_axi_write_data_din = edge_list_ch_47_write_data__din;
  assign edge_list_ch_47_write_data__full_n = edge_list_ch_47__m_axi_write_data_full_n;
  assign edge_list_ch_47__m_axi_write_data_write = edge_list_ch_47_write_data__write;
  assign edge_list_ch_47_write_resp__dout = edge_list_ch_47__m_axi_write_resp_dout;
  assign edge_list_ch_47_write_resp__empty_n = edge_list_ch_47__m_axi_write_resp_empty_n;
  assign edge_list_ch_47__m_axi_write_resp_read = edge_list_ch_47_write_resp__read;
  assign vec_X__m_axi_clk = ap_clk;
  assign m_axi_vec_X_ARADDR = vec_X__m_axi_m_axi_ARADDR;
  assign m_axi_vec_X_ARBURST = vec_X__m_axi_m_axi_ARBURST;
  assign m_axi_vec_X_ARCACHE = vec_X__m_axi_m_axi_ARCACHE;
  assign m_axi_vec_X_ARID = vec_X__m_axi_m_axi_ARID;
  assign m_axi_vec_X_ARLEN = vec_X__m_axi_m_axi_ARLEN;
  assign m_axi_vec_X_ARLOCK = vec_X__m_axi_m_axi_ARLOCK;
  assign m_axi_vec_X_ARPROT = vec_X__m_axi_m_axi_ARPROT;
  assign m_axi_vec_X_ARQOS = vec_X__m_axi_m_axi_ARQOS;
  assign vec_X__m_axi_m_axi_ARREADY = m_axi_vec_X_ARREADY;
  assign m_axi_vec_X_ARSIZE = vec_X__m_axi_m_axi_ARSIZE;
  assign m_axi_vec_X_ARVALID = vec_X__m_axi_m_axi_ARVALID;
  assign m_axi_vec_X_AWADDR = vec_X__m_axi_m_axi_AWADDR;
  assign m_axi_vec_X_AWBURST = vec_X__m_axi_m_axi_AWBURST;
  assign m_axi_vec_X_AWCACHE = vec_X__m_axi_m_axi_AWCACHE;
  assign m_axi_vec_X_AWID = vec_X__m_axi_m_axi_AWID;
  assign m_axi_vec_X_AWLEN = vec_X__m_axi_m_axi_AWLEN;
  assign m_axi_vec_X_AWLOCK = vec_X__m_axi_m_axi_AWLOCK;
  assign m_axi_vec_X_AWPROT = vec_X__m_axi_m_axi_AWPROT;
  assign m_axi_vec_X_AWQOS = vec_X__m_axi_m_axi_AWQOS;
  assign vec_X__m_axi_m_axi_AWREADY = m_axi_vec_X_AWREADY;
  assign m_axi_vec_X_AWSIZE = vec_X__m_axi_m_axi_AWSIZE;
  assign m_axi_vec_X_AWVALID = vec_X__m_axi_m_axi_AWVALID;
  assign vec_X__m_axi_m_axi_BID = m_axi_vec_X_BID;
  assign m_axi_vec_X_BREADY = vec_X__m_axi_m_axi_BREADY;
  assign vec_X__m_axi_m_axi_BRESP = m_axi_vec_X_BRESP;
  assign vec_X__m_axi_m_axi_BVALID = m_axi_vec_X_BVALID;
  assign vec_X__m_axi_m_axi_RDATA = m_axi_vec_X_RDATA;
  assign vec_X__m_axi_m_axi_RID = m_axi_vec_X_RID;
  assign vec_X__m_axi_m_axi_RLAST = m_axi_vec_X_RLAST;
  assign m_axi_vec_X_RREADY = vec_X__m_axi_m_axi_RREADY;
  assign vec_X__m_axi_m_axi_RRESP = m_axi_vec_X_RRESP;
  assign vec_X__m_axi_m_axi_RVALID = m_axi_vec_X_RVALID;
  assign m_axi_vec_X_WDATA = vec_X__m_axi_m_axi_WDATA;
  assign m_axi_vec_X_WLAST = vec_X__m_axi_m_axi_WLAST;
  assign vec_X__m_axi_m_axi_WREADY = m_axi_vec_X_WREADY;
  assign m_axi_vec_X_WSTRB = vec_X__m_axi_m_axi_WSTRB;
  assign m_axi_vec_X_WVALID = vec_X__m_axi_m_axi_WVALID;
  assign vec_X__m_axi_read_addr_din = vec_X_read_addr__din;
  assign vec_X_read_addr__full_n = vec_X__m_axi_read_addr_full_n;
  assign vec_X__m_axi_read_addr_write = vec_X_read_addr__write;
  assign vec_X_read_data__dout = vec_X__m_axi_read_data_dout;
  assign vec_X_read_data__empty_n = vec_X__m_axi_read_data_empty_n;
  assign vec_X__m_axi_read_data_read = vec_X_read_data__read;
  assign vec_X__m_axi_rst = ~ ap_rst_n;
  assign vec_X__m_axi_write_addr_din = vec_X_write_addr__din;
  assign vec_X_write_addr__full_n = vec_X__m_axi_write_addr_full_n;
  assign vec_X__m_axi_write_addr_write = vec_X_write_addr__write;
  assign vec_X__m_axi_write_data_din = vec_X_write_data__din;
  assign vec_X_write_data__full_n = vec_X__m_axi_write_data_full_n;
  assign vec_X__m_axi_write_data_write = vec_X_write_data__write;
  assign vec_X_write_resp__dout = vec_X__m_axi_write_resp_dout;
  assign vec_X_write_resp__empty_n = vec_X__m_axi_write_resp_empty_n;
  assign vec_X__m_axi_write_resp_read = vec_X_write_resp__read;
  assign vec_Y__m_axi_clk = ap_clk;
  assign m_axi_vec_Y_ARADDR = vec_Y__m_axi_m_axi_ARADDR;
  assign m_axi_vec_Y_ARBURST = vec_Y__m_axi_m_axi_ARBURST;
  assign m_axi_vec_Y_ARCACHE = vec_Y__m_axi_m_axi_ARCACHE;
  assign m_axi_vec_Y_ARID = vec_Y__m_axi_m_axi_ARID;
  assign m_axi_vec_Y_ARLEN = vec_Y__m_axi_m_axi_ARLEN;
  assign m_axi_vec_Y_ARLOCK = vec_Y__m_axi_m_axi_ARLOCK;
  assign m_axi_vec_Y_ARPROT = vec_Y__m_axi_m_axi_ARPROT;
  assign m_axi_vec_Y_ARQOS = vec_Y__m_axi_m_axi_ARQOS;
  assign vec_Y__m_axi_m_axi_ARREADY = m_axi_vec_Y_ARREADY;
  assign m_axi_vec_Y_ARSIZE = vec_Y__m_axi_m_axi_ARSIZE;
  assign m_axi_vec_Y_ARVALID = vec_Y__m_axi_m_axi_ARVALID;
  assign m_axi_vec_Y_AWADDR = vec_Y__m_axi_m_axi_AWADDR;
  assign m_axi_vec_Y_AWBURST = vec_Y__m_axi_m_axi_AWBURST;
  assign m_axi_vec_Y_AWCACHE = vec_Y__m_axi_m_axi_AWCACHE;
  assign m_axi_vec_Y_AWID = vec_Y__m_axi_m_axi_AWID;
  assign m_axi_vec_Y_AWLEN = vec_Y__m_axi_m_axi_AWLEN;
  assign m_axi_vec_Y_AWLOCK = vec_Y__m_axi_m_axi_AWLOCK;
  assign m_axi_vec_Y_AWPROT = vec_Y__m_axi_m_axi_AWPROT;
  assign m_axi_vec_Y_AWQOS = vec_Y__m_axi_m_axi_AWQOS;
  assign vec_Y__m_axi_m_axi_AWREADY = m_axi_vec_Y_AWREADY;
  assign m_axi_vec_Y_AWSIZE = vec_Y__m_axi_m_axi_AWSIZE;
  assign m_axi_vec_Y_AWVALID = vec_Y__m_axi_m_axi_AWVALID;
  assign vec_Y__m_axi_m_axi_BID = m_axi_vec_Y_BID;
  assign m_axi_vec_Y_BREADY = vec_Y__m_axi_m_axi_BREADY;
  assign vec_Y__m_axi_m_axi_BRESP = m_axi_vec_Y_BRESP;
  assign vec_Y__m_axi_m_axi_BVALID = m_axi_vec_Y_BVALID;
  assign vec_Y__m_axi_m_axi_RDATA = m_axi_vec_Y_RDATA;
  assign vec_Y__m_axi_m_axi_RID = m_axi_vec_Y_RID;
  assign vec_Y__m_axi_m_axi_RLAST = m_axi_vec_Y_RLAST;
  assign m_axi_vec_Y_RREADY = vec_Y__m_axi_m_axi_RREADY;
  assign vec_Y__m_axi_m_axi_RRESP = m_axi_vec_Y_RRESP;
  assign vec_Y__m_axi_m_axi_RVALID = m_axi_vec_Y_RVALID;
  assign m_axi_vec_Y_WDATA = vec_Y__m_axi_m_axi_WDATA;
  assign m_axi_vec_Y_WLAST = vec_Y__m_axi_m_axi_WLAST;
  assign vec_Y__m_axi_m_axi_WREADY = m_axi_vec_Y_WREADY;
  assign m_axi_vec_Y_WSTRB = vec_Y__m_axi_m_axi_WSTRB;
  assign m_axi_vec_Y_WVALID = vec_Y__m_axi_m_axi_WVALID;
  assign vec_Y__m_axi_read_addr_din = vec_Y_read_addr__din;
  assign vec_Y_read_addr__full_n = vec_Y__m_axi_read_addr_full_n;
  assign vec_Y__m_axi_read_addr_write = vec_Y_read_addr__write;
  assign vec_Y_read_data__dout = vec_Y__m_axi_read_data_dout;
  assign vec_Y_read_data__empty_n = vec_Y__m_axi_read_data_empty_n;
  assign vec_Y__m_axi_read_data_read = vec_Y_read_data__read;
  assign vec_Y__m_axi_rst = ~ ap_rst_n;
  assign vec_Y__m_axi_write_addr_din = vec_Y_write_addr__din;
  assign vec_Y_write_addr__full_n = vec_Y__m_axi_write_addr_full_n;
  assign vec_Y__m_axi_write_addr_write = vec_Y_write_addr__write;
  assign vec_Y__m_axi_write_data_din = vec_Y_write_data__din;
  assign vec_Y_write_data__full_n = vec_Y__m_axi_write_data_full_n;
  assign vec_Y__m_axi_write_data_write = vec_Y_write_data__write;
  assign vec_Y_write_resp__dout = vec_Y__m_axi_write_resp_dout;
  assign vec_Y_write_resp__empty_n = vec_Y__m_axi_write_resp_empty_n;
  assign vec_Y__m_axi_write_resp_read = vec_Y_write_resp__read;
  assign edge_list_ptr__m_axi_clk = ap_clk;
  assign m_axi_edge_list_ptr_ARADDR = edge_list_ptr__m_axi_m_axi_ARADDR;
  assign m_axi_edge_list_ptr_ARBURST = edge_list_ptr__m_axi_m_axi_ARBURST;
  assign m_axi_edge_list_ptr_ARCACHE = edge_list_ptr__m_axi_m_axi_ARCACHE;
  assign m_axi_edge_list_ptr_ARID = edge_list_ptr__m_axi_m_axi_ARID;
  assign m_axi_edge_list_ptr_ARLEN = edge_list_ptr__m_axi_m_axi_ARLEN;
  assign m_axi_edge_list_ptr_ARLOCK = edge_list_ptr__m_axi_m_axi_ARLOCK;
  assign m_axi_edge_list_ptr_ARPROT = edge_list_ptr__m_axi_m_axi_ARPROT;
  assign m_axi_edge_list_ptr_ARQOS = edge_list_ptr__m_axi_m_axi_ARQOS;
  assign edge_list_ptr__m_axi_m_axi_ARREADY = m_axi_edge_list_ptr_ARREADY;
  assign m_axi_edge_list_ptr_ARSIZE = edge_list_ptr__m_axi_m_axi_ARSIZE;
  assign m_axi_edge_list_ptr_ARVALID = edge_list_ptr__m_axi_m_axi_ARVALID;
  assign m_axi_edge_list_ptr_AWADDR = edge_list_ptr__m_axi_m_axi_AWADDR;
  assign m_axi_edge_list_ptr_AWBURST = edge_list_ptr__m_axi_m_axi_AWBURST;
  assign m_axi_edge_list_ptr_AWCACHE = edge_list_ptr__m_axi_m_axi_AWCACHE;
  assign m_axi_edge_list_ptr_AWID = edge_list_ptr__m_axi_m_axi_AWID;
  assign m_axi_edge_list_ptr_AWLEN = edge_list_ptr__m_axi_m_axi_AWLEN;
  assign m_axi_edge_list_ptr_AWLOCK = edge_list_ptr__m_axi_m_axi_AWLOCK;
  assign m_axi_edge_list_ptr_AWPROT = edge_list_ptr__m_axi_m_axi_AWPROT;
  assign m_axi_edge_list_ptr_AWQOS = edge_list_ptr__m_axi_m_axi_AWQOS;
  assign edge_list_ptr__m_axi_m_axi_AWREADY = m_axi_edge_list_ptr_AWREADY;
  assign m_axi_edge_list_ptr_AWSIZE = edge_list_ptr__m_axi_m_axi_AWSIZE;
  assign m_axi_edge_list_ptr_AWVALID = edge_list_ptr__m_axi_m_axi_AWVALID;
  assign edge_list_ptr__m_axi_m_axi_BID = m_axi_edge_list_ptr_BID;
  assign m_axi_edge_list_ptr_BREADY = edge_list_ptr__m_axi_m_axi_BREADY;
  assign edge_list_ptr__m_axi_m_axi_BRESP = m_axi_edge_list_ptr_BRESP;
  assign edge_list_ptr__m_axi_m_axi_BVALID = m_axi_edge_list_ptr_BVALID;
  assign edge_list_ptr__m_axi_m_axi_RDATA = m_axi_edge_list_ptr_RDATA;
  assign edge_list_ptr__m_axi_m_axi_RID = m_axi_edge_list_ptr_RID;
  assign edge_list_ptr__m_axi_m_axi_RLAST = m_axi_edge_list_ptr_RLAST;
  assign m_axi_edge_list_ptr_RREADY = edge_list_ptr__m_axi_m_axi_RREADY;
  assign edge_list_ptr__m_axi_m_axi_RRESP = m_axi_edge_list_ptr_RRESP;
  assign edge_list_ptr__m_axi_m_axi_RVALID = m_axi_edge_list_ptr_RVALID;
  assign m_axi_edge_list_ptr_WDATA = edge_list_ptr__m_axi_m_axi_WDATA;
  assign m_axi_edge_list_ptr_WLAST = edge_list_ptr__m_axi_m_axi_WLAST;
  assign edge_list_ptr__m_axi_m_axi_WREADY = m_axi_edge_list_ptr_WREADY;
  assign m_axi_edge_list_ptr_WSTRB = edge_list_ptr__m_axi_m_axi_WSTRB;
  assign m_axi_edge_list_ptr_WVALID = edge_list_ptr__m_axi_m_axi_WVALID;
  assign edge_list_ptr__m_axi_read_addr_din = edge_list_ptr_read_addr__din;
  assign edge_list_ptr_read_addr__full_n = edge_list_ptr__m_axi_read_addr_full_n;
  assign edge_list_ptr__m_axi_read_addr_write = edge_list_ptr_read_addr__write;
  assign edge_list_ptr_read_data__dout = edge_list_ptr__m_axi_read_data_dout;
  assign edge_list_ptr_read_data__empty_n = edge_list_ptr__m_axi_read_data_empty_n;
  assign edge_list_ptr__m_axi_read_data_read = edge_list_ptr_read_data__read;
  assign edge_list_ptr__m_axi_rst = ~ ap_rst_n;
  assign edge_list_ptr__m_axi_write_addr_din = edge_list_ptr_write_addr__din;
  assign edge_list_ptr_write_addr__full_n = edge_list_ptr__m_axi_write_addr_full_n;
  assign edge_list_ptr__m_axi_write_addr_write = edge_list_ptr_write_addr__write;
  assign edge_list_ptr__m_axi_write_data_din = edge_list_ptr_write_data__din;
  assign edge_list_ptr_write_data__full_n = edge_list_ptr__m_axi_write_data_full_n;
  assign edge_list_ptr__m_axi_write_data_write = edge_list_ptr_write_data__write;
  assign edge_list_ptr_write_resp__dout = edge_list_ptr__m_axi_write_resp_dout;
  assign edge_list_ptr_write_resp__empty_n = edge_list_ptr__m_axi_write_resp_empty_n;
  assign edge_list_ptr__m_axi_write_resp_read = edge_list_ptr_write_resp__read;
  assign vec_Y_out__m_axi_clk = ap_clk;
  assign m_axi_vec_Y_out_ARADDR = vec_Y_out__m_axi_m_axi_ARADDR;
  assign m_axi_vec_Y_out_ARBURST = vec_Y_out__m_axi_m_axi_ARBURST;
  assign m_axi_vec_Y_out_ARCACHE = vec_Y_out__m_axi_m_axi_ARCACHE;
  assign m_axi_vec_Y_out_ARID = vec_Y_out__m_axi_m_axi_ARID;
  assign m_axi_vec_Y_out_ARLEN = vec_Y_out__m_axi_m_axi_ARLEN;
  assign m_axi_vec_Y_out_ARLOCK = vec_Y_out__m_axi_m_axi_ARLOCK;
  assign m_axi_vec_Y_out_ARPROT = vec_Y_out__m_axi_m_axi_ARPROT;
  assign m_axi_vec_Y_out_ARQOS = vec_Y_out__m_axi_m_axi_ARQOS;
  assign vec_Y_out__m_axi_m_axi_ARREADY = m_axi_vec_Y_out_ARREADY;
  assign m_axi_vec_Y_out_ARSIZE = vec_Y_out__m_axi_m_axi_ARSIZE;
  assign m_axi_vec_Y_out_ARVALID = vec_Y_out__m_axi_m_axi_ARVALID;
  assign m_axi_vec_Y_out_AWADDR = vec_Y_out__m_axi_m_axi_AWADDR;
  assign m_axi_vec_Y_out_AWBURST = vec_Y_out__m_axi_m_axi_AWBURST;
  assign m_axi_vec_Y_out_AWCACHE = vec_Y_out__m_axi_m_axi_AWCACHE;
  assign m_axi_vec_Y_out_AWID = vec_Y_out__m_axi_m_axi_AWID;
  assign m_axi_vec_Y_out_AWLEN = vec_Y_out__m_axi_m_axi_AWLEN;
  assign m_axi_vec_Y_out_AWLOCK = vec_Y_out__m_axi_m_axi_AWLOCK;
  assign m_axi_vec_Y_out_AWPROT = vec_Y_out__m_axi_m_axi_AWPROT;
  assign m_axi_vec_Y_out_AWQOS = vec_Y_out__m_axi_m_axi_AWQOS;
  assign vec_Y_out__m_axi_m_axi_AWREADY = m_axi_vec_Y_out_AWREADY;
  assign m_axi_vec_Y_out_AWSIZE = vec_Y_out__m_axi_m_axi_AWSIZE;
  assign m_axi_vec_Y_out_AWVALID = vec_Y_out__m_axi_m_axi_AWVALID;
  assign vec_Y_out__m_axi_m_axi_BID = m_axi_vec_Y_out_BID;
  assign m_axi_vec_Y_out_BREADY = vec_Y_out__m_axi_m_axi_BREADY;
  assign vec_Y_out__m_axi_m_axi_BRESP = m_axi_vec_Y_out_BRESP;
  assign vec_Y_out__m_axi_m_axi_BVALID = m_axi_vec_Y_out_BVALID;
  assign vec_Y_out__m_axi_m_axi_RDATA = m_axi_vec_Y_out_RDATA;
  assign vec_Y_out__m_axi_m_axi_RID = m_axi_vec_Y_out_RID;
  assign vec_Y_out__m_axi_m_axi_RLAST = m_axi_vec_Y_out_RLAST;
  assign m_axi_vec_Y_out_RREADY = vec_Y_out__m_axi_m_axi_RREADY;
  assign vec_Y_out__m_axi_m_axi_RRESP = m_axi_vec_Y_out_RRESP;
  assign vec_Y_out__m_axi_m_axi_RVALID = m_axi_vec_Y_out_RVALID;
  assign m_axi_vec_Y_out_WDATA = vec_Y_out__m_axi_m_axi_WDATA;
  assign m_axi_vec_Y_out_WLAST = vec_Y_out__m_axi_m_axi_WLAST;
  assign vec_Y_out__m_axi_m_axi_WREADY = m_axi_vec_Y_out_WREADY;
  assign m_axi_vec_Y_out_WSTRB = vec_Y_out__m_axi_m_axi_WSTRB;
  assign m_axi_vec_Y_out_WVALID = vec_Y_out__m_axi_m_axi_WVALID;
  assign vec_Y_out__m_axi_read_addr_din = vec_Y_out_read_addr__din;
  assign vec_Y_out_read_addr__full_n = vec_Y_out__m_axi_read_addr_full_n;
  assign vec_Y_out__m_axi_read_addr_write = vec_Y_out_read_addr__write;
  assign vec_Y_out_read_data__dout = vec_Y_out__m_axi_read_data_dout;
  assign vec_Y_out_read_data__empty_n = vec_Y_out__m_axi_read_data_empty_n;
  assign vec_Y_out__m_axi_read_data_read = vec_Y_out_read_data__read;
  assign vec_Y_out__m_axi_rst = ~ ap_rst_n;
  assign vec_Y_out__m_axi_write_addr_din = vec_Y_out_write_addr__din;
  assign vec_Y_out_write_addr__full_n = vec_Y_out__m_axi_write_addr_full_n;
  assign vec_Y_out__m_axi_write_addr_write = vec_Y_out_write_addr__write;
  assign vec_Y_out__m_axi_write_data_din = vec_Y_out_write_data__din;
  assign vec_Y_out_write_data__full_n = vec_Y_out__m_axi_write_data_full_n;
  assign vec_Y_out__m_axi_write_data_write = vec_Y_out_write_data__write;
  assign vec_Y_out_write_resp__dout = vec_Y_out__m_axi_write_resp_dout;
  assign vec_Y_out_write_resp__empty_n = vec_Y_out__m_axi_write_resp_empty_n;
  assign vec_Y_out__m_axi_write_resp_read = vec_Y_out_write_resp__read;
  assign Arbiter_Y_0___M__q0 = __tapa_fsm_unit_Arbiter_Y_0___M__q0;
  assign Arbiter_Y_0___P_N__q0 = __tapa_fsm_unit_Arbiter_Y_0___P_N__q0;
  assign __tapa_fsm_unit_Arbiter_Y_0__ap_done = Arbiter_Y_0__ap_done;
  assign __tapa_fsm_unit_Arbiter_Y_0__ap_idle = Arbiter_Y_0__ap_idle;
  assign __tapa_fsm_unit_Arbiter_Y_0__ap_ready = Arbiter_Y_0__ap_ready;
  assign Arbiter_Y_0__ap_start = __tapa_fsm_unit_Arbiter_Y_0__ap_start;
  assign Arbiter_Y_1___M__q0 = __tapa_fsm_unit_Arbiter_Y_1___M__q0;
  assign Arbiter_Y_1___P_N__q0 = __tapa_fsm_unit_Arbiter_Y_1___P_N__q0;
  assign __tapa_fsm_unit_Arbiter_Y_1__ap_done = Arbiter_Y_1__ap_done;
  assign __tapa_fsm_unit_Arbiter_Y_1__ap_idle = Arbiter_Y_1__ap_idle;
  assign __tapa_fsm_unit_Arbiter_Y_1__ap_ready = Arbiter_Y_1__ap_ready;
  assign Arbiter_Y_1__ap_start = __tapa_fsm_unit_Arbiter_Y_1__ap_start;
  assign Arbiter_Y_2___M__q0 = __tapa_fsm_unit_Arbiter_Y_2___M__q0;
  assign Arbiter_Y_2___P_N__q0 = __tapa_fsm_unit_Arbiter_Y_2___P_N__q0;
  assign __tapa_fsm_unit_Arbiter_Y_2__ap_done = Arbiter_Y_2__ap_done;
  assign __tapa_fsm_unit_Arbiter_Y_2__ap_idle = Arbiter_Y_2__ap_idle;
  assign __tapa_fsm_unit_Arbiter_Y_2__ap_ready = Arbiter_Y_2__ap_ready;
  assign Arbiter_Y_2__ap_start = __tapa_fsm_unit_Arbiter_Y_2__ap_start;
  assign Arbiter_Y_3___M__q0 = __tapa_fsm_unit_Arbiter_Y_3___M__q0;
  assign Arbiter_Y_3___P_N__q0 = __tapa_fsm_unit_Arbiter_Y_3___P_N__q0;
  assign __tapa_fsm_unit_Arbiter_Y_3__ap_done = Arbiter_Y_3__ap_done;
  assign __tapa_fsm_unit_Arbiter_Y_3__ap_idle = Arbiter_Y_3__ap_idle;
  assign __tapa_fsm_unit_Arbiter_Y_3__ap_ready = Arbiter_Y_3__ap_ready;
  assign Arbiter_Y_3__ap_start = __tapa_fsm_unit_Arbiter_Y_3__ap_start;
  assign Arbiter_Y_4___M__q0 = __tapa_fsm_unit_Arbiter_Y_4___M__q0;
  assign Arbiter_Y_4___P_N__q0 = __tapa_fsm_unit_Arbiter_Y_4___P_N__q0;
  assign __tapa_fsm_unit_Arbiter_Y_4__ap_done = Arbiter_Y_4__ap_done;
  assign __tapa_fsm_unit_Arbiter_Y_4__ap_idle = Arbiter_Y_4__ap_idle;
  assign __tapa_fsm_unit_Arbiter_Y_4__ap_ready = Arbiter_Y_4__ap_ready;
  assign Arbiter_Y_4__ap_start = __tapa_fsm_unit_Arbiter_Y_4__ap_start;
  assign Arbiter_Y_5___M__q0 = __tapa_fsm_unit_Arbiter_Y_5___M__q0;
  assign Arbiter_Y_5___P_N__q0 = __tapa_fsm_unit_Arbiter_Y_5___P_N__q0;
  assign __tapa_fsm_unit_Arbiter_Y_5__ap_done = Arbiter_Y_5__ap_done;
  assign __tapa_fsm_unit_Arbiter_Y_5__ap_idle = Arbiter_Y_5__ap_idle;
  assign __tapa_fsm_unit_Arbiter_Y_5__ap_ready = Arbiter_Y_5__ap_ready;
  assign Arbiter_Y_5__ap_start = __tapa_fsm_unit_Arbiter_Y_5__ap_start;
  assign Arbiter_Y_6___M__q0 = __tapa_fsm_unit_Arbiter_Y_6___M__q0;
  assign Arbiter_Y_6___P_N__q0 = __tapa_fsm_unit_Arbiter_Y_6___P_N__q0;
  assign __tapa_fsm_unit_Arbiter_Y_6__ap_done = Arbiter_Y_6__ap_done;
  assign __tapa_fsm_unit_Arbiter_Y_6__ap_idle = Arbiter_Y_6__ap_idle;
  assign __tapa_fsm_unit_Arbiter_Y_6__ap_ready = Arbiter_Y_6__ap_ready;
  assign Arbiter_Y_6__ap_start = __tapa_fsm_unit_Arbiter_Y_6__ap_start;
  assign Arbiter_Y_7___M__q0 = __tapa_fsm_unit_Arbiter_Y_7___M__q0;
  assign Arbiter_Y_7___P_N__q0 = __tapa_fsm_unit_Arbiter_Y_7___P_N__q0;
  assign __tapa_fsm_unit_Arbiter_Y_7__ap_done = Arbiter_Y_7__ap_done;
  assign __tapa_fsm_unit_Arbiter_Y_7__ap_idle = Arbiter_Y_7__ap_idle;
  assign __tapa_fsm_unit_Arbiter_Y_7__ap_ready = Arbiter_Y_7__ap_ready;
  assign Arbiter_Y_7__ap_start = __tapa_fsm_unit_Arbiter_Y_7__ap_start;
  assign FloatvAddFloatv_0__ap_start = __tapa_fsm_unit_FloatvAddFloatv_0__ap_start;
  assign FloatvMultConst_0___M__q0 = __tapa_fsm_unit_FloatvMultConst_0___M__q0;
  assign FloatvMultConst_0___P_N__q0 = __tapa_fsm_unit_FloatvMultConst_0___P_N__q0;
  assign FloatvMultConst_0___alpha_u__q0 = __tapa_fsm_unit_FloatvMultConst_0___alpha_u__q0;
  assign __tapa_fsm_unit_FloatvMultConst_0__ap_done = FloatvMultConst_0__ap_done;
  assign __tapa_fsm_unit_FloatvMultConst_0__ap_idle = FloatvMultConst_0__ap_idle;
  assign __tapa_fsm_unit_FloatvMultConst_0__ap_ready = FloatvMultConst_0__ap_ready;
  assign FloatvMultConst_0__ap_start = __tapa_fsm_unit_FloatvMultConst_0__ap_start;
  assign FloatvMultConst_1___M__q0 = __tapa_fsm_unit_FloatvMultConst_1___M__q0;
  assign FloatvMultConst_1___P_N__q0 = __tapa_fsm_unit_FloatvMultConst_1___P_N__q0;
  assign FloatvMultConst_1___beta_u__q0 = __tapa_fsm_unit_FloatvMultConst_1___beta_u__q0;
  assign __tapa_fsm_unit_FloatvMultConst_1__ap_done = FloatvMultConst_1__ap_done;
  assign __tapa_fsm_unit_FloatvMultConst_1__ap_idle = FloatvMultConst_1__ap_idle;
  assign __tapa_fsm_unit_FloatvMultConst_1__ap_ready = FloatvMultConst_1__ap_ready;
  assign FloatvMultConst_1__ap_start = __tapa_fsm_unit_FloatvMultConst_1__ap_start;
  assign __tapa_fsm_unit_K = K;
  assign __tapa_fsm_unit_M = M;
  assign Merger_Y_0__ap_start = __tapa_fsm_unit_Merger_Y_0__ap_start;
  assign __tapa_fsm_unit_NUM_A_LEN = NUM_A_LEN;
  assign __tapa_fsm_unit_NUM_ITE = NUM_ITE;
  assign __tapa_fsm_unit_PEG_Xvec_0__ap_done = PEG_Xvec_0__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_0__ap_idle = PEG_Xvec_0__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_0__ap_ready = PEG_Xvec_0__ap_ready;
  assign PEG_Xvec_0__ap_start = __tapa_fsm_unit_PEG_Xvec_0__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_10__ap_done = PEG_Xvec_10__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_10__ap_idle = PEG_Xvec_10__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_10__ap_ready = PEG_Xvec_10__ap_ready;
  assign PEG_Xvec_10__ap_start = __tapa_fsm_unit_PEG_Xvec_10__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_11__ap_done = PEG_Xvec_11__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_11__ap_idle = PEG_Xvec_11__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_11__ap_ready = PEG_Xvec_11__ap_ready;
  assign PEG_Xvec_11__ap_start = __tapa_fsm_unit_PEG_Xvec_11__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_12__ap_done = PEG_Xvec_12__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_12__ap_idle = PEG_Xvec_12__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_12__ap_ready = PEG_Xvec_12__ap_ready;
  assign PEG_Xvec_12__ap_start = __tapa_fsm_unit_PEG_Xvec_12__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_13__ap_done = PEG_Xvec_13__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_13__ap_idle = PEG_Xvec_13__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_13__ap_ready = PEG_Xvec_13__ap_ready;
  assign PEG_Xvec_13__ap_start = __tapa_fsm_unit_PEG_Xvec_13__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_14__ap_done = PEG_Xvec_14__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_14__ap_idle = PEG_Xvec_14__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_14__ap_ready = PEG_Xvec_14__ap_ready;
  assign PEG_Xvec_14__ap_start = __tapa_fsm_unit_PEG_Xvec_14__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_15__ap_done = PEG_Xvec_15__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_15__ap_idle = PEG_Xvec_15__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_15__ap_ready = PEG_Xvec_15__ap_ready;
  assign PEG_Xvec_15__ap_start = __tapa_fsm_unit_PEG_Xvec_15__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_16__ap_done = PEG_Xvec_16__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_16__ap_idle = PEG_Xvec_16__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_16__ap_ready = PEG_Xvec_16__ap_ready;
  assign PEG_Xvec_16__ap_start = __tapa_fsm_unit_PEG_Xvec_16__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_17__ap_done = PEG_Xvec_17__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_17__ap_idle = PEG_Xvec_17__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_17__ap_ready = PEG_Xvec_17__ap_ready;
  assign PEG_Xvec_17__ap_start = __tapa_fsm_unit_PEG_Xvec_17__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_18__ap_done = PEG_Xvec_18__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_18__ap_idle = PEG_Xvec_18__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_18__ap_ready = PEG_Xvec_18__ap_ready;
  assign PEG_Xvec_18__ap_start = __tapa_fsm_unit_PEG_Xvec_18__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_19__ap_done = PEG_Xvec_19__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_19__ap_idle = PEG_Xvec_19__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_19__ap_ready = PEG_Xvec_19__ap_ready;
  assign PEG_Xvec_19__ap_start = __tapa_fsm_unit_PEG_Xvec_19__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_1__ap_done = PEG_Xvec_1__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_1__ap_idle = PEG_Xvec_1__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_1__ap_ready = PEG_Xvec_1__ap_ready;
  assign PEG_Xvec_1__ap_start = __tapa_fsm_unit_PEG_Xvec_1__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_20__ap_done = PEG_Xvec_20__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_20__ap_idle = PEG_Xvec_20__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_20__ap_ready = PEG_Xvec_20__ap_ready;
  assign PEG_Xvec_20__ap_start = __tapa_fsm_unit_PEG_Xvec_20__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_21__ap_done = PEG_Xvec_21__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_21__ap_idle = PEG_Xvec_21__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_21__ap_ready = PEG_Xvec_21__ap_ready;
  assign PEG_Xvec_21__ap_start = __tapa_fsm_unit_PEG_Xvec_21__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_22__ap_done = PEG_Xvec_22__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_22__ap_idle = PEG_Xvec_22__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_22__ap_ready = PEG_Xvec_22__ap_ready;
  assign PEG_Xvec_22__ap_start = __tapa_fsm_unit_PEG_Xvec_22__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_23__ap_done = PEG_Xvec_23__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_23__ap_idle = PEG_Xvec_23__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_23__ap_ready = PEG_Xvec_23__ap_ready;
  assign PEG_Xvec_23__ap_start = __tapa_fsm_unit_PEG_Xvec_23__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_24__ap_done = PEG_Xvec_24__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_24__ap_idle = PEG_Xvec_24__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_24__ap_ready = PEG_Xvec_24__ap_ready;
  assign PEG_Xvec_24__ap_start = __tapa_fsm_unit_PEG_Xvec_24__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_25__ap_done = PEG_Xvec_25__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_25__ap_idle = PEG_Xvec_25__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_25__ap_ready = PEG_Xvec_25__ap_ready;
  assign PEG_Xvec_25__ap_start = __tapa_fsm_unit_PEG_Xvec_25__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_26__ap_done = PEG_Xvec_26__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_26__ap_idle = PEG_Xvec_26__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_26__ap_ready = PEG_Xvec_26__ap_ready;
  assign PEG_Xvec_26__ap_start = __tapa_fsm_unit_PEG_Xvec_26__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_27__ap_done = PEG_Xvec_27__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_27__ap_idle = PEG_Xvec_27__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_27__ap_ready = PEG_Xvec_27__ap_ready;
  assign PEG_Xvec_27__ap_start = __tapa_fsm_unit_PEG_Xvec_27__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_28__ap_done = PEG_Xvec_28__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_28__ap_idle = PEG_Xvec_28__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_28__ap_ready = PEG_Xvec_28__ap_ready;
  assign PEG_Xvec_28__ap_start = __tapa_fsm_unit_PEG_Xvec_28__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_29__ap_done = PEG_Xvec_29__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_29__ap_idle = PEG_Xvec_29__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_29__ap_ready = PEG_Xvec_29__ap_ready;
  assign PEG_Xvec_29__ap_start = __tapa_fsm_unit_PEG_Xvec_29__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_2__ap_done = PEG_Xvec_2__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_2__ap_idle = PEG_Xvec_2__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_2__ap_ready = PEG_Xvec_2__ap_ready;
  assign PEG_Xvec_2__ap_start = __tapa_fsm_unit_PEG_Xvec_2__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_30__ap_done = PEG_Xvec_30__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_30__ap_idle = PEG_Xvec_30__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_30__ap_ready = PEG_Xvec_30__ap_ready;
  assign PEG_Xvec_30__ap_start = __tapa_fsm_unit_PEG_Xvec_30__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_31__ap_done = PEG_Xvec_31__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_31__ap_idle = PEG_Xvec_31__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_31__ap_ready = PEG_Xvec_31__ap_ready;
  assign PEG_Xvec_31__ap_start = __tapa_fsm_unit_PEG_Xvec_31__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_32__ap_done = PEG_Xvec_32__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_32__ap_idle = PEG_Xvec_32__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_32__ap_ready = PEG_Xvec_32__ap_ready;
  assign PEG_Xvec_32__ap_start = __tapa_fsm_unit_PEG_Xvec_32__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_33__ap_done = PEG_Xvec_33__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_33__ap_idle = PEG_Xvec_33__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_33__ap_ready = PEG_Xvec_33__ap_ready;
  assign PEG_Xvec_33__ap_start = __tapa_fsm_unit_PEG_Xvec_33__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_34__ap_done = PEG_Xvec_34__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_34__ap_idle = PEG_Xvec_34__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_34__ap_ready = PEG_Xvec_34__ap_ready;
  assign PEG_Xvec_34__ap_start = __tapa_fsm_unit_PEG_Xvec_34__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_35__ap_done = PEG_Xvec_35__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_35__ap_idle = PEG_Xvec_35__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_35__ap_ready = PEG_Xvec_35__ap_ready;
  assign PEG_Xvec_35__ap_start = __tapa_fsm_unit_PEG_Xvec_35__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_36__ap_done = PEG_Xvec_36__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_36__ap_idle = PEG_Xvec_36__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_36__ap_ready = PEG_Xvec_36__ap_ready;
  assign PEG_Xvec_36__ap_start = __tapa_fsm_unit_PEG_Xvec_36__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_37__ap_done = PEG_Xvec_37__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_37__ap_idle = PEG_Xvec_37__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_37__ap_ready = PEG_Xvec_37__ap_ready;
  assign PEG_Xvec_37__ap_start = __tapa_fsm_unit_PEG_Xvec_37__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_38__ap_done = PEG_Xvec_38__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_38__ap_idle = PEG_Xvec_38__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_38__ap_ready = PEG_Xvec_38__ap_ready;
  assign PEG_Xvec_38__ap_start = __tapa_fsm_unit_PEG_Xvec_38__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_39__ap_done = PEG_Xvec_39__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_39__ap_idle = PEG_Xvec_39__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_39__ap_ready = PEG_Xvec_39__ap_ready;
  assign PEG_Xvec_39__ap_start = __tapa_fsm_unit_PEG_Xvec_39__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_3__ap_done = PEG_Xvec_3__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_3__ap_idle = PEG_Xvec_3__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_3__ap_ready = PEG_Xvec_3__ap_ready;
  assign PEG_Xvec_3__ap_start = __tapa_fsm_unit_PEG_Xvec_3__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_40__ap_done = PEG_Xvec_40__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_40__ap_idle = PEG_Xvec_40__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_40__ap_ready = PEG_Xvec_40__ap_ready;
  assign PEG_Xvec_40__ap_start = __tapa_fsm_unit_PEG_Xvec_40__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_41__ap_done = PEG_Xvec_41__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_41__ap_idle = PEG_Xvec_41__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_41__ap_ready = PEG_Xvec_41__ap_ready;
  assign PEG_Xvec_41__ap_start = __tapa_fsm_unit_PEG_Xvec_41__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_42__ap_done = PEG_Xvec_42__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_42__ap_idle = PEG_Xvec_42__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_42__ap_ready = PEG_Xvec_42__ap_ready;
  assign PEG_Xvec_42__ap_start = __tapa_fsm_unit_PEG_Xvec_42__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_43__ap_done = PEG_Xvec_43__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_43__ap_idle = PEG_Xvec_43__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_43__ap_ready = PEG_Xvec_43__ap_ready;
  assign PEG_Xvec_43__ap_start = __tapa_fsm_unit_PEG_Xvec_43__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_44__ap_done = PEG_Xvec_44__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_44__ap_idle = PEG_Xvec_44__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_44__ap_ready = PEG_Xvec_44__ap_ready;
  assign PEG_Xvec_44__ap_start = __tapa_fsm_unit_PEG_Xvec_44__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_45__ap_done = PEG_Xvec_45__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_45__ap_idle = PEG_Xvec_45__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_45__ap_ready = PEG_Xvec_45__ap_ready;
  assign PEG_Xvec_45__ap_start = __tapa_fsm_unit_PEG_Xvec_45__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_46__ap_done = PEG_Xvec_46__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_46__ap_idle = PEG_Xvec_46__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_46__ap_ready = PEG_Xvec_46__ap_ready;
  assign PEG_Xvec_46__ap_start = __tapa_fsm_unit_PEG_Xvec_46__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_47__ap_done = PEG_Xvec_47__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_47__ap_idle = PEG_Xvec_47__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_47__ap_ready = PEG_Xvec_47__ap_ready;
  assign PEG_Xvec_47__ap_start = __tapa_fsm_unit_PEG_Xvec_47__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_4__ap_done = PEG_Xvec_4__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_4__ap_idle = PEG_Xvec_4__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_4__ap_ready = PEG_Xvec_4__ap_ready;
  assign PEG_Xvec_4__ap_start = __tapa_fsm_unit_PEG_Xvec_4__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_5__ap_done = PEG_Xvec_5__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_5__ap_idle = PEG_Xvec_5__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_5__ap_ready = PEG_Xvec_5__ap_ready;
  assign PEG_Xvec_5__ap_start = __tapa_fsm_unit_PEG_Xvec_5__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_6__ap_done = PEG_Xvec_6__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_6__ap_idle = PEG_Xvec_6__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_6__ap_ready = PEG_Xvec_6__ap_ready;
  assign PEG_Xvec_6__ap_start = __tapa_fsm_unit_PEG_Xvec_6__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_7__ap_done = PEG_Xvec_7__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_7__ap_idle = PEG_Xvec_7__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_7__ap_ready = PEG_Xvec_7__ap_ready;
  assign PEG_Xvec_7__ap_start = __tapa_fsm_unit_PEG_Xvec_7__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_8__ap_done = PEG_Xvec_8__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_8__ap_idle = PEG_Xvec_8__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_8__ap_ready = PEG_Xvec_8__ap_ready;
  assign PEG_Xvec_8__ap_start = __tapa_fsm_unit_PEG_Xvec_8__ap_start;
  assign __tapa_fsm_unit_PEG_Xvec_9__ap_done = PEG_Xvec_9__ap_done;
  assign __tapa_fsm_unit_PEG_Xvec_9__ap_idle = PEG_Xvec_9__ap_idle;
  assign __tapa_fsm_unit_PEG_Xvec_9__ap_ready = PEG_Xvec_9__ap_ready;
  assign PEG_Xvec_9__ap_start = __tapa_fsm_unit_PEG_Xvec_9__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_0__ap_done = PEG_Yvec_0__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_0__ap_idle = PEG_Yvec_0__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_0__ap_ready = PEG_Yvec_0__ap_ready;
  assign PEG_Yvec_0__ap_start = __tapa_fsm_unit_PEG_Yvec_0__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_10__ap_done = PEG_Yvec_10__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_10__ap_idle = PEG_Yvec_10__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_10__ap_ready = PEG_Yvec_10__ap_ready;
  assign PEG_Yvec_10__ap_start = __tapa_fsm_unit_PEG_Yvec_10__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_11__ap_done = PEG_Yvec_11__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_11__ap_idle = PEG_Yvec_11__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_11__ap_ready = PEG_Yvec_11__ap_ready;
  assign PEG_Yvec_11__ap_start = __tapa_fsm_unit_PEG_Yvec_11__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_12__ap_done = PEG_Yvec_12__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_12__ap_idle = PEG_Yvec_12__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_12__ap_ready = PEG_Yvec_12__ap_ready;
  assign PEG_Yvec_12__ap_start = __tapa_fsm_unit_PEG_Yvec_12__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_13__ap_done = PEG_Yvec_13__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_13__ap_idle = PEG_Yvec_13__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_13__ap_ready = PEG_Yvec_13__ap_ready;
  assign PEG_Yvec_13__ap_start = __tapa_fsm_unit_PEG_Yvec_13__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_14__ap_done = PEG_Yvec_14__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_14__ap_idle = PEG_Yvec_14__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_14__ap_ready = PEG_Yvec_14__ap_ready;
  assign PEG_Yvec_14__ap_start = __tapa_fsm_unit_PEG_Yvec_14__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_15__ap_done = PEG_Yvec_15__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_15__ap_idle = PEG_Yvec_15__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_15__ap_ready = PEG_Yvec_15__ap_ready;
  assign PEG_Yvec_15__ap_start = __tapa_fsm_unit_PEG_Yvec_15__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_16__ap_done = PEG_Yvec_16__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_16__ap_idle = PEG_Yvec_16__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_16__ap_ready = PEG_Yvec_16__ap_ready;
  assign PEG_Yvec_16__ap_start = __tapa_fsm_unit_PEG_Yvec_16__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_17__ap_done = PEG_Yvec_17__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_17__ap_idle = PEG_Yvec_17__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_17__ap_ready = PEG_Yvec_17__ap_ready;
  assign PEG_Yvec_17__ap_start = __tapa_fsm_unit_PEG_Yvec_17__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_18__ap_done = PEG_Yvec_18__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_18__ap_idle = PEG_Yvec_18__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_18__ap_ready = PEG_Yvec_18__ap_ready;
  assign PEG_Yvec_18__ap_start = __tapa_fsm_unit_PEG_Yvec_18__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_19__ap_done = PEG_Yvec_19__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_19__ap_idle = PEG_Yvec_19__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_19__ap_ready = PEG_Yvec_19__ap_ready;
  assign PEG_Yvec_19__ap_start = __tapa_fsm_unit_PEG_Yvec_19__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_1__ap_done = PEG_Yvec_1__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_1__ap_idle = PEG_Yvec_1__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_1__ap_ready = PEG_Yvec_1__ap_ready;
  assign PEG_Yvec_1__ap_start = __tapa_fsm_unit_PEG_Yvec_1__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_20__ap_done = PEG_Yvec_20__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_20__ap_idle = PEG_Yvec_20__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_20__ap_ready = PEG_Yvec_20__ap_ready;
  assign PEG_Yvec_20__ap_start = __tapa_fsm_unit_PEG_Yvec_20__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_21__ap_done = PEG_Yvec_21__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_21__ap_idle = PEG_Yvec_21__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_21__ap_ready = PEG_Yvec_21__ap_ready;
  assign PEG_Yvec_21__ap_start = __tapa_fsm_unit_PEG_Yvec_21__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_22__ap_done = PEG_Yvec_22__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_22__ap_idle = PEG_Yvec_22__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_22__ap_ready = PEG_Yvec_22__ap_ready;
  assign PEG_Yvec_22__ap_start = __tapa_fsm_unit_PEG_Yvec_22__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_23__ap_done = PEG_Yvec_23__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_23__ap_idle = PEG_Yvec_23__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_23__ap_ready = PEG_Yvec_23__ap_ready;
  assign PEG_Yvec_23__ap_start = __tapa_fsm_unit_PEG_Yvec_23__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_24__ap_done = PEG_Yvec_24__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_24__ap_idle = PEG_Yvec_24__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_24__ap_ready = PEG_Yvec_24__ap_ready;
  assign PEG_Yvec_24__ap_start = __tapa_fsm_unit_PEG_Yvec_24__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_25__ap_done = PEG_Yvec_25__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_25__ap_idle = PEG_Yvec_25__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_25__ap_ready = PEG_Yvec_25__ap_ready;
  assign PEG_Yvec_25__ap_start = __tapa_fsm_unit_PEG_Yvec_25__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_26__ap_done = PEG_Yvec_26__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_26__ap_idle = PEG_Yvec_26__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_26__ap_ready = PEG_Yvec_26__ap_ready;
  assign PEG_Yvec_26__ap_start = __tapa_fsm_unit_PEG_Yvec_26__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_27__ap_done = PEG_Yvec_27__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_27__ap_idle = PEG_Yvec_27__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_27__ap_ready = PEG_Yvec_27__ap_ready;
  assign PEG_Yvec_27__ap_start = __tapa_fsm_unit_PEG_Yvec_27__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_28__ap_done = PEG_Yvec_28__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_28__ap_idle = PEG_Yvec_28__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_28__ap_ready = PEG_Yvec_28__ap_ready;
  assign PEG_Yvec_28__ap_start = __tapa_fsm_unit_PEG_Yvec_28__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_29__ap_done = PEG_Yvec_29__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_29__ap_idle = PEG_Yvec_29__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_29__ap_ready = PEG_Yvec_29__ap_ready;
  assign PEG_Yvec_29__ap_start = __tapa_fsm_unit_PEG_Yvec_29__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_2__ap_done = PEG_Yvec_2__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_2__ap_idle = PEG_Yvec_2__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_2__ap_ready = PEG_Yvec_2__ap_ready;
  assign PEG_Yvec_2__ap_start = __tapa_fsm_unit_PEG_Yvec_2__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_30__ap_done = PEG_Yvec_30__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_30__ap_idle = PEG_Yvec_30__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_30__ap_ready = PEG_Yvec_30__ap_ready;
  assign PEG_Yvec_30__ap_start = __tapa_fsm_unit_PEG_Yvec_30__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_31__ap_done = PEG_Yvec_31__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_31__ap_idle = PEG_Yvec_31__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_31__ap_ready = PEG_Yvec_31__ap_ready;
  assign PEG_Yvec_31__ap_start = __tapa_fsm_unit_PEG_Yvec_31__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_32__ap_done = PEG_Yvec_32__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_32__ap_idle = PEG_Yvec_32__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_32__ap_ready = PEG_Yvec_32__ap_ready;
  assign PEG_Yvec_32__ap_start = __tapa_fsm_unit_PEG_Yvec_32__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_33__ap_done = PEG_Yvec_33__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_33__ap_idle = PEG_Yvec_33__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_33__ap_ready = PEG_Yvec_33__ap_ready;
  assign PEG_Yvec_33__ap_start = __tapa_fsm_unit_PEG_Yvec_33__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_34__ap_done = PEG_Yvec_34__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_34__ap_idle = PEG_Yvec_34__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_34__ap_ready = PEG_Yvec_34__ap_ready;
  assign PEG_Yvec_34__ap_start = __tapa_fsm_unit_PEG_Yvec_34__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_35__ap_done = PEG_Yvec_35__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_35__ap_idle = PEG_Yvec_35__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_35__ap_ready = PEG_Yvec_35__ap_ready;
  assign PEG_Yvec_35__ap_start = __tapa_fsm_unit_PEG_Yvec_35__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_36__ap_done = PEG_Yvec_36__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_36__ap_idle = PEG_Yvec_36__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_36__ap_ready = PEG_Yvec_36__ap_ready;
  assign PEG_Yvec_36__ap_start = __tapa_fsm_unit_PEG_Yvec_36__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_37__ap_done = PEG_Yvec_37__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_37__ap_idle = PEG_Yvec_37__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_37__ap_ready = PEG_Yvec_37__ap_ready;
  assign PEG_Yvec_37__ap_start = __tapa_fsm_unit_PEG_Yvec_37__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_38__ap_done = PEG_Yvec_38__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_38__ap_idle = PEG_Yvec_38__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_38__ap_ready = PEG_Yvec_38__ap_ready;
  assign PEG_Yvec_38__ap_start = __tapa_fsm_unit_PEG_Yvec_38__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_39__ap_done = PEG_Yvec_39__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_39__ap_idle = PEG_Yvec_39__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_39__ap_ready = PEG_Yvec_39__ap_ready;
  assign PEG_Yvec_39__ap_start = __tapa_fsm_unit_PEG_Yvec_39__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_3__ap_done = PEG_Yvec_3__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_3__ap_idle = PEG_Yvec_3__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_3__ap_ready = PEG_Yvec_3__ap_ready;
  assign PEG_Yvec_3__ap_start = __tapa_fsm_unit_PEG_Yvec_3__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_40__ap_done = PEG_Yvec_40__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_40__ap_idle = PEG_Yvec_40__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_40__ap_ready = PEG_Yvec_40__ap_ready;
  assign PEG_Yvec_40__ap_start = __tapa_fsm_unit_PEG_Yvec_40__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_41__ap_done = PEG_Yvec_41__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_41__ap_idle = PEG_Yvec_41__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_41__ap_ready = PEG_Yvec_41__ap_ready;
  assign PEG_Yvec_41__ap_start = __tapa_fsm_unit_PEG_Yvec_41__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_42__ap_done = PEG_Yvec_42__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_42__ap_idle = PEG_Yvec_42__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_42__ap_ready = PEG_Yvec_42__ap_ready;
  assign PEG_Yvec_42__ap_start = __tapa_fsm_unit_PEG_Yvec_42__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_43__ap_done = PEG_Yvec_43__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_43__ap_idle = PEG_Yvec_43__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_43__ap_ready = PEG_Yvec_43__ap_ready;
  assign PEG_Yvec_43__ap_start = __tapa_fsm_unit_PEG_Yvec_43__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_44__ap_done = PEG_Yvec_44__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_44__ap_idle = PEG_Yvec_44__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_44__ap_ready = PEG_Yvec_44__ap_ready;
  assign PEG_Yvec_44__ap_start = __tapa_fsm_unit_PEG_Yvec_44__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_45__ap_done = PEG_Yvec_45__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_45__ap_idle = PEG_Yvec_45__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_45__ap_ready = PEG_Yvec_45__ap_ready;
  assign PEG_Yvec_45__ap_start = __tapa_fsm_unit_PEG_Yvec_45__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_46__ap_done = PEG_Yvec_46__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_46__ap_idle = PEG_Yvec_46__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_46__ap_ready = PEG_Yvec_46__ap_ready;
  assign PEG_Yvec_46__ap_start = __tapa_fsm_unit_PEG_Yvec_46__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_47__ap_done = PEG_Yvec_47__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_47__ap_idle = PEG_Yvec_47__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_47__ap_ready = PEG_Yvec_47__ap_ready;
  assign PEG_Yvec_47__ap_start = __tapa_fsm_unit_PEG_Yvec_47__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_4__ap_done = PEG_Yvec_4__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_4__ap_idle = PEG_Yvec_4__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_4__ap_ready = PEG_Yvec_4__ap_ready;
  assign PEG_Yvec_4__ap_start = __tapa_fsm_unit_PEG_Yvec_4__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_5__ap_done = PEG_Yvec_5__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_5__ap_idle = PEG_Yvec_5__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_5__ap_ready = PEG_Yvec_5__ap_ready;
  assign PEG_Yvec_5__ap_start = __tapa_fsm_unit_PEG_Yvec_5__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_6__ap_done = PEG_Yvec_6__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_6__ap_idle = PEG_Yvec_6__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_6__ap_ready = PEG_Yvec_6__ap_ready;
  assign PEG_Yvec_6__ap_start = __tapa_fsm_unit_PEG_Yvec_6__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_7__ap_done = PEG_Yvec_7__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_7__ap_idle = PEG_Yvec_7__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_7__ap_ready = PEG_Yvec_7__ap_ready;
  assign PEG_Yvec_7__ap_start = __tapa_fsm_unit_PEG_Yvec_7__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_8__ap_done = PEG_Yvec_8__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_8__ap_idle = PEG_Yvec_8__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_8__ap_ready = PEG_Yvec_8__ap_ready;
  assign PEG_Yvec_8__ap_start = __tapa_fsm_unit_PEG_Yvec_8__ap_start;
  assign __tapa_fsm_unit_PEG_Yvec_9__ap_done = PEG_Yvec_9__ap_done;
  assign __tapa_fsm_unit_PEG_Yvec_9__ap_idle = PEG_Yvec_9__ap_idle;
  assign __tapa_fsm_unit_PEG_Yvec_9__ap_ready = PEG_Yvec_9__ap_ready;
  assign PEG_Yvec_9__ap_start = __tapa_fsm_unit_PEG_Yvec_9__ap_start;
  assign __tapa_fsm_unit_P_N = P_N;
  assign __tapa_fsm_unit_alpha_u = alpha_u;
  assign __tapa_fsm_unit_ap_clk = ap_clk;
  assign ap_done = __tapa_fsm_unit_ap_done;
  assign ap_idle = __tapa_fsm_unit_ap_idle;
  assign ap_ready = __tapa_fsm_unit_ap_ready;
  assign __tapa_fsm_unit_ap_rst_n = ap_rst_n;
  assign __tapa_fsm_unit_ap_start = ap_start;
  assign __tapa_fsm_unit_beta_u = beta_u;
  assign black_hole_float_v16_0__ap_start = __tapa_fsm_unit_black_hole_float_v16_0__ap_start;
  assign black_hole_int_0__ap_start = __tapa_fsm_unit_black_hole_int_0__ap_start;
  assign __tapa_fsm_unit_edge_list_ch_0 = edge_list_ch_0;
  assign __tapa_fsm_unit_edge_list_ch_1 = edge_list_ch_1;
  assign __tapa_fsm_unit_edge_list_ch_10 = edge_list_ch_10;
  assign __tapa_fsm_unit_edge_list_ch_11 = edge_list_ch_11;
  assign __tapa_fsm_unit_edge_list_ch_12 = edge_list_ch_12;
  assign __tapa_fsm_unit_edge_list_ch_13 = edge_list_ch_13;
  assign __tapa_fsm_unit_edge_list_ch_14 = edge_list_ch_14;
  assign __tapa_fsm_unit_edge_list_ch_15 = edge_list_ch_15;
  assign __tapa_fsm_unit_edge_list_ch_16 = edge_list_ch_16;
  assign __tapa_fsm_unit_edge_list_ch_17 = edge_list_ch_17;
  assign __tapa_fsm_unit_edge_list_ch_18 = edge_list_ch_18;
  assign __tapa_fsm_unit_edge_list_ch_19 = edge_list_ch_19;
  assign __tapa_fsm_unit_edge_list_ch_2 = edge_list_ch_2;
  assign __tapa_fsm_unit_edge_list_ch_20 = edge_list_ch_20;
  assign __tapa_fsm_unit_edge_list_ch_21 = edge_list_ch_21;
  assign __tapa_fsm_unit_edge_list_ch_22 = edge_list_ch_22;
  assign __tapa_fsm_unit_edge_list_ch_23 = edge_list_ch_23;
  assign __tapa_fsm_unit_edge_list_ch_24 = edge_list_ch_24;
  assign __tapa_fsm_unit_edge_list_ch_25 = edge_list_ch_25;
  assign __tapa_fsm_unit_edge_list_ch_26 = edge_list_ch_26;
  assign __tapa_fsm_unit_edge_list_ch_27 = edge_list_ch_27;
  assign __tapa_fsm_unit_edge_list_ch_28 = edge_list_ch_28;
  assign __tapa_fsm_unit_edge_list_ch_29 = edge_list_ch_29;
  assign __tapa_fsm_unit_edge_list_ch_3 = edge_list_ch_3;
  assign __tapa_fsm_unit_edge_list_ch_30 = edge_list_ch_30;
  assign __tapa_fsm_unit_edge_list_ch_31 = edge_list_ch_31;
  assign __tapa_fsm_unit_edge_list_ch_32 = edge_list_ch_32;
  assign __tapa_fsm_unit_edge_list_ch_33 = edge_list_ch_33;
  assign __tapa_fsm_unit_edge_list_ch_34 = edge_list_ch_34;
  assign __tapa_fsm_unit_edge_list_ch_35 = edge_list_ch_35;
  assign __tapa_fsm_unit_edge_list_ch_36 = edge_list_ch_36;
  assign __tapa_fsm_unit_edge_list_ch_37 = edge_list_ch_37;
  assign __tapa_fsm_unit_edge_list_ch_38 = edge_list_ch_38;
  assign __tapa_fsm_unit_edge_list_ch_39 = edge_list_ch_39;
  assign __tapa_fsm_unit_edge_list_ch_4 = edge_list_ch_4;
  assign __tapa_fsm_unit_edge_list_ch_40 = edge_list_ch_40;
  assign __tapa_fsm_unit_edge_list_ch_41 = edge_list_ch_41;
  assign __tapa_fsm_unit_edge_list_ch_42 = edge_list_ch_42;
  assign __tapa_fsm_unit_edge_list_ch_43 = edge_list_ch_43;
  assign __tapa_fsm_unit_edge_list_ch_44 = edge_list_ch_44;
  assign __tapa_fsm_unit_edge_list_ch_45 = edge_list_ch_45;
  assign __tapa_fsm_unit_edge_list_ch_46 = edge_list_ch_46;
  assign __tapa_fsm_unit_edge_list_ch_47 = edge_list_ch_47;
  assign __tapa_fsm_unit_edge_list_ch_5 = edge_list_ch_5;
  assign __tapa_fsm_unit_edge_list_ch_6 = edge_list_ch_6;
  assign __tapa_fsm_unit_edge_list_ch_7 = edge_list_ch_7;
  assign __tapa_fsm_unit_edge_list_ch_8 = edge_list_ch_8;
  assign __tapa_fsm_unit_edge_list_ch_9 = edge_list_ch_9;
  assign __tapa_fsm_unit_edge_list_ptr = edge_list_ptr;
  assign read_A_0___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_0___NUM_A_LEN__q0;
  assign read_A_0___P_N__q0 = __tapa_fsm_unit_read_A_0___P_N__q0;
  assign read_A_0___edge_list_ch_0__q0 = __tapa_fsm_unit_read_A_0___edge_list_ch_0__q0;
  assign __tapa_fsm_unit_read_A_0__ap_done = read_A_0__ap_done;
  assign __tapa_fsm_unit_read_A_0__ap_idle = read_A_0__ap_idle;
  assign __tapa_fsm_unit_read_A_0__ap_ready = read_A_0__ap_ready;
  assign read_A_0__ap_start = __tapa_fsm_unit_read_A_0__ap_start;
  assign read_A_10___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_10___NUM_A_LEN__q0;
  assign read_A_10___P_N__q0 = __tapa_fsm_unit_read_A_10___P_N__q0;
  assign read_A_10___edge_list_ch_10__q0 = __tapa_fsm_unit_read_A_10___edge_list_ch_10__q0;
  assign __tapa_fsm_unit_read_A_10__ap_done = read_A_10__ap_done;
  assign __tapa_fsm_unit_read_A_10__ap_idle = read_A_10__ap_idle;
  assign __tapa_fsm_unit_read_A_10__ap_ready = read_A_10__ap_ready;
  assign read_A_10__ap_start = __tapa_fsm_unit_read_A_10__ap_start;
  assign read_A_11___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_11___NUM_A_LEN__q0;
  assign read_A_11___P_N__q0 = __tapa_fsm_unit_read_A_11___P_N__q0;
  assign read_A_11___edge_list_ch_11__q0 = __tapa_fsm_unit_read_A_11___edge_list_ch_11__q0;
  assign __tapa_fsm_unit_read_A_11__ap_done = read_A_11__ap_done;
  assign __tapa_fsm_unit_read_A_11__ap_idle = read_A_11__ap_idle;
  assign __tapa_fsm_unit_read_A_11__ap_ready = read_A_11__ap_ready;
  assign read_A_11__ap_start = __tapa_fsm_unit_read_A_11__ap_start;
  assign read_A_12___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_12___NUM_A_LEN__q0;
  assign read_A_12___P_N__q0 = __tapa_fsm_unit_read_A_12___P_N__q0;
  assign read_A_12___edge_list_ch_12__q0 = __tapa_fsm_unit_read_A_12___edge_list_ch_12__q0;
  assign __tapa_fsm_unit_read_A_12__ap_done = read_A_12__ap_done;
  assign __tapa_fsm_unit_read_A_12__ap_idle = read_A_12__ap_idle;
  assign __tapa_fsm_unit_read_A_12__ap_ready = read_A_12__ap_ready;
  assign read_A_12__ap_start = __tapa_fsm_unit_read_A_12__ap_start;
  assign read_A_13___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_13___NUM_A_LEN__q0;
  assign read_A_13___P_N__q0 = __tapa_fsm_unit_read_A_13___P_N__q0;
  assign read_A_13___edge_list_ch_13__q0 = __tapa_fsm_unit_read_A_13___edge_list_ch_13__q0;
  assign __tapa_fsm_unit_read_A_13__ap_done = read_A_13__ap_done;
  assign __tapa_fsm_unit_read_A_13__ap_idle = read_A_13__ap_idle;
  assign __tapa_fsm_unit_read_A_13__ap_ready = read_A_13__ap_ready;
  assign read_A_13__ap_start = __tapa_fsm_unit_read_A_13__ap_start;
  assign read_A_14___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_14___NUM_A_LEN__q0;
  assign read_A_14___P_N__q0 = __tapa_fsm_unit_read_A_14___P_N__q0;
  assign read_A_14___edge_list_ch_14__q0 = __tapa_fsm_unit_read_A_14___edge_list_ch_14__q0;
  assign __tapa_fsm_unit_read_A_14__ap_done = read_A_14__ap_done;
  assign __tapa_fsm_unit_read_A_14__ap_idle = read_A_14__ap_idle;
  assign __tapa_fsm_unit_read_A_14__ap_ready = read_A_14__ap_ready;
  assign read_A_14__ap_start = __tapa_fsm_unit_read_A_14__ap_start;
  assign read_A_15___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_15___NUM_A_LEN__q0;
  assign read_A_15___P_N__q0 = __tapa_fsm_unit_read_A_15___P_N__q0;
  assign read_A_15___edge_list_ch_15__q0 = __tapa_fsm_unit_read_A_15___edge_list_ch_15__q0;
  assign __tapa_fsm_unit_read_A_15__ap_done = read_A_15__ap_done;
  assign __tapa_fsm_unit_read_A_15__ap_idle = read_A_15__ap_idle;
  assign __tapa_fsm_unit_read_A_15__ap_ready = read_A_15__ap_ready;
  assign read_A_15__ap_start = __tapa_fsm_unit_read_A_15__ap_start;
  assign read_A_16___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_16___NUM_A_LEN__q0;
  assign read_A_16___P_N__q0 = __tapa_fsm_unit_read_A_16___P_N__q0;
  assign read_A_16___edge_list_ch_16__q0 = __tapa_fsm_unit_read_A_16___edge_list_ch_16__q0;
  assign __tapa_fsm_unit_read_A_16__ap_done = read_A_16__ap_done;
  assign __tapa_fsm_unit_read_A_16__ap_idle = read_A_16__ap_idle;
  assign __tapa_fsm_unit_read_A_16__ap_ready = read_A_16__ap_ready;
  assign read_A_16__ap_start = __tapa_fsm_unit_read_A_16__ap_start;
  assign read_A_17___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_17___NUM_A_LEN__q0;
  assign read_A_17___P_N__q0 = __tapa_fsm_unit_read_A_17___P_N__q0;
  assign read_A_17___edge_list_ch_17__q0 = __tapa_fsm_unit_read_A_17___edge_list_ch_17__q0;
  assign __tapa_fsm_unit_read_A_17__ap_done = read_A_17__ap_done;
  assign __tapa_fsm_unit_read_A_17__ap_idle = read_A_17__ap_idle;
  assign __tapa_fsm_unit_read_A_17__ap_ready = read_A_17__ap_ready;
  assign read_A_17__ap_start = __tapa_fsm_unit_read_A_17__ap_start;
  assign read_A_18___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_18___NUM_A_LEN__q0;
  assign read_A_18___P_N__q0 = __tapa_fsm_unit_read_A_18___P_N__q0;
  assign read_A_18___edge_list_ch_18__q0 = __tapa_fsm_unit_read_A_18___edge_list_ch_18__q0;
  assign __tapa_fsm_unit_read_A_18__ap_done = read_A_18__ap_done;
  assign __tapa_fsm_unit_read_A_18__ap_idle = read_A_18__ap_idle;
  assign __tapa_fsm_unit_read_A_18__ap_ready = read_A_18__ap_ready;
  assign read_A_18__ap_start = __tapa_fsm_unit_read_A_18__ap_start;
  assign read_A_19___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_19___NUM_A_LEN__q0;
  assign read_A_19___P_N__q0 = __tapa_fsm_unit_read_A_19___P_N__q0;
  assign read_A_19___edge_list_ch_19__q0 = __tapa_fsm_unit_read_A_19___edge_list_ch_19__q0;
  assign __tapa_fsm_unit_read_A_19__ap_done = read_A_19__ap_done;
  assign __tapa_fsm_unit_read_A_19__ap_idle = read_A_19__ap_idle;
  assign __tapa_fsm_unit_read_A_19__ap_ready = read_A_19__ap_ready;
  assign read_A_19__ap_start = __tapa_fsm_unit_read_A_19__ap_start;
  assign read_A_1___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_1___NUM_A_LEN__q0;
  assign read_A_1___P_N__q0 = __tapa_fsm_unit_read_A_1___P_N__q0;
  assign read_A_1___edge_list_ch_1__q0 = __tapa_fsm_unit_read_A_1___edge_list_ch_1__q0;
  assign __tapa_fsm_unit_read_A_1__ap_done = read_A_1__ap_done;
  assign __tapa_fsm_unit_read_A_1__ap_idle = read_A_1__ap_idle;
  assign __tapa_fsm_unit_read_A_1__ap_ready = read_A_1__ap_ready;
  assign read_A_1__ap_start = __tapa_fsm_unit_read_A_1__ap_start;
  assign read_A_20___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_20___NUM_A_LEN__q0;
  assign read_A_20___P_N__q0 = __tapa_fsm_unit_read_A_20___P_N__q0;
  assign read_A_20___edge_list_ch_20__q0 = __tapa_fsm_unit_read_A_20___edge_list_ch_20__q0;
  assign __tapa_fsm_unit_read_A_20__ap_done = read_A_20__ap_done;
  assign __tapa_fsm_unit_read_A_20__ap_idle = read_A_20__ap_idle;
  assign __tapa_fsm_unit_read_A_20__ap_ready = read_A_20__ap_ready;
  assign read_A_20__ap_start = __tapa_fsm_unit_read_A_20__ap_start;
  assign read_A_21___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_21___NUM_A_LEN__q0;
  assign read_A_21___P_N__q0 = __tapa_fsm_unit_read_A_21___P_N__q0;
  assign read_A_21___edge_list_ch_21__q0 = __tapa_fsm_unit_read_A_21___edge_list_ch_21__q0;
  assign __tapa_fsm_unit_read_A_21__ap_done = read_A_21__ap_done;
  assign __tapa_fsm_unit_read_A_21__ap_idle = read_A_21__ap_idle;
  assign __tapa_fsm_unit_read_A_21__ap_ready = read_A_21__ap_ready;
  assign read_A_21__ap_start = __tapa_fsm_unit_read_A_21__ap_start;
  assign read_A_22___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_22___NUM_A_LEN__q0;
  assign read_A_22___P_N__q0 = __tapa_fsm_unit_read_A_22___P_N__q0;
  assign read_A_22___edge_list_ch_22__q0 = __tapa_fsm_unit_read_A_22___edge_list_ch_22__q0;
  assign __tapa_fsm_unit_read_A_22__ap_done = read_A_22__ap_done;
  assign __tapa_fsm_unit_read_A_22__ap_idle = read_A_22__ap_idle;
  assign __tapa_fsm_unit_read_A_22__ap_ready = read_A_22__ap_ready;
  assign read_A_22__ap_start = __tapa_fsm_unit_read_A_22__ap_start;
  assign read_A_23___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_23___NUM_A_LEN__q0;
  assign read_A_23___P_N__q0 = __tapa_fsm_unit_read_A_23___P_N__q0;
  assign read_A_23___edge_list_ch_23__q0 = __tapa_fsm_unit_read_A_23___edge_list_ch_23__q0;
  assign __tapa_fsm_unit_read_A_23__ap_done = read_A_23__ap_done;
  assign __tapa_fsm_unit_read_A_23__ap_idle = read_A_23__ap_idle;
  assign __tapa_fsm_unit_read_A_23__ap_ready = read_A_23__ap_ready;
  assign read_A_23__ap_start = __tapa_fsm_unit_read_A_23__ap_start;
  assign read_A_24___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_24___NUM_A_LEN__q0;
  assign read_A_24___P_N__q0 = __tapa_fsm_unit_read_A_24___P_N__q0;
  assign read_A_24___edge_list_ch_24__q0 = __tapa_fsm_unit_read_A_24___edge_list_ch_24__q0;
  assign __tapa_fsm_unit_read_A_24__ap_done = read_A_24__ap_done;
  assign __tapa_fsm_unit_read_A_24__ap_idle = read_A_24__ap_idle;
  assign __tapa_fsm_unit_read_A_24__ap_ready = read_A_24__ap_ready;
  assign read_A_24__ap_start = __tapa_fsm_unit_read_A_24__ap_start;
  assign read_A_25___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_25___NUM_A_LEN__q0;
  assign read_A_25___P_N__q0 = __tapa_fsm_unit_read_A_25___P_N__q0;
  assign read_A_25___edge_list_ch_25__q0 = __tapa_fsm_unit_read_A_25___edge_list_ch_25__q0;
  assign __tapa_fsm_unit_read_A_25__ap_done = read_A_25__ap_done;
  assign __tapa_fsm_unit_read_A_25__ap_idle = read_A_25__ap_idle;
  assign __tapa_fsm_unit_read_A_25__ap_ready = read_A_25__ap_ready;
  assign read_A_25__ap_start = __tapa_fsm_unit_read_A_25__ap_start;
  assign read_A_26___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_26___NUM_A_LEN__q0;
  assign read_A_26___P_N__q0 = __tapa_fsm_unit_read_A_26___P_N__q0;
  assign read_A_26___edge_list_ch_26__q0 = __tapa_fsm_unit_read_A_26___edge_list_ch_26__q0;
  assign __tapa_fsm_unit_read_A_26__ap_done = read_A_26__ap_done;
  assign __tapa_fsm_unit_read_A_26__ap_idle = read_A_26__ap_idle;
  assign __tapa_fsm_unit_read_A_26__ap_ready = read_A_26__ap_ready;
  assign read_A_26__ap_start = __tapa_fsm_unit_read_A_26__ap_start;
  assign read_A_27___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_27___NUM_A_LEN__q0;
  assign read_A_27___P_N__q0 = __tapa_fsm_unit_read_A_27___P_N__q0;
  assign read_A_27___edge_list_ch_27__q0 = __tapa_fsm_unit_read_A_27___edge_list_ch_27__q0;
  assign __tapa_fsm_unit_read_A_27__ap_done = read_A_27__ap_done;
  assign __tapa_fsm_unit_read_A_27__ap_idle = read_A_27__ap_idle;
  assign __tapa_fsm_unit_read_A_27__ap_ready = read_A_27__ap_ready;
  assign read_A_27__ap_start = __tapa_fsm_unit_read_A_27__ap_start;
  assign read_A_28___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_28___NUM_A_LEN__q0;
  assign read_A_28___P_N__q0 = __tapa_fsm_unit_read_A_28___P_N__q0;
  assign read_A_28___edge_list_ch_28__q0 = __tapa_fsm_unit_read_A_28___edge_list_ch_28__q0;
  assign __tapa_fsm_unit_read_A_28__ap_done = read_A_28__ap_done;
  assign __tapa_fsm_unit_read_A_28__ap_idle = read_A_28__ap_idle;
  assign __tapa_fsm_unit_read_A_28__ap_ready = read_A_28__ap_ready;
  assign read_A_28__ap_start = __tapa_fsm_unit_read_A_28__ap_start;
  assign read_A_29___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_29___NUM_A_LEN__q0;
  assign read_A_29___P_N__q0 = __tapa_fsm_unit_read_A_29___P_N__q0;
  assign read_A_29___edge_list_ch_29__q0 = __tapa_fsm_unit_read_A_29___edge_list_ch_29__q0;
  assign __tapa_fsm_unit_read_A_29__ap_done = read_A_29__ap_done;
  assign __tapa_fsm_unit_read_A_29__ap_idle = read_A_29__ap_idle;
  assign __tapa_fsm_unit_read_A_29__ap_ready = read_A_29__ap_ready;
  assign read_A_29__ap_start = __tapa_fsm_unit_read_A_29__ap_start;
  assign read_A_2___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_2___NUM_A_LEN__q0;
  assign read_A_2___P_N__q0 = __tapa_fsm_unit_read_A_2___P_N__q0;
  assign read_A_2___edge_list_ch_2__q0 = __tapa_fsm_unit_read_A_2___edge_list_ch_2__q0;
  assign __tapa_fsm_unit_read_A_2__ap_done = read_A_2__ap_done;
  assign __tapa_fsm_unit_read_A_2__ap_idle = read_A_2__ap_idle;
  assign __tapa_fsm_unit_read_A_2__ap_ready = read_A_2__ap_ready;
  assign read_A_2__ap_start = __tapa_fsm_unit_read_A_2__ap_start;
  assign read_A_30___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_30___NUM_A_LEN__q0;
  assign read_A_30___P_N__q0 = __tapa_fsm_unit_read_A_30___P_N__q0;
  assign read_A_30___edge_list_ch_30__q0 = __tapa_fsm_unit_read_A_30___edge_list_ch_30__q0;
  assign __tapa_fsm_unit_read_A_30__ap_done = read_A_30__ap_done;
  assign __tapa_fsm_unit_read_A_30__ap_idle = read_A_30__ap_idle;
  assign __tapa_fsm_unit_read_A_30__ap_ready = read_A_30__ap_ready;
  assign read_A_30__ap_start = __tapa_fsm_unit_read_A_30__ap_start;
  assign read_A_31___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_31___NUM_A_LEN__q0;
  assign read_A_31___P_N__q0 = __tapa_fsm_unit_read_A_31___P_N__q0;
  assign read_A_31___edge_list_ch_31__q0 = __tapa_fsm_unit_read_A_31___edge_list_ch_31__q0;
  assign __tapa_fsm_unit_read_A_31__ap_done = read_A_31__ap_done;
  assign __tapa_fsm_unit_read_A_31__ap_idle = read_A_31__ap_idle;
  assign __tapa_fsm_unit_read_A_31__ap_ready = read_A_31__ap_ready;
  assign read_A_31__ap_start = __tapa_fsm_unit_read_A_31__ap_start;
  assign read_A_32___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_32___NUM_A_LEN__q0;
  assign read_A_32___P_N__q0 = __tapa_fsm_unit_read_A_32___P_N__q0;
  assign read_A_32___edge_list_ch_32__q0 = __tapa_fsm_unit_read_A_32___edge_list_ch_32__q0;
  assign __tapa_fsm_unit_read_A_32__ap_done = read_A_32__ap_done;
  assign __tapa_fsm_unit_read_A_32__ap_idle = read_A_32__ap_idle;
  assign __tapa_fsm_unit_read_A_32__ap_ready = read_A_32__ap_ready;
  assign read_A_32__ap_start = __tapa_fsm_unit_read_A_32__ap_start;
  assign read_A_33___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_33___NUM_A_LEN__q0;
  assign read_A_33___P_N__q0 = __tapa_fsm_unit_read_A_33___P_N__q0;
  assign read_A_33___edge_list_ch_33__q0 = __tapa_fsm_unit_read_A_33___edge_list_ch_33__q0;
  assign __tapa_fsm_unit_read_A_33__ap_done = read_A_33__ap_done;
  assign __tapa_fsm_unit_read_A_33__ap_idle = read_A_33__ap_idle;
  assign __tapa_fsm_unit_read_A_33__ap_ready = read_A_33__ap_ready;
  assign read_A_33__ap_start = __tapa_fsm_unit_read_A_33__ap_start;
  assign read_A_34___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_34___NUM_A_LEN__q0;
  assign read_A_34___P_N__q0 = __tapa_fsm_unit_read_A_34___P_N__q0;
  assign read_A_34___edge_list_ch_34__q0 = __tapa_fsm_unit_read_A_34___edge_list_ch_34__q0;
  assign __tapa_fsm_unit_read_A_34__ap_done = read_A_34__ap_done;
  assign __tapa_fsm_unit_read_A_34__ap_idle = read_A_34__ap_idle;
  assign __tapa_fsm_unit_read_A_34__ap_ready = read_A_34__ap_ready;
  assign read_A_34__ap_start = __tapa_fsm_unit_read_A_34__ap_start;
  assign read_A_35___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_35___NUM_A_LEN__q0;
  assign read_A_35___P_N__q0 = __tapa_fsm_unit_read_A_35___P_N__q0;
  assign read_A_35___edge_list_ch_35__q0 = __tapa_fsm_unit_read_A_35___edge_list_ch_35__q0;
  assign __tapa_fsm_unit_read_A_35__ap_done = read_A_35__ap_done;
  assign __tapa_fsm_unit_read_A_35__ap_idle = read_A_35__ap_idle;
  assign __tapa_fsm_unit_read_A_35__ap_ready = read_A_35__ap_ready;
  assign read_A_35__ap_start = __tapa_fsm_unit_read_A_35__ap_start;
  assign read_A_36___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_36___NUM_A_LEN__q0;
  assign read_A_36___P_N__q0 = __tapa_fsm_unit_read_A_36___P_N__q0;
  assign read_A_36___edge_list_ch_36__q0 = __tapa_fsm_unit_read_A_36___edge_list_ch_36__q0;
  assign __tapa_fsm_unit_read_A_36__ap_done = read_A_36__ap_done;
  assign __tapa_fsm_unit_read_A_36__ap_idle = read_A_36__ap_idle;
  assign __tapa_fsm_unit_read_A_36__ap_ready = read_A_36__ap_ready;
  assign read_A_36__ap_start = __tapa_fsm_unit_read_A_36__ap_start;
  assign read_A_37___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_37___NUM_A_LEN__q0;
  assign read_A_37___P_N__q0 = __tapa_fsm_unit_read_A_37___P_N__q0;
  assign read_A_37___edge_list_ch_37__q0 = __tapa_fsm_unit_read_A_37___edge_list_ch_37__q0;
  assign __tapa_fsm_unit_read_A_37__ap_done = read_A_37__ap_done;
  assign __tapa_fsm_unit_read_A_37__ap_idle = read_A_37__ap_idle;
  assign __tapa_fsm_unit_read_A_37__ap_ready = read_A_37__ap_ready;
  assign read_A_37__ap_start = __tapa_fsm_unit_read_A_37__ap_start;
  assign read_A_38___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_38___NUM_A_LEN__q0;
  assign read_A_38___P_N__q0 = __tapa_fsm_unit_read_A_38___P_N__q0;
  assign read_A_38___edge_list_ch_38__q0 = __tapa_fsm_unit_read_A_38___edge_list_ch_38__q0;
  assign __tapa_fsm_unit_read_A_38__ap_done = read_A_38__ap_done;
  assign __tapa_fsm_unit_read_A_38__ap_idle = read_A_38__ap_idle;
  assign __tapa_fsm_unit_read_A_38__ap_ready = read_A_38__ap_ready;
  assign read_A_38__ap_start = __tapa_fsm_unit_read_A_38__ap_start;
  assign read_A_39___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_39___NUM_A_LEN__q0;
  assign read_A_39___P_N__q0 = __tapa_fsm_unit_read_A_39___P_N__q0;
  assign read_A_39___edge_list_ch_39__q0 = __tapa_fsm_unit_read_A_39___edge_list_ch_39__q0;
  assign __tapa_fsm_unit_read_A_39__ap_done = read_A_39__ap_done;
  assign __tapa_fsm_unit_read_A_39__ap_idle = read_A_39__ap_idle;
  assign __tapa_fsm_unit_read_A_39__ap_ready = read_A_39__ap_ready;
  assign read_A_39__ap_start = __tapa_fsm_unit_read_A_39__ap_start;
  assign read_A_3___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_3___NUM_A_LEN__q0;
  assign read_A_3___P_N__q0 = __tapa_fsm_unit_read_A_3___P_N__q0;
  assign read_A_3___edge_list_ch_3__q0 = __tapa_fsm_unit_read_A_3___edge_list_ch_3__q0;
  assign __tapa_fsm_unit_read_A_3__ap_done = read_A_3__ap_done;
  assign __tapa_fsm_unit_read_A_3__ap_idle = read_A_3__ap_idle;
  assign __tapa_fsm_unit_read_A_3__ap_ready = read_A_3__ap_ready;
  assign read_A_3__ap_start = __tapa_fsm_unit_read_A_3__ap_start;
  assign read_A_40___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_40___NUM_A_LEN__q0;
  assign read_A_40___P_N__q0 = __tapa_fsm_unit_read_A_40___P_N__q0;
  assign read_A_40___edge_list_ch_40__q0 = __tapa_fsm_unit_read_A_40___edge_list_ch_40__q0;
  assign __tapa_fsm_unit_read_A_40__ap_done = read_A_40__ap_done;
  assign __tapa_fsm_unit_read_A_40__ap_idle = read_A_40__ap_idle;
  assign __tapa_fsm_unit_read_A_40__ap_ready = read_A_40__ap_ready;
  assign read_A_40__ap_start = __tapa_fsm_unit_read_A_40__ap_start;
  assign read_A_41___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_41___NUM_A_LEN__q0;
  assign read_A_41___P_N__q0 = __tapa_fsm_unit_read_A_41___P_N__q0;
  assign read_A_41___edge_list_ch_41__q0 = __tapa_fsm_unit_read_A_41___edge_list_ch_41__q0;
  assign __tapa_fsm_unit_read_A_41__ap_done = read_A_41__ap_done;
  assign __tapa_fsm_unit_read_A_41__ap_idle = read_A_41__ap_idle;
  assign __tapa_fsm_unit_read_A_41__ap_ready = read_A_41__ap_ready;
  assign read_A_41__ap_start = __tapa_fsm_unit_read_A_41__ap_start;
  assign read_A_42___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_42___NUM_A_LEN__q0;
  assign read_A_42___P_N__q0 = __tapa_fsm_unit_read_A_42___P_N__q0;
  assign read_A_42___edge_list_ch_42__q0 = __tapa_fsm_unit_read_A_42___edge_list_ch_42__q0;
  assign __tapa_fsm_unit_read_A_42__ap_done = read_A_42__ap_done;
  assign __tapa_fsm_unit_read_A_42__ap_idle = read_A_42__ap_idle;
  assign __tapa_fsm_unit_read_A_42__ap_ready = read_A_42__ap_ready;
  assign read_A_42__ap_start = __tapa_fsm_unit_read_A_42__ap_start;
  assign read_A_43___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_43___NUM_A_LEN__q0;
  assign read_A_43___P_N__q0 = __tapa_fsm_unit_read_A_43___P_N__q0;
  assign read_A_43___edge_list_ch_43__q0 = __tapa_fsm_unit_read_A_43___edge_list_ch_43__q0;
  assign __tapa_fsm_unit_read_A_43__ap_done = read_A_43__ap_done;
  assign __tapa_fsm_unit_read_A_43__ap_idle = read_A_43__ap_idle;
  assign __tapa_fsm_unit_read_A_43__ap_ready = read_A_43__ap_ready;
  assign read_A_43__ap_start = __tapa_fsm_unit_read_A_43__ap_start;
  assign read_A_44___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_44___NUM_A_LEN__q0;
  assign read_A_44___P_N__q0 = __tapa_fsm_unit_read_A_44___P_N__q0;
  assign read_A_44___edge_list_ch_44__q0 = __tapa_fsm_unit_read_A_44___edge_list_ch_44__q0;
  assign __tapa_fsm_unit_read_A_44__ap_done = read_A_44__ap_done;
  assign __tapa_fsm_unit_read_A_44__ap_idle = read_A_44__ap_idle;
  assign __tapa_fsm_unit_read_A_44__ap_ready = read_A_44__ap_ready;
  assign read_A_44__ap_start = __tapa_fsm_unit_read_A_44__ap_start;
  assign read_A_45___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_45___NUM_A_LEN__q0;
  assign read_A_45___P_N__q0 = __tapa_fsm_unit_read_A_45___P_N__q0;
  assign read_A_45___edge_list_ch_45__q0 = __tapa_fsm_unit_read_A_45___edge_list_ch_45__q0;
  assign __tapa_fsm_unit_read_A_45__ap_done = read_A_45__ap_done;
  assign __tapa_fsm_unit_read_A_45__ap_idle = read_A_45__ap_idle;
  assign __tapa_fsm_unit_read_A_45__ap_ready = read_A_45__ap_ready;
  assign read_A_45__ap_start = __tapa_fsm_unit_read_A_45__ap_start;
  assign read_A_46___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_46___NUM_A_LEN__q0;
  assign read_A_46___P_N__q0 = __tapa_fsm_unit_read_A_46___P_N__q0;
  assign read_A_46___edge_list_ch_46__q0 = __tapa_fsm_unit_read_A_46___edge_list_ch_46__q0;
  assign __tapa_fsm_unit_read_A_46__ap_done = read_A_46__ap_done;
  assign __tapa_fsm_unit_read_A_46__ap_idle = read_A_46__ap_idle;
  assign __tapa_fsm_unit_read_A_46__ap_ready = read_A_46__ap_ready;
  assign read_A_46__ap_start = __tapa_fsm_unit_read_A_46__ap_start;
  assign read_A_47___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_47___NUM_A_LEN__q0;
  assign read_A_47___P_N__q0 = __tapa_fsm_unit_read_A_47___P_N__q0;
  assign read_A_47___edge_list_ch_47__q0 = __tapa_fsm_unit_read_A_47___edge_list_ch_47__q0;
  assign __tapa_fsm_unit_read_A_47__ap_done = read_A_47__ap_done;
  assign __tapa_fsm_unit_read_A_47__ap_idle = read_A_47__ap_idle;
  assign __tapa_fsm_unit_read_A_47__ap_ready = read_A_47__ap_ready;
  assign read_A_47__ap_start = __tapa_fsm_unit_read_A_47__ap_start;
  assign read_A_4___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_4___NUM_A_LEN__q0;
  assign read_A_4___P_N__q0 = __tapa_fsm_unit_read_A_4___P_N__q0;
  assign read_A_4___edge_list_ch_4__q0 = __tapa_fsm_unit_read_A_4___edge_list_ch_4__q0;
  assign __tapa_fsm_unit_read_A_4__ap_done = read_A_4__ap_done;
  assign __tapa_fsm_unit_read_A_4__ap_idle = read_A_4__ap_idle;
  assign __tapa_fsm_unit_read_A_4__ap_ready = read_A_4__ap_ready;
  assign read_A_4__ap_start = __tapa_fsm_unit_read_A_4__ap_start;
  assign read_A_5___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_5___NUM_A_LEN__q0;
  assign read_A_5___P_N__q0 = __tapa_fsm_unit_read_A_5___P_N__q0;
  assign read_A_5___edge_list_ch_5__q0 = __tapa_fsm_unit_read_A_5___edge_list_ch_5__q0;
  assign __tapa_fsm_unit_read_A_5__ap_done = read_A_5__ap_done;
  assign __tapa_fsm_unit_read_A_5__ap_idle = read_A_5__ap_idle;
  assign __tapa_fsm_unit_read_A_5__ap_ready = read_A_5__ap_ready;
  assign read_A_5__ap_start = __tapa_fsm_unit_read_A_5__ap_start;
  assign read_A_6___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_6___NUM_A_LEN__q0;
  assign read_A_6___P_N__q0 = __tapa_fsm_unit_read_A_6___P_N__q0;
  assign read_A_6___edge_list_ch_6__q0 = __tapa_fsm_unit_read_A_6___edge_list_ch_6__q0;
  assign __tapa_fsm_unit_read_A_6__ap_done = read_A_6__ap_done;
  assign __tapa_fsm_unit_read_A_6__ap_idle = read_A_6__ap_idle;
  assign __tapa_fsm_unit_read_A_6__ap_ready = read_A_6__ap_ready;
  assign read_A_6__ap_start = __tapa_fsm_unit_read_A_6__ap_start;
  assign read_A_7___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_7___NUM_A_LEN__q0;
  assign read_A_7___P_N__q0 = __tapa_fsm_unit_read_A_7___P_N__q0;
  assign read_A_7___edge_list_ch_7__q0 = __tapa_fsm_unit_read_A_7___edge_list_ch_7__q0;
  assign __tapa_fsm_unit_read_A_7__ap_done = read_A_7__ap_done;
  assign __tapa_fsm_unit_read_A_7__ap_idle = read_A_7__ap_idle;
  assign __tapa_fsm_unit_read_A_7__ap_ready = read_A_7__ap_ready;
  assign read_A_7__ap_start = __tapa_fsm_unit_read_A_7__ap_start;
  assign read_A_8___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_8___NUM_A_LEN__q0;
  assign read_A_8___P_N__q0 = __tapa_fsm_unit_read_A_8___P_N__q0;
  assign read_A_8___edge_list_ch_8__q0 = __tapa_fsm_unit_read_A_8___edge_list_ch_8__q0;
  assign __tapa_fsm_unit_read_A_8__ap_done = read_A_8__ap_done;
  assign __tapa_fsm_unit_read_A_8__ap_idle = read_A_8__ap_idle;
  assign __tapa_fsm_unit_read_A_8__ap_ready = read_A_8__ap_ready;
  assign read_A_8__ap_start = __tapa_fsm_unit_read_A_8__ap_start;
  assign read_A_9___NUM_A_LEN__q0 = __tapa_fsm_unit_read_A_9___NUM_A_LEN__q0;
  assign read_A_9___P_N__q0 = __tapa_fsm_unit_read_A_9___P_N__q0;
  assign read_A_9___edge_list_ch_9__q0 = __tapa_fsm_unit_read_A_9___edge_list_ch_9__q0;
  assign __tapa_fsm_unit_read_A_9__ap_done = read_A_9__ap_done;
  assign __tapa_fsm_unit_read_A_9__ap_idle = read_A_9__ap_idle;
  assign __tapa_fsm_unit_read_A_9__ap_ready = read_A_9__ap_ready;
  assign read_A_9__ap_start = __tapa_fsm_unit_read_A_9__ap_start;
  assign read_X_0___K__q0 = __tapa_fsm_unit_read_X_0___K__q0;
  assign read_X_0___P_N__q0 = __tapa_fsm_unit_read_X_0___P_N__q0;
  assign read_X_0___vec_X__q0 = __tapa_fsm_unit_read_X_0___vec_X__q0;
  assign __tapa_fsm_unit_read_X_0__ap_done = read_X_0__ap_done;
  assign __tapa_fsm_unit_read_X_0__ap_idle = read_X_0__ap_idle;
  assign __tapa_fsm_unit_read_X_0__ap_ready = read_X_0__ap_ready;
  assign read_X_0__ap_start = __tapa_fsm_unit_read_X_0__ap_start;
  assign read_Y_0___M__q0 = __tapa_fsm_unit_read_Y_0___M__q0;
  assign read_Y_0___P_N__q0 = __tapa_fsm_unit_read_Y_0___P_N__q0;
  assign read_Y_0___vec_Y__q0 = __tapa_fsm_unit_read_Y_0___vec_Y__q0;
  assign __tapa_fsm_unit_read_Y_0__ap_done = read_Y_0__ap_done;
  assign __tapa_fsm_unit_read_Y_0__ap_idle = read_Y_0__ap_idle;
  assign __tapa_fsm_unit_read_Y_0__ap_ready = read_Y_0__ap_ready;
  assign read_Y_0__ap_start = __tapa_fsm_unit_read_Y_0__ap_start;
  assign read_edge_list_ptr_0___K__q0 = __tapa_fsm_unit_read_edge_list_ptr_0___K__q0;
  assign read_edge_list_ptr_0___M__q0 = __tapa_fsm_unit_read_edge_list_ptr_0___M__q0;
  assign read_edge_list_ptr_0___NUM_ITE__q0 = __tapa_fsm_unit_read_edge_list_ptr_0___NUM_ITE__q0;
  assign read_edge_list_ptr_0___P_N__q0 = __tapa_fsm_unit_read_edge_list_ptr_0___P_N__q0;
  assign read_edge_list_ptr_0___edge_list_ptr__q0 = __tapa_fsm_unit_read_edge_list_ptr_0___edge_list_ptr__q0;
  assign __tapa_fsm_unit_read_edge_list_ptr_0__ap_done = read_edge_list_ptr_0__ap_done;
  assign __tapa_fsm_unit_read_edge_list_ptr_0__ap_idle = read_edge_list_ptr_0__ap_idle;
  assign __tapa_fsm_unit_read_edge_list_ptr_0__ap_ready = read_edge_list_ptr_0__ap_ready;
  assign read_edge_list_ptr_0__ap_start = __tapa_fsm_unit_read_edge_list_ptr_0__ap_start;
  assign __tapa_fsm_unit_vec_X = vec_X;
  assign __tapa_fsm_unit_vec_Y = vec_Y;
  assign __tapa_fsm_unit_vec_Y_out = vec_Y_out;
  assign write_Y_0___M__q0 = __tapa_fsm_unit_write_Y_0___M__q0;
  assign write_Y_0___P_N__q0 = __tapa_fsm_unit_write_Y_0___P_N__q0;
  assign write_Y_0___vec_Y_out__q0 = __tapa_fsm_unit_write_Y_0___vec_Y_out__q0;
  assign __tapa_fsm_unit_write_Y_0__ap_done = write_Y_0__ap_done;
  assign __tapa_fsm_unit_write_Y_0__ap_idle = write_Y_0__ap_idle;
  assign __tapa_fsm_unit_write_Y_0__ap_ready = write_Y_0__ap_ready;
  assign write_Y_0__ap_start = __tapa_fsm_unit_write_Y_0__ap_start;
endmodule