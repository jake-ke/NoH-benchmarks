`timescale 1 ns / 1 ps
module __rs___rs_ap_ctrl_start_ready_pipeline_2_aux #(
    parameter HEAD_LEVEL      = 0,
    parameter BODY_LEVEL      = 2,
    parameter TAIL_LEVEL      = 0,
    parameter __HEAD_REGION   = "",
    parameter __BODY_0_REGION = "",
    parameter __BODY_1_REGION = "",
    parameter __TAIL_REGION   = "",
    parameter GRACE_PERIOD    = ( BODY_LEVEL + HEAD_LEVEL + TAIL_LEVEL ) * 2
) (
    output wire RS_AP_PP_BODY_0_clk,
    output wire RS_AP_PP_BODY_0_reset,
    output wire RS_AP_PP_BODY_1_clk,
    output wire RS_AP_PP_BODY_1_reset,
    output wire RS_AP_PP_HEAD_clk,
    output wire RS_AP_PP_HEAD_reset,
    output wire RS_AP_PP_TAIL_GATE_clk,
    output wire RS_AP_PP_TAIL_GATE_reset,
    output wire RS_AP_PP_TAIL_clk,
    output wire RS_AP_PP_TAIL_reset,
    input wire  clk,
    input wire  reset
);
    
    wire                  body_outbound_0_valid;
    wire                  body_outbound_0_ready;
    
    wire                  body_outbound_1_valid;
    wire                  body_outbound_1_ready;
    
    wire                  body_outbound_2_valid;
    wire                  body_outbound_2_ready;
    
    wire                  tail_gate_valid;
    wire                  tail_gate_ready;
  assign RS_AP_PP_HEAD_clk = clk;
  assign RS_AP_PP_HEAD_reset = reset;
  assign RS_AP_PP_BODY_0_clk = clk;
  assign RS_AP_PP_BODY_0_reset = reset;
  assign RS_AP_PP_BODY_1_clk = clk;
  assign RS_AP_PP_BODY_1_reset = reset;
  assign RS_AP_PP_TAIL_GATE_clk = clk;
  assign RS_AP_PP_TAIL_GATE_reset = reset;
  assign RS_AP_PP_TAIL_clk = clk;
  assign RS_AP_PP_TAIL_reset = reset;
endmodule