`timescale 1 ns / 1 ps
 
(* CORE_GENERATION_INFO = "Knn_Knn,hls_ip_2023_2_2,{HLS_INPUT_TYPE=cxx,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=0,HLS_INPUT_PART=xcvh1582-vsva3697-2MP-e-S,HLS_INPUT_CLOCK=3.330000,HLS_INPUT_ARCH=others,HLS_SYN_CLOCK=1.000000,HLS_SYN_LAT=0,HLS_SYN_TPT=none,HLS_SYN_MEM=0,HLS_SYN_DSP=0,HLS_SYN_FF=2066,HLS_SYN_LUT=3752,HLS_VERSION=2023_2_2}" *)module __rs_Knn_aux #(
    parameter C_S_AXI_CONTROL_DATA_WIDTH  = 32,
    parameter C_S_AXI_CONTROL_ADDR_WIDTH  = 9,
    parameter C_S_AXI_DATA_WIDTH          = 32,
    parameter C_S_AXI_CONTROL_WSTRB_WIDTH = 4,
    parameter C_S_AXI_WSTRB_WIDTH         = 4
) (
    input wire                                           s_axi_control_AWVALID,
    output wire                                          s_axi_control_AWREADY,
    input wire  [    (C_S_AXI_CONTROL_ADDR_WIDTH - 1):0] s_axi_control_AWADDR,
    input wire                                           s_axi_control_WVALID,
    output wire                                          s_axi_control_WREADY,
    input wire  [    (C_S_AXI_CONTROL_DATA_WIDTH - 1):0] s_axi_control_WDATA,
    input wire  [   (C_S_AXI_CONTROL_WSTRB_WIDTH - 1):0] s_axi_control_WSTRB,
    input wire                                           s_axi_control_ARVALID,
    output wire                                          s_axi_control_ARREADY,
    input wire  [    (C_S_AXI_CONTROL_ADDR_WIDTH - 1):0] s_axi_control_ARADDR,
    output wire                                          s_axi_control_RVALID,
    input wire                                           s_axi_control_RREADY,
    output wire [    (C_S_AXI_CONTROL_DATA_WIDTH - 1):0] s_axi_control_RDATA,
    output wire [                                   1:0] s_axi_control_RRESP,
    output wire                                          s_axi_control_BVALID,
    input wire                                           s_axi_control_BREADY,
    output wire [                                   1:0] s_axi_control_BRESP,
    input wire                                           ap_clk,
    input wire                                           ap_rst_n,
    output wire                                          interrupt,
    output wire [                                  63:0] m_axi_L3_out_dist_ARADDR,
    output wire [                                   1:0] m_axi_L3_out_dist_ARBURST,
    output wire [                                   3:0] m_axi_L3_out_dist_ARCACHE,
    output wire [                                   0:0] m_axi_L3_out_dist_ARID,
    output wire [                                   7:0] m_axi_L3_out_dist_ARLEN,
    output wire                                          m_axi_L3_out_dist_ARLOCK,
    output wire [                                   2:0] m_axi_L3_out_dist_ARPROT,
    output wire [                                   3:0] m_axi_L3_out_dist_ARQOS,
    input wire                                           m_axi_L3_out_dist_ARREADY,
    output wire [                                   2:0] m_axi_L3_out_dist_ARSIZE,
    output wire                                          m_axi_L3_out_dist_ARVALID,
    output wire [                                  63:0] m_axi_L3_out_dist_AWADDR,
    output wire [                                   1:0] m_axi_L3_out_dist_AWBURST,
    output wire [                                   3:0] m_axi_L3_out_dist_AWCACHE,
    output wire [                                   0:0] m_axi_L3_out_dist_AWID,
    output wire [                                   7:0] m_axi_L3_out_dist_AWLEN,
    output wire                                          m_axi_L3_out_dist_AWLOCK,
    output wire [                                   2:0] m_axi_L3_out_dist_AWPROT,
    output wire [                                   3:0] m_axi_L3_out_dist_AWQOS,
    input wire                                           m_axi_L3_out_dist_AWREADY,
    output wire [                                   2:0] m_axi_L3_out_dist_AWSIZE,
    output wire                                          m_axi_L3_out_dist_AWVALID,
    input wire  [                                   0:0] m_axi_L3_out_dist_BID,
    output wire                                          m_axi_L3_out_dist_BREADY,
    input wire  [                                   1:0] m_axi_L3_out_dist_BRESP,
    input wire                                           m_axi_L3_out_dist_BVALID,
    input wire  [                                  31:0] m_axi_L3_out_dist_RDATA,
    input wire  [                                   0:0] m_axi_L3_out_dist_RID,
    input wire                                           m_axi_L3_out_dist_RLAST,
    output wire                                          m_axi_L3_out_dist_RREADY,
    input wire  [                                   1:0] m_axi_L3_out_dist_RRESP,
    input wire                                           m_axi_L3_out_dist_RVALID,
    output wire [                                  31:0] m_axi_L3_out_dist_WDATA,
    output wire                                          m_axi_L3_out_dist_WLAST,
    input wire                                           m_axi_L3_out_dist_WREADY,
    output wire [                                   3:0] m_axi_L3_out_dist_WSTRB,
    output wire                                          m_axi_L3_out_dist_WVALID,
    output wire [                                  63:0] m_axi_L3_out_id_ARADDR,
    output wire [                                   1:0] m_axi_L3_out_id_ARBURST,
    output wire [                                   3:0] m_axi_L3_out_id_ARCACHE,
    output wire [                                   0:0] m_axi_L3_out_id_ARID,
    output wire [                                   7:0] m_axi_L3_out_id_ARLEN,
    output wire                                          m_axi_L3_out_id_ARLOCK,
    output wire [                                   2:0] m_axi_L3_out_id_ARPROT,
    output wire [                                   3:0] m_axi_L3_out_id_ARQOS,
    input wire                                           m_axi_L3_out_id_ARREADY,
    output wire [                                   2:0] m_axi_L3_out_id_ARSIZE,
    output wire                                          m_axi_L3_out_id_ARVALID,
    output wire [                                  63:0] m_axi_L3_out_id_AWADDR,
    output wire [                                   1:0] m_axi_L3_out_id_AWBURST,
    output wire [                                   3:0] m_axi_L3_out_id_AWCACHE,
    output wire [                                   0:0] m_axi_L3_out_id_AWID,
    output wire [                                   7:0] m_axi_L3_out_id_AWLEN,
    output wire                                          m_axi_L3_out_id_AWLOCK,
    output wire [                                   2:0] m_axi_L3_out_id_AWPROT,
    output wire [                                   3:0] m_axi_L3_out_id_AWQOS,
    input wire                                           m_axi_L3_out_id_AWREADY,
    output wire [                                   2:0] m_axi_L3_out_id_AWSIZE,
    output wire                                          m_axi_L3_out_id_AWVALID,
    input wire  [                                   0:0] m_axi_L3_out_id_BID,
    output wire                                          m_axi_L3_out_id_BREADY,
    input wire  [                                   1:0] m_axi_L3_out_id_BRESP,
    input wire                                           m_axi_L3_out_id_BVALID,
    input wire  [                                  31:0] m_axi_L3_out_id_RDATA,
    input wire  [                                   0:0] m_axi_L3_out_id_RID,
    input wire                                           m_axi_L3_out_id_RLAST,
    output wire                                          m_axi_L3_out_id_RREADY,
    input wire  [                                   1:0] m_axi_L3_out_id_RRESP,
    input wire                                           m_axi_L3_out_id_RVALID,
    output wire [                                  31:0] m_axi_L3_out_id_WDATA,
    output wire                                          m_axi_L3_out_id_WLAST,
    input wire                                           m_axi_L3_out_id_WREADY,
    output wire [                                   3:0] m_axi_L3_out_id_WSTRB,
    output wire                                          m_axi_L3_out_id_WVALID,
    output wire [                                  63:0] m_axi_in_0_ARADDR,
    output wire [                                   1:0] m_axi_in_0_ARBURST,
    output wire [                                   3:0] m_axi_in_0_ARCACHE,
    output wire [                                   0:0] m_axi_in_0_ARID,
    output wire [                                   7:0] m_axi_in_0_ARLEN,
    output wire                                          m_axi_in_0_ARLOCK,
    output wire [                                   2:0] m_axi_in_0_ARPROT,
    output wire [                                   3:0] m_axi_in_0_ARQOS,
    input wire                                           m_axi_in_0_ARREADY,
    output wire [                                   2:0] m_axi_in_0_ARSIZE,
    output wire                                          m_axi_in_0_ARVALID,
    output wire [                                  63:0] m_axi_in_0_AWADDR,
    output wire [                                   1:0] m_axi_in_0_AWBURST,
    output wire [                                   3:0] m_axi_in_0_AWCACHE,
    output wire [                                   0:0] m_axi_in_0_AWID,
    output wire [                                   7:0] m_axi_in_0_AWLEN,
    output wire                                          m_axi_in_0_AWLOCK,
    output wire [                                   2:0] m_axi_in_0_AWPROT,
    output wire [                                   3:0] m_axi_in_0_AWQOS,
    input wire                                           m_axi_in_0_AWREADY,
    output wire [                                   2:0] m_axi_in_0_AWSIZE,
    output wire                                          m_axi_in_0_AWVALID,
    input wire  [                                   0:0] m_axi_in_0_BID,
    output wire                                          m_axi_in_0_BREADY,
    input wire  [                                   1:0] m_axi_in_0_BRESP,
    input wire                                           m_axi_in_0_BVALID,
    input wire  [                                 255:0] m_axi_in_0_RDATA,
    input wire  [                                   0:0] m_axi_in_0_RID,
    input wire                                           m_axi_in_0_RLAST,
    output wire                                          m_axi_in_0_RREADY,
    input wire  [                                   1:0] m_axi_in_0_RRESP,
    input wire                                           m_axi_in_0_RVALID,
    output wire [                                 255:0] m_axi_in_0_WDATA,
    output wire                                          m_axi_in_0_WLAST,
    input wire                                           m_axi_in_0_WREADY,
    output wire [                                  31:0] m_axi_in_0_WSTRB,
    output wire                                          m_axi_in_0_WVALID,
    output wire [                                  63:0] m_axi_in_1_ARADDR,
    output wire [                                   1:0] m_axi_in_1_ARBURST,
    output wire [                                   3:0] m_axi_in_1_ARCACHE,
    output wire [                                   0:0] m_axi_in_1_ARID,
    output wire [                                   7:0] m_axi_in_1_ARLEN,
    output wire                                          m_axi_in_1_ARLOCK,
    output wire [                                   2:0] m_axi_in_1_ARPROT,
    output wire [                                   3:0] m_axi_in_1_ARQOS,
    input wire                                           m_axi_in_1_ARREADY,
    output wire [                                   2:0] m_axi_in_1_ARSIZE,
    output wire                                          m_axi_in_1_ARVALID,
    output wire [                                  63:0] m_axi_in_1_AWADDR,
    output wire [                                   1:0] m_axi_in_1_AWBURST,
    output wire [                                   3:0] m_axi_in_1_AWCACHE,
    output wire [                                   0:0] m_axi_in_1_AWID,
    output wire [                                   7:0] m_axi_in_1_AWLEN,
    output wire                                          m_axi_in_1_AWLOCK,
    output wire [                                   2:0] m_axi_in_1_AWPROT,
    output wire [                                   3:0] m_axi_in_1_AWQOS,
    input wire                                           m_axi_in_1_AWREADY,
    output wire [                                   2:0] m_axi_in_1_AWSIZE,
    output wire                                          m_axi_in_1_AWVALID,
    input wire  [                                   0:0] m_axi_in_1_BID,
    output wire                                          m_axi_in_1_BREADY,
    input wire  [                                   1:0] m_axi_in_1_BRESP,
    input wire                                           m_axi_in_1_BVALID,
    input wire  [                                 255:0] m_axi_in_1_RDATA,
    input wire  [                                   0:0] m_axi_in_1_RID,
    input wire                                           m_axi_in_1_RLAST,
    output wire                                          m_axi_in_1_RREADY,
    input wire  [                                   1:0] m_axi_in_1_RRESP,
    input wire                                           m_axi_in_1_RVALID,
    output wire [                                 255:0] m_axi_in_1_WDATA,
    output wire                                          m_axi_in_1_WLAST,
    input wire                                           m_axi_in_1_WREADY,
    output wire [                                  31:0] m_axi_in_1_WSTRB,
    output wire                                          m_axi_in_1_WVALID,
    output wire [                                  63:0] m_axi_in_10_ARADDR,
    output wire [                                   1:0] m_axi_in_10_ARBURST,
    output wire [                                   3:0] m_axi_in_10_ARCACHE,
    output wire [                                   0:0] m_axi_in_10_ARID,
    output wire [                                   7:0] m_axi_in_10_ARLEN,
    output wire                                          m_axi_in_10_ARLOCK,
    output wire [                                   2:0] m_axi_in_10_ARPROT,
    output wire [                                   3:0] m_axi_in_10_ARQOS,
    input wire                                           m_axi_in_10_ARREADY,
    output wire [                                   2:0] m_axi_in_10_ARSIZE,
    output wire                                          m_axi_in_10_ARVALID,
    output wire [                                  63:0] m_axi_in_10_AWADDR,
    output wire [                                   1:0] m_axi_in_10_AWBURST,
    output wire [                                   3:0] m_axi_in_10_AWCACHE,
    output wire [                                   0:0] m_axi_in_10_AWID,
    output wire [                                   7:0] m_axi_in_10_AWLEN,
    output wire                                          m_axi_in_10_AWLOCK,
    output wire [                                   2:0] m_axi_in_10_AWPROT,
    output wire [                                   3:0] m_axi_in_10_AWQOS,
    input wire                                           m_axi_in_10_AWREADY,
    output wire [                                   2:0] m_axi_in_10_AWSIZE,
    output wire                                          m_axi_in_10_AWVALID,
    input wire  [                                   0:0] m_axi_in_10_BID,
    output wire                                          m_axi_in_10_BREADY,
    input wire  [                                   1:0] m_axi_in_10_BRESP,
    input wire                                           m_axi_in_10_BVALID,
    input wire  [                                 255:0] m_axi_in_10_RDATA,
    input wire  [                                   0:0] m_axi_in_10_RID,
    input wire                                           m_axi_in_10_RLAST,
    output wire                                          m_axi_in_10_RREADY,
    input wire  [                                   1:0] m_axi_in_10_RRESP,
    input wire                                           m_axi_in_10_RVALID,
    output wire [                                 255:0] m_axi_in_10_WDATA,
    output wire                                          m_axi_in_10_WLAST,
    input wire                                           m_axi_in_10_WREADY,
    output wire [                                  31:0] m_axi_in_10_WSTRB,
    output wire                                          m_axi_in_10_WVALID,
    output wire [                                  63:0] m_axi_in_11_ARADDR,
    output wire [                                   1:0] m_axi_in_11_ARBURST,
    output wire [                                   3:0] m_axi_in_11_ARCACHE,
    output wire [                                   0:0] m_axi_in_11_ARID,
    output wire [                                   7:0] m_axi_in_11_ARLEN,
    output wire                                          m_axi_in_11_ARLOCK,
    output wire [                                   2:0] m_axi_in_11_ARPROT,
    output wire [                                   3:0] m_axi_in_11_ARQOS,
    input wire                                           m_axi_in_11_ARREADY,
    output wire [                                   2:0] m_axi_in_11_ARSIZE,
    output wire                                          m_axi_in_11_ARVALID,
    output wire [                                  63:0] m_axi_in_11_AWADDR,
    output wire [                                   1:0] m_axi_in_11_AWBURST,
    output wire [                                   3:0] m_axi_in_11_AWCACHE,
    output wire [                                   0:0] m_axi_in_11_AWID,
    output wire [                                   7:0] m_axi_in_11_AWLEN,
    output wire                                          m_axi_in_11_AWLOCK,
    output wire [                                   2:0] m_axi_in_11_AWPROT,
    output wire [                                   3:0] m_axi_in_11_AWQOS,
    input wire                                           m_axi_in_11_AWREADY,
    output wire [                                   2:0] m_axi_in_11_AWSIZE,
    output wire                                          m_axi_in_11_AWVALID,
    input wire  [                                   0:0] m_axi_in_11_BID,
    output wire                                          m_axi_in_11_BREADY,
    input wire  [                                   1:0] m_axi_in_11_BRESP,
    input wire                                           m_axi_in_11_BVALID,
    input wire  [                                 255:0] m_axi_in_11_RDATA,
    input wire  [                                   0:0] m_axi_in_11_RID,
    input wire                                           m_axi_in_11_RLAST,
    output wire                                          m_axi_in_11_RREADY,
    input wire  [                                   1:0] m_axi_in_11_RRESP,
    input wire                                           m_axi_in_11_RVALID,
    output wire [                                 255:0] m_axi_in_11_WDATA,
    output wire                                          m_axi_in_11_WLAST,
    input wire                                           m_axi_in_11_WREADY,
    output wire [                                  31:0] m_axi_in_11_WSTRB,
    output wire                                          m_axi_in_11_WVALID,
    output wire [                                  63:0] m_axi_in_12_ARADDR,
    output wire [                                   1:0] m_axi_in_12_ARBURST,
    output wire [                                   3:0] m_axi_in_12_ARCACHE,
    output wire [                                   0:0] m_axi_in_12_ARID,
    output wire [                                   7:0] m_axi_in_12_ARLEN,
    output wire                                          m_axi_in_12_ARLOCK,
    output wire [                                   2:0] m_axi_in_12_ARPROT,
    output wire [                                   3:0] m_axi_in_12_ARQOS,
    input wire                                           m_axi_in_12_ARREADY,
    output wire [                                   2:0] m_axi_in_12_ARSIZE,
    output wire                                          m_axi_in_12_ARVALID,
    output wire [                                  63:0] m_axi_in_12_AWADDR,
    output wire [                                   1:0] m_axi_in_12_AWBURST,
    output wire [                                   3:0] m_axi_in_12_AWCACHE,
    output wire [                                   0:0] m_axi_in_12_AWID,
    output wire [                                   7:0] m_axi_in_12_AWLEN,
    output wire                                          m_axi_in_12_AWLOCK,
    output wire [                                   2:0] m_axi_in_12_AWPROT,
    output wire [                                   3:0] m_axi_in_12_AWQOS,
    input wire                                           m_axi_in_12_AWREADY,
    output wire [                                   2:0] m_axi_in_12_AWSIZE,
    output wire                                          m_axi_in_12_AWVALID,
    input wire  [                                   0:0] m_axi_in_12_BID,
    output wire                                          m_axi_in_12_BREADY,
    input wire  [                                   1:0] m_axi_in_12_BRESP,
    input wire                                           m_axi_in_12_BVALID,
    input wire  [                                 255:0] m_axi_in_12_RDATA,
    input wire  [                                   0:0] m_axi_in_12_RID,
    input wire                                           m_axi_in_12_RLAST,
    output wire                                          m_axi_in_12_RREADY,
    input wire  [                                   1:0] m_axi_in_12_RRESP,
    input wire                                           m_axi_in_12_RVALID,
    output wire [                                 255:0] m_axi_in_12_WDATA,
    output wire                                          m_axi_in_12_WLAST,
    input wire                                           m_axi_in_12_WREADY,
    output wire [                                  31:0] m_axi_in_12_WSTRB,
    output wire                                          m_axi_in_12_WVALID,
    output wire [                                  63:0] m_axi_in_13_ARADDR,
    output wire [                                   1:0] m_axi_in_13_ARBURST,
    output wire [                                   3:0] m_axi_in_13_ARCACHE,
    output wire [                                   0:0] m_axi_in_13_ARID,
    output wire [                                   7:0] m_axi_in_13_ARLEN,
    output wire                                          m_axi_in_13_ARLOCK,
    output wire [                                   2:0] m_axi_in_13_ARPROT,
    output wire [                                   3:0] m_axi_in_13_ARQOS,
    input wire                                           m_axi_in_13_ARREADY,
    output wire [                                   2:0] m_axi_in_13_ARSIZE,
    output wire                                          m_axi_in_13_ARVALID,
    output wire [                                  63:0] m_axi_in_13_AWADDR,
    output wire [                                   1:0] m_axi_in_13_AWBURST,
    output wire [                                   3:0] m_axi_in_13_AWCACHE,
    output wire [                                   0:0] m_axi_in_13_AWID,
    output wire [                                   7:0] m_axi_in_13_AWLEN,
    output wire                                          m_axi_in_13_AWLOCK,
    output wire [                                   2:0] m_axi_in_13_AWPROT,
    output wire [                                   3:0] m_axi_in_13_AWQOS,
    input wire                                           m_axi_in_13_AWREADY,
    output wire [                                   2:0] m_axi_in_13_AWSIZE,
    output wire                                          m_axi_in_13_AWVALID,
    input wire  [                                   0:0] m_axi_in_13_BID,
    output wire                                          m_axi_in_13_BREADY,
    input wire  [                                   1:0] m_axi_in_13_BRESP,
    input wire                                           m_axi_in_13_BVALID,
    input wire  [                                 255:0] m_axi_in_13_RDATA,
    input wire  [                                   0:0] m_axi_in_13_RID,
    input wire                                           m_axi_in_13_RLAST,
    output wire                                          m_axi_in_13_RREADY,
    input wire  [                                   1:0] m_axi_in_13_RRESP,
    input wire                                           m_axi_in_13_RVALID,
    output wire [                                 255:0] m_axi_in_13_WDATA,
    output wire                                          m_axi_in_13_WLAST,
    input wire                                           m_axi_in_13_WREADY,
    output wire [                                  31:0] m_axi_in_13_WSTRB,
    output wire                                          m_axi_in_13_WVALID,
    output wire [                                  63:0] m_axi_in_14_ARADDR,
    output wire [                                   1:0] m_axi_in_14_ARBURST,
    output wire [                                   3:0] m_axi_in_14_ARCACHE,
    output wire [                                   0:0] m_axi_in_14_ARID,
    output wire [                                   7:0] m_axi_in_14_ARLEN,
    output wire                                          m_axi_in_14_ARLOCK,
    output wire [                                   2:0] m_axi_in_14_ARPROT,
    output wire [                                   3:0] m_axi_in_14_ARQOS,
    input wire                                           m_axi_in_14_ARREADY,
    output wire [                                   2:0] m_axi_in_14_ARSIZE,
    output wire                                          m_axi_in_14_ARVALID,
    output wire [                                  63:0] m_axi_in_14_AWADDR,
    output wire [                                   1:0] m_axi_in_14_AWBURST,
    output wire [                                   3:0] m_axi_in_14_AWCACHE,
    output wire [                                   0:0] m_axi_in_14_AWID,
    output wire [                                   7:0] m_axi_in_14_AWLEN,
    output wire                                          m_axi_in_14_AWLOCK,
    output wire [                                   2:0] m_axi_in_14_AWPROT,
    output wire [                                   3:0] m_axi_in_14_AWQOS,
    input wire                                           m_axi_in_14_AWREADY,
    output wire [                                   2:0] m_axi_in_14_AWSIZE,
    output wire                                          m_axi_in_14_AWVALID,
    input wire  [                                   0:0] m_axi_in_14_BID,
    output wire                                          m_axi_in_14_BREADY,
    input wire  [                                   1:0] m_axi_in_14_BRESP,
    input wire                                           m_axi_in_14_BVALID,
    input wire  [                                 255:0] m_axi_in_14_RDATA,
    input wire  [                                   0:0] m_axi_in_14_RID,
    input wire                                           m_axi_in_14_RLAST,
    output wire                                          m_axi_in_14_RREADY,
    input wire  [                                   1:0] m_axi_in_14_RRESP,
    input wire                                           m_axi_in_14_RVALID,
    output wire [                                 255:0] m_axi_in_14_WDATA,
    output wire                                          m_axi_in_14_WLAST,
    input wire                                           m_axi_in_14_WREADY,
    output wire [                                  31:0] m_axi_in_14_WSTRB,
    output wire                                          m_axi_in_14_WVALID,
    output wire [                                  63:0] m_axi_in_15_ARADDR,
    output wire [                                   1:0] m_axi_in_15_ARBURST,
    output wire [                                   3:0] m_axi_in_15_ARCACHE,
    output wire [                                   0:0] m_axi_in_15_ARID,
    output wire [                                   7:0] m_axi_in_15_ARLEN,
    output wire                                          m_axi_in_15_ARLOCK,
    output wire [                                   2:0] m_axi_in_15_ARPROT,
    output wire [                                   3:0] m_axi_in_15_ARQOS,
    input wire                                           m_axi_in_15_ARREADY,
    output wire [                                   2:0] m_axi_in_15_ARSIZE,
    output wire                                          m_axi_in_15_ARVALID,
    output wire [                                  63:0] m_axi_in_15_AWADDR,
    output wire [                                   1:0] m_axi_in_15_AWBURST,
    output wire [                                   3:0] m_axi_in_15_AWCACHE,
    output wire [                                   0:0] m_axi_in_15_AWID,
    output wire [                                   7:0] m_axi_in_15_AWLEN,
    output wire                                          m_axi_in_15_AWLOCK,
    output wire [                                   2:0] m_axi_in_15_AWPROT,
    output wire [                                   3:0] m_axi_in_15_AWQOS,
    input wire                                           m_axi_in_15_AWREADY,
    output wire [                                   2:0] m_axi_in_15_AWSIZE,
    output wire                                          m_axi_in_15_AWVALID,
    input wire  [                                   0:0] m_axi_in_15_BID,
    output wire                                          m_axi_in_15_BREADY,
    input wire  [                                   1:0] m_axi_in_15_BRESP,
    input wire                                           m_axi_in_15_BVALID,
    input wire  [                                 255:0] m_axi_in_15_RDATA,
    input wire  [                                   0:0] m_axi_in_15_RID,
    input wire                                           m_axi_in_15_RLAST,
    output wire                                          m_axi_in_15_RREADY,
    input wire  [                                   1:0] m_axi_in_15_RRESP,
    input wire                                           m_axi_in_15_RVALID,
    output wire [                                 255:0] m_axi_in_15_WDATA,
    output wire                                          m_axi_in_15_WLAST,
    input wire                                           m_axi_in_15_WREADY,
    output wire [                                  31:0] m_axi_in_15_WSTRB,
    output wire                                          m_axi_in_15_WVALID,
    output wire [                                  63:0] m_axi_in_16_ARADDR,
    output wire [                                   1:0] m_axi_in_16_ARBURST,
    output wire [                                   3:0] m_axi_in_16_ARCACHE,
    output wire [                                   0:0] m_axi_in_16_ARID,
    output wire [                                   7:0] m_axi_in_16_ARLEN,
    output wire                                          m_axi_in_16_ARLOCK,
    output wire [                                   2:0] m_axi_in_16_ARPROT,
    output wire [                                   3:0] m_axi_in_16_ARQOS,
    input wire                                           m_axi_in_16_ARREADY,
    output wire [                                   2:0] m_axi_in_16_ARSIZE,
    output wire                                          m_axi_in_16_ARVALID,
    output wire [                                  63:0] m_axi_in_16_AWADDR,
    output wire [                                   1:0] m_axi_in_16_AWBURST,
    output wire [                                   3:0] m_axi_in_16_AWCACHE,
    output wire [                                   0:0] m_axi_in_16_AWID,
    output wire [                                   7:0] m_axi_in_16_AWLEN,
    output wire                                          m_axi_in_16_AWLOCK,
    output wire [                                   2:0] m_axi_in_16_AWPROT,
    output wire [                                   3:0] m_axi_in_16_AWQOS,
    input wire                                           m_axi_in_16_AWREADY,
    output wire [                                   2:0] m_axi_in_16_AWSIZE,
    output wire                                          m_axi_in_16_AWVALID,
    input wire  [                                   0:0] m_axi_in_16_BID,
    output wire                                          m_axi_in_16_BREADY,
    input wire  [                                   1:0] m_axi_in_16_BRESP,
    input wire                                           m_axi_in_16_BVALID,
    input wire  [                                 255:0] m_axi_in_16_RDATA,
    input wire  [                                   0:0] m_axi_in_16_RID,
    input wire                                           m_axi_in_16_RLAST,
    output wire                                          m_axi_in_16_RREADY,
    input wire  [                                   1:0] m_axi_in_16_RRESP,
    input wire                                           m_axi_in_16_RVALID,
    output wire [                                 255:0] m_axi_in_16_WDATA,
    output wire                                          m_axi_in_16_WLAST,
    input wire                                           m_axi_in_16_WREADY,
    output wire [                                  31:0] m_axi_in_16_WSTRB,
    output wire                                          m_axi_in_16_WVALID,
    output wire [                                  63:0] m_axi_in_17_ARADDR,
    output wire [                                   1:0] m_axi_in_17_ARBURST,
    output wire [                                   3:0] m_axi_in_17_ARCACHE,
    output wire [                                   0:0] m_axi_in_17_ARID,
    output wire [                                   7:0] m_axi_in_17_ARLEN,
    output wire                                          m_axi_in_17_ARLOCK,
    output wire [                                   2:0] m_axi_in_17_ARPROT,
    output wire [                                   3:0] m_axi_in_17_ARQOS,
    input wire                                           m_axi_in_17_ARREADY,
    output wire [                                   2:0] m_axi_in_17_ARSIZE,
    output wire                                          m_axi_in_17_ARVALID,
    output wire [                                  63:0] m_axi_in_17_AWADDR,
    output wire [                                   1:0] m_axi_in_17_AWBURST,
    output wire [                                   3:0] m_axi_in_17_AWCACHE,
    output wire [                                   0:0] m_axi_in_17_AWID,
    output wire [                                   7:0] m_axi_in_17_AWLEN,
    output wire                                          m_axi_in_17_AWLOCK,
    output wire [                                   2:0] m_axi_in_17_AWPROT,
    output wire [                                   3:0] m_axi_in_17_AWQOS,
    input wire                                           m_axi_in_17_AWREADY,
    output wire [                                   2:0] m_axi_in_17_AWSIZE,
    output wire                                          m_axi_in_17_AWVALID,
    input wire  [                                   0:0] m_axi_in_17_BID,
    output wire                                          m_axi_in_17_BREADY,
    input wire  [                                   1:0] m_axi_in_17_BRESP,
    input wire                                           m_axi_in_17_BVALID,
    input wire  [                                 255:0] m_axi_in_17_RDATA,
    input wire  [                                   0:0] m_axi_in_17_RID,
    input wire                                           m_axi_in_17_RLAST,
    output wire                                          m_axi_in_17_RREADY,
    input wire  [                                   1:0] m_axi_in_17_RRESP,
    input wire                                           m_axi_in_17_RVALID,
    output wire [                                 255:0] m_axi_in_17_WDATA,
    output wire                                          m_axi_in_17_WLAST,
    input wire                                           m_axi_in_17_WREADY,
    output wire [                                  31:0] m_axi_in_17_WSTRB,
    output wire                                          m_axi_in_17_WVALID,
    output wire [                                  63:0] m_axi_in_18_ARADDR,
    output wire [                                   1:0] m_axi_in_18_ARBURST,
    output wire [                                   3:0] m_axi_in_18_ARCACHE,
    output wire [                                   0:0] m_axi_in_18_ARID,
    output wire [                                   7:0] m_axi_in_18_ARLEN,
    output wire                                          m_axi_in_18_ARLOCK,
    output wire [                                   2:0] m_axi_in_18_ARPROT,
    output wire [                                   3:0] m_axi_in_18_ARQOS,
    input wire                                           m_axi_in_18_ARREADY,
    output wire [                                   2:0] m_axi_in_18_ARSIZE,
    output wire                                          m_axi_in_18_ARVALID,
    output wire [                                  63:0] m_axi_in_18_AWADDR,
    output wire [                                   1:0] m_axi_in_18_AWBURST,
    output wire [                                   3:0] m_axi_in_18_AWCACHE,
    output wire [                                   0:0] m_axi_in_18_AWID,
    output wire [                                   7:0] m_axi_in_18_AWLEN,
    output wire                                          m_axi_in_18_AWLOCK,
    output wire [                                   2:0] m_axi_in_18_AWPROT,
    output wire [                                   3:0] m_axi_in_18_AWQOS,
    input wire                                           m_axi_in_18_AWREADY,
    output wire [                                   2:0] m_axi_in_18_AWSIZE,
    output wire                                          m_axi_in_18_AWVALID,
    input wire  [                                   0:0] m_axi_in_18_BID,
    output wire                                          m_axi_in_18_BREADY,
    input wire  [                                   1:0] m_axi_in_18_BRESP,
    input wire                                           m_axi_in_18_BVALID,
    input wire  [                                 255:0] m_axi_in_18_RDATA,
    input wire  [                                   0:0] m_axi_in_18_RID,
    input wire                                           m_axi_in_18_RLAST,
    output wire                                          m_axi_in_18_RREADY,
    input wire  [                                   1:0] m_axi_in_18_RRESP,
    input wire                                           m_axi_in_18_RVALID,
    output wire [                                 255:0] m_axi_in_18_WDATA,
    output wire                                          m_axi_in_18_WLAST,
    input wire                                           m_axi_in_18_WREADY,
    output wire [                                  31:0] m_axi_in_18_WSTRB,
    output wire                                          m_axi_in_18_WVALID,
    output wire [                                  63:0] m_axi_in_19_ARADDR,
    output wire [                                   1:0] m_axi_in_19_ARBURST,
    output wire [                                   3:0] m_axi_in_19_ARCACHE,
    output wire [                                   0:0] m_axi_in_19_ARID,
    output wire [                                   7:0] m_axi_in_19_ARLEN,
    output wire                                          m_axi_in_19_ARLOCK,
    output wire [                                   2:0] m_axi_in_19_ARPROT,
    output wire [                                   3:0] m_axi_in_19_ARQOS,
    input wire                                           m_axi_in_19_ARREADY,
    output wire [                                   2:0] m_axi_in_19_ARSIZE,
    output wire                                          m_axi_in_19_ARVALID,
    output wire [                                  63:0] m_axi_in_19_AWADDR,
    output wire [                                   1:0] m_axi_in_19_AWBURST,
    output wire [                                   3:0] m_axi_in_19_AWCACHE,
    output wire [                                   0:0] m_axi_in_19_AWID,
    output wire [                                   7:0] m_axi_in_19_AWLEN,
    output wire                                          m_axi_in_19_AWLOCK,
    output wire [                                   2:0] m_axi_in_19_AWPROT,
    output wire [                                   3:0] m_axi_in_19_AWQOS,
    input wire                                           m_axi_in_19_AWREADY,
    output wire [                                   2:0] m_axi_in_19_AWSIZE,
    output wire                                          m_axi_in_19_AWVALID,
    input wire  [                                   0:0] m_axi_in_19_BID,
    output wire                                          m_axi_in_19_BREADY,
    input wire  [                                   1:0] m_axi_in_19_BRESP,
    input wire                                           m_axi_in_19_BVALID,
    input wire  [                                 255:0] m_axi_in_19_RDATA,
    input wire  [                                   0:0] m_axi_in_19_RID,
    input wire                                           m_axi_in_19_RLAST,
    output wire                                          m_axi_in_19_RREADY,
    input wire  [                                   1:0] m_axi_in_19_RRESP,
    input wire                                           m_axi_in_19_RVALID,
    output wire [                                 255:0] m_axi_in_19_WDATA,
    output wire                                          m_axi_in_19_WLAST,
    input wire                                           m_axi_in_19_WREADY,
    output wire [                                  31:0] m_axi_in_19_WSTRB,
    output wire                                          m_axi_in_19_WVALID,
    output wire [                                  63:0] m_axi_in_2_ARADDR,
    output wire [                                   1:0] m_axi_in_2_ARBURST,
    output wire [                                   3:0] m_axi_in_2_ARCACHE,
    output wire [                                   0:0] m_axi_in_2_ARID,
    output wire [                                   7:0] m_axi_in_2_ARLEN,
    output wire                                          m_axi_in_2_ARLOCK,
    output wire [                                   2:0] m_axi_in_2_ARPROT,
    output wire [                                   3:0] m_axi_in_2_ARQOS,
    input wire                                           m_axi_in_2_ARREADY,
    output wire [                                   2:0] m_axi_in_2_ARSIZE,
    output wire                                          m_axi_in_2_ARVALID,
    output wire [                                  63:0] m_axi_in_2_AWADDR,
    output wire [                                   1:0] m_axi_in_2_AWBURST,
    output wire [                                   3:0] m_axi_in_2_AWCACHE,
    output wire [                                   0:0] m_axi_in_2_AWID,
    output wire [                                   7:0] m_axi_in_2_AWLEN,
    output wire                                          m_axi_in_2_AWLOCK,
    output wire [                                   2:0] m_axi_in_2_AWPROT,
    output wire [                                   3:0] m_axi_in_2_AWQOS,
    input wire                                           m_axi_in_2_AWREADY,
    output wire [                                   2:0] m_axi_in_2_AWSIZE,
    output wire                                          m_axi_in_2_AWVALID,
    input wire  [                                   0:0] m_axi_in_2_BID,
    output wire                                          m_axi_in_2_BREADY,
    input wire  [                                   1:0] m_axi_in_2_BRESP,
    input wire                                           m_axi_in_2_BVALID,
    input wire  [                                 255:0] m_axi_in_2_RDATA,
    input wire  [                                   0:0] m_axi_in_2_RID,
    input wire                                           m_axi_in_2_RLAST,
    output wire                                          m_axi_in_2_RREADY,
    input wire  [                                   1:0] m_axi_in_2_RRESP,
    input wire                                           m_axi_in_2_RVALID,
    output wire [                                 255:0] m_axi_in_2_WDATA,
    output wire                                          m_axi_in_2_WLAST,
    input wire                                           m_axi_in_2_WREADY,
    output wire [                                  31:0] m_axi_in_2_WSTRB,
    output wire                                          m_axi_in_2_WVALID,
    output wire [                                  63:0] m_axi_in_20_ARADDR,
    output wire [                                   1:0] m_axi_in_20_ARBURST,
    output wire [                                   3:0] m_axi_in_20_ARCACHE,
    output wire [                                   0:0] m_axi_in_20_ARID,
    output wire [                                   7:0] m_axi_in_20_ARLEN,
    output wire                                          m_axi_in_20_ARLOCK,
    output wire [                                   2:0] m_axi_in_20_ARPROT,
    output wire [                                   3:0] m_axi_in_20_ARQOS,
    input wire                                           m_axi_in_20_ARREADY,
    output wire [                                   2:0] m_axi_in_20_ARSIZE,
    output wire                                          m_axi_in_20_ARVALID,
    output wire [                                  63:0] m_axi_in_20_AWADDR,
    output wire [                                   1:0] m_axi_in_20_AWBURST,
    output wire [                                   3:0] m_axi_in_20_AWCACHE,
    output wire [                                   0:0] m_axi_in_20_AWID,
    output wire [                                   7:0] m_axi_in_20_AWLEN,
    output wire                                          m_axi_in_20_AWLOCK,
    output wire [                                   2:0] m_axi_in_20_AWPROT,
    output wire [                                   3:0] m_axi_in_20_AWQOS,
    input wire                                           m_axi_in_20_AWREADY,
    output wire [                                   2:0] m_axi_in_20_AWSIZE,
    output wire                                          m_axi_in_20_AWVALID,
    input wire  [                                   0:0] m_axi_in_20_BID,
    output wire                                          m_axi_in_20_BREADY,
    input wire  [                                   1:0] m_axi_in_20_BRESP,
    input wire                                           m_axi_in_20_BVALID,
    input wire  [                                 255:0] m_axi_in_20_RDATA,
    input wire  [                                   0:0] m_axi_in_20_RID,
    input wire                                           m_axi_in_20_RLAST,
    output wire                                          m_axi_in_20_RREADY,
    input wire  [                                   1:0] m_axi_in_20_RRESP,
    input wire                                           m_axi_in_20_RVALID,
    output wire [                                 255:0] m_axi_in_20_WDATA,
    output wire                                          m_axi_in_20_WLAST,
    input wire                                           m_axi_in_20_WREADY,
    output wire [                                  31:0] m_axi_in_20_WSTRB,
    output wire                                          m_axi_in_20_WVALID,
    output wire [                                  63:0] m_axi_in_21_ARADDR,
    output wire [                                   1:0] m_axi_in_21_ARBURST,
    output wire [                                   3:0] m_axi_in_21_ARCACHE,
    output wire [                                   0:0] m_axi_in_21_ARID,
    output wire [                                   7:0] m_axi_in_21_ARLEN,
    output wire                                          m_axi_in_21_ARLOCK,
    output wire [                                   2:0] m_axi_in_21_ARPROT,
    output wire [                                   3:0] m_axi_in_21_ARQOS,
    input wire                                           m_axi_in_21_ARREADY,
    output wire [                                   2:0] m_axi_in_21_ARSIZE,
    output wire                                          m_axi_in_21_ARVALID,
    output wire [                                  63:0] m_axi_in_21_AWADDR,
    output wire [                                   1:0] m_axi_in_21_AWBURST,
    output wire [                                   3:0] m_axi_in_21_AWCACHE,
    output wire [                                   0:0] m_axi_in_21_AWID,
    output wire [                                   7:0] m_axi_in_21_AWLEN,
    output wire                                          m_axi_in_21_AWLOCK,
    output wire [                                   2:0] m_axi_in_21_AWPROT,
    output wire [                                   3:0] m_axi_in_21_AWQOS,
    input wire                                           m_axi_in_21_AWREADY,
    output wire [                                   2:0] m_axi_in_21_AWSIZE,
    output wire                                          m_axi_in_21_AWVALID,
    input wire  [                                   0:0] m_axi_in_21_BID,
    output wire                                          m_axi_in_21_BREADY,
    input wire  [                                   1:0] m_axi_in_21_BRESP,
    input wire                                           m_axi_in_21_BVALID,
    input wire  [                                 255:0] m_axi_in_21_RDATA,
    input wire  [                                   0:0] m_axi_in_21_RID,
    input wire                                           m_axi_in_21_RLAST,
    output wire                                          m_axi_in_21_RREADY,
    input wire  [                                   1:0] m_axi_in_21_RRESP,
    input wire                                           m_axi_in_21_RVALID,
    output wire [                                 255:0] m_axi_in_21_WDATA,
    output wire                                          m_axi_in_21_WLAST,
    input wire                                           m_axi_in_21_WREADY,
    output wire [                                  31:0] m_axi_in_21_WSTRB,
    output wire                                          m_axi_in_21_WVALID,
    output wire [                                  63:0] m_axi_in_22_ARADDR,
    output wire [                                   1:0] m_axi_in_22_ARBURST,
    output wire [                                   3:0] m_axi_in_22_ARCACHE,
    output wire [                                   0:0] m_axi_in_22_ARID,
    output wire [                                   7:0] m_axi_in_22_ARLEN,
    output wire                                          m_axi_in_22_ARLOCK,
    output wire [                                   2:0] m_axi_in_22_ARPROT,
    output wire [                                   3:0] m_axi_in_22_ARQOS,
    input wire                                           m_axi_in_22_ARREADY,
    output wire [                                   2:0] m_axi_in_22_ARSIZE,
    output wire                                          m_axi_in_22_ARVALID,
    output wire [                                  63:0] m_axi_in_22_AWADDR,
    output wire [                                   1:0] m_axi_in_22_AWBURST,
    output wire [                                   3:0] m_axi_in_22_AWCACHE,
    output wire [                                   0:0] m_axi_in_22_AWID,
    output wire [                                   7:0] m_axi_in_22_AWLEN,
    output wire                                          m_axi_in_22_AWLOCK,
    output wire [                                   2:0] m_axi_in_22_AWPROT,
    output wire [                                   3:0] m_axi_in_22_AWQOS,
    input wire                                           m_axi_in_22_AWREADY,
    output wire [                                   2:0] m_axi_in_22_AWSIZE,
    output wire                                          m_axi_in_22_AWVALID,
    input wire  [                                   0:0] m_axi_in_22_BID,
    output wire                                          m_axi_in_22_BREADY,
    input wire  [                                   1:0] m_axi_in_22_BRESP,
    input wire                                           m_axi_in_22_BVALID,
    input wire  [                                 255:0] m_axi_in_22_RDATA,
    input wire  [                                   0:0] m_axi_in_22_RID,
    input wire                                           m_axi_in_22_RLAST,
    output wire                                          m_axi_in_22_RREADY,
    input wire  [                                   1:0] m_axi_in_22_RRESP,
    input wire                                           m_axi_in_22_RVALID,
    output wire [                                 255:0] m_axi_in_22_WDATA,
    output wire                                          m_axi_in_22_WLAST,
    input wire                                           m_axi_in_22_WREADY,
    output wire [                                  31:0] m_axi_in_22_WSTRB,
    output wire                                          m_axi_in_22_WVALID,
    output wire [                                  63:0] m_axi_in_23_ARADDR,
    output wire [                                   1:0] m_axi_in_23_ARBURST,
    output wire [                                   3:0] m_axi_in_23_ARCACHE,
    output wire [                                   0:0] m_axi_in_23_ARID,
    output wire [                                   7:0] m_axi_in_23_ARLEN,
    output wire                                          m_axi_in_23_ARLOCK,
    output wire [                                   2:0] m_axi_in_23_ARPROT,
    output wire [                                   3:0] m_axi_in_23_ARQOS,
    input wire                                           m_axi_in_23_ARREADY,
    output wire [                                   2:0] m_axi_in_23_ARSIZE,
    output wire                                          m_axi_in_23_ARVALID,
    output wire [                                  63:0] m_axi_in_23_AWADDR,
    output wire [                                   1:0] m_axi_in_23_AWBURST,
    output wire [                                   3:0] m_axi_in_23_AWCACHE,
    output wire [                                   0:0] m_axi_in_23_AWID,
    output wire [                                   7:0] m_axi_in_23_AWLEN,
    output wire                                          m_axi_in_23_AWLOCK,
    output wire [                                   2:0] m_axi_in_23_AWPROT,
    output wire [                                   3:0] m_axi_in_23_AWQOS,
    input wire                                           m_axi_in_23_AWREADY,
    output wire [                                   2:0] m_axi_in_23_AWSIZE,
    output wire                                          m_axi_in_23_AWVALID,
    input wire  [                                   0:0] m_axi_in_23_BID,
    output wire                                          m_axi_in_23_BREADY,
    input wire  [                                   1:0] m_axi_in_23_BRESP,
    input wire                                           m_axi_in_23_BVALID,
    input wire  [                                 255:0] m_axi_in_23_RDATA,
    input wire  [                                   0:0] m_axi_in_23_RID,
    input wire                                           m_axi_in_23_RLAST,
    output wire                                          m_axi_in_23_RREADY,
    input wire  [                                   1:0] m_axi_in_23_RRESP,
    input wire                                           m_axi_in_23_RVALID,
    output wire [                                 255:0] m_axi_in_23_WDATA,
    output wire                                          m_axi_in_23_WLAST,
    input wire                                           m_axi_in_23_WREADY,
    output wire [                                  31:0] m_axi_in_23_WSTRB,
    output wire                                          m_axi_in_23_WVALID,
    output wire [                                  63:0] m_axi_in_24_ARADDR,
    output wire [                                   1:0] m_axi_in_24_ARBURST,
    output wire [                                   3:0] m_axi_in_24_ARCACHE,
    output wire [                                   0:0] m_axi_in_24_ARID,
    output wire [                                   7:0] m_axi_in_24_ARLEN,
    output wire                                          m_axi_in_24_ARLOCK,
    output wire [                                   2:0] m_axi_in_24_ARPROT,
    output wire [                                   3:0] m_axi_in_24_ARQOS,
    input wire                                           m_axi_in_24_ARREADY,
    output wire [                                   2:0] m_axi_in_24_ARSIZE,
    output wire                                          m_axi_in_24_ARVALID,
    output wire [                                  63:0] m_axi_in_24_AWADDR,
    output wire [                                   1:0] m_axi_in_24_AWBURST,
    output wire [                                   3:0] m_axi_in_24_AWCACHE,
    output wire [                                   0:0] m_axi_in_24_AWID,
    output wire [                                   7:0] m_axi_in_24_AWLEN,
    output wire                                          m_axi_in_24_AWLOCK,
    output wire [                                   2:0] m_axi_in_24_AWPROT,
    output wire [                                   3:0] m_axi_in_24_AWQOS,
    input wire                                           m_axi_in_24_AWREADY,
    output wire [                                   2:0] m_axi_in_24_AWSIZE,
    output wire                                          m_axi_in_24_AWVALID,
    input wire  [                                   0:0] m_axi_in_24_BID,
    output wire                                          m_axi_in_24_BREADY,
    input wire  [                                   1:0] m_axi_in_24_BRESP,
    input wire                                           m_axi_in_24_BVALID,
    input wire  [                                 255:0] m_axi_in_24_RDATA,
    input wire  [                                   0:0] m_axi_in_24_RID,
    input wire                                           m_axi_in_24_RLAST,
    output wire                                          m_axi_in_24_RREADY,
    input wire  [                                   1:0] m_axi_in_24_RRESP,
    input wire                                           m_axi_in_24_RVALID,
    output wire [                                 255:0] m_axi_in_24_WDATA,
    output wire                                          m_axi_in_24_WLAST,
    input wire                                           m_axi_in_24_WREADY,
    output wire [                                  31:0] m_axi_in_24_WSTRB,
    output wire                                          m_axi_in_24_WVALID,
    output wire [                                  63:0] m_axi_in_25_ARADDR,
    output wire [                                   1:0] m_axi_in_25_ARBURST,
    output wire [                                   3:0] m_axi_in_25_ARCACHE,
    output wire [                                   0:0] m_axi_in_25_ARID,
    output wire [                                   7:0] m_axi_in_25_ARLEN,
    output wire                                          m_axi_in_25_ARLOCK,
    output wire [                                   2:0] m_axi_in_25_ARPROT,
    output wire [                                   3:0] m_axi_in_25_ARQOS,
    input wire                                           m_axi_in_25_ARREADY,
    output wire [                                   2:0] m_axi_in_25_ARSIZE,
    output wire                                          m_axi_in_25_ARVALID,
    output wire [                                  63:0] m_axi_in_25_AWADDR,
    output wire [                                   1:0] m_axi_in_25_AWBURST,
    output wire [                                   3:0] m_axi_in_25_AWCACHE,
    output wire [                                   0:0] m_axi_in_25_AWID,
    output wire [                                   7:0] m_axi_in_25_AWLEN,
    output wire                                          m_axi_in_25_AWLOCK,
    output wire [                                   2:0] m_axi_in_25_AWPROT,
    output wire [                                   3:0] m_axi_in_25_AWQOS,
    input wire                                           m_axi_in_25_AWREADY,
    output wire [                                   2:0] m_axi_in_25_AWSIZE,
    output wire                                          m_axi_in_25_AWVALID,
    input wire  [                                   0:0] m_axi_in_25_BID,
    output wire                                          m_axi_in_25_BREADY,
    input wire  [                                   1:0] m_axi_in_25_BRESP,
    input wire                                           m_axi_in_25_BVALID,
    input wire  [                                 255:0] m_axi_in_25_RDATA,
    input wire  [                                   0:0] m_axi_in_25_RID,
    input wire                                           m_axi_in_25_RLAST,
    output wire                                          m_axi_in_25_RREADY,
    input wire  [                                   1:0] m_axi_in_25_RRESP,
    input wire                                           m_axi_in_25_RVALID,
    output wire [                                 255:0] m_axi_in_25_WDATA,
    output wire                                          m_axi_in_25_WLAST,
    input wire                                           m_axi_in_25_WREADY,
    output wire [                                  31:0] m_axi_in_25_WSTRB,
    output wire                                          m_axi_in_25_WVALID,
    output wire [                                  63:0] m_axi_in_26_ARADDR,
    output wire [                                   1:0] m_axi_in_26_ARBURST,
    output wire [                                   3:0] m_axi_in_26_ARCACHE,
    output wire [                                   0:0] m_axi_in_26_ARID,
    output wire [                                   7:0] m_axi_in_26_ARLEN,
    output wire                                          m_axi_in_26_ARLOCK,
    output wire [                                   2:0] m_axi_in_26_ARPROT,
    output wire [                                   3:0] m_axi_in_26_ARQOS,
    input wire                                           m_axi_in_26_ARREADY,
    output wire [                                   2:0] m_axi_in_26_ARSIZE,
    output wire                                          m_axi_in_26_ARVALID,
    output wire [                                  63:0] m_axi_in_26_AWADDR,
    output wire [                                   1:0] m_axi_in_26_AWBURST,
    output wire [                                   3:0] m_axi_in_26_AWCACHE,
    output wire [                                   0:0] m_axi_in_26_AWID,
    output wire [                                   7:0] m_axi_in_26_AWLEN,
    output wire                                          m_axi_in_26_AWLOCK,
    output wire [                                   2:0] m_axi_in_26_AWPROT,
    output wire [                                   3:0] m_axi_in_26_AWQOS,
    input wire                                           m_axi_in_26_AWREADY,
    output wire [                                   2:0] m_axi_in_26_AWSIZE,
    output wire                                          m_axi_in_26_AWVALID,
    input wire  [                                   0:0] m_axi_in_26_BID,
    output wire                                          m_axi_in_26_BREADY,
    input wire  [                                   1:0] m_axi_in_26_BRESP,
    input wire                                           m_axi_in_26_BVALID,
    input wire  [                                 255:0] m_axi_in_26_RDATA,
    input wire  [                                   0:0] m_axi_in_26_RID,
    input wire                                           m_axi_in_26_RLAST,
    output wire                                          m_axi_in_26_RREADY,
    input wire  [                                   1:0] m_axi_in_26_RRESP,
    input wire                                           m_axi_in_26_RVALID,
    output wire [                                 255:0] m_axi_in_26_WDATA,
    output wire                                          m_axi_in_26_WLAST,
    input wire                                           m_axi_in_26_WREADY,
    output wire [                                  31:0] m_axi_in_26_WSTRB,
    output wire                                          m_axi_in_26_WVALID,
    output wire [                                  63:0] m_axi_in_3_ARADDR,
    output wire [                                   1:0] m_axi_in_3_ARBURST,
    output wire [                                   3:0] m_axi_in_3_ARCACHE,
    output wire [                                   0:0] m_axi_in_3_ARID,
    output wire [                                   7:0] m_axi_in_3_ARLEN,
    output wire                                          m_axi_in_3_ARLOCK,
    output wire [                                   2:0] m_axi_in_3_ARPROT,
    output wire [                                   3:0] m_axi_in_3_ARQOS,
    input wire                                           m_axi_in_3_ARREADY,
    output wire [                                   2:0] m_axi_in_3_ARSIZE,
    output wire                                          m_axi_in_3_ARVALID,
    output wire [                                  63:0] m_axi_in_3_AWADDR,
    output wire [                                   1:0] m_axi_in_3_AWBURST,
    output wire [                                   3:0] m_axi_in_3_AWCACHE,
    output wire [                                   0:0] m_axi_in_3_AWID,
    output wire [                                   7:0] m_axi_in_3_AWLEN,
    output wire                                          m_axi_in_3_AWLOCK,
    output wire [                                   2:0] m_axi_in_3_AWPROT,
    output wire [                                   3:0] m_axi_in_3_AWQOS,
    input wire                                           m_axi_in_3_AWREADY,
    output wire [                                   2:0] m_axi_in_3_AWSIZE,
    output wire                                          m_axi_in_3_AWVALID,
    input wire  [                                   0:0] m_axi_in_3_BID,
    output wire                                          m_axi_in_3_BREADY,
    input wire  [                                   1:0] m_axi_in_3_BRESP,
    input wire                                           m_axi_in_3_BVALID,
    input wire  [                                 255:0] m_axi_in_3_RDATA,
    input wire  [                                   0:0] m_axi_in_3_RID,
    input wire                                           m_axi_in_3_RLAST,
    output wire                                          m_axi_in_3_RREADY,
    input wire  [                                   1:0] m_axi_in_3_RRESP,
    input wire                                           m_axi_in_3_RVALID,
    output wire [                                 255:0] m_axi_in_3_WDATA,
    output wire                                          m_axi_in_3_WLAST,
    input wire                                           m_axi_in_3_WREADY,
    output wire [                                  31:0] m_axi_in_3_WSTRB,
    output wire                                          m_axi_in_3_WVALID,
    output wire [                                  63:0] m_axi_in_4_ARADDR,
    output wire [                                   1:0] m_axi_in_4_ARBURST,
    output wire [                                   3:0] m_axi_in_4_ARCACHE,
    output wire [                                   0:0] m_axi_in_4_ARID,
    output wire [                                   7:0] m_axi_in_4_ARLEN,
    output wire                                          m_axi_in_4_ARLOCK,
    output wire [                                   2:0] m_axi_in_4_ARPROT,
    output wire [                                   3:0] m_axi_in_4_ARQOS,
    input wire                                           m_axi_in_4_ARREADY,
    output wire [                                   2:0] m_axi_in_4_ARSIZE,
    output wire                                          m_axi_in_4_ARVALID,
    output wire [                                  63:0] m_axi_in_4_AWADDR,
    output wire [                                   1:0] m_axi_in_4_AWBURST,
    output wire [                                   3:0] m_axi_in_4_AWCACHE,
    output wire [                                   0:0] m_axi_in_4_AWID,
    output wire [                                   7:0] m_axi_in_4_AWLEN,
    output wire                                          m_axi_in_4_AWLOCK,
    output wire [                                   2:0] m_axi_in_4_AWPROT,
    output wire [                                   3:0] m_axi_in_4_AWQOS,
    input wire                                           m_axi_in_4_AWREADY,
    output wire [                                   2:0] m_axi_in_4_AWSIZE,
    output wire                                          m_axi_in_4_AWVALID,
    input wire  [                                   0:0] m_axi_in_4_BID,
    output wire                                          m_axi_in_4_BREADY,
    input wire  [                                   1:0] m_axi_in_4_BRESP,
    input wire                                           m_axi_in_4_BVALID,
    input wire  [                                 255:0] m_axi_in_4_RDATA,
    input wire  [                                   0:0] m_axi_in_4_RID,
    input wire                                           m_axi_in_4_RLAST,
    output wire                                          m_axi_in_4_RREADY,
    input wire  [                                   1:0] m_axi_in_4_RRESP,
    input wire                                           m_axi_in_4_RVALID,
    output wire [                                 255:0] m_axi_in_4_WDATA,
    output wire                                          m_axi_in_4_WLAST,
    input wire                                           m_axi_in_4_WREADY,
    output wire [                                  31:0] m_axi_in_4_WSTRB,
    output wire                                          m_axi_in_4_WVALID,
    output wire [                                  63:0] m_axi_in_5_ARADDR,
    output wire [                                   1:0] m_axi_in_5_ARBURST,
    output wire [                                   3:0] m_axi_in_5_ARCACHE,
    output wire [                                   0:0] m_axi_in_5_ARID,
    output wire [                                   7:0] m_axi_in_5_ARLEN,
    output wire                                          m_axi_in_5_ARLOCK,
    output wire [                                   2:0] m_axi_in_5_ARPROT,
    output wire [                                   3:0] m_axi_in_5_ARQOS,
    input wire                                           m_axi_in_5_ARREADY,
    output wire [                                   2:0] m_axi_in_5_ARSIZE,
    output wire                                          m_axi_in_5_ARVALID,
    output wire [                                  63:0] m_axi_in_5_AWADDR,
    output wire [                                   1:0] m_axi_in_5_AWBURST,
    output wire [                                   3:0] m_axi_in_5_AWCACHE,
    output wire [                                   0:0] m_axi_in_5_AWID,
    output wire [                                   7:0] m_axi_in_5_AWLEN,
    output wire                                          m_axi_in_5_AWLOCK,
    output wire [                                   2:0] m_axi_in_5_AWPROT,
    output wire [                                   3:0] m_axi_in_5_AWQOS,
    input wire                                           m_axi_in_5_AWREADY,
    output wire [                                   2:0] m_axi_in_5_AWSIZE,
    output wire                                          m_axi_in_5_AWVALID,
    input wire  [                                   0:0] m_axi_in_5_BID,
    output wire                                          m_axi_in_5_BREADY,
    input wire  [                                   1:0] m_axi_in_5_BRESP,
    input wire                                           m_axi_in_5_BVALID,
    input wire  [                                 255:0] m_axi_in_5_RDATA,
    input wire  [                                   0:0] m_axi_in_5_RID,
    input wire                                           m_axi_in_5_RLAST,
    output wire                                          m_axi_in_5_RREADY,
    input wire  [                                   1:0] m_axi_in_5_RRESP,
    input wire                                           m_axi_in_5_RVALID,
    output wire [                                 255:0] m_axi_in_5_WDATA,
    output wire                                          m_axi_in_5_WLAST,
    input wire                                           m_axi_in_5_WREADY,
    output wire [                                  31:0] m_axi_in_5_WSTRB,
    output wire                                          m_axi_in_5_WVALID,
    output wire [                                  63:0] m_axi_in_6_ARADDR,
    output wire [                                   1:0] m_axi_in_6_ARBURST,
    output wire [                                   3:0] m_axi_in_6_ARCACHE,
    output wire [                                   0:0] m_axi_in_6_ARID,
    output wire [                                   7:0] m_axi_in_6_ARLEN,
    output wire                                          m_axi_in_6_ARLOCK,
    output wire [                                   2:0] m_axi_in_6_ARPROT,
    output wire [                                   3:0] m_axi_in_6_ARQOS,
    input wire                                           m_axi_in_6_ARREADY,
    output wire [                                   2:0] m_axi_in_6_ARSIZE,
    output wire                                          m_axi_in_6_ARVALID,
    output wire [                                  63:0] m_axi_in_6_AWADDR,
    output wire [                                   1:0] m_axi_in_6_AWBURST,
    output wire [                                   3:0] m_axi_in_6_AWCACHE,
    output wire [                                   0:0] m_axi_in_6_AWID,
    output wire [                                   7:0] m_axi_in_6_AWLEN,
    output wire                                          m_axi_in_6_AWLOCK,
    output wire [                                   2:0] m_axi_in_6_AWPROT,
    output wire [                                   3:0] m_axi_in_6_AWQOS,
    input wire                                           m_axi_in_6_AWREADY,
    output wire [                                   2:0] m_axi_in_6_AWSIZE,
    output wire                                          m_axi_in_6_AWVALID,
    input wire  [                                   0:0] m_axi_in_6_BID,
    output wire                                          m_axi_in_6_BREADY,
    input wire  [                                   1:0] m_axi_in_6_BRESP,
    input wire                                           m_axi_in_6_BVALID,
    input wire  [                                 255:0] m_axi_in_6_RDATA,
    input wire  [                                   0:0] m_axi_in_6_RID,
    input wire                                           m_axi_in_6_RLAST,
    output wire                                          m_axi_in_6_RREADY,
    input wire  [                                   1:0] m_axi_in_6_RRESP,
    input wire                                           m_axi_in_6_RVALID,
    output wire [                                 255:0] m_axi_in_6_WDATA,
    output wire                                          m_axi_in_6_WLAST,
    input wire                                           m_axi_in_6_WREADY,
    output wire [                                  31:0] m_axi_in_6_WSTRB,
    output wire                                          m_axi_in_6_WVALID,
    output wire [                                  63:0] m_axi_in_7_ARADDR,
    output wire [                                   1:0] m_axi_in_7_ARBURST,
    output wire [                                   3:0] m_axi_in_7_ARCACHE,
    output wire [                                   0:0] m_axi_in_7_ARID,
    output wire [                                   7:0] m_axi_in_7_ARLEN,
    output wire                                          m_axi_in_7_ARLOCK,
    output wire [                                   2:0] m_axi_in_7_ARPROT,
    output wire [                                   3:0] m_axi_in_7_ARQOS,
    input wire                                           m_axi_in_7_ARREADY,
    output wire [                                   2:0] m_axi_in_7_ARSIZE,
    output wire                                          m_axi_in_7_ARVALID,
    output wire [                                  63:0] m_axi_in_7_AWADDR,
    output wire [                                   1:0] m_axi_in_7_AWBURST,
    output wire [                                   3:0] m_axi_in_7_AWCACHE,
    output wire [                                   0:0] m_axi_in_7_AWID,
    output wire [                                   7:0] m_axi_in_7_AWLEN,
    output wire                                          m_axi_in_7_AWLOCK,
    output wire [                                   2:0] m_axi_in_7_AWPROT,
    output wire [                                   3:0] m_axi_in_7_AWQOS,
    input wire                                           m_axi_in_7_AWREADY,
    output wire [                                   2:0] m_axi_in_7_AWSIZE,
    output wire                                          m_axi_in_7_AWVALID,
    input wire  [                                   0:0] m_axi_in_7_BID,
    output wire                                          m_axi_in_7_BREADY,
    input wire  [                                   1:0] m_axi_in_7_BRESP,
    input wire                                           m_axi_in_7_BVALID,
    input wire  [                                 255:0] m_axi_in_7_RDATA,
    input wire  [                                   0:0] m_axi_in_7_RID,
    input wire                                           m_axi_in_7_RLAST,
    output wire                                          m_axi_in_7_RREADY,
    input wire  [                                   1:0] m_axi_in_7_RRESP,
    input wire                                           m_axi_in_7_RVALID,
    output wire [                                 255:0] m_axi_in_7_WDATA,
    output wire                                          m_axi_in_7_WLAST,
    input wire                                           m_axi_in_7_WREADY,
    output wire [                                  31:0] m_axi_in_7_WSTRB,
    output wire                                          m_axi_in_7_WVALID,
    output wire [                                  63:0] m_axi_in_8_ARADDR,
    output wire [                                   1:0] m_axi_in_8_ARBURST,
    output wire [                                   3:0] m_axi_in_8_ARCACHE,
    output wire [                                   0:0] m_axi_in_8_ARID,
    output wire [                                   7:0] m_axi_in_8_ARLEN,
    output wire                                          m_axi_in_8_ARLOCK,
    output wire [                                   2:0] m_axi_in_8_ARPROT,
    output wire [                                   3:0] m_axi_in_8_ARQOS,
    input wire                                           m_axi_in_8_ARREADY,
    output wire [                                   2:0] m_axi_in_8_ARSIZE,
    output wire                                          m_axi_in_8_ARVALID,
    output wire [                                  63:0] m_axi_in_8_AWADDR,
    output wire [                                   1:0] m_axi_in_8_AWBURST,
    output wire [                                   3:0] m_axi_in_8_AWCACHE,
    output wire [                                   0:0] m_axi_in_8_AWID,
    output wire [                                   7:0] m_axi_in_8_AWLEN,
    output wire                                          m_axi_in_8_AWLOCK,
    output wire [                                   2:0] m_axi_in_8_AWPROT,
    output wire [                                   3:0] m_axi_in_8_AWQOS,
    input wire                                           m_axi_in_8_AWREADY,
    output wire [                                   2:0] m_axi_in_8_AWSIZE,
    output wire                                          m_axi_in_8_AWVALID,
    input wire  [                                   0:0] m_axi_in_8_BID,
    output wire                                          m_axi_in_8_BREADY,
    input wire  [                                   1:0] m_axi_in_8_BRESP,
    input wire                                           m_axi_in_8_BVALID,
    input wire  [                                 255:0] m_axi_in_8_RDATA,
    input wire  [                                   0:0] m_axi_in_8_RID,
    input wire                                           m_axi_in_8_RLAST,
    output wire                                          m_axi_in_8_RREADY,
    input wire  [                                   1:0] m_axi_in_8_RRESP,
    input wire                                           m_axi_in_8_RVALID,
    output wire [                                 255:0] m_axi_in_8_WDATA,
    output wire                                          m_axi_in_8_WLAST,
    input wire                                           m_axi_in_8_WREADY,
    output wire [                                  31:0] m_axi_in_8_WSTRB,
    output wire                                          m_axi_in_8_WVALID,
    output wire [                                  63:0] m_axi_in_9_ARADDR,
    output wire [                                   1:0] m_axi_in_9_ARBURST,
    output wire [                                   3:0] m_axi_in_9_ARCACHE,
    output wire [                                   0:0] m_axi_in_9_ARID,
    output wire [                                   7:0] m_axi_in_9_ARLEN,
    output wire                                          m_axi_in_9_ARLOCK,
    output wire [                                   2:0] m_axi_in_9_ARPROT,
    output wire [                                   3:0] m_axi_in_9_ARQOS,
    input wire                                           m_axi_in_9_ARREADY,
    output wire [                                   2:0] m_axi_in_9_ARSIZE,
    output wire                                          m_axi_in_9_ARVALID,
    output wire [                                  63:0] m_axi_in_9_AWADDR,
    output wire [                                   1:0] m_axi_in_9_AWBURST,
    output wire [                                   3:0] m_axi_in_9_AWCACHE,
    output wire [                                   0:0] m_axi_in_9_AWID,
    output wire [                                   7:0] m_axi_in_9_AWLEN,
    output wire                                          m_axi_in_9_AWLOCK,
    output wire [                                   2:0] m_axi_in_9_AWPROT,
    output wire [                                   3:0] m_axi_in_9_AWQOS,
    input wire                                           m_axi_in_9_AWREADY,
    output wire [                                   2:0] m_axi_in_9_AWSIZE,
    output wire                                          m_axi_in_9_AWVALID,
    input wire  [                                   0:0] m_axi_in_9_BID,
    output wire                                          m_axi_in_9_BREADY,
    input wire  [                                   1:0] m_axi_in_9_BRESP,
    input wire                                           m_axi_in_9_BVALID,
    input wire  [                                 255:0] m_axi_in_9_RDATA,
    input wire  [                                   0:0] m_axi_in_9_RID,
    input wire                                           m_axi_in_9_RLAST,
    output wire                                          m_axi_in_9_RREADY,
    input wire  [                                   1:0] m_axi_in_9_RRESP,
    input wire                                           m_axi_in_9_RVALID,
    output wire [                                 255:0] m_axi_in_9_WDATA,
    output wire                                          m_axi_in_9_WLAST,
    input wire                                           m_axi_in_9_WREADY,
    output wire [                                  31:0] m_axi_in_9_WSTRB,
    output wire                                          m_axi_in_9_WVALID,
    output wire                                          control_s_axi_U_ACLK,
    output wire                                          control_s_axi_U_ACLK_EN,
    output wire [    (C_S_AXI_CONTROL_ADDR_WIDTH - 1):0] control_s_axi_U_ARADDR,
    output wire                                          control_s_axi_U_ARESET,
    input wire                                           control_s_axi_U_ARREADY,
    output wire                                          control_s_axi_U_ARVALID,
    output wire [    (C_S_AXI_CONTROL_ADDR_WIDTH - 1):0] control_s_axi_U_AWADDR,
    input wire                                           control_s_axi_U_AWREADY,
    output wire                                          control_s_axi_U_AWVALID,
    output wire                                          control_s_axi_U_BREADY,
    input wire  [                                   1:0] control_s_axi_U_BRESP,
    input wire                                           control_s_axi_U_BVALID,
    input wire  [                                  63:0] control_s_axi_U_L3_out_dist,
    input wire  [                                  63:0] control_s_axi_U_L3_out_id,
    input wire  [    (C_S_AXI_CONTROL_DATA_WIDTH - 1):0] control_s_axi_U_RDATA,
    output wire                                          control_s_axi_U_RREADY,
    input wire  [                                   1:0] control_s_axi_U_RRESP,
    input wire                                           control_s_axi_U_RVALID,
    output wire [    (C_S_AXI_CONTROL_DATA_WIDTH - 1):0] control_s_axi_U_WDATA,
    input wire                                           control_s_axi_U_WREADY,
    output wire [(C_S_AXI_CONTROL_DATA_WIDTH / 8 - 1):0] control_s_axi_U_WSTRB,
    output wire                                          control_s_axi_U_WVALID,
    output wire                                          control_s_axi_U_ap_done,
    output wire                                          control_s_axi_U_ap_idle,
    output wire                                          control_s_axi_U_ap_ready,
    input wire                                           control_s_axi_U_ap_start,
    input wire  [                                  63:0] control_s_axi_U_in_0,
    input wire  [                                  63:0] control_s_axi_U_in_1,
    input wire  [                                  63:0] control_s_axi_U_in_10,
    input wire  [                                  63:0] control_s_axi_U_in_11,
    input wire  [                                  63:0] control_s_axi_U_in_12,
    input wire  [                                  63:0] control_s_axi_U_in_13,
    input wire  [                                  63:0] control_s_axi_U_in_14,
    input wire  [                                  63:0] control_s_axi_U_in_15,
    input wire  [                                  63:0] control_s_axi_U_in_16,
    input wire  [                                  63:0] control_s_axi_U_in_17,
    input wire  [                                  63:0] control_s_axi_U_in_18,
    input wire  [                                  63:0] control_s_axi_U_in_19,
    input wire  [                                  63:0] control_s_axi_U_in_2,
    input wire  [                                  63:0] control_s_axi_U_in_20,
    input wire  [                                  63:0] control_s_axi_U_in_21,
    input wire  [                                  63:0] control_s_axi_U_in_22,
    input wire  [                                  63:0] control_s_axi_U_in_23,
    input wire  [                                  63:0] control_s_axi_U_in_24,
    input wire  [                                  63:0] control_s_axi_U_in_25,
    input wire  [                                  63:0] control_s_axi_U_in_26,
    input wire  [                                  63:0] control_s_axi_U_in_3,
    input wire  [                                  63:0] control_s_axi_U_in_4,
    input wire  [                                  63:0] control_s_axi_U_in_5,
    input wire  [                                  63:0] control_s_axi_U_in_6,
    input wire  [                                  63:0] control_s_axi_U_in_7,
    input wire  [                                  63:0] control_s_axi_U_in_8,
    input wire  [                                  63:0] control_s_axi_U_in_9,
    input wire                                           control_s_axi_U_interrupt,
    output wire                                          L1_out_dist_0_clk,
    output wire [                                  65:0] L1_out_dist_0_if_din,
    input wire  [                                  65:0] L1_out_dist_0_if_dout,
    input wire                                           L1_out_dist_0_if_empty_n,
    input wire                                           L1_out_dist_0_if_full_n,
    output wire                                          L1_out_dist_0_if_read,
    output wire                                          L1_out_dist_0_if_read_ce,
    output wire                                          L1_out_dist_0_if_write,
    output wire                                          L1_out_dist_0_if_write_ce,
    output wire                                          L1_out_dist_0_reset,
    output wire                                          L1_out_dist_1_clk,
    output wire [                                  65:0] L1_out_dist_1_if_din,
    input wire  [                                  65:0] L1_out_dist_1_if_dout,
    input wire                                           L1_out_dist_1_if_empty_n,
    input wire                                           L1_out_dist_1_if_full_n,
    output wire                                          L1_out_dist_1_if_read,
    output wire                                          L1_out_dist_1_if_read_ce,
    output wire                                          L1_out_dist_1_if_write,
    output wire                                          L1_out_dist_1_if_write_ce,
    output wire                                          L1_out_dist_1_reset,
    output wire                                          L1_out_dist_2_clk,
    output wire [                                  65:0] L1_out_dist_2_if_din,
    input wire  [                                  65:0] L1_out_dist_2_if_dout,
    input wire                                           L1_out_dist_2_if_empty_n,
    input wire                                           L1_out_dist_2_if_full_n,
    output wire                                          L1_out_dist_2_if_read,
    output wire                                          L1_out_dist_2_if_read_ce,
    output wire                                          L1_out_dist_2_if_write,
    output wire                                          L1_out_dist_2_if_write_ce,
    output wire                                          L1_out_dist_2_reset,
    output wire                                          L1_out_dist_3_clk,
    output wire [                                  65:0] L1_out_dist_3_if_din,
    input wire  [                                  65:0] L1_out_dist_3_if_dout,
    input wire                                           L1_out_dist_3_if_empty_n,
    input wire                                           L1_out_dist_3_if_full_n,
    output wire                                          L1_out_dist_3_if_read,
    output wire                                          L1_out_dist_3_if_read_ce,
    output wire                                          L1_out_dist_3_if_write,
    output wire                                          L1_out_dist_3_if_write_ce,
    output wire                                          L1_out_dist_3_reset,
    output wire                                          L1_out_dist_4_clk,
    output wire [                                  65:0] L1_out_dist_4_if_din,
    input wire  [                                  65:0] L1_out_dist_4_if_dout,
    input wire                                           L1_out_dist_4_if_empty_n,
    input wire                                           L1_out_dist_4_if_full_n,
    output wire                                          L1_out_dist_4_if_read,
    output wire                                          L1_out_dist_4_if_read_ce,
    output wire                                          L1_out_dist_4_if_write,
    output wire                                          L1_out_dist_4_if_write_ce,
    output wire                                          L1_out_dist_4_reset,
    output wire                                          L1_out_dist_5_clk,
    output wire [                                  65:0] L1_out_dist_5_if_din,
    input wire  [                                  65:0] L1_out_dist_5_if_dout,
    input wire                                           L1_out_dist_5_if_empty_n,
    input wire                                           L1_out_dist_5_if_full_n,
    output wire                                          L1_out_dist_5_if_read,
    output wire                                          L1_out_dist_5_if_read_ce,
    output wire                                          L1_out_dist_5_if_write,
    output wire                                          L1_out_dist_5_if_write_ce,
    output wire                                          L1_out_dist_5_reset,
    output wire                                          L1_out_dist_6_clk,
    output wire [                                  65:0] L1_out_dist_6_if_din,
    input wire  [                                  65:0] L1_out_dist_6_if_dout,
    input wire                                           L1_out_dist_6_if_empty_n,
    input wire                                           L1_out_dist_6_if_full_n,
    output wire                                          L1_out_dist_6_if_read,
    output wire                                          L1_out_dist_6_if_read_ce,
    output wire                                          L1_out_dist_6_if_write,
    output wire                                          L1_out_dist_6_if_write_ce,
    output wire                                          L1_out_dist_6_reset,
    output wire                                          L1_out_dist_7_clk,
    output wire [                                  65:0] L1_out_dist_7_if_din,
    input wire  [                                  65:0] L1_out_dist_7_if_dout,
    input wire                                           L1_out_dist_7_if_empty_n,
    input wire                                           L1_out_dist_7_if_full_n,
    output wire                                          L1_out_dist_7_if_read,
    output wire                                          L1_out_dist_7_if_read_ce,
    output wire                                          L1_out_dist_7_if_write,
    output wire                                          L1_out_dist_7_if_write_ce,
    output wire                                          L1_out_dist_7_reset,
    output wire                                          L1_out_dist_8_clk,
    output wire [                                  65:0] L1_out_dist_8_if_din,
    input wire  [                                  65:0] L1_out_dist_8_if_dout,
    input wire                                           L1_out_dist_8_if_empty_n,
    input wire                                           L1_out_dist_8_if_full_n,
    output wire                                          L1_out_dist_8_if_read,
    output wire                                          L1_out_dist_8_if_read_ce,
    output wire                                          L1_out_dist_8_if_write,
    output wire                                          L1_out_dist_8_if_write_ce,
    output wire                                          L1_out_dist_8_reset,
    output wire                                          L1_out_id_0_clk,
    output wire [                                  65:0] L1_out_id_0_if_din,
    input wire  [                                  65:0] L1_out_id_0_if_dout,
    input wire                                           L1_out_id_0_if_empty_n,
    input wire                                           L1_out_id_0_if_full_n,
    output wire                                          L1_out_id_0_if_read,
    output wire                                          L1_out_id_0_if_read_ce,
    output wire                                          L1_out_id_0_if_write,
    output wire                                          L1_out_id_0_if_write_ce,
    output wire                                          L1_out_id_0_reset,
    output wire                                          L1_out_id_1_clk,
    output wire [                                  65:0] L1_out_id_1_if_din,
    input wire  [                                  65:0] L1_out_id_1_if_dout,
    input wire                                           L1_out_id_1_if_empty_n,
    input wire                                           L1_out_id_1_if_full_n,
    output wire                                          L1_out_id_1_if_read,
    output wire                                          L1_out_id_1_if_read_ce,
    output wire                                          L1_out_id_1_if_write,
    output wire                                          L1_out_id_1_if_write_ce,
    output wire                                          L1_out_id_1_reset,
    output wire                                          L1_out_id_2_clk,
    output wire [                                  65:0] L1_out_id_2_if_din,
    input wire  [                                  65:0] L1_out_id_2_if_dout,
    input wire                                           L1_out_id_2_if_empty_n,
    input wire                                           L1_out_id_2_if_full_n,
    output wire                                          L1_out_id_2_if_read,
    output wire                                          L1_out_id_2_if_read_ce,
    output wire                                          L1_out_id_2_if_write,
    output wire                                          L1_out_id_2_if_write_ce,
    output wire                                          L1_out_id_2_reset,
    output wire                                          L1_out_id_3_clk,
    output wire [                                  65:0] L1_out_id_3_if_din,
    input wire  [                                  65:0] L1_out_id_3_if_dout,
    input wire                                           L1_out_id_3_if_empty_n,
    input wire                                           L1_out_id_3_if_full_n,
    output wire                                          L1_out_id_3_if_read,
    output wire                                          L1_out_id_3_if_read_ce,
    output wire                                          L1_out_id_3_if_write,
    output wire                                          L1_out_id_3_if_write_ce,
    output wire                                          L1_out_id_3_reset,
    output wire                                          L1_out_id_4_clk,
    output wire [                                  65:0] L1_out_id_4_if_din,
    input wire  [                                  65:0] L1_out_id_4_if_dout,
    input wire                                           L1_out_id_4_if_empty_n,
    input wire                                           L1_out_id_4_if_full_n,
    output wire                                          L1_out_id_4_if_read,
    output wire                                          L1_out_id_4_if_read_ce,
    output wire                                          L1_out_id_4_if_write,
    output wire                                          L1_out_id_4_if_write_ce,
    output wire                                          L1_out_id_4_reset,
    output wire                                          L1_out_id_5_clk,
    output wire [                                  65:0] L1_out_id_5_if_din,
    input wire  [                                  65:0] L1_out_id_5_if_dout,
    input wire                                           L1_out_id_5_if_empty_n,
    input wire                                           L1_out_id_5_if_full_n,
    output wire                                          L1_out_id_5_if_read,
    output wire                                          L1_out_id_5_if_read_ce,
    output wire                                          L1_out_id_5_if_write,
    output wire                                          L1_out_id_5_if_write_ce,
    output wire                                          L1_out_id_5_reset,
    output wire                                          L1_out_id_6_clk,
    output wire [                                  65:0] L1_out_id_6_if_din,
    input wire  [                                  65:0] L1_out_id_6_if_dout,
    input wire                                           L1_out_id_6_if_empty_n,
    input wire                                           L1_out_id_6_if_full_n,
    output wire                                          L1_out_id_6_if_read,
    output wire                                          L1_out_id_6_if_read_ce,
    output wire                                          L1_out_id_6_if_write,
    output wire                                          L1_out_id_6_if_write_ce,
    output wire                                          L1_out_id_6_reset,
    output wire                                          L1_out_id_7_clk,
    output wire [                                  65:0] L1_out_id_7_if_din,
    input wire  [                                  65:0] L1_out_id_7_if_dout,
    input wire                                           L1_out_id_7_if_empty_n,
    input wire                                           L1_out_id_7_if_full_n,
    output wire                                          L1_out_id_7_if_read,
    output wire                                          L1_out_id_7_if_read_ce,
    output wire                                          L1_out_id_7_if_write,
    output wire                                          L1_out_id_7_if_write_ce,
    output wire                                          L1_out_id_7_reset,
    output wire                                          L1_out_id_8_clk,
    output wire [                                  65:0] L1_out_id_8_if_din,
    input wire  [                                  65:0] L1_out_id_8_if_dout,
    input wire                                           L1_out_id_8_if_empty_n,
    input wire                                           L1_out_id_8_if_full_n,
    output wire                                          L1_out_id_8_if_read,
    output wire                                          L1_out_id_8_if_read_ce,
    output wire                                          L1_out_id_8_if_write,
    output wire                                          L1_out_id_8_if_write_ce,
    output wire                                          L1_out_id_8_reset,
    output wire                                          L2_out_dist0_clk,
    output wire [                                  65:0] L2_out_dist0_if_din,
    input wire  [                                  65:0] L2_out_dist0_if_dout,
    input wire                                           L2_out_dist0_if_empty_n,
    input wire                                           L2_out_dist0_if_full_n,
    output wire                                          L2_out_dist0_if_read,
    output wire                                          L2_out_dist0_if_read_ce,
    output wire                                          L2_out_dist0_if_write,
    output wire                                          L2_out_dist0_if_write_ce,
    output wire                                          L2_out_dist0_reset,
    output wire                                          L2_out_dist1_clk,
    output wire [                                  65:0] L2_out_dist1_if_din,
    input wire  [                                  65:0] L2_out_dist1_if_dout,
    input wire                                           L2_out_dist1_if_empty_n,
    input wire                                           L2_out_dist1_if_full_n,
    output wire                                          L2_out_dist1_if_read,
    output wire                                          L2_out_dist1_if_read_ce,
    output wire                                          L2_out_dist1_if_write,
    output wire                                          L2_out_dist1_if_write_ce,
    output wire                                          L2_out_dist1_reset,
    output wire                                          L2_out_dist2_clk,
    output wire [                                  65:0] L2_out_dist2_if_din,
    input wire  [                                  65:0] L2_out_dist2_if_dout,
    input wire                                           L2_out_dist2_if_empty_n,
    input wire                                           L2_out_dist2_if_full_n,
    output wire                                          L2_out_dist2_if_read,
    output wire                                          L2_out_dist2_if_read_ce,
    output wire                                          L2_out_dist2_if_write,
    output wire                                          L2_out_dist2_if_write_ce,
    output wire                                          L2_out_dist2_reset,
    output wire                                          L2_out_id0_clk,
    output wire [                                  65:0] L2_out_id0_if_din,
    input wire  [                                  65:0] L2_out_id0_if_dout,
    input wire                                           L2_out_id0_if_empty_n,
    input wire                                           L2_out_id0_if_full_n,
    output wire                                          L2_out_id0_if_read,
    output wire                                          L2_out_id0_if_read_ce,
    output wire                                          L2_out_id0_if_write,
    output wire                                          L2_out_id0_if_write_ce,
    output wire                                          L2_out_id0_reset,
    output wire                                          L2_out_id1_clk,
    output wire [                                  65:0] L2_out_id1_if_din,
    input wire  [                                  65:0] L2_out_id1_if_dout,
    input wire                                           L2_out_id1_if_empty_n,
    input wire                                           L2_out_id1_if_full_n,
    output wire                                          L2_out_id1_if_read,
    output wire                                          L2_out_id1_if_read_ce,
    output wire                                          L2_out_id1_if_write,
    output wire                                          L2_out_id1_if_write_ce,
    output wire                                          L2_out_id1_reset,
    output wire                                          L2_out_id2_clk,
    output wire [                                  65:0] L2_out_id2_if_din,
    input wire  [                                  65:0] L2_out_id2_if_dout,
    input wire                                           L2_out_id2_if_empty_n,
    input wire                                           L2_out_id2_if_full_n,
    output wire                                          L2_out_id2_if_read,
    output wire                                          L2_out_id2_if_read_ce,
    output wire                                          L2_out_id2_if_write,
    output wire                                          L2_out_id2_if_write_ce,
    output wire                                          L2_out_id2_reset,
    output wire                                          L3_out_dist_stream_clk,
    output wire [                                  65:0] L3_out_dist_stream_if_din,
    input wire  [                                  65:0] L3_out_dist_stream_if_dout,
    input wire                                           L3_out_dist_stream_if_empty_n,
    input wire                                           L3_out_dist_stream_if_full_n,
    output wire                                          L3_out_dist_stream_if_read,
    output wire                                          L3_out_dist_stream_if_read_ce,
    output wire                                          L3_out_dist_stream_if_write,
    output wire                                          L3_out_dist_stream_if_write_ce,
    output wire                                          L3_out_dist_stream_reset,
    output wire                                          L3_out_id_stream_clk,
    output wire [                                  65:0] L3_out_id_stream_if_din,
    input wire  [                                  65:0] L3_out_id_stream_if_dout,
    input wire                                           L3_out_id_stream_if_empty_n,
    input wire                                           L3_out_id_stream_if_full_n,
    output wire                                          L3_out_id_stream_if_read,
    output wire                                          L3_out_id_stream_if_read_ce,
    output wire                                          L3_out_id_stream_if_write,
    output wire                                          L3_out_id_stream_if_write_ce,
    output wire                                          L3_out_id_stream_reset,
    output wire                                          out_dist_0_clk,
    output wire [                                  65:0] out_dist_0_if_din,
    input wire  [                                  65:0] out_dist_0_if_dout,
    input wire                                           out_dist_0_if_empty_n,
    input wire                                           out_dist_0_if_full_n,
    output wire                                          out_dist_0_if_read,
    output wire                                          out_dist_0_if_read_ce,
    output wire                                          out_dist_0_if_write,
    output wire                                          out_dist_0_if_write_ce,
    output wire                                          out_dist_0_reset,
    output wire                                          out_dist_10_clk,
    output wire [                                  65:0] out_dist_10_if_din,
    input wire  [                                  65:0] out_dist_10_if_dout,
    input wire                                           out_dist_10_if_empty_n,
    input wire                                           out_dist_10_if_full_n,
    output wire                                          out_dist_10_if_read,
    output wire                                          out_dist_10_if_read_ce,
    output wire                                          out_dist_10_if_write,
    output wire                                          out_dist_10_if_write_ce,
    output wire                                          out_dist_10_reset,
    output wire                                          out_dist_11_clk,
    output wire [                                  65:0] out_dist_11_if_din,
    input wire  [                                  65:0] out_dist_11_if_dout,
    input wire                                           out_dist_11_if_empty_n,
    input wire                                           out_dist_11_if_full_n,
    output wire                                          out_dist_11_if_read,
    output wire                                          out_dist_11_if_read_ce,
    output wire                                          out_dist_11_if_write,
    output wire                                          out_dist_11_if_write_ce,
    output wire                                          out_dist_11_reset,
    output wire                                          out_dist_12_clk,
    output wire [                                  65:0] out_dist_12_if_din,
    input wire  [                                  65:0] out_dist_12_if_dout,
    input wire                                           out_dist_12_if_empty_n,
    input wire                                           out_dist_12_if_full_n,
    output wire                                          out_dist_12_if_read,
    output wire                                          out_dist_12_if_read_ce,
    output wire                                          out_dist_12_if_write,
    output wire                                          out_dist_12_if_write_ce,
    output wire                                          out_dist_12_reset,
    output wire                                          out_dist_13_clk,
    output wire [                                  65:0] out_dist_13_if_din,
    input wire  [                                  65:0] out_dist_13_if_dout,
    input wire                                           out_dist_13_if_empty_n,
    input wire                                           out_dist_13_if_full_n,
    output wire                                          out_dist_13_if_read,
    output wire                                          out_dist_13_if_read_ce,
    output wire                                          out_dist_13_if_write,
    output wire                                          out_dist_13_if_write_ce,
    output wire                                          out_dist_13_reset,
    output wire                                          out_dist_14_clk,
    output wire [                                  65:0] out_dist_14_if_din,
    input wire  [                                  65:0] out_dist_14_if_dout,
    input wire                                           out_dist_14_if_empty_n,
    input wire                                           out_dist_14_if_full_n,
    output wire                                          out_dist_14_if_read,
    output wire                                          out_dist_14_if_read_ce,
    output wire                                          out_dist_14_if_write,
    output wire                                          out_dist_14_if_write_ce,
    output wire                                          out_dist_14_reset,
    output wire                                          out_dist_15_clk,
    output wire [                                  65:0] out_dist_15_if_din,
    input wire  [                                  65:0] out_dist_15_if_dout,
    input wire                                           out_dist_15_if_empty_n,
    input wire                                           out_dist_15_if_full_n,
    output wire                                          out_dist_15_if_read,
    output wire                                          out_dist_15_if_read_ce,
    output wire                                          out_dist_15_if_write,
    output wire                                          out_dist_15_if_write_ce,
    output wire                                          out_dist_15_reset,
    output wire                                          out_dist_16_clk,
    output wire [                                  65:0] out_dist_16_if_din,
    input wire  [                                  65:0] out_dist_16_if_dout,
    input wire                                           out_dist_16_if_empty_n,
    input wire                                           out_dist_16_if_full_n,
    output wire                                          out_dist_16_if_read,
    output wire                                          out_dist_16_if_read_ce,
    output wire                                          out_dist_16_if_write,
    output wire                                          out_dist_16_if_write_ce,
    output wire                                          out_dist_16_reset,
    output wire                                          out_dist_17_clk,
    output wire [                                  65:0] out_dist_17_if_din,
    input wire  [                                  65:0] out_dist_17_if_dout,
    input wire                                           out_dist_17_if_empty_n,
    input wire                                           out_dist_17_if_full_n,
    output wire                                          out_dist_17_if_read,
    output wire                                          out_dist_17_if_read_ce,
    output wire                                          out_dist_17_if_write,
    output wire                                          out_dist_17_if_write_ce,
    output wire                                          out_dist_17_reset,
    output wire                                          out_dist_18_clk,
    output wire [                                  65:0] out_dist_18_if_din,
    input wire  [                                  65:0] out_dist_18_if_dout,
    input wire                                           out_dist_18_if_empty_n,
    input wire                                           out_dist_18_if_full_n,
    output wire                                          out_dist_18_if_read,
    output wire                                          out_dist_18_if_read_ce,
    output wire                                          out_dist_18_if_write,
    output wire                                          out_dist_18_if_write_ce,
    output wire                                          out_dist_18_reset,
    output wire                                          out_dist_19_clk,
    output wire [                                  65:0] out_dist_19_if_din,
    input wire  [                                  65:0] out_dist_19_if_dout,
    input wire                                           out_dist_19_if_empty_n,
    input wire                                           out_dist_19_if_full_n,
    output wire                                          out_dist_19_if_read,
    output wire                                          out_dist_19_if_read_ce,
    output wire                                          out_dist_19_if_write,
    output wire                                          out_dist_19_if_write_ce,
    output wire                                          out_dist_19_reset,
    output wire                                          out_dist_1_clk,
    output wire [                                  65:0] out_dist_1_if_din,
    input wire  [                                  65:0] out_dist_1_if_dout,
    input wire                                           out_dist_1_if_empty_n,
    input wire                                           out_dist_1_if_full_n,
    output wire                                          out_dist_1_if_read,
    output wire                                          out_dist_1_if_read_ce,
    output wire                                          out_dist_1_if_write,
    output wire                                          out_dist_1_if_write_ce,
    output wire                                          out_dist_1_reset,
    output wire                                          out_dist_20_clk,
    output wire [                                  65:0] out_dist_20_if_din,
    input wire  [                                  65:0] out_dist_20_if_dout,
    input wire                                           out_dist_20_if_empty_n,
    input wire                                           out_dist_20_if_full_n,
    output wire                                          out_dist_20_if_read,
    output wire                                          out_dist_20_if_read_ce,
    output wire                                          out_dist_20_if_write,
    output wire                                          out_dist_20_if_write_ce,
    output wire                                          out_dist_20_reset,
    output wire                                          out_dist_21_clk,
    output wire [                                  65:0] out_dist_21_if_din,
    input wire  [                                  65:0] out_dist_21_if_dout,
    input wire                                           out_dist_21_if_empty_n,
    input wire                                           out_dist_21_if_full_n,
    output wire                                          out_dist_21_if_read,
    output wire                                          out_dist_21_if_read_ce,
    output wire                                          out_dist_21_if_write,
    output wire                                          out_dist_21_if_write_ce,
    output wire                                          out_dist_21_reset,
    output wire                                          out_dist_22_clk,
    output wire [                                  65:0] out_dist_22_if_din,
    input wire  [                                  65:0] out_dist_22_if_dout,
    input wire                                           out_dist_22_if_empty_n,
    input wire                                           out_dist_22_if_full_n,
    output wire                                          out_dist_22_if_read,
    output wire                                          out_dist_22_if_read_ce,
    output wire                                          out_dist_22_if_write,
    output wire                                          out_dist_22_if_write_ce,
    output wire                                          out_dist_22_reset,
    output wire                                          out_dist_23_clk,
    output wire [                                  65:0] out_dist_23_if_din,
    input wire  [                                  65:0] out_dist_23_if_dout,
    input wire                                           out_dist_23_if_empty_n,
    input wire                                           out_dist_23_if_full_n,
    output wire                                          out_dist_23_if_read,
    output wire                                          out_dist_23_if_read_ce,
    output wire                                          out_dist_23_if_write,
    output wire                                          out_dist_23_if_write_ce,
    output wire                                          out_dist_23_reset,
    output wire                                          out_dist_24_clk,
    output wire [                                  65:0] out_dist_24_if_din,
    input wire  [                                  65:0] out_dist_24_if_dout,
    input wire                                           out_dist_24_if_empty_n,
    input wire                                           out_dist_24_if_full_n,
    output wire                                          out_dist_24_if_read,
    output wire                                          out_dist_24_if_read_ce,
    output wire                                          out_dist_24_if_write,
    output wire                                          out_dist_24_if_write_ce,
    output wire                                          out_dist_24_reset,
    output wire                                          out_dist_25_clk,
    output wire [                                  65:0] out_dist_25_if_din,
    input wire  [                                  65:0] out_dist_25_if_dout,
    input wire                                           out_dist_25_if_empty_n,
    input wire                                           out_dist_25_if_full_n,
    output wire                                          out_dist_25_if_read,
    output wire                                          out_dist_25_if_read_ce,
    output wire                                          out_dist_25_if_write,
    output wire                                          out_dist_25_if_write_ce,
    output wire                                          out_dist_25_reset,
    output wire                                          out_dist_26_clk,
    output wire [                                  65:0] out_dist_26_if_din,
    input wire  [                                  65:0] out_dist_26_if_dout,
    input wire                                           out_dist_26_if_empty_n,
    input wire                                           out_dist_26_if_full_n,
    output wire                                          out_dist_26_if_read,
    output wire                                          out_dist_26_if_read_ce,
    output wire                                          out_dist_26_if_write,
    output wire                                          out_dist_26_if_write_ce,
    output wire                                          out_dist_26_reset,
    output wire                                          out_dist_2_clk,
    output wire [                                  65:0] out_dist_2_if_din,
    input wire  [                                  65:0] out_dist_2_if_dout,
    input wire                                           out_dist_2_if_empty_n,
    input wire                                           out_dist_2_if_full_n,
    output wire                                          out_dist_2_if_read,
    output wire                                          out_dist_2_if_read_ce,
    output wire                                          out_dist_2_if_write,
    output wire                                          out_dist_2_if_write_ce,
    output wire                                          out_dist_2_reset,
    output wire                                          out_dist_3_clk,
    output wire [                                  65:0] out_dist_3_if_din,
    input wire  [                                  65:0] out_dist_3_if_dout,
    input wire                                           out_dist_3_if_empty_n,
    input wire                                           out_dist_3_if_full_n,
    output wire                                          out_dist_3_if_read,
    output wire                                          out_dist_3_if_read_ce,
    output wire                                          out_dist_3_if_write,
    output wire                                          out_dist_3_if_write_ce,
    output wire                                          out_dist_3_reset,
    output wire                                          out_dist_4_clk,
    output wire [                                  65:0] out_dist_4_if_din,
    input wire  [                                  65:0] out_dist_4_if_dout,
    input wire                                           out_dist_4_if_empty_n,
    input wire                                           out_dist_4_if_full_n,
    output wire                                          out_dist_4_if_read,
    output wire                                          out_dist_4_if_read_ce,
    output wire                                          out_dist_4_if_write,
    output wire                                          out_dist_4_if_write_ce,
    output wire                                          out_dist_4_reset,
    output wire                                          out_dist_5_clk,
    output wire [                                  65:0] out_dist_5_if_din,
    input wire  [                                  65:0] out_dist_5_if_dout,
    input wire                                           out_dist_5_if_empty_n,
    input wire                                           out_dist_5_if_full_n,
    output wire                                          out_dist_5_if_read,
    output wire                                          out_dist_5_if_read_ce,
    output wire                                          out_dist_5_if_write,
    output wire                                          out_dist_5_if_write_ce,
    output wire                                          out_dist_5_reset,
    output wire                                          out_dist_6_clk,
    output wire [                                  65:0] out_dist_6_if_din,
    input wire  [                                  65:0] out_dist_6_if_dout,
    input wire                                           out_dist_6_if_empty_n,
    input wire                                           out_dist_6_if_full_n,
    output wire                                          out_dist_6_if_read,
    output wire                                          out_dist_6_if_read_ce,
    output wire                                          out_dist_6_if_write,
    output wire                                          out_dist_6_if_write_ce,
    output wire                                          out_dist_6_reset,
    output wire                                          out_dist_7_clk,
    output wire [                                  65:0] out_dist_7_if_din,
    input wire  [                                  65:0] out_dist_7_if_dout,
    input wire                                           out_dist_7_if_empty_n,
    input wire                                           out_dist_7_if_full_n,
    output wire                                          out_dist_7_if_read,
    output wire                                          out_dist_7_if_read_ce,
    output wire                                          out_dist_7_if_write,
    output wire                                          out_dist_7_if_write_ce,
    output wire                                          out_dist_7_reset,
    output wire                                          out_dist_8_clk,
    output wire [                                  65:0] out_dist_8_if_din,
    input wire  [                                  65:0] out_dist_8_if_dout,
    input wire                                           out_dist_8_if_empty_n,
    input wire                                           out_dist_8_if_full_n,
    output wire                                          out_dist_8_if_read,
    output wire                                          out_dist_8_if_read_ce,
    output wire                                          out_dist_8_if_write,
    output wire                                          out_dist_8_if_write_ce,
    output wire                                          out_dist_8_reset,
    output wire                                          out_dist_9_clk,
    output wire [                                  65:0] out_dist_9_if_din,
    input wire  [                                  65:0] out_dist_9_if_dout,
    input wire                                           out_dist_9_if_empty_n,
    input wire                                           out_dist_9_if_full_n,
    output wire                                          out_dist_9_if_read,
    output wire                                          out_dist_9_if_read_ce,
    output wire                                          out_dist_9_if_write,
    output wire                                          out_dist_9_if_write_ce,
    output wire                                          out_dist_9_reset,
    output wire                                          out_id_0_clk,
    output wire [                                  65:0] out_id_0_if_din,
    input wire  [                                  65:0] out_id_0_if_dout,
    input wire                                           out_id_0_if_empty_n,
    input wire                                           out_id_0_if_full_n,
    output wire                                          out_id_0_if_read,
    output wire                                          out_id_0_if_read_ce,
    output wire                                          out_id_0_if_write,
    output wire                                          out_id_0_if_write_ce,
    output wire                                          out_id_0_reset,
    output wire                                          out_id_10_clk,
    output wire [                                  65:0] out_id_10_if_din,
    input wire  [                                  65:0] out_id_10_if_dout,
    input wire                                           out_id_10_if_empty_n,
    input wire                                           out_id_10_if_full_n,
    output wire                                          out_id_10_if_read,
    output wire                                          out_id_10_if_read_ce,
    output wire                                          out_id_10_if_write,
    output wire                                          out_id_10_if_write_ce,
    output wire                                          out_id_10_reset,
    output wire                                          out_id_11_clk,
    output wire [                                  65:0] out_id_11_if_din,
    input wire  [                                  65:0] out_id_11_if_dout,
    input wire                                           out_id_11_if_empty_n,
    input wire                                           out_id_11_if_full_n,
    output wire                                          out_id_11_if_read,
    output wire                                          out_id_11_if_read_ce,
    output wire                                          out_id_11_if_write,
    output wire                                          out_id_11_if_write_ce,
    output wire                                          out_id_11_reset,
    output wire                                          out_id_12_clk,
    output wire [                                  65:0] out_id_12_if_din,
    input wire  [                                  65:0] out_id_12_if_dout,
    input wire                                           out_id_12_if_empty_n,
    input wire                                           out_id_12_if_full_n,
    output wire                                          out_id_12_if_read,
    output wire                                          out_id_12_if_read_ce,
    output wire                                          out_id_12_if_write,
    output wire                                          out_id_12_if_write_ce,
    output wire                                          out_id_12_reset,
    output wire                                          out_id_13_clk,
    output wire [                                  65:0] out_id_13_if_din,
    input wire  [                                  65:0] out_id_13_if_dout,
    input wire                                           out_id_13_if_empty_n,
    input wire                                           out_id_13_if_full_n,
    output wire                                          out_id_13_if_read,
    output wire                                          out_id_13_if_read_ce,
    output wire                                          out_id_13_if_write,
    output wire                                          out_id_13_if_write_ce,
    output wire                                          out_id_13_reset,
    output wire                                          out_id_14_clk,
    output wire [                                  65:0] out_id_14_if_din,
    input wire  [                                  65:0] out_id_14_if_dout,
    input wire                                           out_id_14_if_empty_n,
    input wire                                           out_id_14_if_full_n,
    output wire                                          out_id_14_if_read,
    output wire                                          out_id_14_if_read_ce,
    output wire                                          out_id_14_if_write,
    output wire                                          out_id_14_if_write_ce,
    output wire                                          out_id_14_reset,
    output wire                                          out_id_15_clk,
    output wire [                                  65:0] out_id_15_if_din,
    input wire  [                                  65:0] out_id_15_if_dout,
    input wire                                           out_id_15_if_empty_n,
    input wire                                           out_id_15_if_full_n,
    output wire                                          out_id_15_if_read,
    output wire                                          out_id_15_if_read_ce,
    output wire                                          out_id_15_if_write,
    output wire                                          out_id_15_if_write_ce,
    output wire                                          out_id_15_reset,
    output wire                                          out_id_16_clk,
    output wire [                                  65:0] out_id_16_if_din,
    input wire  [                                  65:0] out_id_16_if_dout,
    input wire                                           out_id_16_if_empty_n,
    input wire                                           out_id_16_if_full_n,
    output wire                                          out_id_16_if_read,
    output wire                                          out_id_16_if_read_ce,
    output wire                                          out_id_16_if_write,
    output wire                                          out_id_16_if_write_ce,
    output wire                                          out_id_16_reset,
    output wire                                          out_id_17_clk,
    output wire [                                  65:0] out_id_17_if_din,
    input wire  [                                  65:0] out_id_17_if_dout,
    input wire                                           out_id_17_if_empty_n,
    input wire                                           out_id_17_if_full_n,
    output wire                                          out_id_17_if_read,
    output wire                                          out_id_17_if_read_ce,
    output wire                                          out_id_17_if_write,
    output wire                                          out_id_17_if_write_ce,
    output wire                                          out_id_17_reset,
    output wire                                          out_id_18_clk,
    output wire [                                  65:0] out_id_18_if_din,
    input wire  [                                  65:0] out_id_18_if_dout,
    input wire                                           out_id_18_if_empty_n,
    input wire                                           out_id_18_if_full_n,
    output wire                                          out_id_18_if_read,
    output wire                                          out_id_18_if_read_ce,
    output wire                                          out_id_18_if_write,
    output wire                                          out_id_18_if_write_ce,
    output wire                                          out_id_18_reset,
    output wire                                          out_id_19_clk,
    output wire [                                  65:0] out_id_19_if_din,
    input wire  [                                  65:0] out_id_19_if_dout,
    input wire                                           out_id_19_if_empty_n,
    input wire                                           out_id_19_if_full_n,
    output wire                                          out_id_19_if_read,
    output wire                                          out_id_19_if_read_ce,
    output wire                                          out_id_19_if_write,
    output wire                                          out_id_19_if_write_ce,
    output wire                                          out_id_19_reset,
    output wire                                          out_id_1_clk,
    output wire [                                  65:0] out_id_1_if_din,
    input wire  [                                  65:0] out_id_1_if_dout,
    input wire                                           out_id_1_if_empty_n,
    input wire                                           out_id_1_if_full_n,
    output wire                                          out_id_1_if_read,
    output wire                                          out_id_1_if_read_ce,
    output wire                                          out_id_1_if_write,
    output wire                                          out_id_1_if_write_ce,
    output wire                                          out_id_1_reset,
    output wire                                          out_id_20_clk,
    output wire [                                  65:0] out_id_20_if_din,
    input wire  [                                  65:0] out_id_20_if_dout,
    input wire                                           out_id_20_if_empty_n,
    input wire                                           out_id_20_if_full_n,
    output wire                                          out_id_20_if_read,
    output wire                                          out_id_20_if_read_ce,
    output wire                                          out_id_20_if_write,
    output wire                                          out_id_20_if_write_ce,
    output wire                                          out_id_20_reset,
    output wire                                          out_id_21_clk,
    output wire [                                  65:0] out_id_21_if_din,
    input wire  [                                  65:0] out_id_21_if_dout,
    input wire                                           out_id_21_if_empty_n,
    input wire                                           out_id_21_if_full_n,
    output wire                                          out_id_21_if_read,
    output wire                                          out_id_21_if_read_ce,
    output wire                                          out_id_21_if_write,
    output wire                                          out_id_21_if_write_ce,
    output wire                                          out_id_21_reset,
    output wire                                          out_id_22_clk,
    output wire [                                  65:0] out_id_22_if_din,
    input wire  [                                  65:0] out_id_22_if_dout,
    input wire                                           out_id_22_if_empty_n,
    input wire                                           out_id_22_if_full_n,
    output wire                                          out_id_22_if_read,
    output wire                                          out_id_22_if_read_ce,
    output wire                                          out_id_22_if_write,
    output wire                                          out_id_22_if_write_ce,
    output wire                                          out_id_22_reset,
    output wire                                          out_id_23_clk,
    output wire [                                  65:0] out_id_23_if_din,
    input wire  [                                  65:0] out_id_23_if_dout,
    input wire                                           out_id_23_if_empty_n,
    input wire                                           out_id_23_if_full_n,
    output wire                                          out_id_23_if_read,
    output wire                                          out_id_23_if_read_ce,
    output wire                                          out_id_23_if_write,
    output wire                                          out_id_23_if_write_ce,
    output wire                                          out_id_23_reset,
    output wire                                          out_id_24_clk,
    output wire [                                  65:0] out_id_24_if_din,
    input wire  [                                  65:0] out_id_24_if_dout,
    input wire                                           out_id_24_if_empty_n,
    input wire                                           out_id_24_if_full_n,
    output wire                                          out_id_24_if_read,
    output wire                                          out_id_24_if_read_ce,
    output wire                                          out_id_24_if_write,
    output wire                                          out_id_24_if_write_ce,
    output wire                                          out_id_24_reset,
    output wire                                          out_id_25_clk,
    output wire [                                  65:0] out_id_25_if_din,
    input wire  [                                  65:0] out_id_25_if_dout,
    input wire                                           out_id_25_if_empty_n,
    input wire                                           out_id_25_if_full_n,
    output wire                                          out_id_25_if_read,
    output wire                                          out_id_25_if_read_ce,
    output wire                                          out_id_25_if_write,
    output wire                                          out_id_25_if_write_ce,
    output wire                                          out_id_25_reset,
    output wire                                          out_id_26_clk,
    output wire [                                  65:0] out_id_26_if_din,
    input wire  [                                  65:0] out_id_26_if_dout,
    input wire                                           out_id_26_if_empty_n,
    input wire                                           out_id_26_if_full_n,
    output wire                                          out_id_26_if_read,
    output wire                                          out_id_26_if_read_ce,
    output wire                                          out_id_26_if_write,
    output wire                                          out_id_26_if_write_ce,
    output wire                                          out_id_26_reset,
    output wire                                          out_id_2_clk,
    output wire [                                  65:0] out_id_2_if_din,
    input wire  [                                  65:0] out_id_2_if_dout,
    input wire                                           out_id_2_if_empty_n,
    input wire                                           out_id_2_if_full_n,
    output wire                                          out_id_2_if_read,
    output wire                                          out_id_2_if_read_ce,
    output wire                                          out_id_2_if_write,
    output wire                                          out_id_2_if_write_ce,
    output wire                                          out_id_2_reset,
    output wire                                          out_id_3_clk,
    output wire [                                  65:0] out_id_3_if_din,
    input wire  [                                  65:0] out_id_3_if_dout,
    input wire                                           out_id_3_if_empty_n,
    input wire                                           out_id_3_if_full_n,
    output wire                                          out_id_3_if_read,
    output wire                                          out_id_3_if_read_ce,
    output wire                                          out_id_3_if_write,
    output wire                                          out_id_3_if_write_ce,
    output wire                                          out_id_3_reset,
    output wire                                          out_id_4_clk,
    output wire [                                  65:0] out_id_4_if_din,
    input wire  [                                  65:0] out_id_4_if_dout,
    input wire                                           out_id_4_if_empty_n,
    input wire                                           out_id_4_if_full_n,
    output wire                                          out_id_4_if_read,
    output wire                                          out_id_4_if_read_ce,
    output wire                                          out_id_4_if_write,
    output wire                                          out_id_4_if_write_ce,
    output wire                                          out_id_4_reset,
    output wire                                          out_id_5_clk,
    output wire [                                  65:0] out_id_5_if_din,
    input wire  [                                  65:0] out_id_5_if_dout,
    input wire                                           out_id_5_if_empty_n,
    input wire                                           out_id_5_if_full_n,
    output wire                                          out_id_5_if_read,
    output wire                                          out_id_5_if_read_ce,
    output wire                                          out_id_5_if_write,
    output wire                                          out_id_5_if_write_ce,
    output wire                                          out_id_5_reset,
    output wire                                          out_id_6_clk,
    output wire [                                  65:0] out_id_6_if_din,
    input wire  [                                  65:0] out_id_6_if_dout,
    input wire                                           out_id_6_if_empty_n,
    input wire                                           out_id_6_if_full_n,
    output wire                                          out_id_6_if_read,
    output wire                                          out_id_6_if_read_ce,
    output wire                                          out_id_6_if_write,
    output wire                                          out_id_6_if_write_ce,
    output wire                                          out_id_6_reset,
    output wire                                          out_id_7_clk,
    output wire [                                  65:0] out_id_7_if_din,
    input wire  [                                  65:0] out_id_7_if_dout,
    input wire                                           out_id_7_if_empty_n,
    input wire                                           out_id_7_if_full_n,
    output wire                                          out_id_7_if_read,
    output wire                                          out_id_7_if_read_ce,
    output wire                                          out_id_7_if_write,
    output wire                                          out_id_7_if_write_ce,
    output wire                                          out_id_7_reset,
    output wire                                          out_id_8_clk,
    output wire [                                  65:0] out_id_8_if_din,
    input wire  [                                  65:0] out_id_8_if_dout,
    input wire                                           out_id_8_if_empty_n,
    input wire                                           out_id_8_if_full_n,
    output wire                                          out_id_8_if_read,
    output wire                                          out_id_8_if_read_ce,
    output wire                                          out_id_8_if_write,
    output wire                                          out_id_8_if_write_ce,
    output wire                                          out_id_8_reset,
    output wire                                          out_id_9_clk,
    output wire [                                  65:0] out_id_9_if_din,
    input wire  [                                  65:0] out_id_9_if_dout,
    input wire                                           out_id_9_if_empty_n,
    input wire                                           out_id_9_if_full_n,
    output wire                                          out_id_9_if_read,
    output wire                                          out_id_9_if_read_ce,
    output wire                                          out_id_9_if_write,
    output wire                                          out_id_9_if_write_ce,
    output wire                                          out_id_9_reset,
    output wire                                          krnl_globalSort_L1_L2_0_ap_clk,
    input wire                                           krnl_globalSort_L1_L2_0_ap_done,
    input wire                                           krnl_globalSort_L1_L2_0_ap_idle,
    input wire                                           krnl_globalSort_L1_L2_0_ap_ready,
    output wire                                          krnl_globalSort_L1_L2_0_ap_rst_n,
    output wire                                          krnl_globalSort_L1_L2_0_ap_start,
    output wire [                                  65:0] krnl_globalSort_L1_L2_0_in_dist0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_0_in_dist0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_0_in_dist0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_0_in_dist0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_0_in_dist0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_0_in_dist0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_0_in_dist1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_0_in_dist1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_0_in_dist1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_0_in_dist1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_0_in_dist1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_0_in_dist1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_0_in_dist2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_0_in_dist2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_0_in_dist2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_0_in_dist2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_0_in_dist2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_0_in_dist2_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_0_in_id0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_0_in_id0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_0_in_id0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_0_in_id0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_0_in_id0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_0_in_id0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_0_in_id1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_0_in_id1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_0_in_id1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_0_in_id1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_0_in_id1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_0_in_id1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_0_in_id2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_0_in_id2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_0_in_id2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_0_in_id2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_0_in_id2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_0_in_id2_s_read,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_0_out_dist_din,
    output wire                                          krnl_globalSort_L1_L2_0_out_dist_full_n,
    input wire                                           krnl_globalSort_L1_L2_0_out_dist_write,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_0_out_id_din,
    output wire                                          krnl_globalSort_L1_L2_0_out_id_full_n,
    input wire                                           krnl_globalSort_L1_L2_0_out_id_write,
    output wire                                          krnl_globalSort_L1_L2_1_ap_clk,
    input wire                                           krnl_globalSort_L1_L2_1_ap_done,
    input wire                                           krnl_globalSort_L1_L2_1_ap_idle,
    input wire                                           krnl_globalSort_L1_L2_1_ap_ready,
    output wire                                          krnl_globalSort_L1_L2_1_ap_rst_n,
    output wire                                          krnl_globalSort_L1_L2_1_ap_start,
    output wire [                                  65:0] krnl_globalSort_L1_L2_1_in_dist0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_1_in_dist0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_1_in_dist0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_1_in_dist0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_1_in_dist0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_1_in_dist0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_1_in_dist1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_1_in_dist1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_1_in_dist1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_1_in_dist1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_1_in_dist1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_1_in_dist1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_1_in_dist2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_1_in_dist2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_1_in_dist2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_1_in_dist2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_1_in_dist2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_1_in_dist2_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_1_in_id0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_1_in_id0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_1_in_id0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_1_in_id0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_1_in_id0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_1_in_id0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_1_in_id1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_1_in_id1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_1_in_id1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_1_in_id1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_1_in_id1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_1_in_id1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_1_in_id2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_1_in_id2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_1_in_id2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_1_in_id2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_1_in_id2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_1_in_id2_s_read,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_1_out_dist_din,
    output wire                                          krnl_globalSort_L1_L2_1_out_dist_full_n,
    input wire                                           krnl_globalSort_L1_L2_1_out_dist_write,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_1_out_id_din,
    output wire                                          krnl_globalSort_L1_L2_1_out_id_full_n,
    input wire                                           krnl_globalSort_L1_L2_1_out_id_write,
    output wire                                          krnl_globalSort_L1_L2_2_ap_clk,
    input wire                                           krnl_globalSort_L1_L2_2_ap_done,
    input wire                                           krnl_globalSort_L1_L2_2_ap_idle,
    input wire                                           krnl_globalSort_L1_L2_2_ap_ready,
    output wire                                          krnl_globalSort_L1_L2_2_ap_rst_n,
    output wire                                          krnl_globalSort_L1_L2_2_ap_start,
    output wire [                                  65:0] krnl_globalSort_L1_L2_2_in_dist0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_2_in_dist0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_2_in_dist0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_2_in_dist0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_2_in_dist0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_2_in_dist0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_2_in_dist1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_2_in_dist1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_2_in_dist1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_2_in_dist1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_2_in_dist1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_2_in_dist1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_2_in_dist2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_2_in_dist2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_2_in_dist2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_2_in_dist2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_2_in_dist2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_2_in_dist2_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_2_in_id0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_2_in_id0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_2_in_id0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_2_in_id0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_2_in_id0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_2_in_id0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_2_in_id1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_2_in_id1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_2_in_id1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_2_in_id1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_2_in_id1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_2_in_id1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_2_in_id2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_2_in_id2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_2_in_id2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_2_in_id2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_2_in_id2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_2_in_id2_s_read,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_2_out_dist_din,
    output wire                                          krnl_globalSort_L1_L2_2_out_dist_full_n,
    input wire                                           krnl_globalSort_L1_L2_2_out_dist_write,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_2_out_id_din,
    output wire                                          krnl_globalSort_L1_L2_2_out_id_full_n,
    input wire                                           krnl_globalSort_L1_L2_2_out_id_write,
    output wire                                          krnl_globalSort_L1_L2_3_ap_clk,
    input wire                                           krnl_globalSort_L1_L2_3_ap_done,
    input wire                                           krnl_globalSort_L1_L2_3_ap_idle,
    input wire                                           krnl_globalSort_L1_L2_3_ap_ready,
    output wire                                          krnl_globalSort_L1_L2_3_ap_rst_n,
    output wire                                          krnl_globalSort_L1_L2_3_ap_start,
    output wire [                                  65:0] krnl_globalSort_L1_L2_3_in_dist0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_3_in_dist0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_3_in_dist0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_3_in_dist0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_3_in_dist0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_3_in_dist0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_3_in_dist1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_3_in_dist1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_3_in_dist1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_3_in_dist1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_3_in_dist1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_3_in_dist1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_3_in_dist2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_3_in_dist2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_3_in_dist2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_3_in_dist2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_3_in_dist2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_3_in_dist2_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_3_in_id0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_3_in_id0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_3_in_id0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_3_in_id0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_3_in_id0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_3_in_id0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_3_in_id1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_3_in_id1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_3_in_id1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_3_in_id1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_3_in_id1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_3_in_id1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_3_in_id2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_3_in_id2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_3_in_id2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_3_in_id2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_3_in_id2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_3_in_id2_s_read,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_3_out_dist_din,
    output wire                                          krnl_globalSort_L1_L2_3_out_dist_full_n,
    input wire                                           krnl_globalSort_L1_L2_3_out_dist_write,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_3_out_id_din,
    output wire                                          krnl_globalSort_L1_L2_3_out_id_full_n,
    input wire                                           krnl_globalSort_L1_L2_3_out_id_write,
    output wire                                          krnl_globalSort_L1_L2_4_ap_clk,
    input wire                                           krnl_globalSort_L1_L2_4_ap_done,
    input wire                                           krnl_globalSort_L1_L2_4_ap_idle,
    input wire                                           krnl_globalSort_L1_L2_4_ap_ready,
    output wire                                          krnl_globalSort_L1_L2_4_ap_rst_n,
    output wire                                          krnl_globalSort_L1_L2_4_ap_start,
    output wire [                                  65:0] krnl_globalSort_L1_L2_4_in_dist0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_4_in_dist0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_4_in_dist0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_4_in_dist0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_4_in_dist0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_4_in_dist0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_4_in_dist1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_4_in_dist1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_4_in_dist1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_4_in_dist1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_4_in_dist1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_4_in_dist1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_4_in_dist2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_4_in_dist2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_4_in_dist2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_4_in_dist2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_4_in_dist2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_4_in_dist2_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_4_in_id0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_4_in_id0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_4_in_id0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_4_in_id0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_4_in_id0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_4_in_id0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_4_in_id1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_4_in_id1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_4_in_id1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_4_in_id1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_4_in_id1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_4_in_id1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_4_in_id2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_4_in_id2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_4_in_id2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_4_in_id2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_4_in_id2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_4_in_id2_s_read,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_4_out_dist_din,
    output wire                                          krnl_globalSort_L1_L2_4_out_dist_full_n,
    input wire                                           krnl_globalSort_L1_L2_4_out_dist_write,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_4_out_id_din,
    output wire                                          krnl_globalSort_L1_L2_4_out_id_full_n,
    input wire                                           krnl_globalSort_L1_L2_4_out_id_write,
    output wire                                          krnl_globalSort_L1_L2_5_ap_clk,
    input wire                                           krnl_globalSort_L1_L2_5_ap_done,
    input wire                                           krnl_globalSort_L1_L2_5_ap_idle,
    input wire                                           krnl_globalSort_L1_L2_5_ap_ready,
    output wire                                          krnl_globalSort_L1_L2_5_ap_rst_n,
    output wire                                          krnl_globalSort_L1_L2_5_ap_start,
    output wire [                                  65:0] krnl_globalSort_L1_L2_5_in_dist0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_5_in_dist0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_5_in_dist0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_5_in_dist0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_5_in_dist0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_5_in_dist0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_5_in_dist1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_5_in_dist1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_5_in_dist1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_5_in_dist1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_5_in_dist1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_5_in_dist1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_5_in_dist2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_5_in_dist2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_5_in_dist2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_5_in_dist2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_5_in_dist2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_5_in_dist2_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_5_in_id0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_5_in_id0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_5_in_id0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_5_in_id0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_5_in_id0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_5_in_id0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_5_in_id1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_5_in_id1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_5_in_id1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_5_in_id1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_5_in_id1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_5_in_id1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_5_in_id2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_5_in_id2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_5_in_id2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_5_in_id2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_5_in_id2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_5_in_id2_s_read,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_5_out_dist_din,
    output wire                                          krnl_globalSort_L1_L2_5_out_dist_full_n,
    input wire                                           krnl_globalSort_L1_L2_5_out_dist_write,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_5_out_id_din,
    output wire                                          krnl_globalSort_L1_L2_5_out_id_full_n,
    input wire                                           krnl_globalSort_L1_L2_5_out_id_write,
    output wire                                          krnl_globalSort_L1_L2_6_ap_clk,
    input wire                                           krnl_globalSort_L1_L2_6_ap_done,
    input wire                                           krnl_globalSort_L1_L2_6_ap_idle,
    input wire                                           krnl_globalSort_L1_L2_6_ap_ready,
    output wire                                          krnl_globalSort_L1_L2_6_ap_rst_n,
    output wire                                          krnl_globalSort_L1_L2_6_ap_start,
    output wire [                                  65:0] krnl_globalSort_L1_L2_6_in_dist0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_6_in_dist0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_6_in_dist0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_6_in_dist0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_6_in_dist0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_6_in_dist0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_6_in_dist1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_6_in_dist1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_6_in_dist1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_6_in_dist1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_6_in_dist1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_6_in_dist1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_6_in_dist2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_6_in_dist2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_6_in_dist2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_6_in_dist2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_6_in_dist2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_6_in_dist2_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_6_in_id0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_6_in_id0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_6_in_id0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_6_in_id0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_6_in_id0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_6_in_id0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_6_in_id1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_6_in_id1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_6_in_id1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_6_in_id1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_6_in_id1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_6_in_id1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_6_in_id2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_6_in_id2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_6_in_id2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_6_in_id2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_6_in_id2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_6_in_id2_s_read,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_6_out_dist_din,
    output wire                                          krnl_globalSort_L1_L2_6_out_dist_full_n,
    input wire                                           krnl_globalSort_L1_L2_6_out_dist_write,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_6_out_id_din,
    output wire                                          krnl_globalSort_L1_L2_6_out_id_full_n,
    input wire                                           krnl_globalSort_L1_L2_6_out_id_write,
    output wire                                          krnl_globalSort_L1_L2_7_ap_clk,
    input wire                                           krnl_globalSort_L1_L2_7_ap_done,
    input wire                                           krnl_globalSort_L1_L2_7_ap_idle,
    input wire                                           krnl_globalSort_L1_L2_7_ap_ready,
    output wire                                          krnl_globalSort_L1_L2_7_ap_rst_n,
    output wire                                          krnl_globalSort_L1_L2_7_ap_start,
    output wire [                                  65:0] krnl_globalSort_L1_L2_7_in_dist0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_7_in_dist0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_7_in_dist0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_7_in_dist0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_7_in_dist0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_7_in_dist0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_7_in_dist1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_7_in_dist1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_7_in_dist1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_7_in_dist1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_7_in_dist1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_7_in_dist1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_7_in_dist2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_7_in_dist2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_7_in_dist2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_7_in_dist2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_7_in_dist2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_7_in_dist2_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_7_in_id0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_7_in_id0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_7_in_id0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_7_in_id0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_7_in_id0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_7_in_id0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_7_in_id1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_7_in_id1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_7_in_id1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_7_in_id1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_7_in_id1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_7_in_id1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_7_in_id2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_7_in_id2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_7_in_id2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_7_in_id2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_7_in_id2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_7_in_id2_s_read,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_7_out_dist_din,
    output wire                                          krnl_globalSort_L1_L2_7_out_dist_full_n,
    input wire                                           krnl_globalSort_L1_L2_7_out_dist_write,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_7_out_id_din,
    output wire                                          krnl_globalSort_L1_L2_7_out_id_full_n,
    input wire                                           krnl_globalSort_L1_L2_7_out_id_write,
    output wire                                          krnl_globalSort_L1_L2_8_ap_clk,
    input wire                                           krnl_globalSort_L1_L2_8_ap_done,
    input wire                                           krnl_globalSort_L1_L2_8_ap_idle,
    input wire                                           krnl_globalSort_L1_L2_8_ap_ready,
    output wire                                          krnl_globalSort_L1_L2_8_ap_rst_n,
    output wire                                          krnl_globalSort_L1_L2_8_ap_start,
    output wire [                                  65:0] krnl_globalSort_L1_L2_8_in_dist0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_8_in_dist0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_8_in_dist0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_8_in_dist0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_8_in_dist0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_8_in_dist0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_8_in_dist1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_8_in_dist1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_8_in_dist1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_8_in_dist1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_8_in_dist1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_8_in_dist1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_8_in_dist2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_8_in_dist2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_8_in_dist2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_8_in_dist2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_8_in_dist2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_8_in_dist2_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_8_in_id0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_8_in_id0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_8_in_id0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_8_in_id0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_8_in_id0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_8_in_id0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_8_in_id1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_8_in_id1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_8_in_id1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_8_in_id1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_8_in_id1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_8_in_id1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_8_in_id2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_8_in_id2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_8_in_id2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_8_in_id2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_8_in_id2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_8_in_id2_s_read,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_8_out_dist_din,
    output wire                                          krnl_globalSort_L1_L2_8_out_dist_full_n,
    input wire                                           krnl_globalSort_L1_L2_8_out_dist_write,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_8_out_id_din,
    output wire                                          krnl_globalSort_L1_L2_8_out_id_full_n,
    input wire                                           krnl_globalSort_L1_L2_8_out_id_write,
    output wire                                          krnl_globalSort_L1_L2_9_ap_clk,
    input wire                                           krnl_globalSort_L1_L2_9_ap_done,
    input wire                                           krnl_globalSort_L1_L2_9_ap_idle,
    input wire                                           krnl_globalSort_L1_L2_9_ap_ready,
    output wire                                          krnl_globalSort_L1_L2_9_ap_rst_n,
    output wire                                          krnl_globalSort_L1_L2_9_ap_start,
    output wire [                                  65:0] krnl_globalSort_L1_L2_9_in_dist0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_9_in_dist0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_9_in_dist0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_9_in_dist0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_9_in_dist0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_9_in_dist0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_9_in_dist1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_9_in_dist1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_9_in_dist1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_9_in_dist1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_9_in_dist1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_9_in_dist1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_9_in_dist2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_9_in_dist2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_9_in_dist2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_9_in_dist2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_9_in_dist2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_9_in_dist2_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_9_in_id0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_9_in_id0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_9_in_id0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_9_in_id0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_9_in_id0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_9_in_id0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_9_in_id1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_9_in_id1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_9_in_id1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_9_in_id1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_9_in_id1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_9_in_id1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_9_in_id2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_9_in_id2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_9_in_id2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_9_in_id2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_9_in_id2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_9_in_id2_s_read,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_9_out_dist_din,
    output wire                                          krnl_globalSort_L1_L2_9_out_dist_full_n,
    input wire                                           krnl_globalSort_L1_L2_9_out_dist_write,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_9_out_id_din,
    output wire                                          krnl_globalSort_L1_L2_9_out_id_full_n,
    input wire                                           krnl_globalSort_L1_L2_9_out_id_write,
    output wire                                          krnl_globalSort_L1_L2_10_ap_clk,
    input wire                                           krnl_globalSort_L1_L2_10_ap_done,
    input wire                                           krnl_globalSort_L1_L2_10_ap_idle,
    input wire                                           krnl_globalSort_L1_L2_10_ap_ready,
    output wire                                          krnl_globalSort_L1_L2_10_ap_rst_n,
    output wire                                          krnl_globalSort_L1_L2_10_ap_start,
    output wire [                                  65:0] krnl_globalSort_L1_L2_10_in_dist0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_10_in_dist0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_10_in_dist0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_10_in_dist0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_10_in_dist0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_10_in_dist0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_10_in_dist1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_10_in_dist1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_10_in_dist1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_10_in_dist1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_10_in_dist1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_10_in_dist1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_10_in_dist2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_10_in_dist2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_10_in_dist2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_10_in_dist2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_10_in_dist2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_10_in_dist2_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_10_in_id0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_10_in_id0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_10_in_id0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_10_in_id0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_10_in_id0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_10_in_id0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_10_in_id1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_10_in_id1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_10_in_id1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_10_in_id1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_10_in_id1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_10_in_id1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_10_in_id2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_10_in_id2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_10_in_id2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_10_in_id2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_10_in_id2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_10_in_id2_s_read,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_10_out_dist_din,
    output wire                                          krnl_globalSort_L1_L2_10_out_dist_full_n,
    input wire                                           krnl_globalSort_L1_L2_10_out_dist_write,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_10_out_id_din,
    output wire                                          krnl_globalSort_L1_L2_10_out_id_full_n,
    input wire                                           krnl_globalSort_L1_L2_10_out_id_write,
    output wire                                          krnl_globalSort_L1_L2_11_ap_clk,
    input wire                                           krnl_globalSort_L1_L2_11_ap_done,
    input wire                                           krnl_globalSort_L1_L2_11_ap_idle,
    input wire                                           krnl_globalSort_L1_L2_11_ap_ready,
    output wire                                          krnl_globalSort_L1_L2_11_ap_rst_n,
    output wire                                          krnl_globalSort_L1_L2_11_ap_start,
    output wire [                                  65:0] krnl_globalSort_L1_L2_11_in_dist0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_11_in_dist0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_11_in_dist0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_11_in_dist0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_11_in_dist0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_11_in_dist0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_11_in_dist1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_11_in_dist1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_11_in_dist1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_11_in_dist1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_11_in_dist1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_11_in_dist1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_11_in_dist2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_11_in_dist2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_11_in_dist2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_11_in_dist2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_11_in_dist2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_11_in_dist2_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_11_in_id0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_11_in_id0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_11_in_id0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_11_in_id0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_11_in_id0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_11_in_id0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_11_in_id1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_11_in_id1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_11_in_id1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_11_in_id1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_11_in_id1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_11_in_id1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_11_in_id2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_11_in_id2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_11_in_id2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_11_in_id2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_11_in_id2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_11_in_id2_s_read,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_11_out_dist_din,
    output wire                                          krnl_globalSort_L1_L2_11_out_dist_full_n,
    input wire                                           krnl_globalSort_L1_L2_11_out_dist_write,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_11_out_id_din,
    output wire                                          krnl_globalSort_L1_L2_11_out_id_full_n,
    input wire                                           krnl_globalSort_L1_L2_11_out_id_write,
    output wire                                          krnl_globalSort_L1_L2_12_ap_clk,
    input wire                                           krnl_globalSort_L1_L2_12_ap_done,
    input wire                                           krnl_globalSort_L1_L2_12_ap_idle,
    input wire                                           krnl_globalSort_L1_L2_12_ap_ready,
    output wire                                          krnl_globalSort_L1_L2_12_ap_rst_n,
    output wire                                          krnl_globalSort_L1_L2_12_ap_start,
    output wire [                                  65:0] krnl_globalSort_L1_L2_12_in_dist0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_12_in_dist0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_12_in_dist0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_12_in_dist0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_12_in_dist0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_12_in_dist0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_12_in_dist1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_12_in_dist1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_12_in_dist1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_12_in_dist1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_12_in_dist1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_12_in_dist1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_12_in_dist2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_12_in_dist2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_12_in_dist2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_12_in_dist2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_12_in_dist2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_12_in_dist2_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_12_in_id0_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_12_in_id0_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_12_in_id0_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_12_in_id0_s_dout,
    output wire                                          krnl_globalSort_L1_L2_12_in_id0_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_12_in_id0_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_12_in_id1_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_12_in_id1_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_12_in_id1_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_12_in_id1_s_dout,
    output wire                                          krnl_globalSort_L1_L2_12_in_id1_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_12_in_id1_s_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_12_in_id2_peek_dout,
    output wire                                          krnl_globalSort_L1_L2_12_in_id2_peek_empty_n,
    input wire                                           krnl_globalSort_L1_L2_12_in_id2_peek_read,
    output wire [                                  65:0] krnl_globalSort_L1_L2_12_in_id2_s_dout,
    output wire                                          krnl_globalSort_L1_L2_12_in_id2_s_empty_n,
    input wire                                           krnl_globalSort_L1_L2_12_in_id2_s_read,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_12_out_dist_din,
    output wire                                          krnl_globalSort_L1_L2_12_out_dist_full_n,
    input wire                                           krnl_globalSort_L1_L2_12_out_dist_write,
    input wire  [                                  65:0] krnl_globalSort_L1_L2_12_out_id_din,
    output wire                                          krnl_globalSort_L1_L2_12_out_id_full_n,
    input wire                                           krnl_globalSort_L1_L2_12_out_id_write,
    output wire                                          krnl_output_dist_id_0_ap_clk,
    input wire                                           krnl_output_dist_id_0_ap_done,
    input wire                                           krnl_output_dist_id_0_ap_idle,
    input wire                                           krnl_output_dist_id_0_ap_ready,
    output wire                                          krnl_output_dist_id_0_ap_rst_n,
    output wire                                          krnl_output_dist_id_0_ap_start,
    output wire [                                  65:0] krnl_output_dist_id_0_in_dist_peek_dout,
    output wire                                          krnl_output_dist_id_0_in_dist_peek_empty_n,
    input wire                                           krnl_output_dist_id_0_in_dist_peek_read,
    output wire [                                  65:0] krnl_output_dist_id_0_in_dist_s_dout,
    output wire                                          krnl_output_dist_id_0_in_dist_s_empty_n,
    input wire                                           krnl_output_dist_id_0_in_dist_s_read,
    output wire [                                  65:0] krnl_output_dist_id_0_in_id_peek_dout,
    output wire                                          krnl_output_dist_id_0_in_id_peek_empty_n,
    input wire                                           krnl_output_dist_id_0_in_id_peek_read,
    output wire [                                  65:0] krnl_output_dist_id_0_in_id_s_dout,
    output wire                                          krnl_output_dist_id_0_in_id_s_empty_n,
    input wire                                           krnl_output_dist_id_0_in_id_s_read,
    output wire [                                  63:0] krnl_output_dist_id_0_output_knnDist_read_addr_offset,
    input wire  [                                  63:0] krnl_output_dist_id_0_output_knnDist_read_addr_s_din,
    output wire                                          krnl_output_dist_id_0_output_knnDist_read_addr_s_full_n,
    input wire                                           krnl_output_dist_id_0_output_knnDist_read_addr_s_write,
    output wire [                                  32:0] krnl_output_dist_id_0_output_knnDist_read_data_peek_dout,
    output wire                                          krnl_output_dist_id_0_output_knnDist_read_data_peek_empty_n,
    input wire                                           krnl_output_dist_id_0_output_knnDist_read_data_peek_read,
    output wire [                                  32:0] krnl_output_dist_id_0_output_knnDist_read_data_s_dout,
    output wire                                          krnl_output_dist_id_0_output_knnDist_read_data_s_empty_n,
    input wire                                           krnl_output_dist_id_0_output_knnDist_read_data_s_read,
    output wire [                                  63:0] krnl_output_dist_id_0_output_knnDist_write_addr_offset,
    input wire  [                                  63:0] krnl_output_dist_id_0_output_knnDist_write_addr_s_din,
    output wire                                          krnl_output_dist_id_0_output_knnDist_write_addr_s_full_n,
    input wire                                           krnl_output_dist_id_0_output_knnDist_write_addr_s_write,
    input wire  [                                  32:0] krnl_output_dist_id_0_output_knnDist_write_data_din,
    output wire                                          krnl_output_dist_id_0_output_knnDist_write_data_full_n,
    input wire                                           krnl_output_dist_id_0_output_knnDist_write_data_write,
    output wire [                                   8:0] krnl_output_dist_id_0_output_knnDist_write_resp_peek_dout,
    output wire                                          krnl_output_dist_id_0_output_knnDist_write_resp_peek_empty_n,
    input wire                                           krnl_output_dist_id_0_output_knnDist_write_resp_peek_read,
    output wire [                                   8:0] krnl_output_dist_id_0_output_knnDist_write_resp_s_dout,
    output wire                                          krnl_output_dist_id_0_output_knnDist_write_resp_s_empty_n,
    input wire                                           krnl_output_dist_id_0_output_knnDist_write_resp_s_read,
    output wire [                                  63:0] krnl_output_dist_id_0_output_knnId_read_addr_offset,
    input wire  [                                  63:0] krnl_output_dist_id_0_output_knnId_read_addr_s_din,
    output wire                                          krnl_output_dist_id_0_output_knnId_read_addr_s_full_n,
    input wire                                           krnl_output_dist_id_0_output_knnId_read_addr_s_write,
    output wire [                                  32:0] krnl_output_dist_id_0_output_knnId_read_data_peek_dout,
    output wire                                          krnl_output_dist_id_0_output_knnId_read_data_peek_empty_n,
    input wire                                           krnl_output_dist_id_0_output_knnId_read_data_peek_read,
    output wire [                                  32:0] krnl_output_dist_id_0_output_knnId_read_data_s_dout,
    output wire                                          krnl_output_dist_id_0_output_knnId_read_data_s_empty_n,
    input wire                                           krnl_output_dist_id_0_output_knnId_read_data_s_read,
    output wire [                                  63:0] krnl_output_dist_id_0_output_knnId_write_addr_offset,
    input wire  [                                  63:0] krnl_output_dist_id_0_output_knnId_write_addr_s_din,
    output wire                                          krnl_output_dist_id_0_output_knnId_write_addr_s_full_n,
    input wire                                           krnl_output_dist_id_0_output_knnId_write_addr_s_write,
    input wire  [                                  32:0] krnl_output_dist_id_0_output_knnId_write_data_din,
    output wire                                          krnl_output_dist_id_0_output_knnId_write_data_full_n,
    input wire                                           krnl_output_dist_id_0_output_knnId_write_data_write,
    output wire [                                   8:0] krnl_output_dist_id_0_output_knnId_write_resp_peek_dout,
    output wire                                          krnl_output_dist_id_0_output_knnId_write_resp_peek_empty_n,
    input wire                                           krnl_output_dist_id_0_output_knnId_write_resp_peek_read,
    output wire [                                   8:0] krnl_output_dist_id_0_output_knnId_write_resp_s_dout,
    output wire                                          krnl_output_dist_id_0_output_knnId_write_resp_s_empty_n,
    input wire                                           krnl_output_dist_id_0_output_knnId_write_resp_s_read,
    output wire                                          krnl_partialKnn_wrapper_0_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_0_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_0_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_0_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_0_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_0_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_0_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_0_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_0_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_0_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_0_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_0_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_0_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_0_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_0_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_0_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_0_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_0_0_searchSpace_0_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_0_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_0_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_0_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_0_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_0_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_0_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_0_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_0_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_0_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_0_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_0_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_0_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_0_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_0_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_0_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_0_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_0_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_0_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_1_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_1_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_1_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_1_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_1_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_1_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_1_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_1_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_1_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_1_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_1_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_1_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_1_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_1_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_1_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_1_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_1_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_1_0_searchSpace_0_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_1_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_1_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_1_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_1_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_1_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_1_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_1_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_1_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_1_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_1_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_1_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_1_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_1_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_1_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_1_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_1_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_1_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_1_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_10_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_10_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_10_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_10_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_10_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_10_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_10_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_10_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_10_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_10_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_10_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_10_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_10_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_10_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_10_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_10_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_10_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_10_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_10_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_10_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_10_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_10_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_10_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_10_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_10_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_10_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_10_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_10_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_10_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_10_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_10_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_10_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_10_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_10_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_10_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_10_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_11_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_11_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_11_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_11_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_11_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_11_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_11_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_11_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_11_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_11_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_11_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_11_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_11_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_11_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_11_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_11_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_11_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_11_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_11_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_11_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_11_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_11_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_11_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_11_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_11_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_11_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_11_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_11_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_11_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_11_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_11_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_11_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_11_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_11_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_11_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_11_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_12_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_12_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_12_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_12_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_12_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_12_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_12_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_12_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_12_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_12_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_12_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_12_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_12_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_12_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_12_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_12_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_12_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_12_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_12_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_12_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_12_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_12_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_12_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_12_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_12_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_12_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_12_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_12_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_12_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_12_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_12_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_12_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_12_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_12_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_12_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_12_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_13_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_13_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_13_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_13_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_13_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_13_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_13_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_13_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_13_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_13_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_13_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_13_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_13_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_13_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_13_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_13_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_13_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_13_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_13_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_13_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_13_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_13_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_13_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_13_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_13_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_13_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_13_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_13_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_13_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_13_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_13_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_13_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_13_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_13_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_13_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_13_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_14_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_14_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_14_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_14_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_14_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_14_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_14_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_14_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_14_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_14_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_14_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_14_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_14_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_14_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_14_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_14_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_14_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_14_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_14_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_14_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_14_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_14_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_14_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_14_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_14_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_14_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_14_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_14_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_14_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_14_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_14_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_14_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_14_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_14_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_14_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_14_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_15_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_15_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_15_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_15_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_15_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_15_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_15_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_15_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_15_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_15_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_15_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_15_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_15_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_15_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_15_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_15_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_15_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_15_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_15_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_15_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_15_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_15_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_15_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_15_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_15_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_15_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_15_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_15_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_15_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_15_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_15_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_15_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_15_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_15_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_15_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_15_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_16_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_16_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_16_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_16_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_16_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_16_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_16_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_16_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_16_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_16_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_16_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_16_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_16_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_16_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_16_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_16_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_16_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_16_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_16_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_16_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_16_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_16_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_16_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_16_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_16_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_16_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_16_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_16_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_16_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_16_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_16_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_16_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_16_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_16_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_16_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_16_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_17_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_17_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_17_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_17_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_17_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_17_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_17_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_17_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_17_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_17_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_17_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_17_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_17_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_17_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_17_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_17_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_17_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_17_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_17_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_17_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_17_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_17_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_17_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_17_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_17_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_17_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_17_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_17_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_17_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_17_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_17_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_17_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_17_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_17_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_17_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_17_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_18_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_18_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_18_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_18_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_18_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_18_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_18_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_18_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_18_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_18_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_18_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_18_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_18_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_18_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_18_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_18_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_18_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_18_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_18_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_18_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_18_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_18_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_18_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_18_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_18_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_18_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_18_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_18_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_18_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_18_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_18_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_18_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_18_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_18_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_18_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_18_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_19_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_19_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_19_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_19_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_19_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_19_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_19_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_19_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_19_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_19_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_19_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_19_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_19_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_19_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_19_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_19_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_19_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_19_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_19_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_19_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_19_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_19_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_19_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_19_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_19_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_19_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_19_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_19_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_19_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_19_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_19_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_19_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_19_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_19_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_19_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_19_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_2_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_2_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_2_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_2_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_2_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_2_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_2_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_2_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_2_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_2_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_2_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_2_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_2_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_2_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_2_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_2_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_2_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_2_0_searchSpace_0_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_2_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_2_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_2_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_2_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_2_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_2_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_2_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_2_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_2_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_2_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_2_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_2_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_2_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_2_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_2_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_2_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_2_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_2_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_20_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_20_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_20_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_20_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_20_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_20_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_20_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_20_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_20_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_20_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_20_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_20_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_20_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_20_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_20_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_20_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_20_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_20_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_20_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_20_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_20_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_20_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_20_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_20_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_20_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_20_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_20_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_20_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_20_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_20_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_20_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_20_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_20_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_20_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_20_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_20_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_21_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_21_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_21_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_21_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_21_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_21_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_21_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_21_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_21_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_21_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_21_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_21_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_21_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_21_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_21_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_21_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_21_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_21_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_21_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_21_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_21_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_21_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_21_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_21_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_21_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_21_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_21_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_21_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_21_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_21_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_21_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_21_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_21_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_21_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_21_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_21_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_22_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_22_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_22_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_22_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_22_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_22_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_22_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_22_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_22_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_22_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_22_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_22_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_22_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_22_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_22_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_22_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_22_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_22_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_22_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_22_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_22_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_22_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_22_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_22_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_22_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_22_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_22_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_22_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_22_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_22_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_22_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_22_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_22_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_22_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_22_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_22_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_23_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_23_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_23_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_23_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_23_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_23_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_23_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_23_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_23_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_23_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_23_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_23_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_23_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_23_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_23_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_23_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_23_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_23_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_23_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_23_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_23_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_23_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_23_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_23_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_23_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_23_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_23_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_23_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_23_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_23_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_23_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_23_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_23_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_23_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_23_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_23_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_24_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_24_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_24_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_24_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_24_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_24_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_24_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_24_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_24_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_24_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_24_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_24_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_24_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_24_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_24_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_24_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_24_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_24_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_24_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_24_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_24_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_24_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_24_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_24_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_24_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_24_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_24_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_24_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_24_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_24_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_24_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_24_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_24_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_24_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_24_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_24_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_25_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_25_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_25_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_25_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_25_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_25_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_25_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_25_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_25_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_25_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_25_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_25_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_25_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_25_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_25_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_25_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_25_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_25_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_25_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_25_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_25_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_25_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_25_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_25_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_25_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_25_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_25_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_25_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_25_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_25_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_25_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_25_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_25_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_25_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_25_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_25_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_26_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_26_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_26_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_26_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_26_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_26_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_26_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_26_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_26_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_26_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_26_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_26_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_26_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_26_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_26_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_26_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_26_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_26_0_searchSpace_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_26_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_26_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_26_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_26_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_26_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_26_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_26_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_26_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_26_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_26_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_26_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_26_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_26_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_26_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_26_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_26_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_26_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_26_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_3_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_3_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_3_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_3_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_3_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_3_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_3_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_3_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_3_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_3_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_3_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_3_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_3_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_3_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_3_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_3_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_3_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_3_0_searchSpace_0_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_3_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_3_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_3_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_3_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_3_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_3_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_3_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_3_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_3_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_3_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_3_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_3_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_3_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_3_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_3_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_3_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_3_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_3_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_4_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_4_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_4_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_4_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_4_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_4_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_4_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_4_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_4_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_4_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_4_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_4_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_4_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_4_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_4_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_4_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_4_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_4_0_searchSpace_0_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_4_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_4_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_4_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_4_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_4_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_4_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_4_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_4_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_4_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_4_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_4_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_4_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_4_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_4_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_4_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_4_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_4_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_4_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_5_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_5_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_5_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_5_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_5_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_5_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_5_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_5_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_5_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_5_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_5_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_5_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_5_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_5_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_5_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_5_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_5_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_5_0_searchSpace_0_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_5_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_5_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_5_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_5_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_5_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_5_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_5_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_5_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_5_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_5_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_5_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_5_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_5_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_5_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_5_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_5_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_5_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_5_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_6_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_6_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_6_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_6_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_6_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_6_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_6_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_6_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_6_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_6_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_6_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_6_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_6_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_6_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_6_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_6_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_6_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_6_0_searchSpace_0_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_6_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_6_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_6_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_6_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_6_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_6_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_6_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_6_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_6_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_6_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_6_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_6_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_6_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_6_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_6_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_6_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_6_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_6_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_7_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_7_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_7_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_7_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_7_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_7_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_7_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_7_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_7_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_7_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_7_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_7_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_7_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_7_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_7_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_7_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_7_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_7_0_searchSpace_0_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_7_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_7_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_7_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_7_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_7_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_7_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_7_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_7_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_7_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_7_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_7_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_7_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_7_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_7_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_7_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_7_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_7_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_7_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_8_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_8_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_8_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_8_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_8_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_8_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_8_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_8_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_8_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_8_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_8_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_8_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_8_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_8_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_8_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_8_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_8_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_8_0_searchSpace_0_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_8_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_8_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_8_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_8_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_8_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_8_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_8_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_8_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_8_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_8_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_8_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_8_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_8_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_8_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_8_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_8_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_8_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_8_0_start_id_0,
    output wire                                          krnl_partialKnn_wrapper_9_0_ap_clk,
    input wire                                           krnl_partialKnn_wrapper_9_0_ap_done,
    input wire                                           krnl_partialKnn_wrapper_9_0_ap_idle,
    input wire                                           krnl_partialKnn_wrapper_9_0_ap_ready,
    output wire                                          krnl_partialKnn_wrapper_9_0_ap_rst_n,
    output wire                                          krnl_partialKnn_wrapper_9_0_ap_start,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_9_0_out_dist_din,
    output wire                                          krnl_partialKnn_wrapper_9_0_out_dist_full_n,
    input wire                                           krnl_partialKnn_wrapper_9_0_out_dist_write,
    input wire  [                                  65:0] krnl_partialKnn_wrapper_9_0_out_id_din,
    output wire                                          krnl_partialKnn_wrapper_9_0_out_id_full_n,
    input wire                                           krnl_partialKnn_wrapper_9_0_out_id_write,
    output wire [                                  63:0] krnl_partialKnn_wrapper_9_0_searchSpace_0_read_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_9_0_searchSpace_0_read_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_9_0_searchSpace_0_read_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_9_0_searchSpace_0_read_addr_s_write,
    output wire [                                 256:0] krnl_partialKnn_wrapper_9_0_searchSpace_0_read_data_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_9_0_searchSpace_0_read_data_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_9_0_searchSpace_0_read_data_peek_read,
    output wire [                                 256:0] krnl_partialKnn_wrapper_9_0_searchSpace_0_read_data_s_dout,
    output wire                                          krnl_partialKnn_wrapper_9_0_searchSpace_0_read_data_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_9_0_searchSpace_0_read_data_s_read,
    output wire [                                  63:0] krnl_partialKnn_wrapper_9_0_searchSpace_0_write_addr_offset,
    input wire  [                                  63:0] krnl_partialKnn_wrapper_9_0_searchSpace_0_write_addr_s_din,
    output wire                                          krnl_partialKnn_wrapper_9_0_searchSpace_0_write_addr_s_full_n,
    input wire                                           krnl_partialKnn_wrapper_9_0_searchSpace_0_write_addr_s_write,
    input wire  [                                 256:0] krnl_partialKnn_wrapper_9_0_searchSpace_0_write_data_din,
    output wire                                          krnl_partialKnn_wrapper_9_0_searchSpace_0_write_data_full_n,
    input wire                                           krnl_partialKnn_wrapper_9_0_searchSpace_0_write_data_write,
    output wire [                                   8:0] krnl_partialKnn_wrapper_9_0_searchSpace_0_write_resp_peek_dout,
    output wire                                          krnl_partialKnn_wrapper_9_0_searchSpace_write_resp_peek_empty_n,
    input wire                                           krnl_partialKnn_wrapper_9_0_searchSpace_0_write_resp_peek_read,
    output wire [                                   8:0] krnl_partialKnn_wrapper_9_0_searchSpace_0_write_resp_s_dout,
    output wire                                          krnl_partialKnn_wrapper_9_0_searchSpace_0_write_resp_s_empty_n,
    input wire                                           krnl_partialKnn_wrapper_9_0_searchSpace_0_write_resp_s_read,
    output wire [                                  31:0] krnl_partialKnn_wrapper_9_0_start_id_0,
    output wire                                          L3_out_dist__m_axi_clk,
    input wire  [                                  63:0] L3_out_dist__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] L3_out_dist__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] L3_out_dist__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] L3_out_dist__m_axi_m_axi_ARID,
    input wire  [                                   7:0] L3_out_dist__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] L3_out_dist__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] L3_out_dist__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] L3_out_dist__m_axi_m_axi_ARQOS,
    output wire                                          L3_out_dist__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] L3_out_dist__m_axi_m_axi_ARSIZE,
    input wire                                           L3_out_dist__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] L3_out_dist__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] L3_out_dist__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] L3_out_dist__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] L3_out_dist__m_axi_m_axi_AWID,
    input wire  [                                   7:0] L3_out_dist__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] L3_out_dist__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] L3_out_dist__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] L3_out_dist__m_axi_m_axi_AWQOS,
    output wire                                          L3_out_dist__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] L3_out_dist__m_axi_m_axi_AWSIZE,
    input wire                                           L3_out_dist__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] L3_out_dist__m_axi_m_axi_BID,
    input wire                                           L3_out_dist__m_axi_m_axi_BREADY,
    output wire [                                   1:0] L3_out_dist__m_axi_m_axi_BRESP,
    output wire                                          L3_out_dist__m_axi_m_axi_BVALID,
    output wire [                                  31:0] L3_out_dist__m_axi_m_axi_RDATA,
    output wire [                                   0:0] L3_out_dist__m_axi_m_axi_RID,
    output wire                                          L3_out_dist__m_axi_m_axi_RLAST,
    input wire                                           L3_out_dist__m_axi_m_axi_RREADY,
    output wire [                                   1:0] L3_out_dist__m_axi_m_axi_RRESP,
    output wire                                          L3_out_dist__m_axi_m_axi_RVALID,
    input wire  [                                  31:0] L3_out_dist__m_axi_m_axi_WDATA,
    input wire                                           L3_out_dist__m_axi_m_axi_WLAST,
    output wire                                          L3_out_dist__m_axi_m_axi_WREADY,
    input wire  [                                   3:0] L3_out_dist__m_axi_m_axi_WSTRB,
    input wire                                           L3_out_dist__m_axi_m_axi_WVALID,
    output wire [                                  63:0] L3_out_dist__m_axi_read_addr_din,
    input wire                                           L3_out_dist__m_axi_read_addr_full_n,
    output wire                                          L3_out_dist__m_axi_read_addr_write,
    input wire  [                                  31:0] L3_out_dist__m_axi_read_data_dout,
    input wire                                           L3_out_dist__m_axi_read_data_empty_n,
    output wire                                          L3_out_dist__m_axi_read_data_read,
    output wire                                          L3_out_dist__m_axi_rst,
    output wire [                                  63:0] L3_out_dist__m_axi_write_addr_din,
    input wire                                           L3_out_dist__m_axi_write_addr_full_n,
    output wire                                          L3_out_dist__m_axi_write_addr_write,
    output wire [                                  31:0] L3_out_dist__m_axi_write_data_din,
    input wire                                           L3_out_dist__m_axi_write_data_full_n,
    output wire                                          L3_out_dist__m_axi_write_data_write,
    input wire  [                                   7:0] L3_out_dist__m_axi_write_resp_dout,
    input wire                                           L3_out_dist__m_axi_write_resp_empty_n,
    output wire                                          L3_out_dist__m_axi_write_resp_read,
    output wire                                          L3_out_id__m_axi_clk,
    input wire  [                                  63:0] L3_out_id__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] L3_out_id__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] L3_out_id__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] L3_out_id__m_axi_m_axi_ARID,
    input wire  [                                   7:0] L3_out_id__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] L3_out_id__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] L3_out_id__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] L3_out_id__m_axi_m_axi_ARQOS,
    output wire                                          L3_out_id__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] L3_out_id__m_axi_m_axi_ARSIZE,
    input wire                                           L3_out_id__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] L3_out_id__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] L3_out_id__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] L3_out_id__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] L3_out_id__m_axi_m_axi_AWID,
    input wire  [                                   7:0] L3_out_id__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] L3_out_id__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] L3_out_id__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] L3_out_id__m_axi_m_axi_AWQOS,
    output wire                                          L3_out_id__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] L3_out_id__m_axi_m_axi_AWSIZE,
    input wire                                           L3_out_id__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] L3_out_id__m_axi_m_axi_BID,
    input wire                                           L3_out_id__m_axi_m_axi_BREADY,
    output wire [                                   1:0] L3_out_id__m_axi_m_axi_BRESP,
    output wire                                          L3_out_id__m_axi_m_axi_BVALID,
    output wire [                                  31:0] L3_out_id__m_axi_m_axi_RDATA,
    output wire [                                   0:0] L3_out_id__m_axi_m_axi_RID,
    output wire                                          L3_out_id__m_axi_m_axi_RLAST,
    input wire                                           L3_out_id__m_axi_m_axi_RREADY,
    output wire [                                   1:0] L3_out_id__m_axi_m_axi_RRESP,
    output wire                                          L3_out_id__m_axi_m_axi_RVALID,
    input wire  [                                  31:0] L3_out_id__m_axi_m_axi_WDATA,
    input wire                                           L3_out_id__m_axi_m_axi_WLAST,
    output wire                                          L3_out_id__m_axi_m_axi_WREADY,
    input wire  [                                   3:0] L3_out_id__m_axi_m_axi_WSTRB,
    input wire                                           L3_out_id__m_axi_m_axi_WVALID,
    output wire [                                  63:0] L3_out_id__m_axi_read_addr_din,
    input wire                                           L3_out_id__m_axi_read_addr_full_n,
    output wire                                          L3_out_id__m_axi_read_addr_write,
    input wire  [                                  31:0] L3_out_id__m_axi_read_data_dout,
    input wire                                           L3_out_id__m_axi_read_data_empty_n,
    output wire                                          L3_out_id__m_axi_read_data_read,
    output wire                                          L3_out_id__m_axi_rst,
    output wire [                                  63:0] L3_out_id__m_axi_write_addr_din,
    input wire                                           L3_out_id__m_axi_write_addr_full_n,
    output wire                                          L3_out_id__m_axi_write_addr_write,
    output wire [                                  31:0] L3_out_id__m_axi_write_data_din,
    input wire                                           L3_out_id__m_axi_write_data_full_n,
    output wire                                          L3_out_id__m_axi_write_data_write,
    input wire  [                                   7:0] L3_out_id__m_axi_write_resp_dout,
    input wire                                           L3_out_id__m_axi_write_resp_empty_n,
    output wire                                          L3_out_id__m_axi_write_resp_read,
    output wire                                          in_0__m_axi_clk,
    input wire  [                                  63:0] in_0__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_0__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_0__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_0__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_0__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_0__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_0__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_0__m_axi_m_axi_ARQOS,
    output wire                                          in_0__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_0__m_axi_m_axi_ARSIZE,
    input wire                                           in_0__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_0__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_0__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_0__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_0__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_0__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_0__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_0__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_0__m_axi_m_axi_AWQOS,
    output wire                                          in_0__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_0__m_axi_m_axi_AWSIZE,
    input wire                                           in_0__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_0__m_axi_m_axi_BID,
    input wire                                           in_0__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_0__m_axi_m_axi_BRESP,
    output wire                                          in_0__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_0__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_0__m_axi_m_axi_RID,
    output wire                                          in_0__m_axi_m_axi_RLAST,
    input wire                                           in_0__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_0__m_axi_m_axi_RRESP,
    output wire                                          in_0__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_0__m_axi_m_axi_WDATA,
    input wire                                           in_0__m_axi_m_axi_WLAST,
    output wire                                          in_0__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_0__m_axi_m_axi_WSTRB,
    input wire                                           in_0__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_0__m_axi_read_addr_din,
    input wire                                           in_0__m_axi_read_addr_full_n,
    output wire                                          in_0__m_axi_read_addr_write,
    input wire  [                                 255:0] in_0__m_axi_read_data_dout,
    input wire                                           in_0__m_axi_read_data_empty_n,
    output wire                                          in_0__m_axi_read_data_read,
    output wire                                          in_0__m_axi_rst,
    output wire [                                  63:0] in_0__m_axi_write_addr_din,
    input wire                                           in_0__m_axi_write_addr_full_n,
    output wire                                          in_0__m_axi_write_addr_write,
    output wire [                                 255:0] in_0__m_axi_write_data_din,
    input wire                                           in_0__m_axi_write_data_full_n,
    output wire                                          in_0__m_axi_write_data_write,
    input wire  [                                   7:0] in_0__m_axi_write_resp_dout,
    input wire                                           in_0__m_axi_write_resp_empty_n,
    output wire                                          in_0__m_axi_write_resp_read,
    output wire                                          in_1__m_axi_clk,
    input wire  [                                  63:0] in_1__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_1__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_1__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_1__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_1__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_1__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_1__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_1__m_axi_m_axi_ARQOS,
    output wire                                          in_1__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_1__m_axi_m_axi_ARSIZE,
    input wire                                           in_1__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_1__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_1__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_1__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_1__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_1__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_1__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_1__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_1__m_axi_m_axi_AWQOS,
    output wire                                          in_1__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_1__m_axi_m_axi_AWSIZE,
    input wire                                           in_1__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_1__m_axi_m_axi_BID,
    input wire                                           in_1__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_1__m_axi_m_axi_BRESP,
    output wire                                          in_1__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_1__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_1__m_axi_m_axi_RID,
    output wire                                          in_1__m_axi_m_axi_RLAST,
    input wire                                           in_1__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_1__m_axi_m_axi_RRESP,
    output wire                                          in_1__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_1__m_axi_m_axi_WDATA,
    input wire                                           in_1__m_axi_m_axi_WLAST,
    output wire                                          in_1__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_1__m_axi_m_axi_WSTRB,
    input wire                                           in_1__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_1__m_axi_read_addr_din,
    input wire                                           in_1__m_axi_read_addr_full_n,
    output wire                                          in_1__m_axi_read_addr_write,
    input wire  [                                 255:0] in_1__m_axi_read_data_dout,
    input wire                                           in_1__m_axi_read_data_empty_n,
    output wire                                          in_1__m_axi_read_data_read,
    output wire                                          in_1__m_axi_rst,
    output wire [                                  63:0] in_1__m_axi_write_addr_din,
    input wire                                           in_1__m_axi_write_addr_full_n,
    output wire                                          in_1__m_axi_write_addr_write,
    output wire [                                 255:0] in_1__m_axi_write_data_din,
    input wire                                           in_1__m_axi_write_data_full_n,
    output wire                                          in_1__m_axi_write_data_write,
    input wire  [                                   7:0] in_1__m_axi_write_resp_dout,
    input wire                                           in_1__m_axi_write_resp_empty_n,
    output wire                                          in_1__m_axi_write_resp_read,
    output wire                                          in_10__m_axi_clk,
    input wire  [                                  63:0] in_10__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_10__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_10__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_10__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_10__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_10__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_10__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_10__m_axi_m_axi_ARQOS,
    output wire                                          in_10__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_10__m_axi_m_axi_ARSIZE,
    input wire                                           in_10__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_10__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_10__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_10__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_10__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_10__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_10__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_10__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_10__m_axi_m_axi_AWQOS,
    output wire                                          in_10__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_10__m_axi_m_axi_AWSIZE,
    input wire                                           in_10__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_10__m_axi_m_axi_BID,
    input wire                                           in_10__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_10__m_axi_m_axi_BRESP,
    output wire                                          in_10__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_10__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_10__m_axi_m_axi_RID,
    output wire                                          in_10__m_axi_m_axi_RLAST,
    input wire                                           in_10__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_10__m_axi_m_axi_RRESP,
    output wire                                          in_10__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_10__m_axi_m_axi_WDATA,
    input wire                                           in_10__m_axi_m_axi_WLAST,
    output wire                                          in_10__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_10__m_axi_m_axi_WSTRB,
    input wire                                           in_10__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_10__m_axi_read_addr_din,
    input wire                                           in_10__m_axi_read_addr_full_n,
    output wire                                          in_10__m_axi_read_addr_write,
    input wire  [                                 255:0] in_10__m_axi_read_data_dout,
    input wire                                           in_10__m_axi_read_data_empty_n,
    output wire                                          in_10__m_axi_read_data_read,
    output wire                                          in_10__m_axi_rst,
    output wire [                                  63:0] in_10__m_axi_write_addr_din,
    input wire                                           in_10__m_axi_write_addr_full_n,
    output wire                                          in_10__m_axi_write_addr_write,
    output wire [                                 255:0] in_10__m_axi_write_data_din,
    input wire                                           in_10__m_axi_write_data_full_n,
    output wire                                          in_10__m_axi_write_data_write,
    input wire  [                                   7:0] in_10__m_axi_write_resp_dout,
    input wire                                           in_10__m_axi_write_resp_empty_n,
    output wire                                          in_10__m_axi_write_resp_read,
    output wire                                          in_11__m_axi_clk,
    input wire  [                                  63:0] in_11__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_11__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_11__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_11__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_11__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_11__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_11__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_11__m_axi_m_axi_ARQOS,
    output wire                                          in_11__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_11__m_axi_m_axi_ARSIZE,
    input wire                                           in_11__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_11__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_11__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_11__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_11__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_11__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_11__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_11__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_11__m_axi_m_axi_AWQOS,
    output wire                                          in_11__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_11__m_axi_m_axi_AWSIZE,
    input wire                                           in_11__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_11__m_axi_m_axi_BID,
    input wire                                           in_11__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_11__m_axi_m_axi_BRESP,
    output wire                                          in_11__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_11__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_11__m_axi_m_axi_RID,
    output wire                                          in_11__m_axi_m_axi_RLAST,
    input wire                                           in_11__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_11__m_axi_m_axi_RRESP,
    output wire                                          in_11__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_11__m_axi_m_axi_WDATA,
    input wire                                           in_11__m_axi_m_axi_WLAST,
    output wire                                          in_11__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_11__m_axi_m_axi_WSTRB,
    input wire                                           in_11__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_11__m_axi_read_addr_din,
    input wire                                           in_11__m_axi_read_addr_full_n,
    output wire                                          in_11__m_axi_read_addr_write,
    input wire  [                                 255:0] in_11__m_axi_read_data_dout,
    input wire                                           in_11__m_axi_read_data_empty_n,
    output wire                                          in_11__m_axi_read_data_read,
    output wire                                          in_11__m_axi_rst,
    output wire [                                  63:0] in_11__m_axi_write_addr_din,
    input wire                                           in_11__m_axi_write_addr_full_n,
    output wire                                          in_11__m_axi_write_addr_write,
    output wire [                                 255:0] in_11__m_axi_write_data_din,
    input wire                                           in_11__m_axi_write_data_full_n,
    output wire                                          in_11__m_axi_write_data_write,
    input wire  [                                   7:0] in_11__m_axi_write_resp_dout,
    input wire                                           in_11__m_axi_write_resp_empty_n,
    output wire                                          in_11__m_axi_write_resp_read,
    output wire                                          in_12__m_axi_clk,
    input wire  [                                  63:0] in_12__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_12__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_12__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_12__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_12__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_12__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_12__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_12__m_axi_m_axi_ARQOS,
    output wire                                          in_12__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_12__m_axi_m_axi_ARSIZE,
    input wire                                           in_12__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_12__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_12__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_12__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_12__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_12__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_12__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_12__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_12__m_axi_m_axi_AWQOS,
    output wire                                          in_12__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_12__m_axi_m_axi_AWSIZE,
    input wire                                           in_12__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_12__m_axi_m_axi_BID,
    input wire                                           in_12__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_12__m_axi_m_axi_BRESP,
    output wire                                          in_12__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_12__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_12__m_axi_m_axi_RID,
    output wire                                          in_12__m_axi_m_axi_RLAST,
    input wire                                           in_12__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_12__m_axi_m_axi_RRESP,
    output wire                                          in_12__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_12__m_axi_m_axi_WDATA,
    input wire                                           in_12__m_axi_m_axi_WLAST,
    output wire                                          in_12__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_12__m_axi_m_axi_WSTRB,
    input wire                                           in_12__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_12__m_axi_read_addr_din,
    input wire                                           in_12__m_axi_read_addr_full_n,
    output wire                                          in_12__m_axi_read_addr_write,
    input wire  [                                 255:0] in_12__m_axi_read_data_dout,
    input wire                                           in_12__m_axi_read_data_empty_n,
    output wire                                          in_12__m_axi_read_data_read,
    output wire                                          in_12__m_axi_rst,
    output wire [                                  63:0] in_12__m_axi_write_addr_din,
    input wire                                           in_12__m_axi_write_addr_full_n,
    output wire                                          in_12__m_axi_write_addr_write,
    output wire [                                 255:0] in_12__m_axi_write_data_din,
    input wire                                           in_12__m_axi_write_data_full_n,
    output wire                                          in_12__m_axi_write_data_write,
    input wire  [                                   7:0] in_12__m_axi_write_resp_dout,
    input wire                                           in_12__m_axi_write_resp_empty_n,
    output wire                                          in_12__m_axi_write_resp_read,
    output wire                                          in_13__m_axi_clk,
    input wire  [                                  63:0] in_13__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_13__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_13__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_13__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_13__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_13__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_13__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_13__m_axi_m_axi_ARQOS,
    output wire                                          in_13__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_13__m_axi_m_axi_ARSIZE,
    input wire                                           in_13__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_13__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_13__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_13__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_13__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_13__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_13__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_13__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_13__m_axi_m_axi_AWQOS,
    output wire                                          in_13__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_13__m_axi_m_axi_AWSIZE,
    input wire                                           in_13__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_13__m_axi_m_axi_BID,
    input wire                                           in_13__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_13__m_axi_m_axi_BRESP,
    output wire                                          in_13__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_13__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_13__m_axi_m_axi_RID,
    output wire                                          in_13__m_axi_m_axi_RLAST,
    input wire                                           in_13__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_13__m_axi_m_axi_RRESP,
    output wire                                          in_13__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_13__m_axi_m_axi_WDATA,
    input wire                                           in_13__m_axi_m_axi_WLAST,
    output wire                                          in_13__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_13__m_axi_m_axi_WSTRB,
    input wire                                           in_13__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_13__m_axi_read_addr_din,
    input wire                                           in_13__m_axi_read_addr_full_n,
    output wire                                          in_13__m_axi_read_addr_write,
    input wire  [                                 255:0] in_13__m_axi_read_data_dout,
    input wire                                           in_13__m_axi_read_data_empty_n,
    output wire                                          in_13__m_axi_read_data_read,
    output wire                                          in_13__m_axi_rst,
    output wire [                                  63:0] in_13__m_axi_write_addr_din,
    input wire                                           in_13__m_axi_write_addr_full_n,
    output wire                                          in_13__m_axi_write_addr_write,
    output wire [                                 255:0] in_13__m_axi_write_data_din,
    input wire                                           in_13__m_axi_write_data_full_n,
    output wire                                          in_13__m_axi_write_data_write,
    input wire  [                                   7:0] in_13__m_axi_write_resp_dout,
    input wire                                           in_13__m_axi_write_resp_empty_n,
    output wire                                          in_13__m_axi_write_resp_read,
    output wire                                          in_14__m_axi_clk,
    input wire  [                                  63:0] in_14__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_14__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_14__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_14__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_14__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_14__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_14__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_14__m_axi_m_axi_ARQOS,
    output wire                                          in_14__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_14__m_axi_m_axi_ARSIZE,
    input wire                                           in_14__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_14__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_14__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_14__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_14__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_14__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_14__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_14__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_14__m_axi_m_axi_AWQOS,
    output wire                                          in_14__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_14__m_axi_m_axi_AWSIZE,
    input wire                                           in_14__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_14__m_axi_m_axi_BID,
    input wire                                           in_14__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_14__m_axi_m_axi_BRESP,
    output wire                                          in_14__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_14__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_14__m_axi_m_axi_RID,
    output wire                                          in_14__m_axi_m_axi_RLAST,
    input wire                                           in_14__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_14__m_axi_m_axi_RRESP,
    output wire                                          in_14__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_14__m_axi_m_axi_WDATA,
    input wire                                           in_14__m_axi_m_axi_WLAST,
    output wire                                          in_14__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_14__m_axi_m_axi_WSTRB,
    input wire                                           in_14__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_14__m_axi_read_addr_din,
    input wire                                           in_14__m_axi_read_addr_full_n,
    output wire                                          in_14__m_axi_read_addr_write,
    input wire  [                                 255:0] in_14__m_axi_read_data_dout,
    input wire                                           in_14__m_axi_read_data_empty_n,
    output wire                                          in_14__m_axi_read_data_read,
    output wire                                          in_14__m_axi_rst,
    output wire [                                  63:0] in_14__m_axi_write_addr_din,
    input wire                                           in_14__m_axi_write_addr_full_n,
    output wire                                          in_14__m_axi_write_addr_write,
    output wire [                                 255:0] in_14__m_axi_write_data_din,
    input wire                                           in_14__m_axi_write_data_full_n,
    output wire                                          in_14__m_axi_write_data_write,
    input wire  [                                   7:0] in_14__m_axi_write_resp_dout,
    input wire                                           in_14__m_axi_write_resp_empty_n,
    output wire                                          in_14__m_axi_write_resp_read,
    output wire                                          in_15__m_axi_clk,
    input wire  [                                  63:0] in_15__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_15__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_15__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_15__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_15__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_15__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_15__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_15__m_axi_m_axi_ARQOS,
    output wire                                          in_15__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_15__m_axi_m_axi_ARSIZE,
    input wire                                           in_15__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_15__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_15__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_15__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_15__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_15__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_15__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_15__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_15__m_axi_m_axi_AWQOS,
    output wire                                          in_15__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_15__m_axi_m_axi_AWSIZE,
    input wire                                           in_15__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_15__m_axi_m_axi_BID,
    input wire                                           in_15__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_15__m_axi_m_axi_BRESP,
    output wire                                          in_15__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_15__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_15__m_axi_m_axi_RID,
    output wire                                          in_15__m_axi_m_axi_RLAST,
    input wire                                           in_15__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_15__m_axi_m_axi_RRESP,
    output wire                                          in_15__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_15__m_axi_m_axi_WDATA,
    input wire                                           in_15__m_axi_m_axi_WLAST,
    output wire                                          in_15__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_15__m_axi_m_axi_WSTRB,
    input wire                                           in_15__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_15__m_axi_read_addr_din,
    input wire                                           in_15__m_axi_read_addr_full_n,
    output wire                                          in_15__m_axi_read_addr_write,
    input wire  [                                 255:0] in_15__m_axi_read_data_dout,
    input wire                                           in_15__m_axi_read_data_empty_n,
    output wire                                          in_15__m_axi_read_data_read,
    output wire                                          in_15__m_axi_rst,
    output wire [                                  63:0] in_15__m_axi_write_addr_din,
    input wire                                           in_15__m_axi_write_addr_full_n,
    output wire                                          in_15__m_axi_write_addr_write,
    output wire [                                 255:0] in_15__m_axi_write_data_din,
    input wire                                           in_15__m_axi_write_data_full_n,
    output wire                                          in_15__m_axi_write_data_write,
    input wire  [                                   7:0] in_15__m_axi_write_resp_dout,
    input wire                                           in_15__m_axi_write_resp_empty_n,
    output wire                                          in_15__m_axi_write_resp_read,
    output wire                                          in_16__m_axi_clk,
    input wire  [                                  63:0] in_16__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_16__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_16__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_16__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_16__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_16__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_16__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_16__m_axi_m_axi_ARQOS,
    output wire                                          in_16__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_16__m_axi_m_axi_ARSIZE,
    input wire                                           in_16__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_16__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_16__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_16__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_16__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_16__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_16__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_16__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_16__m_axi_m_axi_AWQOS,
    output wire                                          in_16__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_16__m_axi_m_axi_AWSIZE,
    input wire                                           in_16__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_16__m_axi_m_axi_BID,
    input wire                                           in_16__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_16__m_axi_m_axi_BRESP,
    output wire                                          in_16__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_16__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_16__m_axi_m_axi_RID,
    output wire                                          in_16__m_axi_m_axi_RLAST,
    input wire                                           in_16__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_16__m_axi_m_axi_RRESP,
    output wire                                          in_16__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_16__m_axi_m_axi_WDATA,
    input wire                                           in_16__m_axi_m_axi_WLAST,
    output wire                                          in_16__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_16__m_axi_m_axi_WSTRB,
    input wire                                           in_16__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_16__m_axi_read_addr_din,
    input wire                                           in_16__m_axi_read_addr_full_n,
    output wire                                          in_16__m_axi_read_addr_write,
    input wire  [                                 255:0] in_16__m_axi_read_data_dout,
    input wire                                           in_16__m_axi_read_data_empty_n,
    output wire                                          in_16__m_axi_read_data_read,
    output wire                                          in_16__m_axi_rst,
    output wire [                                  63:0] in_16__m_axi_write_addr_din,
    input wire                                           in_16__m_axi_write_addr_full_n,
    output wire                                          in_16__m_axi_write_addr_write,
    output wire [                                 255:0] in_16__m_axi_write_data_din,
    input wire                                           in_16__m_axi_write_data_full_n,
    output wire                                          in_16__m_axi_write_data_write,
    input wire  [                                   7:0] in_16__m_axi_write_resp_dout,
    input wire                                           in_16__m_axi_write_resp_empty_n,
    output wire                                          in_16__m_axi_write_resp_read,
    output wire                                          in_17__m_axi_clk,
    input wire  [                                  63:0] in_17__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_17__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_17__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_17__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_17__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_17__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_17__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_17__m_axi_m_axi_ARQOS,
    output wire                                          in_17__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_17__m_axi_m_axi_ARSIZE,
    input wire                                           in_17__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_17__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_17__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_17__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_17__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_17__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_17__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_17__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_17__m_axi_m_axi_AWQOS,
    output wire                                          in_17__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_17__m_axi_m_axi_AWSIZE,
    input wire                                           in_17__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_17__m_axi_m_axi_BID,
    input wire                                           in_17__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_17__m_axi_m_axi_BRESP,
    output wire                                          in_17__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_17__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_17__m_axi_m_axi_RID,
    output wire                                          in_17__m_axi_m_axi_RLAST,
    input wire                                           in_17__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_17__m_axi_m_axi_RRESP,
    output wire                                          in_17__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_17__m_axi_m_axi_WDATA,
    input wire                                           in_17__m_axi_m_axi_WLAST,
    output wire                                          in_17__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_17__m_axi_m_axi_WSTRB,
    input wire                                           in_17__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_17__m_axi_read_addr_din,
    input wire                                           in_17__m_axi_read_addr_full_n,
    output wire                                          in_17__m_axi_read_addr_write,
    input wire  [                                 255:0] in_17__m_axi_read_data_dout,
    input wire                                           in_17__m_axi_read_data_empty_n,
    output wire                                          in_17__m_axi_read_data_read,
    output wire                                          in_17__m_axi_rst,
    output wire [                                  63:0] in_17__m_axi_write_addr_din,
    input wire                                           in_17__m_axi_write_addr_full_n,
    output wire                                          in_17__m_axi_write_addr_write,
    output wire [                                 255:0] in_17__m_axi_write_data_din,
    input wire                                           in_17__m_axi_write_data_full_n,
    output wire                                          in_17__m_axi_write_data_write,
    input wire  [                                   7:0] in_17__m_axi_write_resp_dout,
    input wire                                           in_17__m_axi_write_resp_empty_n,
    output wire                                          in_17__m_axi_write_resp_read,
    output wire                                          in_18__m_axi_clk,
    input wire  [                                  63:0] in_18__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_18__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_18__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_18__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_18__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_18__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_18__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_18__m_axi_m_axi_ARQOS,
    output wire                                          in_18__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_18__m_axi_m_axi_ARSIZE,
    input wire                                           in_18__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_18__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_18__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_18__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_18__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_18__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_18__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_18__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_18__m_axi_m_axi_AWQOS,
    output wire                                          in_18__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_18__m_axi_m_axi_AWSIZE,
    input wire                                           in_18__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_18__m_axi_m_axi_BID,
    input wire                                           in_18__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_18__m_axi_m_axi_BRESP,
    output wire                                          in_18__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_18__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_18__m_axi_m_axi_RID,
    output wire                                          in_18__m_axi_m_axi_RLAST,
    input wire                                           in_18__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_18__m_axi_m_axi_RRESP,
    output wire                                          in_18__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_18__m_axi_m_axi_WDATA,
    input wire                                           in_18__m_axi_m_axi_WLAST,
    output wire                                          in_18__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_18__m_axi_m_axi_WSTRB,
    input wire                                           in_18__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_18__m_axi_read_addr_din,
    input wire                                           in_18__m_axi_read_addr_full_n,
    output wire                                          in_18__m_axi_read_addr_write,
    input wire  [                                 255:0] in_18__m_axi_read_data_dout,
    input wire                                           in_18__m_axi_read_data_empty_n,
    output wire                                          in_18__m_axi_read_data_read,
    output wire                                          in_18__m_axi_rst,
    output wire [                                  63:0] in_18__m_axi_write_addr_din,
    input wire                                           in_18__m_axi_write_addr_full_n,
    output wire                                          in_18__m_axi_write_addr_write,
    output wire [                                 255:0] in_18__m_axi_write_data_din,
    input wire                                           in_18__m_axi_write_data_full_n,
    output wire                                          in_18__m_axi_write_data_write,
    input wire  [                                   7:0] in_18__m_axi_write_resp_dout,
    input wire                                           in_18__m_axi_write_resp_empty_n,
    output wire                                          in_18__m_axi_write_resp_read,
    output wire                                          in_19__m_axi_clk,
    input wire  [                                  63:0] in_19__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_19__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_19__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_19__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_19__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_19__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_19__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_19__m_axi_m_axi_ARQOS,
    output wire                                          in_19__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_19__m_axi_m_axi_ARSIZE,
    input wire                                           in_19__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_19__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_19__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_19__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_19__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_19__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_19__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_19__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_19__m_axi_m_axi_AWQOS,
    output wire                                          in_19__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_19__m_axi_m_axi_AWSIZE,
    input wire                                           in_19__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_19__m_axi_m_axi_BID,
    input wire                                           in_19__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_19__m_axi_m_axi_BRESP,
    output wire                                          in_19__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_19__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_19__m_axi_m_axi_RID,
    output wire                                          in_19__m_axi_m_axi_RLAST,
    input wire                                           in_19__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_19__m_axi_m_axi_RRESP,
    output wire                                          in_19__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_19__m_axi_m_axi_WDATA,
    input wire                                           in_19__m_axi_m_axi_WLAST,
    output wire                                          in_19__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_19__m_axi_m_axi_WSTRB,
    input wire                                           in_19__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_19__m_axi_read_addr_din,
    input wire                                           in_19__m_axi_read_addr_full_n,
    output wire                                          in_19__m_axi_read_addr_write,
    input wire  [                                 255:0] in_19__m_axi_read_data_dout,
    input wire                                           in_19__m_axi_read_data_empty_n,
    output wire                                          in_19__m_axi_read_data_read,
    output wire                                          in_19__m_axi_rst,
    output wire [                                  63:0] in_19__m_axi_write_addr_din,
    input wire                                           in_19__m_axi_write_addr_full_n,
    output wire                                          in_19__m_axi_write_addr_write,
    output wire [                                 255:0] in_19__m_axi_write_data_din,
    input wire                                           in_19__m_axi_write_data_full_n,
    output wire                                          in_19__m_axi_write_data_write,
    input wire  [                                   7:0] in_19__m_axi_write_resp_dout,
    input wire                                           in_19__m_axi_write_resp_empty_n,
    output wire                                          in_19__m_axi_write_resp_read,
    output wire                                          in_2__m_axi_clk,
    input wire  [                                  63:0] in_2__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_2__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_2__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_2__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_2__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_2__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_2__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_2__m_axi_m_axi_ARQOS,
    output wire                                          in_2__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_2__m_axi_m_axi_ARSIZE,
    input wire                                           in_2__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_2__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_2__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_2__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_2__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_2__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_2__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_2__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_2__m_axi_m_axi_AWQOS,
    output wire                                          in_2__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_2__m_axi_m_axi_AWSIZE,
    input wire                                           in_2__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_2__m_axi_m_axi_BID,
    input wire                                           in_2__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_2__m_axi_m_axi_BRESP,
    output wire                                          in_2__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_2__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_2__m_axi_m_axi_RID,
    output wire                                          in_2__m_axi_m_axi_RLAST,
    input wire                                           in_2__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_2__m_axi_m_axi_RRESP,
    output wire                                          in_2__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_2__m_axi_m_axi_WDATA,
    input wire                                           in_2__m_axi_m_axi_WLAST,
    output wire                                          in_2__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_2__m_axi_m_axi_WSTRB,
    input wire                                           in_2__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_2__m_axi_read_addr_din,
    input wire                                           in_2__m_axi_read_addr_full_n,
    output wire                                          in_2__m_axi_read_addr_write,
    input wire  [                                 255:0] in_2__m_axi_read_data_dout,
    input wire                                           in_2__m_axi_read_data_empty_n,
    output wire                                          in_2__m_axi_read_data_read,
    output wire                                          in_2__m_axi_rst,
    output wire [                                  63:0] in_2__m_axi_write_addr_din,
    input wire                                           in_2__m_axi_write_addr_full_n,
    output wire                                          in_2__m_axi_write_addr_write,
    output wire [                                 255:0] in_2__m_axi_write_data_din,
    input wire                                           in_2__m_axi_write_data_full_n,
    output wire                                          in_2__m_axi_write_data_write,
    input wire  [                                   7:0] in_2__m_axi_write_resp_dout,
    input wire                                           in_2__m_axi_write_resp_empty_n,
    output wire                                          in_2__m_axi_write_resp_read,
    output wire                                          in_20__m_axi_clk,
    input wire  [                                  63:0] in_20__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_20__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_20__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_20__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_20__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_20__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_20__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_20__m_axi_m_axi_ARQOS,
    output wire                                          in_20__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_20__m_axi_m_axi_ARSIZE,
    input wire                                           in_20__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_20__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_20__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_20__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_20__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_20__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_20__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_20__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_20__m_axi_m_axi_AWQOS,
    output wire                                          in_20__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_20__m_axi_m_axi_AWSIZE,
    input wire                                           in_20__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_20__m_axi_m_axi_BID,
    input wire                                           in_20__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_20__m_axi_m_axi_BRESP,
    output wire                                          in_20__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_20__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_20__m_axi_m_axi_RID,
    output wire                                          in_20__m_axi_m_axi_RLAST,
    input wire                                           in_20__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_20__m_axi_m_axi_RRESP,
    output wire                                          in_20__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_20__m_axi_m_axi_WDATA,
    input wire                                           in_20__m_axi_m_axi_WLAST,
    output wire                                          in_20__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_20__m_axi_m_axi_WSTRB,
    input wire                                           in_20__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_20__m_axi_read_addr_din,
    input wire                                           in_20__m_axi_read_addr_full_n,
    output wire                                          in_20__m_axi_read_addr_write,
    input wire  [                                 255:0] in_20__m_axi_read_data_dout,
    input wire                                           in_20__m_axi_read_data_empty_n,
    output wire                                          in_20__m_axi_read_data_read,
    output wire                                          in_20__m_axi_rst,
    output wire [                                  63:0] in_20__m_axi_write_addr_din,
    input wire                                           in_20__m_axi_write_addr_full_n,
    output wire                                          in_20__m_axi_write_addr_write,
    output wire [                                 255:0] in_20__m_axi_write_data_din,
    input wire                                           in_20__m_axi_write_data_full_n,
    output wire                                          in_20__m_axi_write_data_write,
    input wire  [                                   7:0] in_20__m_axi_write_resp_dout,
    input wire                                           in_20__m_axi_write_resp_empty_n,
    output wire                                          in_20__m_axi_write_resp_read,
    output wire                                          in_21__m_axi_clk,
    input wire  [                                  63:0] in_21__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_21__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_21__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_21__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_21__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_21__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_21__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_21__m_axi_m_axi_ARQOS,
    output wire                                          in_21__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_21__m_axi_m_axi_ARSIZE,
    input wire                                           in_21__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_21__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_21__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_21__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_21__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_21__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_21__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_21__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_21__m_axi_m_axi_AWQOS,
    output wire                                          in_21__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_21__m_axi_m_axi_AWSIZE,
    input wire                                           in_21__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_21__m_axi_m_axi_BID,
    input wire                                           in_21__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_21__m_axi_m_axi_BRESP,
    output wire                                          in_21__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_21__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_21__m_axi_m_axi_RID,
    output wire                                          in_21__m_axi_m_axi_RLAST,
    input wire                                           in_21__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_21__m_axi_m_axi_RRESP,
    output wire                                          in_21__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_21__m_axi_m_axi_WDATA,
    input wire                                           in_21__m_axi_m_axi_WLAST,
    output wire                                          in_21__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_21__m_axi_m_axi_WSTRB,
    input wire                                           in_21__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_21__m_axi_read_addr_din,
    input wire                                           in_21__m_axi_read_addr_full_n,
    output wire                                          in_21__m_axi_read_addr_write,
    input wire  [                                 255:0] in_21__m_axi_read_data_dout,
    input wire                                           in_21__m_axi_read_data_empty_n,
    output wire                                          in_21__m_axi_read_data_read,
    output wire                                          in_21__m_axi_rst,
    output wire [                                  63:0] in_21__m_axi_write_addr_din,
    input wire                                           in_21__m_axi_write_addr_full_n,
    output wire                                          in_21__m_axi_write_addr_write,
    output wire [                                 255:0] in_21__m_axi_write_data_din,
    input wire                                           in_21__m_axi_write_data_full_n,
    output wire                                          in_21__m_axi_write_data_write,
    input wire  [                                   7:0] in_21__m_axi_write_resp_dout,
    input wire                                           in_21__m_axi_write_resp_empty_n,
    output wire                                          in_21__m_axi_write_resp_read,
    output wire                                          in_22__m_axi_clk,
    input wire  [                                  63:0] in_22__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_22__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_22__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_22__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_22__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_22__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_22__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_22__m_axi_m_axi_ARQOS,
    output wire                                          in_22__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_22__m_axi_m_axi_ARSIZE,
    input wire                                           in_22__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_22__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_22__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_22__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_22__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_22__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_22__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_22__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_22__m_axi_m_axi_AWQOS,
    output wire                                          in_22__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_22__m_axi_m_axi_AWSIZE,
    input wire                                           in_22__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_22__m_axi_m_axi_BID,
    input wire                                           in_22__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_22__m_axi_m_axi_BRESP,
    output wire                                          in_22__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_22__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_22__m_axi_m_axi_RID,
    output wire                                          in_22__m_axi_m_axi_RLAST,
    input wire                                           in_22__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_22__m_axi_m_axi_RRESP,
    output wire                                          in_22__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_22__m_axi_m_axi_WDATA,
    input wire                                           in_22__m_axi_m_axi_WLAST,
    output wire                                          in_22__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_22__m_axi_m_axi_WSTRB,
    input wire                                           in_22__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_22__m_axi_read_addr_din,
    input wire                                           in_22__m_axi_read_addr_full_n,
    output wire                                          in_22__m_axi_read_addr_write,
    input wire  [                                 255:0] in_22__m_axi_read_data_dout,
    input wire                                           in_22__m_axi_read_data_empty_n,
    output wire                                          in_22__m_axi_read_data_read,
    output wire                                          in_22__m_axi_rst,
    output wire [                                  63:0] in_22__m_axi_write_addr_din,
    input wire                                           in_22__m_axi_write_addr_full_n,
    output wire                                          in_22__m_axi_write_addr_write,
    output wire [                                 255:0] in_22__m_axi_write_data_din,
    input wire                                           in_22__m_axi_write_data_full_n,
    output wire                                          in_22__m_axi_write_data_write,
    input wire  [                                   7:0] in_22__m_axi_write_resp_dout,
    input wire                                           in_22__m_axi_write_resp_empty_n,
    output wire                                          in_22__m_axi_write_resp_read,
    output wire                                          in_23__m_axi_clk,
    input wire  [                                  63:0] in_23__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_23__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_23__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_23__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_23__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_23__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_23__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_23__m_axi_m_axi_ARQOS,
    output wire                                          in_23__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_23__m_axi_m_axi_ARSIZE,
    input wire                                           in_23__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_23__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_23__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_23__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_23__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_23__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_23__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_23__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_23__m_axi_m_axi_AWQOS,
    output wire                                          in_23__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_23__m_axi_m_axi_AWSIZE,
    input wire                                           in_23__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_23__m_axi_m_axi_BID,
    input wire                                           in_23__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_23__m_axi_m_axi_BRESP,
    output wire                                          in_23__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_23__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_23__m_axi_m_axi_RID,
    output wire                                          in_23__m_axi_m_axi_RLAST,
    input wire                                           in_23__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_23__m_axi_m_axi_RRESP,
    output wire                                          in_23__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_23__m_axi_m_axi_WDATA,
    input wire                                           in_23__m_axi_m_axi_WLAST,
    output wire                                          in_23__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_23__m_axi_m_axi_WSTRB,
    input wire                                           in_23__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_23__m_axi_read_addr_din,
    input wire                                           in_23__m_axi_read_addr_full_n,
    output wire                                          in_23__m_axi_read_addr_write,
    input wire  [                                 255:0] in_23__m_axi_read_data_dout,
    input wire                                           in_23__m_axi_read_data_empty_n,
    output wire                                          in_23__m_axi_read_data_read,
    output wire                                          in_23__m_axi_rst,
    output wire [                                  63:0] in_23__m_axi_write_addr_din,
    input wire                                           in_23__m_axi_write_addr_full_n,
    output wire                                          in_23__m_axi_write_addr_write,
    output wire [                                 255:0] in_23__m_axi_write_data_din,
    input wire                                           in_23__m_axi_write_data_full_n,
    output wire                                          in_23__m_axi_write_data_write,
    input wire  [                                   7:0] in_23__m_axi_write_resp_dout,
    input wire                                           in_23__m_axi_write_resp_empty_n,
    output wire                                          in_23__m_axi_write_resp_read,
    output wire                                          in_24__m_axi_clk,
    input wire  [                                  63:0] in_24__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_24__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_24__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_24__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_24__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_24__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_24__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_24__m_axi_m_axi_ARQOS,
    output wire                                          in_24__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_24__m_axi_m_axi_ARSIZE,
    input wire                                           in_24__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_24__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_24__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_24__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_24__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_24__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_24__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_24__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_24__m_axi_m_axi_AWQOS,
    output wire                                          in_24__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_24__m_axi_m_axi_AWSIZE,
    input wire                                           in_24__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_24__m_axi_m_axi_BID,
    input wire                                           in_24__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_24__m_axi_m_axi_BRESP,
    output wire                                          in_24__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_24__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_24__m_axi_m_axi_RID,
    output wire                                          in_24__m_axi_m_axi_RLAST,
    input wire                                           in_24__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_24__m_axi_m_axi_RRESP,
    output wire                                          in_24__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_24__m_axi_m_axi_WDATA,
    input wire                                           in_24__m_axi_m_axi_WLAST,
    output wire                                          in_24__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_24__m_axi_m_axi_WSTRB,
    input wire                                           in_24__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_24__m_axi_read_addr_din,
    input wire                                           in_24__m_axi_read_addr_full_n,
    output wire                                          in_24__m_axi_read_addr_write,
    input wire  [                                 255:0] in_24__m_axi_read_data_dout,
    input wire                                           in_24__m_axi_read_data_empty_n,
    output wire                                          in_24__m_axi_read_data_read,
    output wire                                          in_24__m_axi_rst,
    output wire [                                  63:0] in_24__m_axi_write_addr_din,
    input wire                                           in_24__m_axi_write_addr_full_n,
    output wire                                          in_24__m_axi_write_addr_write,
    output wire [                                 255:0] in_24__m_axi_write_data_din,
    input wire                                           in_24__m_axi_write_data_full_n,
    output wire                                          in_24__m_axi_write_data_write,
    input wire  [                                   7:0] in_24__m_axi_write_resp_dout,
    input wire                                           in_24__m_axi_write_resp_empty_n,
    output wire                                          in_24__m_axi_write_resp_read,
    output wire                                          in_25__m_axi_clk,
    input wire  [                                  63:0] in_25__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_25__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_25__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_25__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_25__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_25__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_25__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_25__m_axi_m_axi_ARQOS,
    output wire                                          in_25__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_25__m_axi_m_axi_ARSIZE,
    input wire                                           in_25__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_25__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_25__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_25__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_25__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_25__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_25__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_25__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_25__m_axi_m_axi_AWQOS,
    output wire                                          in_25__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_25__m_axi_m_axi_AWSIZE,
    input wire                                           in_25__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_25__m_axi_m_axi_BID,
    input wire                                           in_25__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_25__m_axi_m_axi_BRESP,
    output wire                                          in_25__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_25__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_25__m_axi_m_axi_RID,
    output wire                                          in_25__m_axi_m_axi_RLAST,
    input wire                                           in_25__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_25__m_axi_m_axi_RRESP,
    output wire                                          in_25__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_25__m_axi_m_axi_WDATA,
    input wire                                           in_25__m_axi_m_axi_WLAST,
    output wire                                          in_25__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_25__m_axi_m_axi_WSTRB,
    input wire                                           in_25__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_25__m_axi_read_addr_din,
    input wire                                           in_25__m_axi_read_addr_full_n,
    output wire                                          in_25__m_axi_read_addr_write,
    input wire  [                                 255:0] in_25__m_axi_read_data_dout,
    input wire                                           in_25__m_axi_read_data_empty_n,
    output wire                                          in_25__m_axi_read_data_read,
    output wire                                          in_25__m_axi_rst,
    output wire [                                  63:0] in_25__m_axi_write_addr_din,
    input wire                                           in_25__m_axi_write_addr_full_n,
    output wire                                          in_25__m_axi_write_addr_write,
    output wire [                                 255:0] in_25__m_axi_write_data_din,
    input wire                                           in_25__m_axi_write_data_full_n,
    output wire                                          in_25__m_axi_write_data_write,
    input wire  [                                   7:0] in_25__m_axi_write_resp_dout,
    input wire                                           in_25__m_axi_write_resp_empty_n,
    output wire                                          in_25__m_axi_write_resp_read,
    output wire                                          in_26__m_axi_clk,
    input wire  [                                  63:0] in_26__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_26__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_26__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_26__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_26__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_26__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_26__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_26__m_axi_m_axi_ARQOS,
    output wire                                          in_26__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_26__m_axi_m_axi_ARSIZE,
    input wire                                           in_26__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_26__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_26__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_26__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_26__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_26__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_26__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_26__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_26__m_axi_m_axi_AWQOS,
    output wire                                          in_26__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_26__m_axi_m_axi_AWSIZE,
    input wire                                           in_26__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_26__m_axi_m_axi_BID,
    input wire                                           in_26__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_26__m_axi_m_axi_BRESP,
    output wire                                          in_26__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_26__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_26__m_axi_m_axi_RID,
    output wire                                          in_26__m_axi_m_axi_RLAST,
    input wire                                           in_26__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_26__m_axi_m_axi_RRESP,
    output wire                                          in_26__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_26__m_axi_m_axi_WDATA,
    input wire                                           in_26__m_axi_m_axi_WLAST,
    output wire                                          in_26__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_26__m_axi_m_axi_WSTRB,
    input wire                                           in_26__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_26__m_axi_read_addr_din,
    input wire                                           in_26__m_axi_read_addr_full_n,
    output wire                                          in_26__m_axi_read_addr_write,
    input wire  [                                 255:0] in_26__m_axi_read_data_dout,
    input wire                                           in_26__m_axi_read_data_empty_n,
    output wire                                          in_26__m_axi_read_data_read,
    output wire                                          in_26__m_axi_rst,
    output wire [                                  63:0] in_26__m_axi_write_addr_din,
    input wire                                           in_26__m_axi_write_addr_full_n,
    output wire                                          in_26__m_axi_write_addr_write,
    output wire [                                 255:0] in_26__m_axi_write_data_din,
    input wire                                           in_26__m_axi_write_data_full_n,
    output wire                                          in_26__m_axi_write_data_write,
    input wire  [                                   7:0] in_26__m_axi_write_resp_dout,
    input wire                                           in_26__m_axi_write_resp_empty_n,
    output wire                                          in_26__m_axi_write_resp_read,
    output wire                                          in_3__m_axi_clk,
    input wire  [                                  63:0] in_3__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_3__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_3__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_3__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_3__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_3__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_3__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_3__m_axi_m_axi_ARQOS,
    output wire                                          in_3__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_3__m_axi_m_axi_ARSIZE,
    input wire                                           in_3__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_3__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_3__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_3__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_3__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_3__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_3__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_3__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_3__m_axi_m_axi_AWQOS,
    output wire                                          in_3__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_3__m_axi_m_axi_AWSIZE,
    input wire                                           in_3__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_3__m_axi_m_axi_BID,
    input wire                                           in_3__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_3__m_axi_m_axi_BRESP,
    output wire                                          in_3__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_3__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_3__m_axi_m_axi_RID,
    output wire                                          in_3__m_axi_m_axi_RLAST,
    input wire                                           in_3__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_3__m_axi_m_axi_RRESP,
    output wire                                          in_3__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_3__m_axi_m_axi_WDATA,
    input wire                                           in_3__m_axi_m_axi_WLAST,
    output wire                                          in_3__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_3__m_axi_m_axi_WSTRB,
    input wire                                           in_3__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_3__m_axi_read_addr_din,
    input wire                                           in_3__m_axi_read_addr_full_n,
    output wire                                          in_3__m_axi_read_addr_write,
    input wire  [                                 255:0] in_3__m_axi_read_data_dout,
    input wire                                           in_3__m_axi_read_data_empty_n,
    output wire                                          in_3__m_axi_read_data_read,
    output wire                                          in_3__m_axi_rst,
    output wire [                                  63:0] in_3__m_axi_write_addr_din,
    input wire                                           in_3__m_axi_write_addr_full_n,
    output wire                                          in_3__m_axi_write_addr_write,
    output wire [                                 255:0] in_3__m_axi_write_data_din,
    input wire                                           in_3__m_axi_write_data_full_n,
    output wire                                          in_3__m_axi_write_data_write,
    input wire  [                                   7:0] in_3__m_axi_write_resp_dout,
    input wire                                           in_3__m_axi_write_resp_empty_n,
    output wire                                          in_3__m_axi_write_resp_read,
    output wire                                          in_4__m_axi_clk,
    input wire  [                                  63:0] in_4__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_4__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_4__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_4__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_4__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_4__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_4__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_4__m_axi_m_axi_ARQOS,
    output wire                                          in_4__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_4__m_axi_m_axi_ARSIZE,
    input wire                                           in_4__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_4__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_4__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_4__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_4__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_4__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_4__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_4__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_4__m_axi_m_axi_AWQOS,
    output wire                                          in_4__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_4__m_axi_m_axi_AWSIZE,
    input wire                                           in_4__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_4__m_axi_m_axi_BID,
    input wire                                           in_4__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_4__m_axi_m_axi_BRESP,
    output wire                                          in_4__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_4__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_4__m_axi_m_axi_RID,
    output wire                                          in_4__m_axi_m_axi_RLAST,
    input wire                                           in_4__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_4__m_axi_m_axi_RRESP,
    output wire                                          in_4__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_4__m_axi_m_axi_WDATA,
    input wire                                           in_4__m_axi_m_axi_WLAST,
    output wire                                          in_4__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_4__m_axi_m_axi_WSTRB,
    input wire                                           in_4__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_4__m_axi_read_addr_din,
    input wire                                           in_4__m_axi_read_addr_full_n,
    output wire                                          in_4__m_axi_read_addr_write,
    input wire  [                                 255:0] in_4__m_axi_read_data_dout,
    input wire                                           in_4__m_axi_read_data_empty_n,
    output wire                                          in_4__m_axi_read_data_read,
    output wire                                          in_4__m_axi_rst,
    output wire [                                  63:0] in_4__m_axi_write_addr_din,
    input wire                                           in_4__m_axi_write_addr_full_n,
    output wire                                          in_4__m_axi_write_addr_write,
    output wire [                                 255:0] in_4__m_axi_write_data_din,
    input wire                                           in_4__m_axi_write_data_full_n,
    output wire                                          in_4__m_axi_write_data_write,
    input wire  [                                   7:0] in_4__m_axi_write_resp_dout,
    input wire                                           in_4__m_axi_write_resp_empty_n,
    output wire                                          in_4__m_axi_write_resp_read,
    output wire                                          in_5__m_axi_clk,
    input wire  [                                  63:0] in_5__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_5__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_5__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_5__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_5__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_5__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_5__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_5__m_axi_m_axi_ARQOS,
    output wire                                          in_5__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_5__m_axi_m_axi_ARSIZE,
    input wire                                           in_5__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_5__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_5__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_5__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_5__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_5__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_5__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_5__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_5__m_axi_m_axi_AWQOS,
    output wire                                          in_5__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_5__m_axi_m_axi_AWSIZE,
    input wire                                           in_5__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_5__m_axi_m_axi_BID,
    input wire                                           in_5__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_5__m_axi_m_axi_BRESP,
    output wire                                          in_5__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_5__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_5__m_axi_m_axi_RID,
    output wire                                          in_5__m_axi_m_axi_RLAST,
    input wire                                           in_5__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_5__m_axi_m_axi_RRESP,
    output wire                                          in_5__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_5__m_axi_m_axi_WDATA,
    input wire                                           in_5__m_axi_m_axi_WLAST,
    output wire                                          in_5__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_5__m_axi_m_axi_WSTRB,
    input wire                                           in_5__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_5__m_axi_read_addr_din,
    input wire                                           in_5__m_axi_read_addr_full_n,
    output wire                                          in_5__m_axi_read_addr_write,
    input wire  [                                 255:0] in_5__m_axi_read_data_dout,
    input wire                                           in_5__m_axi_read_data_empty_n,
    output wire                                          in_5__m_axi_read_data_read,
    output wire                                          in_5__m_axi_rst,
    output wire [                                  63:0] in_5__m_axi_write_addr_din,
    input wire                                           in_5__m_axi_write_addr_full_n,
    output wire                                          in_5__m_axi_write_addr_write,
    output wire [                                 255:0] in_5__m_axi_write_data_din,
    input wire                                           in_5__m_axi_write_data_full_n,
    output wire                                          in_5__m_axi_write_data_write,
    input wire  [                                   7:0] in_5__m_axi_write_resp_dout,
    input wire                                           in_5__m_axi_write_resp_empty_n,
    output wire                                          in_5__m_axi_write_resp_read,
    output wire                                          in_6__m_axi_clk,
    input wire  [                                  63:0] in_6__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_6__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_6__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_6__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_6__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_6__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_6__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_6__m_axi_m_axi_ARQOS,
    output wire                                          in_6__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_6__m_axi_m_axi_ARSIZE,
    input wire                                           in_6__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_6__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_6__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_6__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_6__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_6__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_6__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_6__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_6__m_axi_m_axi_AWQOS,
    output wire                                          in_6__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_6__m_axi_m_axi_AWSIZE,
    input wire                                           in_6__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_6__m_axi_m_axi_BID,
    input wire                                           in_6__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_6__m_axi_m_axi_BRESP,
    output wire                                          in_6__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_6__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_6__m_axi_m_axi_RID,
    output wire                                          in_6__m_axi_m_axi_RLAST,
    input wire                                           in_6__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_6__m_axi_m_axi_RRESP,
    output wire                                          in_6__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_6__m_axi_m_axi_WDATA,
    input wire                                           in_6__m_axi_m_axi_WLAST,
    output wire                                          in_6__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_6__m_axi_m_axi_WSTRB,
    input wire                                           in_6__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_6__m_axi_read_addr_din,
    input wire                                           in_6__m_axi_read_addr_full_n,
    output wire                                          in_6__m_axi_read_addr_write,
    input wire  [                                 255:0] in_6__m_axi_read_data_dout,
    input wire                                           in_6__m_axi_read_data_empty_n,
    output wire                                          in_6__m_axi_read_data_read,
    output wire                                          in_6__m_axi_rst,
    output wire [                                  63:0] in_6__m_axi_write_addr_din,
    input wire                                           in_6__m_axi_write_addr_full_n,
    output wire                                          in_6__m_axi_write_addr_write,
    output wire [                                 255:0] in_6__m_axi_write_data_din,
    input wire                                           in_6__m_axi_write_data_full_n,
    output wire                                          in_6__m_axi_write_data_write,
    input wire  [                                   7:0] in_6__m_axi_write_resp_dout,
    input wire                                           in_6__m_axi_write_resp_empty_n,
    output wire                                          in_6__m_axi_write_resp_read,
    output wire                                          in_7__m_axi_clk,
    input wire  [                                  63:0] in_7__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_7__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_7__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_7__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_7__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_7__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_7__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_7__m_axi_m_axi_ARQOS,
    output wire                                          in_7__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_7__m_axi_m_axi_ARSIZE,
    input wire                                           in_7__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_7__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_7__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_7__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_7__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_7__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_7__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_7__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_7__m_axi_m_axi_AWQOS,
    output wire                                          in_7__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_7__m_axi_m_axi_AWSIZE,
    input wire                                           in_7__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_7__m_axi_m_axi_BID,
    input wire                                           in_7__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_7__m_axi_m_axi_BRESP,
    output wire                                          in_7__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_7__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_7__m_axi_m_axi_RID,
    output wire                                          in_7__m_axi_m_axi_RLAST,
    input wire                                           in_7__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_7__m_axi_m_axi_RRESP,
    output wire                                          in_7__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_7__m_axi_m_axi_WDATA,
    input wire                                           in_7__m_axi_m_axi_WLAST,
    output wire                                          in_7__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_7__m_axi_m_axi_WSTRB,
    input wire                                           in_7__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_7__m_axi_read_addr_din,
    input wire                                           in_7__m_axi_read_addr_full_n,
    output wire                                          in_7__m_axi_read_addr_write,
    input wire  [                                 255:0] in_7__m_axi_read_data_dout,
    input wire                                           in_7__m_axi_read_data_empty_n,
    output wire                                          in_7__m_axi_read_data_read,
    output wire                                          in_7__m_axi_rst,
    output wire [                                  63:0] in_7__m_axi_write_addr_din,
    input wire                                           in_7__m_axi_write_addr_full_n,
    output wire                                          in_7__m_axi_write_addr_write,
    output wire [                                 255:0] in_7__m_axi_write_data_din,
    input wire                                           in_7__m_axi_write_data_full_n,
    output wire                                          in_7__m_axi_write_data_write,
    input wire  [                                   7:0] in_7__m_axi_write_resp_dout,
    input wire                                           in_7__m_axi_write_resp_empty_n,
    output wire                                          in_7__m_axi_write_resp_read,
    output wire                                          in_8__m_axi_clk,
    input wire  [                                  63:0] in_8__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_8__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_8__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_8__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_8__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_8__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_8__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_8__m_axi_m_axi_ARQOS,
    output wire                                          in_8__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_8__m_axi_m_axi_ARSIZE,
    input wire                                           in_8__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_8__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_8__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_8__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_8__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_8__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_8__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_8__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_8__m_axi_m_axi_AWQOS,
    output wire                                          in_8__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_8__m_axi_m_axi_AWSIZE,
    input wire                                           in_8__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_8__m_axi_m_axi_BID,
    input wire                                           in_8__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_8__m_axi_m_axi_BRESP,
    output wire                                          in_8__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_8__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_8__m_axi_m_axi_RID,
    output wire                                          in_8__m_axi_m_axi_RLAST,
    input wire                                           in_8__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_8__m_axi_m_axi_RRESP,
    output wire                                          in_8__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_8__m_axi_m_axi_WDATA,
    input wire                                           in_8__m_axi_m_axi_WLAST,
    output wire                                          in_8__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_8__m_axi_m_axi_WSTRB,
    input wire                                           in_8__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_8__m_axi_read_addr_din,
    input wire                                           in_8__m_axi_read_addr_full_n,
    output wire                                          in_8__m_axi_read_addr_write,
    input wire  [                                 255:0] in_8__m_axi_read_data_dout,
    input wire                                           in_8__m_axi_read_data_empty_n,
    output wire                                          in_8__m_axi_read_data_read,
    output wire                                          in_8__m_axi_rst,
    output wire [                                  63:0] in_8__m_axi_write_addr_din,
    input wire                                           in_8__m_axi_write_addr_full_n,
    output wire                                          in_8__m_axi_write_addr_write,
    output wire [                                 255:0] in_8__m_axi_write_data_din,
    input wire                                           in_8__m_axi_write_data_full_n,
    output wire                                          in_8__m_axi_write_data_write,
    input wire  [                                   7:0] in_8__m_axi_write_resp_dout,
    input wire                                           in_8__m_axi_write_resp_empty_n,
    output wire                                          in_8__m_axi_write_resp_read,
    output wire                                          in_9__m_axi_clk,
    input wire  [                                  63:0] in_9__m_axi_m_axi_ARADDR,
    input wire  [                                   1:0] in_9__m_axi_m_axi_ARBURST,
    input wire  [                                   3:0] in_9__m_axi_m_axi_ARCACHE,
    input wire  [                                   0:0] in_9__m_axi_m_axi_ARID,
    input wire  [                                   7:0] in_9__m_axi_m_axi_ARLEN,
    input wire  [                                   0:0] in_9__m_axi_m_axi_ARLOCK,
    input wire  [                                   2:0] in_9__m_axi_m_axi_ARPROT,
    input wire  [                                   3:0] in_9__m_axi_m_axi_ARQOS,
    output wire                                          in_9__m_axi_m_axi_ARREADY,
    input wire  [                                   2:0] in_9__m_axi_m_axi_ARSIZE,
    input wire                                           in_9__m_axi_m_axi_ARVALID,
    input wire  [                                  63:0] in_9__m_axi_m_axi_AWADDR,
    input wire  [                                   1:0] in_9__m_axi_m_axi_AWBURST,
    input wire  [                                   3:0] in_9__m_axi_m_axi_AWCACHE,
    input wire  [                                   0:0] in_9__m_axi_m_axi_AWID,
    input wire  [                                   7:0] in_9__m_axi_m_axi_AWLEN,
    input wire  [                                   0:0] in_9__m_axi_m_axi_AWLOCK,
    input wire  [                                   2:0] in_9__m_axi_m_axi_AWPROT,
    input wire  [                                   3:0] in_9__m_axi_m_axi_AWQOS,
    output wire                                          in_9__m_axi_m_axi_AWREADY,
    input wire  [                                   2:0] in_9__m_axi_m_axi_AWSIZE,
    input wire                                           in_9__m_axi_m_axi_AWVALID,
    output wire [                                   0:0] in_9__m_axi_m_axi_BID,
    input wire                                           in_9__m_axi_m_axi_BREADY,
    output wire [                                   1:0] in_9__m_axi_m_axi_BRESP,
    output wire                                          in_9__m_axi_m_axi_BVALID,
    output wire [                                 255:0] in_9__m_axi_m_axi_RDATA,
    output wire [                                   0:0] in_9__m_axi_m_axi_RID,
    output wire                                          in_9__m_axi_m_axi_RLAST,
    input wire                                           in_9__m_axi_m_axi_RREADY,
    output wire [                                   1:0] in_9__m_axi_m_axi_RRESP,
    output wire                                          in_9__m_axi_m_axi_RVALID,
    input wire  [                                 255:0] in_9__m_axi_m_axi_WDATA,
    input wire                                           in_9__m_axi_m_axi_WLAST,
    output wire                                          in_9__m_axi_m_axi_WREADY,
    input wire  [                                  31:0] in_9__m_axi_m_axi_WSTRB,
    input wire                                           in_9__m_axi_m_axi_WVALID,
    output wire [                                  63:0] in_9__m_axi_read_addr_din,
    input wire                                           in_9__m_axi_read_addr_full_n,
    output wire                                          in_9__m_axi_read_addr_write,
    input wire  [                                 255:0] in_9__m_axi_read_data_dout,
    input wire                                           in_9__m_axi_read_data_empty_n,
    output wire                                          in_9__m_axi_read_data_read,
    output wire                                          in_9__m_axi_rst,
    output wire [                                  63:0] in_9__m_axi_write_addr_din,
    input wire                                           in_9__m_axi_write_addr_full_n,
    output wire                                          in_9__m_axi_write_addr_write,
    output wire [                                 255:0] in_9__m_axi_write_data_din,
    input wire                                           in_9__m_axi_write_data_full_n,
    output wire                                          in_9__m_axi_write_data_write,
    input wire  [                                   7:0] in_9__m_axi_write_resp_dout,
    input wire                                           in_9__m_axi_write_resp_empty_n,
    output wire                                          in_9__m_axi_write_resp_read,
    output wire [                                  63:0] __tapa_fsm_unit_L3_out_dist,
    output wire [                                  63:0] __tapa_fsm_unit_L3_out_id,
    output wire                                          __tapa_fsm_unit_ap_clk,
    input wire                                           __tapa_fsm_unit_ap_done,
    input wire                                           __tapa_fsm_unit_ap_idle,
    input wire                                           __tapa_fsm_unit_ap_ready,
    output wire                                          __tapa_fsm_unit_ap_rst_n,
    output wire                                          __tapa_fsm_unit_ap_start,
    output wire [                                  63:0] __tapa_fsm_unit_in_0,
    output wire [                                  63:0] __tapa_fsm_unit_in_1,
    output wire [                                  63:0] __tapa_fsm_unit_in_10,
    output wire [                                  63:0] __tapa_fsm_unit_in_11,
    output wire [                                  63:0] __tapa_fsm_unit_in_12,
    output wire [                                  63:0] __tapa_fsm_unit_in_13,
    output wire [                                  63:0] __tapa_fsm_unit_in_14,
    output wire [                                  63:0] __tapa_fsm_unit_in_15,
    output wire [                                  63:0] __tapa_fsm_unit_in_16,
    output wire [                                  63:0] __tapa_fsm_unit_in_17,
    output wire [                                  63:0] __tapa_fsm_unit_in_18,
    output wire [                                  63:0] __tapa_fsm_unit_in_19,
    output wire [                                  63:0] __tapa_fsm_unit_in_2,
    output wire [                                  63:0] __tapa_fsm_unit_in_20,
    output wire [                                  63:0] __tapa_fsm_unit_in_21,
    output wire [                                  63:0] __tapa_fsm_unit_in_22,
    output wire [                                  63:0] __tapa_fsm_unit_in_23,
    output wire [                                  63:0] __tapa_fsm_unit_in_24,
    output wire [                                  63:0] __tapa_fsm_unit_in_25,
    output wire [                                  63:0] __tapa_fsm_unit_in_26,
    output wire [                                  63:0] __tapa_fsm_unit_in_3,
    output wire [                                  63:0] __tapa_fsm_unit_in_4,
    output wire [                                  63:0] __tapa_fsm_unit_in_5,
    output wire [                                  63:0] __tapa_fsm_unit_in_6,
    output wire [                                  63:0] __tapa_fsm_unit_in_7,
    output wire [                                  63:0] __tapa_fsm_unit_in_8,
    output wire [                                  63:0] __tapa_fsm_unit_in_9,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_globalSort_L1_L2_0__ap_start,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_10__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_10__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_10__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_globalSort_L1_L2_10__ap_start,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_11__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_11__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_11__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_globalSort_L1_L2_11__ap_start,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_12__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_12__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_12__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_globalSort_L1_L2_12__ap_start,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_1__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_1__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_1__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_globalSort_L1_L2_1__ap_start,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_2__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_2__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_2__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_globalSort_L1_L2_2__ap_start,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_3__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_3__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_3__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_globalSort_L1_L2_3__ap_start,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_4__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_4__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_4__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_globalSort_L1_L2_4__ap_start,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_5__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_5__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_5__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_globalSort_L1_L2_5__ap_start,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_6__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_6__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_6__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_globalSort_L1_L2_6__ap_start,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_7__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_7__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_7__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_globalSort_L1_L2_7__ap_start,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_8__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_8__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_8__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_globalSort_L1_L2_8__ap_start,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_9__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_9__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_globalSort_L1_L2_9__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_globalSort_L1_L2_9__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_output_dist_id_0___L3_out_dist__q0,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_output_dist_id_0___L3_out_id__q0,
    output wire                                          __tapa_fsm_unit_krnl_output_dist_id_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_output_dist_id_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_output_dist_id_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_output_dist_id_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_0_0___in_0__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_0_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_0_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_0_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_0_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_10_0___in_10__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_10_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_10_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_10_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_10_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_11_0___in_11__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_11_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_11_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_11_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_11_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_12_0___in_12__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_12_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_12_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_12_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_12_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_13_0___in_13__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_13_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_13_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_13_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_13_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_14_0___in_14__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_14_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_14_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_14_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_14_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_15_0___in_15__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_15_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_15_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_15_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_15_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_16_0___in_16__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_16_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_16_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_16_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_16_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_17_0___in_17__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_17_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_17_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_17_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_17_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_18_0___in_18__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_18_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_18_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_18_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_18_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_19_0___in_19__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_19_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_19_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_19_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_19_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_1_0___in_1__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_1_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_1_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_1_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_1_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_20_0___in_20__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_20_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_20_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_20_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_20_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_21_0___in_21__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_21_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_21_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_21_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_21_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_22_0___in_22__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_22_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_22_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_22_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_22_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_23_0___in_23__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_23_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_23_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_23_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_23_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_24_0___in_24__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_24_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_24_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_24_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_24_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_25_0___in_25__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_25_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_25_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_25_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_25_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_26_0___in_26__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_26_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_26_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_26_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_26_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_2_0___in_2__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_2_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_2_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_2_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_2_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_3_0___in_3__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_3_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_3_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_3_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_3_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_4_0___in_4__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_4_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_4_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_4_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_4_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_5_0___in_5__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_5_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_5_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_5_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_5_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_6_0___in_6__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_6_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_6_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_6_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_6_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_7_0___in_7__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_7_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_7_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_7_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_7_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_8_0___in_8__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_8_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_8_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_8_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_8_0__ap_start,
    input wire  [                                  63:0] __tapa_fsm_unit_krnl_partialKnn_wrapper_9_0___in_9__q0,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_9_0__ap_done,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_9_0__ap_idle,
    output wire                                          __tapa_fsm_unit_krnl_partialKnn_wrapper_9_0__ap_ready,
    input wire                                           __tapa_fsm_unit_krnl_partialKnn_wrapper_9_0__ap_start
);
  wire ap_start;
  wire [63:0] in_0;
  wire [63:0] in_1;
  wire [63:0] in_2;
  wire [63:0] in_3;
  wire [63:0] in_4;
  wire [63:0] in_5;
  wire [63:0] in_6;
  wire [63:0] in_7;
  wire [63:0] in_8;
  wire [63:0] in_9;
  wire [63:0] in_10;
  wire [63:0] in_11;
  wire [63:0] in_12;
  wire [63:0] in_13;
  wire [63:0] in_14;
  wire [63:0] in_15;
  wire [63:0] in_16;
  wire [63:0] in_17;
  wire [63:0] in_18;
  wire [63:0] in_19;
  wire [63:0] in_20;
  wire [63:0] in_21;
  wire [63:0] in_22;
  wire [63:0] in_23;
  wire [63:0] in_24;
  wire [63:0] in_25;
  wire [63:0] in_26;
  wire [63:0] L3_out_dist;
  wire [63:0] L3_out_id;
  wire [65:0] L1_out_dist_0__dout;
  wire L1_out_dist_0__empty_n;
  wire L1_out_dist_0__read;
  wire [65:0] L1_out_dist_0__din;
  wire L1_out_dist_0__full_n;
  wire L1_out_dist_0__write;
  wire [65:0] L1_out_dist_1__dout;
  wire L1_out_dist_1__empty_n;
  wire L1_out_dist_1__read;
  wire [65:0] L1_out_dist_1__din;
  wire L1_out_dist_1__full_n;
  wire L1_out_dist_1__write;
  wire [65:0] L1_out_dist_2__dout;
  wire L1_out_dist_2__empty_n;
  wire L1_out_dist_2__read;
  wire [65:0] L1_out_dist_2__din;
  wire L1_out_dist_2__full_n;
  wire L1_out_dist_2__write;
  wire [65:0] L1_out_dist_3__dout;
  wire L1_out_dist_3__empty_n;
  wire L1_out_dist_3__read;
  wire [65:0] L1_out_dist_3__din;
  wire L1_out_dist_3__full_n;
  wire L1_out_dist_3__write;
  wire [65:0] L1_out_dist_4__dout;
  wire L1_out_dist_4__empty_n;
  wire L1_out_dist_4__read;
  wire [65:0] L1_out_dist_4__din;
  wire L1_out_dist_4__full_n;
  wire L1_out_dist_4__write;
  wire [65:0] L1_out_dist_5__dout;
  wire L1_out_dist_5__empty_n;
  wire L1_out_dist_5__read;
  wire [65:0] L1_out_dist_5__din;
  wire L1_out_dist_5__full_n;
  wire L1_out_dist_5__write;
  wire [65:0] L1_out_dist_6__dout;
  wire L1_out_dist_6__empty_n;
  wire L1_out_dist_6__read;
  wire [65:0] L1_out_dist_6__din;
  wire L1_out_dist_6__full_n;
  wire L1_out_dist_6__write;
  wire [65:0] L1_out_dist_7__dout;
  wire L1_out_dist_7__empty_n;
  wire L1_out_dist_7__read;
  wire [65:0] L1_out_dist_7__din;
  wire L1_out_dist_7__full_n;
  wire L1_out_dist_7__write;
  wire [65:0] L1_out_dist_8__dout;
  wire L1_out_dist_8__empty_n;
  wire L1_out_dist_8__read;
  wire [65:0] L1_out_dist_8__din;
  wire L1_out_dist_8__full_n;
  wire L1_out_dist_8__write;
  wire [65:0] L1_out_id_0__dout;
  wire L1_out_id_0__empty_n;
  wire L1_out_id_0__read;
  wire [65:0] L1_out_id_0__din;
  wire L1_out_id_0__full_n;
  wire L1_out_id_0__write;
  wire [65:0] L1_out_id_1__dout;
  wire L1_out_id_1__empty_n;
  wire L1_out_id_1__read;
  wire [65:0] L1_out_id_1__din;
  wire L1_out_id_1__full_n;
  wire L1_out_id_1__write;
  wire [65:0] L1_out_id_2__dout;
  wire L1_out_id_2__empty_n;
  wire L1_out_id_2__read;
  wire [65:0] L1_out_id_2__din;
  wire L1_out_id_2__full_n;
  wire L1_out_id_2__write;
  wire [65:0] L1_out_id_3__dout;
  wire L1_out_id_3__empty_n;
  wire L1_out_id_3__read;
  wire [65:0] L1_out_id_3__din;
  wire L1_out_id_3__full_n;
  wire L1_out_id_3__write;
  wire [65:0] L1_out_id_4__dout;
  wire L1_out_id_4__empty_n;
  wire L1_out_id_4__read;
  wire [65:0] L1_out_id_4__din;
  wire L1_out_id_4__full_n;
  wire L1_out_id_4__write;
  wire [65:0] L1_out_id_5__dout;
  wire L1_out_id_5__empty_n;
  wire L1_out_id_5__read;
  wire [65:0] L1_out_id_5__din;
  wire L1_out_id_5__full_n;
  wire L1_out_id_5__write;
  wire [65:0] L1_out_id_6__dout;
  wire L1_out_id_6__empty_n;
  wire L1_out_id_6__read;
  wire [65:0] L1_out_id_6__din;
  wire L1_out_id_6__full_n;
  wire L1_out_id_6__write;
  wire [65:0] L1_out_id_7__dout;
  wire L1_out_id_7__empty_n;
  wire L1_out_id_7__read;
  wire [65:0] L1_out_id_7__din;
  wire L1_out_id_7__full_n;
  wire L1_out_id_7__write;
  wire [65:0] L1_out_id_8__dout;
  wire L1_out_id_8__empty_n;
  wire L1_out_id_8__read;
  wire [65:0] L1_out_id_8__din;
  wire L1_out_id_8__full_n;
  wire L1_out_id_8__write;
  wire [65:0] L2_out_dist0__dout;
  wire L2_out_dist0__empty_n;
  wire L2_out_dist0__read;
  wire [65:0] L2_out_dist0__din;
  wire L2_out_dist0__full_n;
  wire L2_out_dist0__write;
  wire [65:0] L2_out_dist1__dout;
  wire L2_out_dist1__empty_n;
  wire L2_out_dist1__read;
  wire [65:0] L2_out_dist1__din;
  wire L2_out_dist1__full_n;
  wire L2_out_dist1__write;
  wire [65:0] L2_out_dist2__dout;
  wire L2_out_dist2__empty_n;
  wire L2_out_dist2__read;
  wire [65:0] L2_out_dist2__din;
  wire L2_out_dist2__full_n;
  wire L2_out_dist2__write;
  wire [65:0] L2_out_id0__dout;
  wire L2_out_id0__empty_n;
  wire L2_out_id0__read;
  wire [65:0] L2_out_id0__din;
  wire L2_out_id0__full_n;
  wire L2_out_id0__write;
  wire [65:0] L2_out_id1__dout;
  wire L2_out_id1__empty_n;
  wire L2_out_id1__read;
  wire [65:0] L2_out_id1__din;
  wire L2_out_id1__full_n;
  wire L2_out_id1__write;
  wire [65:0] L2_out_id2__dout;
  wire L2_out_id2__empty_n;
  wire L2_out_id2__read;
  wire [65:0] L2_out_id2__din;
  wire L2_out_id2__full_n;
  wire L2_out_id2__write;
  wire [65:0] L3_out_dist_stream__dout;
  wire L3_out_dist_stream__empty_n;
  wire L3_out_dist_stream__read;
  wire [65:0] L3_out_dist_stream__din;
  wire L3_out_dist_stream__full_n;
  wire L3_out_dist_stream__write;
  wire [65:0] L3_out_id_stream__dout;
  wire L3_out_id_stream__empty_n;
  wire L3_out_id_stream__read;
  wire [65:0] L3_out_id_stream__din;
  wire L3_out_id_stream__full_n;
  wire L3_out_id_stream__write;
  wire [65:0] out_dist_0__dout;
  wire out_dist_0__empty_n;
  wire out_dist_0__read;
  wire [65:0] out_dist_0__din;
  wire out_dist_0__full_n;
  wire out_dist_0__write;
  wire [65:0] out_dist_10__dout;
  wire out_dist_10__empty_n;
  wire out_dist_10__read;
  wire [65:0] out_dist_10__din;
  wire out_dist_10__full_n;
  wire out_dist_10__write;
  wire [65:0] out_dist_11__dout;
  wire out_dist_11__empty_n;
  wire out_dist_11__read;
  wire [65:0] out_dist_11__din;
  wire out_dist_11__full_n;
  wire out_dist_11__write;
  wire [65:0] out_dist_12__dout;
  wire out_dist_12__empty_n;
  wire out_dist_12__read;
  wire [65:0] out_dist_12__din;
  wire out_dist_12__full_n;
  wire out_dist_12__write;
  wire [65:0] out_dist_13__dout;
  wire out_dist_13__empty_n;
  wire out_dist_13__read;
  wire [65:0] out_dist_13__din;
  wire out_dist_13__full_n;
  wire out_dist_13__write;
  wire [65:0] out_dist_14__dout;
  wire out_dist_14__empty_n;
  wire out_dist_14__read;
  wire [65:0] out_dist_14__din;
  wire out_dist_14__full_n;
  wire out_dist_14__write;
  wire [65:0] out_dist_15__dout;
  wire out_dist_15__empty_n;
  wire out_dist_15__read;
  wire [65:0] out_dist_15__din;
  wire out_dist_15__full_n;
  wire out_dist_15__write;
  wire [65:0] out_dist_16__dout;
  wire out_dist_16__empty_n;
  wire out_dist_16__read;
  wire [65:0] out_dist_16__din;
  wire out_dist_16__full_n;
  wire out_dist_16__write;
  wire [65:0] out_dist_17__dout;
  wire out_dist_17__empty_n;
  wire out_dist_17__read;
  wire [65:0] out_dist_17__din;
  wire out_dist_17__full_n;
  wire out_dist_17__write;
  wire [65:0] out_dist_18__dout;
  wire out_dist_18__empty_n;
  wire out_dist_18__read;
  wire [65:0] out_dist_18__din;
  wire out_dist_18__full_n;
  wire out_dist_18__write;
  wire [65:0] out_dist_19__dout;
  wire out_dist_19__empty_n;
  wire out_dist_19__read;
  wire [65:0] out_dist_19__din;
  wire out_dist_19__full_n;
  wire out_dist_19__write;
  wire [65:0] out_dist_1__dout;
  wire out_dist_1__empty_n;
  wire out_dist_1__read;
  wire [65:0] out_dist_1__din;
  wire out_dist_1__full_n;
  wire out_dist_1__write;
  wire [65:0] out_dist_20__dout;
  wire out_dist_20__empty_n;
  wire out_dist_20__read;
  wire [65:0] out_dist_20__din;
  wire out_dist_20__full_n;
  wire out_dist_20__write;
  wire [65:0] out_dist_21__dout;
  wire out_dist_21__empty_n;
  wire out_dist_21__read;
  wire [65:0] out_dist_21__din;
  wire out_dist_21__full_n;
  wire out_dist_21__write;
  wire [65:0] out_dist_22__dout;
  wire out_dist_22__empty_n;
  wire out_dist_22__read;
  wire [65:0] out_dist_22__din;
  wire out_dist_22__full_n;
  wire out_dist_22__write;
  wire [65:0] out_dist_23__dout;
  wire out_dist_23__empty_n;
  wire out_dist_23__read;
  wire [65:0] out_dist_23__din;
  wire out_dist_23__full_n;
  wire out_dist_23__write;
  wire [65:0] out_dist_24__dout;
  wire out_dist_24__empty_n;
  wire out_dist_24__read;
  wire [65:0] out_dist_24__din;
  wire out_dist_24__full_n;
  wire out_dist_24__write;
  wire [65:0] out_dist_25__dout;
  wire out_dist_25__empty_n;
  wire out_dist_25__read;
  wire [65:0] out_dist_25__din;
  wire out_dist_25__full_n;
  wire out_dist_25__write;
  wire [65:0] out_dist_26__dout;
  wire out_dist_26__empty_n;
  wire out_dist_26__read;
  wire [65:0] out_dist_26__din;
  wire out_dist_26__full_n;
  wire out_dist_26__write;
  wire [65:0] out_dist_2__dout;
  wire out_dist_2__empty_n;
  wire out_dist_2__read;
  wire [65:0] out_dist_2__din;
  wire out_dist_2__full_n;
  wire out_dist_2__write;
  wire [65:0] out_dist_3__dout;
  wire out_dist_3__empty_n;
  wire out_dist_3__read;
  wire [65:0] out_dist_3__din;
  wire out_dist_3__full_n;
  wire out_dist_3__write;
  wire [65:0] out_dist_4__dout;
  wire out_dist_4__empty_n;
  wire out_dist_4__read;
  wire [65:0] out_dist_4__din;
  wire out_dist_4__full_n;
  wire out_dist_4__write;
  wire [65:0] out_dist_5__dout;
  wire out_dist_5__empty_n;
  wire out_dist_5__read;
  wire [65:0] out_dist_5__din;
  wire out_dist_5__full_n;
  wire out_dist_5__write;
  wire [65:0] out_dist_6__dout;
  wire out_dist_6__empty_n;
  wire out_dist_6__read;
  wire [65:0] out_dist_6__din;
  wire out_dist_6__full_n;
  wire out_dist_6__write;
  wire [65:0] out_dist_7__dout;
  wire out_dist_7__empty_n;
  wire out_dist_7__read;
  wire [65:0] out_dist_7__din;
  wire out_dist_7__full_n;
  wire out_dist_7__write;
  wire [65:0] out_dist_8__dout;
  wire out_dist_8__empty_n;
  wire out_dist_8__read;
  wire [65:0] out_dist_8__din;
  wire out_dist_8__full_n;
  wire out_dist_8__write;
  wire [65:0] out_dist_9__dout;
  wire out_dist_9__empty_n;
  wire out_dist_9__read;
  wire [65:0] out_dist_9__din;
  wire out_dist_9__full_n;
  wire out_dist_9__write;
  wire [65:0] out_id_0__dout;
  wire out_id_0__empty_n;
  wire out_id_0__read;
  wire [65:0] out_id_0__din;
  wire out_id_0__full_n;
  wire out_id_0__write;
  wire [65:0] out_id_10__dout;
  wire out_id_10__empty_n;
  wire out_id_10__read;
  wire [65:0] out_id_10__din;
  wire out_id_10__full_n;
  wire out_id_10__write;
  wire [65:0] out_id_11__dout;
  wire out_id_11__empty_n;
  wire out_id_11__read;
  wire [65:0] out_id_11__din;
  wire out_id_11__full_n;
  wire out_id_11__write;
  wire [65:0] out_id_12__dout;
  wire out_id_12__empty_n;
  wire out_id_12__read;
  wire [65:0] out_id_12__din;
  wire out_id_12__full_n;
  wire out_id_12__write;
  wire [65:0] out_id_13__dout;
  wire out_id_13__empty_n;
  wire out_id_13__read;
  wire [65:0] out_id_13__din;
  wire out_id_13__full_n;
  wire out_id_13__write;
  wire [65:0] out_id_14__dout;
  wire out_id_14__empty_n;
  wire out_id_14__read;
  wire [65:0] out_id_14__din;
  wire out_id_14__full_n;
  wire out_id_14__write;
  wire [65:0] out_id_15__dout;
  wire out_id_15__empty_n;
  wire out_id_15__read;
  wire [65:0] out_id_15__din;
  wire out_id_15__full_n;
  wire out_id_15__write;
  wire [65:0] out_id_16__dout;
  wire out_id_16__empty_n;
  wire out_id_16__read;
  wire [65:0] out_id_16__din;
  wire out_id_16__full_n;
  wire out_id_16__write;
  wire [65:0] out_id_17__dout;
  wire out_id_17__empty_n;
  wire out_id_17__read;
  wire [65:0] out_id_17__din;
  wire out_id_17__full_n;
  wire out_id_17__write;
  wire [65:0] out_id_18__dout;
  wire out_id_18__empty_n;
  wire out_id_18__read;
  wire [65:0] out_id_18__din;
  wire out_id_18__full_n;
  wire out_id_18__write;
  wire [65:0] out_id_19__dout;
  wire out_id_19__empty_n;
  wire out_id_19__read;
  wire [65:0] out_id_19__din;
  wire out_id_19__full_n;
  wire out_id_19__write;
  wire [65:0] out_id_1__dout;
  wire out_id_1__empty_n;
  wire out_id_1__read;
  wire [65:0] out_id_1__din;
  wire out_id_1__full_n;
  wire out_id_1__write;
  wire [65:0] out_id_20__dout;
  wire out_id_20__empty_n;
  wire out_id_20__read;
  wire [65:0] out_id_20__din;
  wire out_id_20__full_n;
  wire out_id_20__write;
  wire [65:0] out_id_21__dout;
  wire out_id_21__empty_n;
  wire out_id_21__read;
  wire [65:0] out_id_21__din;
  wire out_id_21__full_n;
  wire out_id_21__write;
  wire [65:0] out_id_22__dout;
  wire out_id_22__empty_n;
  wire out_id_22__read;
  wire [65:0] out_id_22__din;
  wire out_id_22__full_n;
  wire out_id_22__write;
  wire [65:0] out_id_23__dout;
  wire out_id_23__empty_n;
  wire out_id_23__read;
  wire [65:0] out_id_23__din;
  wire out_id_23__full_n;
  wire out_id_23__write;
  wire [65:0] out_id_24__dout;
  wire out_id_24__empty_n;
  wire out_id_24__read;
  wire [65:0] out_id_24__din;
  wire out_id_24__full_n;
  wire out_id_24__write;
  wire [65:0] out_id_25__dout;
  wire out_id_25__empty_n;
  wire out_id_25__read;
  wire [65:0] out_id_25__din;
  wire out_id_25__full_n;
  wire out_id_25__write;
  wire [65:0] out_id_26__dout;
  wire out_id_26__empty_n;
  wire out_id_26__read;
  wire [65:0] out_id_26__din;
  wire out_id_26__full_n;
  wire out_id_26__write;
  wire [65:0] out_id_2__dout;
  wire out_id_2__empty_n;
  wire out_id_2__read;
  wire [65:0] out_id_2__din;
  wire out_id_2__full_n;
  wire out_id_2__write;
  wire [65:0] out_id_3__dout;
  wire out_id_3__empty_n;
  wire out_id_3__read;
  wire [65:0] out_id_3__din;
  wire out_id_3__full_n;
  wire out_id_3__write;
  wire [65:0] out_id_4__dout;
  wire out_id_4__empty_n;
  wire out_id_4__read;
  wire [65:0] out_id_4__din;
  wire out_id_4__full_n;
  wire out_id_4__write;
  wire [65:0] out_id_5__dout;
  wire out_id_5__empty_n;
  wire out_id_5__read;
  wire [65:0] out_id_5__din;
  wire out_id_5__full_n;
  wire out_id_5__write;
  wire [65:0] out_id_6__dout;
  wire out_id_6__empty_n;
  wire out_id_6__read;
  wire [65:0] out_id_6__din;
  wire out_id_6__full_n;
  wire out_id_6__write;
  wire [65:0] out_id_7__dout;
  wire out_id_7__empty_n;
  wire out_id_7__read;
  wire [65:0] out_id_7__din;
  wire out_id_7__full_n;
  wire out_id_7__write;
  wire [65:0] out_id_8__dout;
  wire out_id_8__empty_n;
  wire out_id_8__read;
  wire [65:0] out_id_8__din;
  wire out_id_8__full_n;
  wire out_id_8__write;
  wire [65:0] out_id_9__dout;
  wire out_id_9__empty_n;
  wire out_id_9__read;
  wire [65:0] out_id_9__din;
  wire out_id_9__full_n;
  wire out_id_9__write;
  wire krnl_globalSort_L1_L2_0__ap_start;
  wire krnl_globalSort_L1_L2_0__ap_ready;
  wire krnl_globalSort_L1_L2_0__ap_done;
  wire krnl_globalSort_L1_L2_0__ap_idle;
  wire krnl_globalSort_L1_L2_1__ap_start;
  wire krnl_globalSort_L1_L2_1__ap_ready;
  wire krnl_globalSort_L1_L2_1__ap_done;
  wire krnl_globalSort_L1_L2_1__ap_idle;
  wire krnl_globalSort_L1_L2_2__ap_start;
  wire krnl_globalSort_L1_L2_2__ap_ready;
  wire krnl_globalSort_L1_L2_2__ap_done;
  wire krnl_globalSort_L1_L2_2__ap_idle;
  wire krnl_globalSort_L1_L2_3__ap_start;
  wire krnl_globalSort_L1_L2_3__ap_ready;
  wire krnl_globalSort_L1_L2_3__ap_done;
  wire krnl_globalSort_L1_L2_3__ap_idle;
  wire krnl_globalSort_L1_L2_4__ap_start;
  wire krnl_globalSort_L1_L2_4__ap_ready;
  wire krnl_globalSort_L1_L2_4__ap_done;
  wire krnl_globalSort_L1_L2_4__ap_idle;
  wire krnl_globalSort_L1_L2_5__ap_start;
  wire krnl_globalSort_L1_L2_5__ap_ready;
  wire krnl_globalSort_L1_L2_5__ap_done;
  wire krnl_globalSort_L1_L2_5__ap_idle;
  wire krnl_globalSort_L1_L2_6__ap_start;
  wire krnl_globalSort_L1_L2_6__ap_ready;
  wire krnl_globalSort_L1_L2_6__ap_done;
  wire krnl_globalSort_L1_L2_6__ap_idle;
  wire krnl_globalSort_L1_L2_7__ap_start;
  wire krnl_globalSort_L1_L2_7__ap_ready;
  wire krnl_globalSort_L1_L2_7__ap_done;
  wire krnl_globalSort_L1_L2_7__ap_idle;
  wire krnl_globalSort_L1_L2_8__ap_start;
  wire krnl_globalSort_L1_L2_8__ap_ready;
  wire krnl_globalSort_L1_L2_8__ap_done;
  wire krnl_globalSort_L1_L2_8__ap_idle;
  wire krnl_globalSort_L1_L2_9__ap_start;
  wire krnl_globalSort_L1_L2_9__ap_ready;
  wire krnl_globalSort_L1_L2_9__ap_done;
  wire krnl_globalSort_L1_L2_9__ap_idle;
  wire krnl_globalSort_L1_L2_10__ap_start;
  wire krnl_globalSort_L1_L2_10__ap_ready;
  wire krnl_globalSort_L1_L2_10__ap_done;
  wire krnl_globalSort_L1_L2_10__ap_idle;
  wire krnl_globalSort_L1_L2_11__ap_start;
  wire krnl_globalSort_L1_L2_11__ap_ready;
  wire krnl_globalSort_L1_L2_11__ap_done;
  wire krnl_globalSort_L1_L2_11__ap_idle;
  wire krnl_globalSort_L1_L2_12__ap_start;
  wire krnl_globalSort_L1_L2_12__ap_ready;
  wire krnl_globalSort_L1_L2_12__ap_done;
  wire krnl_globalSort_L1_L2_12__ap_idle;
  wire [63:0] krnl_output_dist_id_0___L3_out_dist__q0;
  wire [63:0] L3_out_dist_read_addr__din;
  wire L3_out_dist_read_addr__full_n;
  wire L3_out_dist_read_addr__write;
  wire [31:0] L3_out_dist_read_data__dout;
  wire L3_out_dist_read_data__empty_n;
  wire L3_out_dist_read_data__read;
  wire [63:0] L3_out_dist_write_addr__din;
  wire L3_out_dist_write_addr__full_n;
  wire L3_out_dist_write_addr__write;
  wire [31:0] L3_out_dist_write_data__din;
  wire L3_out_dist_write_data__full_n;
  wire L3_out_dist_write_data__write;
  wire [7:0] L3_out_dist_write_resp__dout;
  wire L3_out_dist_write_resp__empty_n;
  wire L3_out_dist_write_resp__read;
  wire [63:0] krnl_output_dist_id_0___L3_out_id__q0;
  wire [63:0] L3_out_id_read_addr__din;
  wire L3_out_id_read_addr__full_n;
  wire L3_out_id_read_addr__write;
  wire [31:0] L3_out_id_read_data__dout;
  wire L3_out_id_read_data__empty_n;
  wire L3_out_id_read_data__read;
  wire [63:0] L3_out_id_write_addr__din;
  wire L3_out_id_write_addr__full_n;
  wire L3_out_id_write_addr__write;
  wire [31:0] L3_out_id_write_data__din;
  wire L3_out_id_write_data__full_n;
  wire L3_out_id_write_data__write;
  wire [7:0] L3_out_id_write_resp__dout;
  wire L3_out_id_write_resp__empty_n;
  wire L3_out_id_write_resp__read;
  wire krnl_output_dist_id_0__ap_start;
  wire krnl_output_dist_id_0__ap_ready;
  wire krnl_output_dist_id_0__ap_done;
  wire krnl_output_dist_id_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_0_0___in_0__q0;
  wire [63:0] in_0_read_addr__din;
  wire in_0_read_addr__full_n;
  wire in_0_read_addr__write;
  wire [255:0] in_0_read_data__dout;
  wire in_0_read_data__empty_n;
  wire in_0_read_data__read;
  wire [63:0] in_0_write_addr__din;
  wire in_0_write_addr__full_n;
  wire in_0_write_addr__write;
  wire [255:0] in_0_write_data__din;
  wire in_0_write_data__full_n;
  wire in_0_write_data__write;
  wire [7:0] in_0_write_resp__dout;
  wire in_0_write_resp__empty_n;
  wire in_0_write_resp__read;
  wire krnl_partialKnn_wrapper_0_0__ap_start;
  wire krnl_partialKnn_wrapper_0_0__ap_ready;
  wire krnl_partialKnn_wrapper_0_0__ap_done;
  wire krnl_partialKnn_wrapper_0_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_1_0___in_1__q0;
  wire [63:0] in_1_read_addr__din;
  wire in_1_read_addr__full_n;
  wire in_1_read_addr__write;
  wire [255:0] in_1_read_data__dout;
  wire in_1_read_data__empty_n;
  wire in_1_read_data__read;
  wire [63:0] in_1_write_addr__din;
  wire in_1_write_addr__full_n;
  wire in_1_write_addr__write;
  wire [255:0] in_1_write_data__din;
  wire in_1_write_data__full_n;
  wire in_1_write_data__write;
  wire [7:0] in_1_write_resp__dout;
  wire in_1_write_resp__empty_n;
  wire in_1_write_resp__read;
  wire krnl_partialKnn_wrapper_1_0__ap_start;
  wire krnl_partialKnn_wrapper_1_0__ap_ready;
  wire krnl_partialKnn_wrapper_1_0__ap_done;
  wire krnl_partialKnn_wrapper_1_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_10_0___in_10__q0;
  wire [63:0] in_10_read_addr__din;
  wire in_10_read_addr__full_n;
  wire in_10_read_addr__write;
  wire [255:0] in_10_read_data__dout;
  wire in_10_read_data__empty_n;
  wire in_10_read_data__read;
  wire [63:0] in_10_write_addr__din;
  wire in_10_write_addr__full_n;
  wire in_10_write_addr__write;
  wire [255:0] in_10_write_data__din;
  wire in_10_write_data__full_n;
  wire in_10_write_data__write;
  wire [7:0] in_10_write_resp__dout;
  wire in_10_write_resp__empty_n;
  wire in_10_write_resp__read;
  wire krnl_partialKnn_wrapper_10_0__ap_start;
  wire krnl_partialKnn_wrapper_10_0__ap_ready;
  wire krnl_partialKnn_wrapper_10_0__ap_done;
  wire krnl_partialKnn_wrapper_10_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_11_0___in_11__q0;
  wire [63:0] in_11_read_addr__din;
  wire in_11_read_addr__full_n;
  wire in_11_read_addr__write;
  wire [255:0] in_11_read_data__dout;
  wire in_11_read_data__empty_n;
  wire in_11_read_data__read;
  wire [63:0] in_11_write_addr__din;
  wire in_11_write_addr__full_n;
  wire in_11_write_addr__write;
  wire [255:0] in_11_write_data__din;
  wire in_11_write_data__full_n;
  wire in_11_write_data__write;
  wire [7:0] in_11_write_resp__dout;
  wire in_11_write_resp__empty_n;
  wire in_11_write_resp__read;
  wire krnl_partialKnn_wrapper_11_0__ap_start;
  wire krnl_partialKnn_wrapper_11_0__ap_ready;
  wire krnl_partialKnn_wrapper_11_0__ap_done;
  wire krnl_partialKnn_wrapper_11_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_12_0___in_12__q0;
  wire [63:0] in_12_read_addr__din;
  wire in_12_read_addr__full_n;
  wire in_12_read_addr__write;
  wire [255:0] in_12_read_data__dout;
  wire in_12_read_data__empty_n;
  wire in_12_read_data__read;
  wire [63:0] in_12_write_addr__din;
  wire in_12_write_addr__full_n;
  wire in_12_write_addr__write;
  wire [255:0] in_12_write_data__din;
  wire in_12_write_data__full_n;
  wire in_12_write_data__write;
  wire [7:0] in_12_write_resp__dout;
  wire in_12_write_resp__empty_n;
  wire in_12_write_resp__read;
  wire krnl_partialKnn_wrapper_12_0__ap_start;
  wire krnl_partialKnn_wrapper_12_0__ap_ready;
  wire krnl_partialKnn_wrapper_12_0__ap_done;
  wire krnl_partialKnn_wrapper_12_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_13_0___in_13__q0;
  wire [63:0] in_13_read_addr__din;
  wire in_13_read_addr__full_n;
  wire in_13_read_addr__write;
  wire [255:0] in_13_read_data__dout;
  wire in_13_read_data__empty_n;
  wire in_13_read_data__read;
  wire [63:0] in_13_write_addr__din;
  wire in_13_write_addr__full_n;
  wire in_13_write_addr__write;
  wire [255:0] in_13_write_data__din;
  wire in_13_write_data__full_n;
  wire in_13_write_data__write;
  wire [7:0] in_13_write_resp__dout;
  wire in_13_write_resp__empty_n;
  wire in_13_write_resp__read;
  wire krnl_partialKnn_wrapper_13_0__ap_start;
  wire krnl_partialKnn_wrapper_13_0__ap_ready;
  wire krnl_partialKnn_wrapper_13_0__ap_done;
  wire krnl_partialKnn_wrapper_13_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_14_0___in_14__q0;
  wire [63:0] in_14_read_addr__din;
  wire in_14_read_addr__full_n;
  wire in_14_read_addr__write;
  wire [255:0] in_14_read_data__dout;
  wire in_14_read_data__empty_n;
  wire in_14_read_data__read;
  wire [63:0] in_14_write_addr__din;
  wire in_14_write_addr__full_n;
  wire in_14_write_addr__write;
  wire [255:0] in_14_write_data__din;
  wire in_14_write_data__full_n;
  wire in_14_write_data__write;
  wire [7:0] in_14_write_resp__dout;
  wire in_14_write_resp__empty_n;
  wire in_14_write_resp__read;
  wire krnl_partialKnn_wrapper_14_0__ap_start;
  wire krnl_partialKnn_wrapper_14_0__ap_ready;
  wire krnl_partialKnn_wrapper_14_0__ap_done;
  wire krnl_partialKnn_wrapper_14_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_15_0___in_15__q0;
  wire [63:0] in_15_read_addr__din;
  wire in_15_read_addr__full_n;
  wire in_15_read_addr__write;
  wire [255:0] in_15_read_data__dout;
  wire in_15_read_data__empty_n;
  wire in_15_read_data__read;
  wire [63:0] in_15_write_addr__din;
  wire in_15_write_addr__full_n;
  wire in_15_write_addr__write;
  wire [255:0] in_15_write_data__din;
  wire in_15_write_data__full_n;
  wire in_15_write_data__write;
  wire [7:0] in_15_write_resp__dout;
  wire in_15_write_resp__empty_n;
  wire in_15_write_resp__read;
  wire krnl_partialKnn_wrapper_15_0__ap_start;
  wire krnl_partialKnn_wrapper_15_0__ap_ready;
  wire krnl_partialKnn_wrapper_15_0__ap_done;
  wire krnl_partialKnn_wrapper_15_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_16_0___in_16__q0;
  wire [63:0] in_16_read_addr__din;
  wire in_16_read_addr__full_n;
  wire in_16_read_addr__write;
  wire [255:0] in_16_read_data__dout;
  wire in_16_read_data__empty_n;
  wire in_16_read_data__read;
  wire [63:0] in_16_write_addr__din;
  wire in_16_write_addr__full_n;
  wire in_16_write_addr__write;
  wire [255:0] in_16_write_data__din;
  wire in_16_write_data__full_n;
  wire in_16_write_data__write;
  wire [7:0] in_16_write_resp__dout;
  wire in_16_write_resp__empty_n;
  wire in_16_write_resp__read;
  wire krnl_partialKnn_wrapper_16_0__ap_start;
  wire krnl_partialKnn_wrapper_16_0__ap_ready;
  wire krnl_partialKnn_wrapper_16_0__ap_done;
  wire krnl_partialKnn_wrapper_16_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_17_0___in_17__q0;
  wire [63:0] in_17_read_addr__din;
  wire in_17_read_addr__full_n;
  wire in_17_read_addr__write;
  wire [255:0] in_17_read_data__dout;
  wire in_17_read_data__empty_n;
  wire in_17_read_data__read;
  wire [63:0] in_17_write_addr__din;
  wire in_17_write_addr__full_n;
  wire in_17_write_addr__write;
  wire [255:0] in_17_write_data__din;
  wire in_17_write_data__full_n;
  wire in_17_write_data__write;
  wire [7:0] in_17_write_resp__dout;
  wire in_17_write_resp__empty_n;
  wire in_17_write_resp__read;
  wire krnl_partialKnn_wrapper_17_0__ap_start;
  wire krnl_partialKnn_wrapper_17_0__ap_ready;
  wire krnl_partialKnn_wrapper_17_0__ap_done;
  wire krnl_partialKnn_wrapper_17_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_18_0___in_18__q0;
  wire [63:0] in_18_read_addr__din;
  wire in_18_read_addr__full_n;
  wire in_18_read_addr__write;
  wire [255:0] in_18_read_data__dout;
  wire in_18_read_data__empty_n;
  wire in_18_read_data__read;
  wire [63:0] in_18_write_addr__din;
  wire in_18_write_addr__full_n;
  wire in_18_write_addr__write;
  wire [255:0] in_18_write_data__din;
  wire in_18_write_data__full_n;
  wire in_18_write_data__write;
  wire [7:0] in_18_write_resp__dout;
  wire in_18_write_resp__empty_n;
  wire in_18_write_resp__read;
  wire krnl_partialKnn_wrapper_18_0__ap_start;
  wire krnl_partialKnn_wrapper_18_0__ap_ready;
  wire krnl_partialKnn_wrapper_18_0__ap_done;
  wire krnl_partialKnn_wrapper_18_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_19_0___in_19__q0;
  wire [63:0] in_19_read_addr__din;
  wire in_19_read_addr__full_n;
  wire in_19_read_addr__write;
  wire [255:0] in_19_read_data__dout;
  wire in_19_read_data__empty_n;
  wire in_19_read_data__read;
  wire [63:0] in_19_write_addr__din;
  wire in_19_write_addr__full_n;
  wire in_19_write_addr__write;
  wire [255:0] in_19_write_data__din;
  wire in_19_write_data__full_n;
  wire in_19_write_data__write;
  wire [7:0] in_19_write_resp__dout;
  wire in_19_write_resp__empty_n;
  wire in_19_write_resp__read;
  wire krnl_partialKnn_wrapper_19_0__ap_start;
  wire krnl_partialKnn_wrapper_19_0__ap_ready;
  wire krnl_partialKnn_wrapper_19_0__ap_done;
  wire krnl_partialKnn_wrapper_19_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_2_0___in_2__q0;
  wire [63:0] in_2_read_addr__din;
  wire in_2_read_addr__full_n;
  wire in_2_read_addr__write;
  wire [255:0] in_2_read_data__dout;
  wire in_2_read_data__empty_n;
  wire in_2_read_data__read;
  wire [63:0] in_2_write_addr__din;
  wire in_2_write_addr__full_n;
  wire in_2_write_addr__write;
  wire [255:0] in_2_write_data__din;
  wire in_2_write_data__full_n;
  wire in_2_write_data__write;
  wire [7:0] in_2_write_resp__dout;
  wire in_2_write_resp__empty_n;
  wire in_2_write_resp__read;
  wire krnl_partialKnn_wrapper_2_0__ap_start;
  wire krnl_partialKnn_wrapper_2_0__ap_ready;
  wire krnl_partialKnn_wrapper_2_0__ap_done;
  wire krnl_partialKnn_wrapper_2_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_20_0___in_20__q0;
  wire [63:0] in_20_read_addr__din;
  wire in_20_read_addr__full_n;
  wire in_20_read_addr__write;
  wire [255:0] in_20_read_data__dout;
  wire in_20_read_data__empty_n;
  wire in_20_read_data__read;
  wire [63:0] in_20_write_addr__din;
  wire in_20_write_addr__full_n;
  wire in_20_write_addr__write;
  wire [255:0] in_20_write_data__din;
  wire in_20_write_data__full_n;
  wire in_20_write_data__write;
  wire [7:0] in_20_write_resp__dout;
  wire in_20_write_resp__empty_n;
  wire in_20_write_resp__read;
  wire krnl_partialKnn_wrapper_20_0__ap_start;
  wire krnl_partialKnn_wrapper_20_0__ap_ready;
  wire krnl_partialKnn_wrapper_20_0__ap_done;
  wire krnl_partialKnn_wrapper_20_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_21_0___in_21__q0;
  wire [63:0] in_21_read_addr__din;
  wire in_21_read_addr__full_n;
  wire in_21_read_addr__write;
  wire [255:0] in_21_read_data__dout;
  wire in_21_read_data__empty_n;
  wire in_21_read_data__read;
  wire [63:0] in_21_write_addr__din;
  wire in_21_write_addr__full_n;
  wire in_21_write_addr__write;
  wire [255:0] in_21_write_data__din;
  wire in_21_write_data__full_n;
  wire in_21_write_data__write;
  wire [7:0] in_21_write_resp__dout;
  wire in_21_write_resp__empty_n;
  wire in_21_write_resp__read;
  wire krnl_partialKnn_wrapper_21_0__ap_start;
  wire krnl_partialKnn_wrapper_21_0__ap_ready;
  wire krnl_partialKnn_wrapper_21_0__ap_done;
  wire krnl_partialKnn_wrapper_21_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_22_0___in_22__q0;
  wire [63:0] in_22_read_addr__din;
  wire in_22_read_addr__full_n;
  wire in_22_read_addr__write;
  wire [255:0] in_22_read_data__dout;
  wire in_22_read_data__empty_n;
  wire in_22_read_data__read;
  wire [63:0] in_22_write_addr__din;
  wire in_22_write_addr__full_n;
  wire in_22_write_addr__write;
  wire [255:0] in_22_write_data__din;
  wire in_22_write_data__full_n;
  wire in_22_write_data__write;
  wire [7:0] in_22_write_resp__dout;
  wire in_22_write_resp__empty_n;
  wire in_22_write_resp__read;
  wire krnl_partialKnn_wrapper_22_0__ap_start;
  wire krnl_partialKnn_wrapper_22_0__ap_ready;
  wire krnl_partialKnn_wrapper_22_0__ap_done;
  wire krnl_partialKnn_wrapper_22_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_23_0___in_23__q0;
  wire [63:0] in_23_read_addr__din;
  wire in_23_read_addr__full_n;
  wire in_23_read_addr__write;
  wire [255:0] in_23_read_data__dout;
  wire in_23_read_data__empty_n;
  wire in_23_read_data__read;
  wire [63:0] in_23_write_addr__din;
  wire in_23_write_addr__full_n;
  wire in_23_write_addr__write;
  wire [255:0] in_23_write_data__din;
  wire in_23_write_data__full_n;
  wire in_23_write_data__write;
  wire [7:0] in_23_write_resp__dout;
  wire in_23_write_resp__empty_n;
  wire in_23_write_resp__read;
  wire krnl_partialKnn_wrapper_23_0__ap_start;
  wire krnl_partialKnn_wrapper_23_0__ap_ready;
  wire krnl_partialKnn_wrapper_23_0__ap_done;
  wire krnl_partialKnn_wrapper_23_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_24_0___in_24__q0;
  wire [63:0] in_24_read_addr__din;
  wire in_24_read_addr__full_n;
  wire in_24_read_addr__write;
  wire [255:0] in_24_read_data__dout;
  wire in_24_read_data__empty_n;
  wire in_24_read_data__read;
  wire [63:0] in_24_write_addr__din;
  wire in_24_write_addr__full_n;
  wire in_24_write_addr__write;
  wire [255:0] in_24_write_data__din;
  wire in_24_write_data__full_n;
  wire in_24_write_data__write;
  wire [7:0] in_24_write_resp__dout;
  wire in_24_write_resp__empty_n;
  wire in_24_write_resp__read;
  wire krnl_partialKnn_wrapper_24_0__ap_start;
  wire krnl_partialKnn_wrapper_24_0__ap_ready;
  wire krnl_partialKnn_wrapper_24_0__ap_done;
  wire krnl_partialKnn_wrapper_24_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_25_0___in_25__q0;
  wire [63:0] in_25_read_addr__din;
  wire in_25_read_addr__full_n;
  wire in_25_read_addr__write;
  wire [255:0] in_25_read_data__dout;
  wire in_25_read_data__empty_n;
  wire in_25_read_data__read;
  wire [63:0] in_25_write_addr__din;
  wire in_25_write_addr__full_n;
  wire in_25_write_addr__write;
  wire [255:0] in_25_write_data__din;
  wire in_25_write_data__full_n;
  wire in_25_write_data__write;
  wire [7:0] in_25_write_resp__dout;
  wire in_25_write_resp__empty_n;
  wire in_25_write_resp__read;
  wire krnl_partialKnn_wrapper_25_0__ap_start;
  wire krnl_partialKnn_wrapper_25_0__ap_ready;
  wire krnl_partialKnn_wrapper_25_0__ap_done;
  wire krnl_partialKnn_wrapper_25_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_26_0___in_26__q0;
  wire [63:0] in_26_read_addr__din;
  wire in_26_read_addr__full_n;
  wire in_26_read_addr__write;
  wire [255:0] in_26_read_data__dout;
  wire in_26_read_data__empty_n;
  wire in_26_read_data__read;
  wire [63:0] in_26_write_addr__din;
  wire in_26_write_addr__full_n;
  wire in_26_write_addr__write;
  wire [255:0] in_26_write_data__din;
  wire in_26_write_data__full_n;
  wire in_26_write_data__write;
  wire [7:0] in_26_write_resp__dout;
  wire in_26_write_resp__empty_n;
  wire in_26_write_resp__read;
  wire krnl_partialKnn_wrapper_26_0__ap_start;
  wire krnl_partialKnn_wrapper_26_0__ap_ready;
  wire krnl_partialKnn_wrapper_26_0__ap_done;
  wire krnl_partialKnn_wrapper_26_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_3_0___in_3__q0;
  wire [63:0] in_3_read_addr__din;
  wire in_3_read_addr__full_n;
  wire in_3_read_addr__write;
  wire [255:0] in_3_read_data__dout;
  wire in_3_read_data__empty_n;
  wire in_3_read_data__read;
  wire [63:0] in_3_write_addr__din;
  wire in_3_write_addr__full_n;
  wire in_3_write_addr__write;
  wire [255:0] in_3_write_data__din;
  wire in_3_write_data__full_n;
  wire in_3_write_data__write;
  wire [7:0] in_3_write_resp__dout;
  wire in_3_write_resp__empty_n;
  wire in_3_write_resp__read;
  wire krnl_partialKnn_wrapper_3_0__ap_start;
  wire krnl_partialKnn_wrapper_3_0__ap_ready;
  wire krnl_partialKnn_wrapper_3_0__ap_done;
  wire krnl_partialKnn_wrapper_3_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_4_0___in_4__q0;
  wire [63:0] in_4_read_addr__din;
  wire in_4_read_addr__full_n;
  wire in_4_read_addr__write;
  wire [255:0] in_4_read_data__dout;
  wire in_4_read_data__empty_n;
  wire in_4_read_data__read;
  wire [63:0] in_4_write_addr__din;
  wire in_4_write_addr__full_n;
  wire in_4_write_addr__write;
  wire [255:0] in_4_write_data__din;
  wire in_4_write_data__full_n;
  wire in_4_write_data__write;
  wire [7:0] in_4_write_resp__dout;
  wire in_4_write_resp__empty_n;
  wire in_4_write_resp__read;
  wire krnl_partialKnn_wrapper_4_0__ap_start;
  wire krnl_partialKnn_wrapper_4_0__ap_ready;
  wire krnl_partialKnn_wrapper_4_0__ap_done;
  wire krnl_partialKnn_wrapper_4_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_5_0___in_5__q0;
  wire [63:0] in_5_read_addr__din;
  wire in_5_read_addr__full_n;
  wire in_5_read_addr__write;
  wire [255:0] in_5_read_data__dout;
  wire in_5_read_data__empty_n;
  wire in_5_read_data__read;
  wire [63:0] in_5_write_addr__din;
  wire in_5_write_addr__full_n;
  wire in_5_write_addr__write;
  wire [255:0] in_5_write_data__din;
  wire in_5_write_data__full_n;
  wire in_5_write_data__write;
  wire [7:0] in_5_write_resp__dout;
  wire in_5_write_resp__empty_n;
  wire in_5_write_resp__read;
  wire krnl_partialKnn_wrapper_5_0__ap_start;
  wire krnl_partialKnn_wrapper_5_0__ap_ready;
  wire krnl_partialKnn_wrapper_5_0__ap_done;
  wire krnl_partialKnn_wrapper_5_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_6_0___in_6__q0;
  wire [63:0] in_6_read_addr__din;
  wire in_6_read_addr__full_n;
  wire in_6_read_addr__write;
  wire [255:0] in_6_read_data__dout;
  wire in_6_read_data__empty_n;
  wire in_6_read_data__read;
  wire [63:0] in_6_write_addr__din;
  wire in_6_write_addr__full_n;
  wire in_6_write_addr__write;
  wire [255:0] in_6_write_data__din;
  wire in_6_write_data__full_n;
  wire in_6_write_data__write;
  wire [7:0] in_6_write_resp__dout;
  wire in_6_write_resp__empty_n;
  wire in_6_write_resp__read;
  wire krnl_partialKnn_wrapper_6_0__ap_start;
  wire krnl_partialKnn_wrapper_6_0__ap_ready;
  wire krnl_partialKnn_wrapper_6_0__ap_done;
  wire krnl_partialKnn_wrapper_6_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_7_0___in_7__q0;
  wire [63:0] in_7_read_addr__din;
  wire in_7_read_addr__full_n;
  wire in_7_read_addr__write;
  wire [255:0] in_7_read_data__dout;
  wire in_7_read_data__empty_n;
  wire in_7_read_data__read;
  wire [63:0] in_7_write_addr__din;
  wire in_7_write_addr__full_n;
  wire in_7_write_addr__write;
  wire [255:0] in_7_write_data__din;
  wire in_7_write_data__full_n;
  wire in_7_write_data__write;
  wire [7:0] in_7_write_resp__dout;
  wire in_7_write_resp__empty_n;
  wire in_7_write_resp__read;
  wire krnl_partialKnn_wrapper_7_0__ap_start;
  wire krnl_partialKnn_wrapper_7_0__ap_ready;
  wire krnl_partialKnn_wrapper_7_0__ap_done;
  wire krnl_partialKnn_wrapper_7_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_8_0___in_8__q0;
  wire [63:0] in_8_read_addr__din;
  wire in_8_read_addr__full_n;
  wire in_8_read_addr__write;
  wire [255:0] in_8_read_data__dout;
  wire in_8_read_data__empty_n;
  wire in_8_read_data__read;
  wire [63:0] in_8_write_addr__din;
  wire in_8_write_addr__full_n;
  wire in_8_write_addr__write;
  wire [255:0] in_8_write_data__din;
  wire in_8_write_data__full_n;
  wire in_8_write_data__write;
  wire [7:0] in_8_write_resp__dout;
  wire in_8_write_resp__empty_n;
  wire in_8_write_resp__read;
  wire krnl_partialKnn_wrapper_8_0__ap_start;
  wire krnl_partialKnn_wrapper_8_0__ap_ready;
  wire krnl_partialKnn_wrapper_8_0__ap_done;
  wire krnl_partialKnn_wrapper_8_0__ap_idle;
  wire [63:0] krnl_partialKnn_wrapper_9_0___in_9__q0;
  wire [63:0] in_9_read_addr__din;
  wire in_9_read_addr__full_n;
  wire in_9_read_addr__write;
  wire [255:0] in_9_read_data__dout;
  wire in_9_read_data__empty_n;
  wire in_9_read_data__read;
  wire [63:0] in_9_write_addr__din;
  wire in_9_write_addr__full_n;
  wire in_9_write_addr__write;
  wire [255:0] in_9_write_data__din;
  wire in_9_write_data__full_n;
  wire in_9_write_data__write;
  wire [7:0] in_9_write_resp__dout;
  wire in_9_write_resp__empty_n;
  wire in_9_write_resp__read;
  wire krnl_partialKnn_wrapper_9_0__ap_start;
  wire krnl_partialKnn_wrapper_9_0__ap_ready;
  wire krnl_partialKnn_wrapper_9_0__ap_done;
  wire krnl_partialKnn_wrapper_9_0__ap_idle;
  wire ap_rst_n_inv;
  wire ap_done;
  wire ap_idle;
  wire ap_ready;
  assign ap_rst_n_inv = (~ap_rst_n);
  assign control_s_axi_U_ACLK = ap_clk;
  assign control_s_axi_U_ACLK_EN = 1'b1;
  assign control_s_axi_U_ARADDR = s_axi_control_ARADDR;
  assign control_s_axi_U_ARESET = ap_rst_n_inv;
  assign s_axi_control_ARREADY = control_s_axi_U_ARREADY;
  assign control_s_axi_U_ARVALID = s_axi_control_ARVALID;
  assign control_s_axi_U_AWADDR = s_axi_control_AWADDR;
  assign s_axi_control_AWREADY = control_s_axi_U_AWREADY;
  assign control_s_axi_U_AWVALID = s_axi_control_AWVALID;
  assign control_s_axi_U_BREADY = s_axi_control_BREADY;
  assign s_axi_control_BRESP = control_s_axi_U_BRESP;
  assign s_axi_control_BVALID = control_s_axi_U_BVALID;
  assign L3_out_dist = control_s_axi_U_L3_out_dist;
  assign L3_out_id = control_s_axi_U_L3_out_id;
  assign s_axi_control_RDATA = control_s_axi_U_RDATA;
  assign control_s_axi_U_RREADY = s_axi_control_RREADY;
  assign s_axi_control_RRESP = control_s_axi_U_RRESP;
  assign s_axi_control_RVALID = control_s_axi_U_RVALID;
  assign control_s_axi_U_WDATA = s_axi_control_WDATA;
  assign s_axi_control_WREADY = control_s_axi_U_WREADY;
  assign control_s_axi_U_WSTRB = s_axi_control_WSTRB;
  assign control_s_axi_U_WVALID = s_axi_control_WVALID;
  assign control_s_axi_U_ap_done = ap_done;
  assign control_s_axi_U_ap_idle = ap_idle;
  assign control_s_axi_U_ap_ready = ap_ready;
  assign ap_start = control_s_axi_U_ap_start;
  assign in_0 = control_s_axi_U_in_0;
  assign in_1 = control_s_axi_U_in_1;
  assign in_10 = control_s_axi_U_in_10;
  assign in_11 = control_s_axi_U_in_11;
  assign in_12 = control_s_axi_U_in_12;
  assign in_13 = control_s_axi_U_in_13;
  assign in_14 = control_s_axi_U_in_14;
  assign in_15 = control_s_axi_U_in_15;
  assign in_16 = control_s_axi_U_in_16;
  assign in_17 = control_s_axi_U_in_17;
  assign in_18 = control_s_axi_U_in_18;
  assign in_19 = control_s_axi_U_in_19;
  assign in_2 = control_s_axi_U_in_2;
  assign in_20 = control_s_axi_U_in_20;
  assign in_21 = control_s_axi_U_in_21;
  assign in_22 = control_s_axi_U_in_22;
  assign in_23 = control_s_axi_U_in_23;
  assign in_24 = control_s_axi_U_in_24;
  assign in_25 = control_s_axi_U_in_25;
  assign in_26 = control_s_axi_U_in_26;
  assign in_3 = control_s_axi_U_in_3;
  assign in_4 = control_s_axi_U_in_4;
  assign in_5 = control_s_axi_U_in_5;
  assign in_6 = control_s_axi_U_in_6;
  assign in_7 = control_s_axi_U_in_7;
  assign in_8 = control_s_axi_U_in_8;
  assign in_9 = control_s_axi_U_in_9;
  assign interrupt = control_s_axi_U_interrupt;
  assign L1_out_dist_0_clk = ap_clk;
  assign L1_out_dist_0_if_din = L1_out_dist_0__din;
  assign L1_out_dist_0__dout = L1_out_dist_0_if_dout;
  assign L1_out_dist_0__empty_n = L1_out_dist_0_if_empty_n;
  assign L1_out_dist_0__full_n = L1_out_dist_0_if_full_n;
  assign L1_out_dist_0_if_read = L1_out_dist_0__read;
  assign L1_out_dist_0_if_read_ce = 1'b1;
  assign L1_out_dist_0_if_write = L1_out_dist_0__write;
  assign L1_out_dist_0_if_write_ce = 1'b1;
  assign L1_out_dist_0_reset = ~ ap_rst_n;
  assign L1_out_dist_1_clk = ap_clk;
  assign L1_out_dist_1_if_din = L1_out_dist_1__din;
  assign L1_out_dist_1__dout = L1_out_dist_1_if_dout;
  assign L1_out_dist_1__empty_n = L1_out_dist_1_if_empty_n;
  assign L1_out_dist_1__full_n = L1_out_dist_1_if_full_n;
  assign L1_out_dist_1_if_read = L1_out_dist_1__read;
  assign L1_out_dist_1_if_read_ce = 1'b1;
  assign L1_out_dist_1_if_write = L1_out_dist_1__write;
  assign L1_out_dist_1_if_write_ce = 1'b1;
  assign L1_out_dist_1_reset = ~ ap_rst_n;
  assign L1_out_dist_2_clk = ap_clk;
  assign L1_out_dist_2_if_din = L1_out_dist_2__din;
  assign L1_out_dist_2__dout = L1_out_dist_2_if_dout;
  assign L1_out_dist_2__empty_n = L1_out_dist_2_if_empty_n;
  assign L1_out_dist_2__full_n = L1_out_dist_2_if_full_n;
  assign L1_out_dist_2_if_read = L1_out_dist_2__read;
  assign L1_out_dist_2_if_read_ce = 1'b1;
  assign L1_out_dist_2_if_write = L1_out_dist_2__write;
  assign L1_out_dist_2_if_write_ce = 1'b1;
  assign L1_out_dist_2_reset = ~ ap_rst_n;
  assign L1_out_dist_3_clk = ap_clk;
  assign L1_out_dist_3_if_din = L1_out_dist_3__din;
  assign L1_out_dist_3__dout = L1_out_dist_3_if_dout;
  assign L1_out_dist_3__empty_n = L1_out_dist_3_if_empty_n;
  assign L1_out_dist_3__full_n = L1_out_dist_3_if_full_n;
  assign L1_out_dist_3_if_read = L1_out_dist_3__read;
  assign L1_out_dist_3_if_read_ce = 1'b1;
  assign L1_out_dist_3_if_write = L1_out_dist_3__write;
  assign L1_out_dist_3_if_write_ce = 1'b1;
  assign L1_out_dist_3_reset = ~ ap_rst_n;
  assign L1_out_dist_4_clk = ap_clk;
  assign L1_out_dist_4_if_din = L1_out_dist_4__din;
  assign L1_out_dist_4__dout = L1_out_dist_4_if_dout;
  assign L1_out_dist_4__empty_n = L1_out_dist_4_if_empty_n;
  assign L1_out_dist_4__full_n = L1_out_dist_4_if_full_n;
  assign L1_out_dist_4_if_read = L1_out_dist_4__read;
  assign L1_out_dist_4_if_read_ce = 1'b1;
  assign L1_out_dist_4_if_write = L1_out_dist_4__write;
  assign L1_out_dist_4_if_write_ce = 1'b1;
  assign L1_out_dist_4_reset = ~ ap_rst_n;
  assign L1_out_dist_5_clk = ap_clk;
  assign L1_out_dist_5_if_din = L1_out_dist_5__din;
  assign L1_out_dist_5__dout = L1_out_dist_5_if_dout;
  assign L1_out_dist_5__empty_n = L1_out_dist_5_if_empty_n;
  assign L1_out_dist_5__full_n = L1_out_dist_5_if_full_n;
  assign L1_out_dist_5_if_read = L1_out_dist_5__read;
  assign L1_out_dist_5_if_read_ce = 1'b1;
  assign L1_out_dist_5_if_write = L1_out_dist_5__write;
  assign L1_out_dist_5_if_write_ce = 1'b1;
  assign L1_out_dist_5_reset = ~ ap_rst_n;
  assign L1_out_dist_6_clk = ap_clk;
  assign L1_out_dist_6_if_din = L1_out_dist_6__din;
  assign L1_out_dist_6__dout = L1_out_dist_6_if_dout;
  assign L1_out_dist_6__empty_n = L1_out_dist_6_if_empty_n;
  assign L1_out_dist_6__full_n = L1_out_dist_6_if_full_n;
  assign L1_out_dist_6_if_read = L1_out_dist_6__read;
  assign L1_out_dist_6_if_read_ce = 1'b1;
  assign L1_out_dist_6_if_write = L1_out_dist_6__write;
  assign L1_out_dist_6_if_write_ce = 1'b1;
  assign L1_out_dist_6_reset = ~ ap_rst_n;
  assign L1_out_dist_7_clk = ap_clk;
  assign L1_out_dist_7_if_din = L1_out_dist_7__din;
  assign L1_out_dist_7__dout = L1_out_dist_7_if_dout;
  assign L1_out_dist_7__empty_n = L1_out_dist_7_if_empty_n;
  assign L1_out_dist_7__full_n = L1_out_dist_7_if_full_n;
  assign L1_out_dist_7_if_read = L1_out_dist_7__read;
  assign L1_out_dist_7_if_read_ce = 1'b1;
  assign L1_out_dist_7_if_write = L1_out_dist_7__write;
  assign L1_out_dist_7_if_write_ce = 1'b1;
  assign L1_out_dist_7_reset = ~ ap_rst_n;
  assign L1_out_dist_8_clk = ap_clk;
  assign L1_out_dist_8_if_din = L1_out_dist_8__din;
  assign L1_out_dist_8__dout = L1_out_dist_8_if_dout;
  assign L1_out_dist_8__empty_n = L1_out_dist_8_if_empty_n;
  assign L1_out_dist_8__full_n = L1_out_dist_8_if_full_n;
  assign L1_out_dist_8_if_read = L1_out_dist_8__read;
  assign L1_out_dist_8_if_read_ce = 1'b1;
  assign L1_out_dist_8_if_write = L1_out_dist_8__write;
  assign L1_out_dist_8_if_write_ce = 1'b1;
  assign L1_out_dist_8_reset = ~ ap_rst_n;
  assign L1_out_id_0_clk = ap_clk;
  assign L1_out_id_0_if_din = L1_out_id_0__din;
  assign L1_out_id_0__dout = L1_out_id_0_if_dout;
  assign L1_out_id_0__empty_n = L1_out_id_0_if_empty_n;
  assign L1_out_id_0__full_n = L1_out_id_0_if_full_n;
  assign L1_out_id_0_if_read = L1_out_id_0__read;
  assign L1_out_id_0_if_read_ce = 1'b1;
  assign L1_out_id_0_if_write = L1_out_id_0__write;
  assign L1_out_id_0_if_write_ce = 1'b1;
  assign L1_out_id_0_reset = ~ ap_rst_n;
  assign L1_out_id_1_clk = ap_clk;
  assign L1_out_id_1_if_din = L1_out_id_1__din;
  assign L1_out_id_1__dout = L1_out_id_1_if_dout;
  assign L1_out_id_1__empty_n = L1_out_id_1_if_empty_n;
  assign L1_out_id_1__full_n = L1_out_id_1_if_full_n;
  assign L1_out_id_1_if_read = L1_out_id_1__read;
  assign L1_out_id_1_if_read_ce = 1'b1;
  assign L1_out_id_1_if_write = L1_out_id_1__write;
  assign L1_out_id_1_if_write_ce = 1'b1;
  assign L1_out_id_1_reset = ~ ap_rst_n;
  assign L1_out_id_2_clk = ap_clk;
  assign L1_out_id_2_if_din = L1_out_id_2__din;
  assign L1_out_id_2__dout = L1_out_id_2_if_dout;
  assign L1_out_id_2__empty_n = L1_out_id_2_if_empty_n;
  assign L1_out_id_2__full_n = L1_out_id_2_if_full_n;
  assign L1_out_id_2_if_read = L1_out_id_2__read;
  assign L1_out_id_2_if_read_ce = 1'b1;
  assign L1_out_id_2_if_write = L1_out_id_2__write;
  assign L1_out_id_2_if_write_ce = 1'b1;
  assign L1_out_id_2_reset = ~ ap_rst_n;
  assign L1_out_id_3_clk = ap_clk;
  assign L1_out_id_3_if_din = L1_out_id_3__din;
  assign L1_out_id_3__dout = L1_out_id_3_if_dout;
  assign L1_out_id_3__empty_n = L1_out_id_3_if_empty_n;
  assign L1_out_id_3__full_n = L1_out_id_3_if_full_n;
  assign L1_out_id_3_if_read = L1_out_id_3__read;
  assign L1_out_id_3_if_read_ce = 1'b1;
  assign L1_out_id_3_if_write = L1_out_id_3__write;
  assign L1_out_id_3_if_write_ce = 1'b1;
  assign L1_out_id_3_reset = ~ ap_rst_n;
  assign L1_out_id_4_clk = ap_clk;
  assign L1_out_id_4_if_din = L1_out_id_4__din;
  assign L1_out_id_4__dout = L1_out_id_4_if_dout;
  assign L1_out_id_4__empty_n = L1_out_id_4_if_empty_n;
  assign L1_out_id_4__full_n = L1_out_id_4_if_full_n;
  assign L1_out_id_4_if_read = L1_out_id_4__read;
  assign L1_out_id_4_if_read_ce = 1'b1;
  assign L1_out_id_4_if_write = L1_out_id_4__write;
  assign L1_out_id_4_if_write_ce = 1'b1;
  assign L1_out_id_4_reset = ~ ap_rst_n;
  assign L1_out_id_5_clk = ap_clk;
  assign L1_out_id_5_if_din = L1_out_id_5__din;
  assign L1_out_id_5__dout = L1_out_id_5_if_dout;
  assign L1_out_id_5__empty_n = L1_out_id_5_if_empty_n;
  assign L1_out_id_5__full_n = L1_out_id_5_if_full_n;
  assign L1_out_id_5_if_read = L1_out_id_5__read;
  assign L1_out_id_5_if_read_ce = 1'b1;
  assign L1_out_id_5_if_write = L1_out_id_5__write;
  assign L1_out_id_5_if_write_ce = 1'b1;
  assign L1_out_id_5_reset = ~ ap_rst_n;
  assign L1_out_id_6_clk = ap_clk;
  assign L1_out_id_6_if_din = L1_out_id_6__din;
  assign L1_out_id_6__dout = L1_out_id_6_if_dout;
  assign L1_out_id_6__empty_n = L1_out_id_6_if_empty_n;
  assign L1_out_id_6__full_n = L1_out_id_6_if_full_n;
  assign L1_out_id_6_if_read = L1_out_id_6__read;
  assign L1_out_id_6_if_read_ce = 1'b1;
  assign L1_out_id_6_if_write = L1_out_id_6__write;
  assign L1_out_id_6_if_write_ce = 1'b1;
  assign L1_out_id_6_reset = ~ ap_rst_n;
  assign L1_out_id_7_clk = ap_clk;
  assign L1_out_id_7_if_din = L1_out_id_7__din;
  assign L1_out_id_7__dout = L1_out_id_7_if_dout;
  assign L1_out_id_7__empty_n = L1_out_id_7_if_empty_n;
  assign L1_out_id_7__full_n = L1_out_id_7_if_full_n;
  assign L1_out_id_7_if_read = L1_out_id_7__read;
  assign L1_out_id_7_if_read_ce = 1'b1;
  assign L1_out_id_7_if_write = L1_out_id_7__write;
  assign L1_out_id_7_if_write_ce = 1'b1;
  assign L1_out_id_7_reset = ~ ap_rst_n;
  assign L1_out_id_8_clk = ap_clk;
  assign L1_out_id_8_if_din = L1_out_id_8__din;
  assign L1_out_id_8__dout = L1_out_id_8_if_dout;
  assign L1_out_id_8__empty_n = L1_out_id_8_if_empty_n;
  assign L1_out_id_8__full_n = L1_out_id_8_if_full_n;
  assign L1_out_id_8_if_read = L1_out_id_8__read;
  assign L1_out_id_8_if_read_ce = 1'b1;
  assign L1_out_id_8_if_write = L1_out_id_8__write;
  assign L1_out_id_8_if_write_ce = 1'b1;
  assign L1_out_id_8_reset = ~ ap_rst_n;
  assign L2_out_dist0_clk = ap_clk;
  assign L2_out_dist0_if_din = L2_out_dist0__din;
  assign L2_out_dist0__dout = L2_out_dist0_if_dout;
  assign L2_out_dist0__empty_n = L2_out_dist0_if_empty_n;
  assign L2_out_dist0__full_n = L2_out_dist0_if_full_n;
  assign L2_out_dist0_if_read = L2_out_dist0__read;
  assign L2_out_dist0_if_read_ce = 1'b1;
  assign L2_out_dist0_if_write = L2_out_dist0__write;
  assign L2_out_dist0_if_write_ce = 1'b1;
  assign L2_out_dist0_reset = ~ ap_rst_n;
  assign L2_out_dist1_clk = ap_clk;
  assign L2_out_dist1_if_din = L2_out_dist1__din;
  assign L2_out_dist1__dout = L2_out_dist1_if_dout;
  assign L2_out_dist1__empty_n = L2_out_dist1_if_empty_n;
  assign L2_out_dist1__full_n = L2_out_dist1_if_full_n;
  assign L2_out_dist1_if_read = L2_out_dist1__read;
  assign L2_out_dist1_if_read_ce = 1'b1;
  assign L2_out_dist1_if_write = L2_out_dist1__write;
  assign L2_out_dist1_if_write_ce = 1'b1;
  assign L2_out_dist1_reset = ~ ap_rst_n;
  assign L2_out_dist2_clk = ap_clk;
  assign L2_out_dist2_if_din = L2_out_dist2__din;
  assign L2_out_dist2__dout = L2_out_dist2_if_dout;
  assign L2_out_dist2__empty_n = L2_out_dist2_if_empty_n;
  assign L2_out_dist2__full_n = L2_out_dist2_if_full_n;
  assign L2_out_dist2_if_read = L2_out_dist2__read;
  assign L2_out_dist2_if_read_ce = 1'b1;
  assign L2_out_dist2_if_write = L2_out_dist2__write;
  assign L2_out_dist2_if_write_ce = 1'b1;
  assign L2_out_dist2_reset = ~ ap_rst_n;
  assign L2_out_id0_clk = ap_clk;
  assign L2_out_id0_if_din = L2_out_id0__din;
  assign L2_out_id0__dout = L2_out_id0_if_dout;
  assign L2_out_id0__empty_n = L2_out_id0_if_empty_n;
  assign L2_out_id0__full_n = L2_out_id0_if_full_n;
  assign L2_out_id0_if_read = L2_out_id0__read;
  assign L2_out_id0_if_read_ce = 1'b1;
  assign L2_out_id0_if_write = L2_out_id0__write;
  assign L2_out_id0_if_write_ce = 1'b1;
  assign L2_out_id0_reset = ~ ap_rst_n;
  assign L2_out_id1_clk = ap_clk;
  assign L2_out_id1_if_din = L2_out_id1__din;
  assign L2_out_id1__dout = L2_out_id1_if_dout;
  assign L2_out_id1__empty_n = L2_out_id1_if_empty_n;
  assign L2_out_id1__full_n = L2_out_id1_if_full_n;
  assign L2_out_id1_if_read = L2_out_id1__read;
  assign L2_out_id1_if_read_ce = 1'b1;
  assign L2_out_id1_if_write = L2_out_id1__write;
  assign L2_out_id1_if_write_ce = 1'b1;
  assign L2_out_id1_reset = ~ ap_rst_n;
  assign L2_out_id2_clk = ap_clk;
  assign L2_out_id2_if_din = L2_out_id2__din;
  assign L2_out_id2__dout = L2_out_id2_if_dout;
  assign L2_out_id2__empty_n = L2_out_id2_if_empty_n;
  assign L2_out_id2__full_n = L2_out_id2_if_full_n;
  assign L2_out_id2_if_read = L2_out_id2__read;
  assign L2_out_id2_if_read_ce = 1'b1;
  assign L2_out_id2_if_write = L2_out_id2__write;
  assign L2_out_id2_if_write_ce = 1'b1;
  assign L2_out_id2_reset = ~ ap_rst_n;
  assign L3_out_dist_stream_clk = ap_clk;
  assign L3_out_dist_stream_if_din = L3_out_dist_stream__din;
  assign L3_out_dist_stream__dout = L3_out_dist_stream_if_dout;
  assign L3_out_dist_stream__empty_n = L3_out_dist_stream_if_empty_n;
  assign L3_out_dist_stream__full_n = L3_out_dist_stream_if_full_n;
  assign L3_out_dist_stream_if_read = L3_out_dist_stream__read;
  assign L3_out_dist_stream_if_read_ce = 1'b1;
  assign L3_out_dist_stream_if_write = L3_out_dist_stream__write;
  assign L3_out_dist_stream_if_write_ce = 1'b1;
  assign L3_out_dist_stream_reset = ~ ap_rst_n;
  assign L3_out_id_stream_clk = ap_clk;
  assign L3_out_id_stream_if_din = L3_out_id_stream__din;
  assign L3_out_id_stream__dout = L3_out_id_stream_if_dout;
  assign L3_out_id_stream__empty_n = L3_out_id_stream_if_empty_n;
  assign L3_out_id_stream__full_n = L3_out_id_stream_if_full_n;
  assign L3_out_id_stream_if_read = L3_out_id_stream__read;
  assign L3_out_id_stream_if_read_ce = 1'b1;
  assign L3_out_id_stream_if_write = L3_out_id_stream__write;
  assign L3_out_id_stream_if_write_ce = 1'b1;
  assign L3_out_id_stream_reset = ~ ap_rst_n;
  assign out_dist_0_clk = ap_clk;
  assign out_dist_0_if_din = out_dist_0__din;
  assign out_dist_0__dout = out_dist_0_if_dout;
  assign out_dist_0__empty_n = out_dist_0_if_empty_n;
  assign out_dist_0__full_n = out_dist_0_if_full_n;
  assign out_dist_0_if_read = out_dist_0__read;
  assign out_dist_0_if_read_ce = 1'b1;
  assign out_dist_0_if_write = out_dist_0__write;
  assign out_dist_0_if_write_ce = 1'b1;
  assign out_dist_0_reset = ~ ap_rst_n;
  assign out_dist_10_clk = ap_clk;
  assign out_dist_10_if_din = out_dist_10__din;
  assign out_dist_10__dout = out_dist_10_if_dout;
  assign out_dist_10__empty_n = out_dist_10_if_empty_n;
  assign out_dist_10__full_n = out_dist_10_if_full_n;
  assign out_dist_10_if_read = out_dist_10__read;
  assign out_dist_10_if_read_ce = 1'b1;
  assign out_dist_10_if_write = out_dist_10__write;
  assign out_dist_10_if_write_ce = 1'b1;
  assign out_dist_10_reset = ~ ap_rst_n;
  assign out_dist_11_clk = ap_clk;
  assign out_dist_11_if_din = out_dist_11__din;
  assign out_dist_11__dout = out_dist_11_if_dout;
  assign out_dist_11__empty_n = out_dist_11_if_empty_n;
  assign out_dist_11__full_n = out_dist_11_if_full_n;
  assign out_dist_11_if_read = out_dist_11__read;
  assign out_dist_11_if_read_ce = 1'b1;
  assign out_dist_11_if_write = out_dist_11__write;
  assign out_dist_11_if_write_ce = 1'b1;
  assign out_dist_11_reset = ~ ap_rst_n;
  assign out_dist_12_clk = ap_clk;
  assign out_dist_12_if_din = out_dist_12__din;
  assign out_dist_12__dout = out_dist_12_if_dout;
  assign out_dist_12__empty_n = out_dist_12_if_empty_n;
  assign out_dist_12__full_n = out_dist_12_if_full_n;
  assign out_dist_12_if_read = out_dist_12__read;
  assign out_dist_12_if_read_ce = 1'b1;
  assign out_dist_12_if_write = out_dist_12__write;
  assign out_dist_12_if_write_ce = 1'b1;
  assign out_dist_12_reset = ~ ap_rst_n;
  assign out_dist_13_clk = ap_clk;
  assign out_dist_13_if_din = out_dist_13__din;
  assign out_dist_13__dout = out_dist_13_if_dout;
  assign out_dist_13__empty_n = out_dist_13_if_empty_n;
  assign out_dist_13__full_n = out_dist_13_if_full_n;
  assign out_dist_13_if_read = out_dist_13__read;
  assign out_dist_13_if_read_ce = 1'b1;
  assign out_dist_13_if_write = out_dist_13__write;
  assign out_dist_13_if_write_ce = 1'b1;
  assign out_dist_13_reset = ~ ap_rst_n;
  assign out_dist_14_clk = ap_clk;
  assign out_dist_14_if_din = out_dist_14__din;
  assign out_dist_14__dout = out_dist_14_if_dout;
  assign out_dist_14__empty_n = out_dist_14_if_empty_n;
  assign out_dist_14__full_n = out_dist_14_if_full_n;
  assign out_dist_14_if_read = out_dist_14__read;
  assign out_dist_14_if_read_ce = 1'b1;
  assign out_dist_14_if_write = out_dist_14__write;
  assign out_dist_14_if_write_ce = 1'b1;
  assign out_dist_14_reset = ~ ap_rst_n;
  assign out_dist_15_clk = ap_clk;
  assign out_dist_15_if_din = out_dist_15__din;
  assign out_dist_15__dout = out_dist_15_if_dout;
  assign out_dist_15__empty_n = out_dist_15_if_empty_n;
  assign out_dist_15__full_n = out_dist_15_if_full_n;
  assign out_dist_15_if_read = out_dist_15__read;
  assign out_dist_15_if_read_ce = 1'b1;
  assign out_dist_15_if_write = out_dist_15__write;
  assign out_dist_15_if_write_ce = 1'b1;
  assign out_dist_15_reset = ~ ap_rst_n;
  assign out_dist_16_clk = ap_clk;
  assign out_dist_16_if_din = out_dist_16__din;
  assign out_dist_16__dout = out_dist_16_if_dout;
  assign out_dist_16__empty_n = out_dist_16_if_empty_n;
  assign out_dist_16__full_n = out_dist_16_if_full_n;
  assign out_dist_16_if_read = out_dist_16__read;
  assign out_dist_16_if_read_ce = 1'b1;
  assign out_dist_16_if_write = out_dist_16__write;
  assign out_dist_16_if_write_ce = 1'b1;
  assign out_dist_16_reset = ~ ap_rst_n;
  assign out_dist_17_clk = ap_clk;
  assign out_dist_17_if_din = out_dist_17__din;
  assign out_dist_17__dout = out_dist_17_if_dout;
  assign out_dist_17__empty_n = out_dist_17_if_empty_n;
  assign out_dist_17__full_n = out_dist_17_if_full_n;
  assign out_dist_17_if_read = out_dist_17__read;
  assign out_dist_17_if_read_ce = 1'b1;
  assign out_dist_17_if_write = out_dist_17__write;
  assign out_dist_17_if_write_ce = 1'b1;
  assign out_dist_17_reset = ~ ap_rst_n;
  assign out_dist_18_clk = ap_clk;
  assign out_dist_18_if_din = out_dist_18__din;
  assign out_dist_18__dout = out_dist_18_if_dout;
  assign out_dist_18__empty_n = out_dist_18_if_empty_n;
  assign out_dist_18__full_n = out_dist_18_if_full_n;
  assign out_dist_18_if_read = out_dist_18__read;
  assign out_dist_18_if_read_ce = 1'b1;
  assign out_dist_18_if_write = out_dist_18__write;
  assign out_dist_18_if_write_ce = 1'b1;
  assign out_dist_18_reset = ~ ap_rst_n;
  assign out_dist_19_clk = ap_clk;
  assign out_dist_19_if_din = out_dist_19__din;
  assign out_dist_19__dout = out_dist_19_if_dout;
  assign out_dist_19__empty_n = out_dist_19_if_empty_n;
  assign out_dist_19__full_n = out_dist_19_if_full_n;
  assign out_dist_19_if_read = out_dist_19__read;
  assign out_dist_19_if_read_ce = 1'b1;
  assign out_dist_19_if_write = out_dist_19__write;
  assign out_dist_19_if_write_ce = 1'b1;
  assign out_dist_19_reset = ~ ap_rst_n;
  assign out_dist_1_clk = ap_clk;
  assign out_dist_1_if_din = out_dist_1__din;
  assign out_dist_1__dout = out_dist_1_if_dout;
  assign out_dist_1__empty_n = out_dist_1_if_empty_n;
  assign out_dist_1__full_n = out_dist_1_if_full_n;
  assign out_dist_1_if_read = out_dist_1__read;
  assign out_dist_1_if_read_ce = 1'b1;
  assign out_dist_1_if_write = out_dist_1__write;
  assign out_dist_1_if_write_ce = 1'b1;
  assign out_dist_1_reset = ~ ap_rst_n;
  assign out_dist_20_clk = ap_clk;
  assign out_dist_20_if_din = out_dist_20__din;
  assign out_dist_20__dout = out_dist_20_if_dout;
  assign out_dist_20__empty_n = out_dist_20_if_empty_n;
  assign out_dist_20__full_n = out_dist_20_if_full_n;
  assign out_dist_20_if_read = out_dist_20__read;
  assign out_dist_20_if_read_ce = 1'b1;
  assign out_dist_20_if_write = out_dist_20__write;
  assign out_dist_20_if_write_ce = 1'b1;
  assign out_dist_20_reset = ~ ap_rst_n;
  assign out_dist_21_clk = ap_clk;
  assign out_dist_21_if_din = out_dist_21__din;
  assign out_dist_21__dout = out_dist_21_if_dout;
  assign out_dist_21__empty_n = out_dist_21_if_empty_n;
  assign out_dist_21__full_n = out_dist_21_if_full_n;
  assign out_dist_21_if_read = out_dist_21__read;
  assign out_dist_21_if_read_ce = 1'b1;
  assign out_dist_21_if_write = out_dist_21__write;
  assign out_dist_21_if_write_ce = 1'b1;
  assign out_dist_21_reset = ~ ap_rst_n;
  assign out_dist_22_clk = ap_clk;
  assign out_dist_22_if_din = out_dist_22__din;
  assign out_dist_22__dout = out_dist_22_if_dout;
  assign out_dist_22__empty_n = out_dist_22_if_empty_n;
  assign out_dist_22__full_n = out_dist_22_if_full_n;
  assign out_dist_22_if_read = out_dist_22__read;
  assign out_dist_22_if_read_ce = 1'b1;
  assign out_dist_22_if_write = out_dist_22__write;
  assign out_dist_22_if_write_ce = 1'b1;
  assign out_dist_22_reset = ~ ap_rst_n;
  assign out_dist_23_clk = ap_clk;
  assign out_dist_23_if_din = out_dist_23__din;
  assign out_dist_23__dout = out_dist_23_if_dout;
  assign out_dist_23__empty_n = out_dist_23_if_empty_n;
  assign out_dist_23__full_n = out_dist_23_if_full_n;
  assign out_dist_23_if_read = out_dist_23__read;
  assign out_dist_23_if_read_ce = 1'b1;
  assign out_dist_23_if_write = out_dist_23__write;
  assign out_dist_23_if_write_ce = 1'b1;
  assign out_dist_23_reset = ~ ap_rst_n;
  assign out_dist_24_clk = ap_clk;
  assign out_dist_24_if_din = out_dist_24__din;
  assign out_dist_24__dout = out_dist_24_if_dout;
  assign out_dist_24__empty_n = out_dist_24_if_empty_n;
  assign out_dist_24__full_n = out_dist_24_if_full_n;
  assign out_dist_24_if_read = out_dist_24__read;
  assign out_dist_24_if_read_ce = 1'b1;
  assign out_dist_24_if_write = out_dist_24__write;
  assign out_dist_24_if_write_ce = 1'b1;
  assign out_dist_24_reset = ~ ap_rst_n;
  assign out_dist_25_clk = ap_clk;
  assign out_dist_25_if_din = out_dist_25__din;
  assign out_dist_25__dout = out_dist_25_if_dout;
  assign out_dist_25__empty_n = out_dist_25_if_empty_n;
  assign out_dist_25__full_n = out_dist_25_if_full_n;
  assign out_dist_25_if_read = out_dist_25__read;
  assign out_dist_25_if_read_ce = 1'b1;
  assign out_dist_25_if_write = out_dist_25__write;
  assign out_dist_25_if_write_ce = 1'b1;
  assign out_dist_25_reset = ~ ap_rst_n;
  assign out_dist_26_clk = ap_clk;
  assign out_dist_26_if_din = out_dist_26__din;
  assign out_dist_26__dout = out_dist_26_if_dout;
  assign out_dist_26__empty_n = out_dist_26_if_empty_n;
  assign out_dist_26__full_n = out_dist_26_if_full_n;
  assign out_dist_26_if_read = out_dist_26__read;
  assign out_dist_26_if_read_ce = 1'b1;
  assign out_dist_26_if_write = out_dist_26__write;
  assign out_dist_26_if_write_ce = 1'b1;
  assign out_dist_26_reset = ~ ap_rst_n;
  assign out_dist_2_clk = ap_clk;
  assign out_dist_2_if_din = out_dist_2__din;
  assign out_dist_2__dout = out_dist_2_if_dout;
  assign out_dist_2__empty_n = out_dist_2_if_empty_n;
  assign out_dist_2__full_n = out_dist_2_if_full_n;
  assign out_dist_2_if_read = out_dist_2__read;
  assign out_dist_2_if_read_ce = 1'b1;
  assign out_dist_2_if_write = out_dist_2__write;
  assign out_dist_2_if_write_ce = 1'b1;
  assign out_dist_2_reset = ~ ap_rst_n;
  assign out_dist_3_clk = ap_clk;
  assign out_dist_3_if_din = out_dist_3__din;
  assign out_dist_3__dout = out_dist_3_if_dout;
  assign out_dist_3__empty_n = out_dist_3_if_empty_n;
  assign out_dist_3__full_n = out_dist_3_if_full_n;
  assign out_dist_3_if_read = out_dist_3__read;
  assign out_dist_3_if_read_ce = 1'b1;
  assign out_dist_3_if_write = out_dist_3__write;
  assign out_dist_3_if_write_ce = 1'b1;
  assign out_dist_3_reset = ~ ap_rst_n;
  assign out_dist_4_clk = ap_clk;
  assign out_dist_4_if_din = out_dist_4__din;
  assign out_dist_4__dout = out_dist_4_if_dout;
  assign out_dist_4__empty_n = out_dist_4_if_empty_n;
  assign out_dist_4__full_n = out_dist_4_if_full_n;
  assign out_dist_4_if_read = out_dist_4__read;
  assign out_dist_4_if_read_ce = 1'b1;
  assign out_dist_4_if_write = out_dist_4__write;
  assign out_dist_4_if_write_ce = 1'b1;
  assign out_dist_4_reset = ~ ap_rst_n;
  assign out_dist_5_clk = ap_clk;
  assign out_dist_5_if_din = out_dist_5__din;
  assign out_dist_5__dout = out_dist_5_if_dout;
  assign out_dist_5__empty_n = out_dist_5_if_empty_n;
  assign out_dist_5__full_n = out_dist_5_if_full_n;
  assign out_dist_5_if_read = out_dist_5__read;
  assign out_dist_5_if_read_ce = 1'b1;
  assign out_dist_5_if_write = out_dist_5__write;
  assign out_dist_5_if_write_ce = 1'b1;
  assign out_dist_5_reset = ~ ap_rst_n;
  assign out_dist_6_clk = ap_clk;
  assign out_dist_6_if_din = out_dist_6__din;
  assign out_dist_6__dout = out_dist_6_if_dout;
  assign out_dist_6__empty_n = out_dist_6_if_empty_n;
  assign out_dist_6__full_n = out_dist_6_if_full_n;
  assign out_dist_6_if_read = out_dist_6__read;
  assign out_dist_6_if_read_ce = 1'b1;
  assign out_dist_6_if_write = out_dist_6__write;
  assign out_dist_6_if_write_ce = 1'b1;
  assign out_dist_6_reset = ~ ap_rst_n;
  assign out_dist_7_clk = ap_clk;
  assign out_dist_7_if_din = out_dist_7__din;
  assign out_dist_7__dout = out_dist_7_if_dout;
  assign out_dist_7__empty_n = out_dist_7_if_empty_n;
  assign out_dist_7__full_n = out_dist_7_if_full_n;
  assign out_dist_7_if_read = out_dist_7__read;
  assign out_dist_7_if_read_ce = 1'b1;
  assign out_dist_7_if_write = out_dist_7__write;
  assign out_dist_7_if_write_ce = 1'b1;
  assign out_dist_7_reset = ~ ap_rst_n;
  assign out_dist_8_clk = ap_clk;
  assign out_dist_8_if_din = out_dist_8__din;
  assign out_dist_8__dout = out_dist_8_if_dout;
  assign out_dist_8__empty_n = out_dist_8_if_empty_n;
  assign out_dist_8__full_n = out_dist_8_if_full_n;
  assign out_dist_8_if_read = out_dist_8__read;
  assign out_dist_8_if_read_ce = 1'b1;
  assign out_dist_8_if_write = out_dist_8__write;
  assign out_dist_8_if_write_ce = 1'b1;
  assign out_dist_8_reset = ~ ap_rst_n;
  assign out_dist_9_clk = ap_clk;
  assign out_dist_9_if_din = out_dist_9__din;
  assign out_dist_9__dout = out_dist_9_if_dout;
  assign out_dist_9__empty_n = out_dist_9_if_empty_n;
  assign out_dist_9__full_n = out_dist_9_if_full_n;
  assign out_dist_9_if_read = out_dist_9__read;
  assign out_dist_9_if_read_ce = 1'b1;
  assign out_dist_9_if_write = out_dist_9__write;
  assign out_dist_9_if_write_ce = 1'b1;
  assign out_dist_9_reset = ~ ap_rst_n;
  assign out_id_0_clk = ap_clk;
  assign out_id_0_if_din = out_id_0__din;
  assign out_id_0__dout = out_id_0_if_dout;
  assign out_id_0__empty_n = out_id_0_if_empty_n;
  assign out_id_0__full_n = out_id_0_if_full_n;
  assign out_id_0_if_read = out_id_0__read;
  assign out_id_0_if_read_ce = 1'b1;
  assign out_id_0_if_write = out_id_0__write;
  assign out_id_0_if_write_ce = 1'b1;
  assign out_id_0_reset = ~ ap_rst_n;
  assign out_id_10_clk = ap_clk;
  assign out_id_10_if_din = out_id_10__din;
  assign out_id_10__dout = out_id_10_if_dout;
  assign out_id_10__empty_n = out_id_10_if_empty_n;
  assign out_id_10__full_n = out_id_10_if_full_n;
  assign out_id_10_if_read = out_id_10__read;
  assign out_id_10_if_read_ce = 1'b1;
  assign out_id_10_if_write = out_id_10__write;
  assign out_id_10_if_write_ce = 1'b1;
  assign out_id_10_reset = ~ ap_rst_n;
  assign out_id_11_clk = ap_clk;
  assign out_id_11_if_din = out_id_11__din;
  assign out_id_11__dout = out_id_11_if_dout;
  assign out_id_11__empty_n = out_id_11_if_empty_n;
  assign out_id_11__full_n = out_id_11_if_full_n;
  assign out_id_11_if_read = out_id_11__read;
  assign out_id_11_if_read_ce = 1'b1;
  assign out_id_11_if_write = out_id_11__write;
  assign out_id_11_if_write_ce = 1'b1;
  assign out_id_11_reset = ~ ap_rst_n;
  assign out_id_12_clk = ap_clk;
  assign out_id_12_if_din = out_id_12__din;
  assign out_id_12__dout = out_id_12_if_dout;
  assign out_id_12__empty_n = out_id_12_if_empty_n;
  assign out_id_12__full_n = out_id_12_if_full_n;
  assign out_id_12_if_read = out_id_12__read;
  assign out_id_12_if_read_ce = 1'b1;
  assign out_id_12_if_write = out_id_12__write;
  assign out_id_12_if_write_ce = 1'b1;
  assign out_id_12_reset = ~ ap_rst_n;
  assign out_id_13_clk = ap_clk;
  assign out_id_13_if_din = out_id_13__din;
  assign out_id_13__dout = out_id_13_if_dout;
  assign out_id_13__empty_n = out_id_13_if_empty_n;
  assign out_id_13__full_n = out_id_13_if_full_n;
  assign out_id_13_if_read = out_id_13__read;
  assign out_id_13_if_read_ce = 1'b1;
  assign out_id_13_if_write = out_id_13__write;
  assign out_id_13_if_write_ce = 1'b1;
  assign out_id_13_reset = ~ ap_rst_n;
  assign out_id_14_clk = ap_clk;
  assign out_id_14_if_din = out_id_14__din;
  assign out_id_14__dout = out_id_14_if_dout;
  assign out_id_14__empty_n = out_id_14_if_empty_n;
  assign out_id_14__full_n = out_id_14_if_full_n;
  assign out_id_14_if_read = out_id_14__read;
  assign out_id_14_if_read_ce = 1'b1;
  assign out_id_14_if_write = out_id_14__write;
  assign out_id_14_if_write_ce = 1'b1;
  assign out_id_14_reset = ~ ap_rst_n;
  assign out_id_15_clk = ap_clk;
  assign out_id_15_if_din = out_id_15__din;
  assign out_id_15__dout = out_id_15_if_dout;
  assign out_id_15__empty_n = out_id_15_if_empty_n;
  assign out_id_15__full_n = out_id_15_if_full_n;
  assign out_id_15_if_read = out_id_15__read;
  assign out_id_15_if_read_ce = 1'b1;
  assign out_id_15_if_write = out_id_15__write;
  assign out_id_15_if_write_ce = 1'b1;
  assign out_id_15_reset = ~ ap_rst_n;
  assign out_id_16_clk = ap_clk;
  assign out_id_16_if_din = out_id_16__din;
  assign out_id_16__dout = out_id_16_if_dout;
  assign out_id_16__empty_n = out_id_16_if_empty_n;
  assign out_id_16__full_n = out_id_16_if_full_n;
  assign out_id_16_if_read = out_id_16__read;
  assign out_id_16_if_read_ce = 1'b1;
  assign out_id_16_if_write = out_id_16__write;
  assign out_id_16_if_write_ce = 1'b1;
  assign out_id_16_reset = ~ ap_rst_n;
  assign out_id_17_clk = ap_clk;
  assign out_id_17_if_din = out_id_17__din;
  assign out_id_17__dout = out_id_17_if_dout;
  assign out_id_17__empty_n = out_id_17_if_empty_n;
  assign out_id_17__full_n = out_id_17_if_full_n;
  assign out_id_17_if_read = out_id_17__read;
  assign out_id_17_if_read_ce = 1'b1;
  assign out_id_17_if_write = out_id_17__write;
  assign out_id_17_if_write_ce = 1'b1;
  assign out_id_17_reset = ~ ap_rst_n;
  assign out_id_18_clk = ap_clk;
  assign out_id_18_if_din = out_id_18__din;
  assign out_id_18__dout = out_id_18_if_dout;
  assign out_id_18__empty_n = out_id_18_if_empty_n;
  assign out_id_18__full_n = out_id_18_if_full_n;
  assign out_id_18_if_read = out_id_18__read;
  assign out_id_18_if_read_ce = 1'b1;
  assign out_id_18_if_write = out_id_18__write;
  assign out_id_18_if_write_ce = 1'b1;
  assign out_id_18_reset = ~ ap_rst_n;
  assign out_id_19_clk = ap_clk;
  assign out_id_19_if_din = out_id_19__din;
  assign out_id_19__dout = out_id_19_if_dout;
  assign out_id_19__empty_n = out_id_19_if_empty_n;
  assign out_id_19__full_n = out_id_19_if_full_n;
  assign out_id_19_if_read = out_id_19__read;
  assign out_id_19_if_read_ce = 1'b1;
  assign out_id_19_if_write = out_id_19__write;
  assign out_id_19_if_write_ce = 1'b1;
  assign out_id_19_reset = ~ ap_rst_n;
  assign out_id_1_clk = ap_clk;
  assign out_id_1_if_din = out_id_1__din;
  assign out_id_1__dout = out_id_1_if_dout;
  assign out_id_1__empty_n = out_id_1_if_empty_n;
  assign out_id_1__full_n = out_id_1_if_full_n;
  assign out_id_1_if_read = out_id_1__read;
  assign out_id_1_if_read_ce = 1'b1;
  assign out_id_1_if_write = out_id_1__write;
  assign out_id_1_if_write_ce = 1'b1;
  assign out_id_1_reset = ~ ap_rst_n;
  assign out_id_20_clk = ap_clk;
  assign out_id_20_if_din = out_id_20__din;
  assign out_id_20__dout = out_id_20_if_dout;
  assign out_id_20__empty_n = out_id_20_if_empty_n;
  assign out_id_20__full_n = out_id_20_if_full_n;
  assign out_id_20_if_read = out_id_20__read;
  assign out_id_20_if_read_ce = 1'b1;
  assign out_id_20_if_write = out_id_20__write;
  assign out_id_20_if_write_ce = 1'b1;
  assign out_id_20_reset = ~ ap_rst_n;
  assign out_id_21_clk = ap_clk;
  assign out_id_21_if_din = out_id_21__din;
  assign out_id_21__dout = out_id_21_if_dout;
  assign out_id_21__empty_n = out_id_21_if_empty_n;
  assign out_id_21__full_n = out_id_21_if_full_n;
  assign out_id_21_if_read = out_id_21__read;
  assign out_id_21_if_read_ce = 1'b1;
  assign out_id_21_if_write = out_id_21__write;
  assign out_id_21_if_write_ce = 1'b1;
  assign out_id_21_reset = ~ ap_rst_n;
  assign out_id_22_clk = ap_clk;
  assign out_id_22_if_din = out_id_22__din;
  assign out_id_22__dout = out_id_22_if_dout;
  assign out_id_22__empty_n = out_id_22_if_empty_n;
  assign out_id_22__full_n = out_id_22_if_full_n;
  assign out_id_22_if_read = out_id_22__read;
  assign out_id_22_if_read_ce = 1'b1;
  assign out_id_22_if_write = out_id_22__write;
  assign out_id_22_if_write_ce = 1'b1;
  assign out_id_22_reset = ~ ap_rst_n;
  assign out_id_23_clk = ap_clk;
  assign out_id_23_if_din = out_id_23__din;
  assign out_id_23__dout = out_id_23_if_dout;
  assign out_id_23__empty_n = out_id_23_if_empty_n;
  assign out_id_23__full_n = out_id_23_if_full_n;
  assign out_id_23_if_read = out_id_23__read;
  assign out_id_23_if_read_ce = 1'b1;
  assign out_id_23_if_write = out_id_23__write;
  assign out_id_23_if_write_ce = 1'b1;
  assign out_id_23_reset = ~ ap_rst_n;
  assign out_id_24_clk = ap_clk;
  assign out_id_24_if_din = out_id_24__din;
  assign out_id_24__dout = out_id_24_if_dout;
  assign out_id_24__empty_n = out_id_24_if_empty_n;
  assign out_id_24__full_n = out_id_24_if_full_n;
  assign out_id_24_if_read = out_id_24__read;
  assign out_id_24_if_read_ce = 1'b1;
  assign out_id_24_if_write = out_id_24__write;
  assign out_id_24_if_write_ce = 1'b1;
  assign out_id_24_reset = ~ ap_rst_n;
  assign out_id_25_clk = ap_clk;
  assign out_id_25_if_din = out_id_25__din;
  assign out_id_25__dout = out_id_25_if_dout;
  assign out_id_25__empty_n = out_id_25_if_empty_n;
  assign out_id_25__full_n = out_id_25_if_full_n;
  assign out_id_25_if_read = out_id_25__read;
  assign out_id_25_if_read_ce = 1'b1;
  assign out_id_25_if_write = out_id_25__write;
  assign out_id_25_if_write_ce = 1'b1;
  assign out_id_25_reset = ~ ap_rst_n;
  assign out_id_26_clk = ap_clk;
  assign out_id_26_if_din = out_id_26__din;
  assign out_id_26__dout = out_id_26_if_dout;
  assign out_id_26__empty_n = out_id_26_if_empty_n;
  assign out_id_26__full_n = out_id_26_if_full_n;
  assign out_id_26_if_read = out_id_26__read;
  assign out_id_26_if_read_ce = 1'b1;
  assign out_id_26_if_write = out_id_26__write;
  assign out_id_26_if_write_ce = 1'b1;
  assign out_id_26_reset = ~ ap_rst_n;
  assign out_id_2_clk = ap_clk;
  assign out_id_2_if_din = out_id_2__din;
  assign out_id_2__dout = out_id_2_if_dout;
  assign out_id_2__empty_n = out_id_2_if_empty_n;
  assign out_id_2__full_n = out_id_2_if_full_n;
  assign out_id_2_if_read = out_id_2__read;
  assign out_id_2_if_read_ce = 1'b1;
  assign out_id_2_if_write = out_id_2__write;
  assign out_id_2_if_write_ce = 1'b1;
  assign out_id_2_reset = ~ ap_rst_n;
  assign out_id_3_clk = ap_clk;
  assign out_id_3_if_din = out_id_3__din;
  assign out_id_3__dout = out_id_3_if_dout;
  assign out_id_3__empty_n = out_id_3_if_empty_n;
  assign out_id_3__full_n = out_id_3_if_full_n;
  assign out_id_3_if_read = out_id_3__read;
  assign out_id_3_if_read_ce = 1'b1;
  assign out_id_3_if_write = out_id_3__write;
  assign out_id_3_if_write_ce = 1'b1;
  assign out_id_3_reset = ~ ap_rst_n;
  assign out_id_4_clk = ap_clk;
  assign out_id_4_if_din = out_id_4__din;
  assign out_id_4__dout = out_id_4_if_dout;
  assign out_id_4__empty_n = out_id_4_if_empty_n;
  assign out_id_4__full_n = out_id_4_if_full_n;
  assign out_id_4_if_read = out_id_4__read;
  assign out_id_4_if_read_ce = 1'b1;
  assign out_id_4_if_write = out_id_4__write;
  assign out_id_4_if_write_ce = 1'b1;
  assign out_id_4_reset = ~ ap_rst_n;
  assign out_id_5_clk = ap_clk;
  assign out_id_5_if_din = out_id_5__din;
  assign out_id_5__dout = out_id_5_if_dout;
  assign out_id_5__empty_n = out_id_5_if_empty_n;
  assign out_id_5__full_n = out_id_5_if_full_n;
  assign out_id_5_if_read = out_id_5__read;
  assign out_id_5_if_read_ce = 1'b1;
  assign out_id_5_if_write = out_id_5__write;
  assign out_id_5_if_write_ce = 1'b1;
  assign out_id_5_reset = ~ ap_rst_n;
  assign out_id_6_clk = ap_clk;
  assign out_id_6_if_din = out_id_6__din;
  assign out_id_6__dout = out_id_6_if_dout;
  assign out_id_6__empty_n = out_id_6_if_empty_n;
  assign out_id_6__full_n = out_id_6_if_full_n;
  assign out_id_6_if_read = out_id_6__read;
  assign out_id_6_if_read_ce = 1'b1;
  assign out_id_6_if_write = out_id_6__write;
  assign out_id_6_if_write_ce = 1'b1;
  assign out_id_6_reset = ~ ap_rst_n;
  assign out_id_7_clk = ap_clk;
  assign out_id_7_if_din = out_id_7__din;
  assign out_id_7__dout = out_id_7_if_dout;
  assign out_id_7__empty_n = out_id_7_if_empty_n;
  assign out_id_7__full_n = out_id_7_if_full_n;
  assign out_id_7_if_read = out_id_7__read;
  assign out_id_7_if_read_ce = 1'b1;
  assign out_id_7_if_write = out_id_7__write;
  assign out_id_7_if_write_ce = 1'b1;
  assign out_id_7_reset = ~ ap_rst_n;
  assign out_id_8_clk = ap_clk;
  assign out_id_8_if_din = out_id_8__din;
  assign out_id_8__dout = out_id_8_if_dout;
  assign out_id_8__empty_n = out_id_8_if_empty_n;
  assign out_id_8__full_n = out_id_8_if_full_n;
  assign out_id_8_if_read = out_id_8__read;
  assign out_id_8_if_read_ce = 1'b1;
  assign out_id_8_if_write = out_id_8__write;
  assign out_id_8_if_write_ce = 1'b1;
  assign out_id_8_reset = ~ ap_rst_n;
  assign out_id_9_clk = ap_clk;
  assign out_id_9_if_din = out_id_9__din;
  assign out_id_9__dout = out_id_9_if_dout;
  assign out_id_9__empty_n = out_id_9_if_empty_n;
  assign out_id_9__full_n = out_id_9_if_full_n;
  assign out_id_9_if_read = out_id_9__read;
  assign out_id_9_if_read_ce = 1'b1;
  assign out_id_9_if_write = out_id_9__write;
  assign out_id_9_if_write_ce = 1'b1;
  assign out_id_9_reset = ~ ap_rst_n;
  assign krnl_globalSort_L1_L2_0_ap_clk = ap_clk;
  assign krnl_globalSort_L1_L2_0__ap_done = krnl_globalSort_L1_L2_0_ap_done;
  assign krnl_globalSort_L1_L2_0__ap_idle = krnl_globalSort_L1_L2_0_ap_idle;
  assign krnl_globalSort_L1_L2_0__ap_ready = krnl_globalSort_L1_L2_0_ap_ready;
  assign krnl_globalSort_L1_L2_0_ap_rst_n = ap_rst_n;
  assign krnl_globalSort_L1_L2_0_ap_start = krnl_globalSort_L1_L2_0__ap_start;
  assign krnl_globalSort_L1_L2_0_in_dist0_peek_dout = out_dist_0__dout;
  assign krnl_globalSort_L1_L2_0_in_dist0_peek_empty_n = out_dist_0__empty_n;
  assign krnl_globalSort_L1_L2_0_in_dist0_s_dout = out_dist_0__dout;
  assign krnl_globalSort_L1_L2_0_in_dist0_s_empty_n = out_dist_0__empty_n;
  assign out_dist_0__read = krnl_globalSort_L1_L2_0_in_dist0_s_read;
  assign krnl_globalSort_L1_L2_0_in_dist1_peek_dout = out_dist_1__dout;
  assign krnl_globalSort_L1_L2_0_in_dist1_peek_empty_n = out_dist_1__empty_n;
  assign krnl_globalSort_L1_L2_0_in_dist1_s_dout = out_dist_1__dout;
  assign krnl_globalSort_L1_L2_0_in_dist1_s_empty_n = out_dist_1__empty_n;
  assign out_dist_1__read = krnl_globalSort_L1_L2_0_in_dist1_s_read;
  assign krnl_globalSort_L1_L2_0_in_dist2_peek_dout = out_dist_2__dout;
  assign krnl_globalSort_L1_L2_0_in_dist2_peek_empty_n = out_dist_2__empty_n;
  assign krnl_globalSort_L1_L2_0_in_dist2_s_dout = out_dist_2__dout;
  assign krnl_globalSort_L1_L2_0_in_dist2_s_empty_n = out_dist_2__empty_n;
  assign out_dist_2__read = krnl_globalSort_L1_L2_0_in_dist2_s_read;
  assign krnl_globalSort_L1_L2_0_in_id0_peek_dout = out_id_0__dout;
  assign krnl_globalSort_L1_L2_0_in_id0_peek_empty_n = out_id_0__empty_n;
  assign krnl_globalSort_L1_L2_0_in_id0_s_dout = out_id_0__dout;
  assign krnl_globalSort_L1_L2_0_in_id0_s_empty_n = out_id_0__empty_n;
  assign out_id_0__read = krnl_globalSort_L1_L2_0_in_id0_s_read;
  assign krnl_globalSort_L1_L2_0_in_id1_peek_dout = out_id_1__dout;
  assign krnl_globalSort_L1_L2_0_in_id1_peek_empty_n = out_id_1__empty_n;
  assign krnl_globalSort_L1_L2_0_in_id1_s_dout = out_id_1__dout;
  assign krnl_globalSort_L1_L2_0_in_id1_s_empty_n = out_id_1__empty_n;
  assign out_id_1__read = krnl_globalSort_L1_L2_0_in_id1_s_read;
  assign krnl_globalSort_L1_L2_0_in_id2_peek_dout = out_id_2__dout;
  assign krnl_globalSort_L1_L2_0_in_id2_peek_empty_n = out_id_2__empty_n;
  assign krnl_globalSort_L1_L2_0_in_id2_s_dout = out_id_2__dout;
  assign krnl_globalSort_L1_L2_0_in_id2_s_empty_n = out_id_2__empty_n;
  assign out_id_2__read = krnl_globalSort_L1_L2_0_in_id2_s_read;
  assign L1_out_dist_0__din = krnl_globalSort_L1_L2_0_out_dist_din;
  assign krnl_globalSort_L1_L2_0_out_dist_full_n = L1_out_dist_0__full_n;
  assign L1_out_dist_0__write = krnl_globalSort_L1_L2_0_out_dist_write;
  assign L1_out_id_0__din = krnl_globalSort_L1_L2_0_out_id_din;
  assign krnl_globalSort_L1_L2_0_out_id_full_n = L1_out_id_0__full_n;
  assign L1_out_id_0__write = krnl_globalSort_L1_L2_0_out_id_write;
  assign krnl_globalSort_L1_L2_1_ap_clk = ap_clk;
  assign krnl_globalSort_L1_L2_1__ap_done = krnl_globalSort_L1_L2_1_ap_done;
  assign krnl_globalSort_L1_L2_1__ap_idle = krnl_globalSort_L1_L2_1_ap_idle;
  assign krnl_globalSort_L1_L2_1__ap_ready = krnl_globalSort_L1_L2_1_ap_ready;
  assign krnl_globalSort_L1_L2_1_ap_rst_n = ap_rst_n;
  assign krnl_globalSort_L1_L2_1_ap_start = krnl_globalSort_L1_L2_1__ap_start;
  assign krnl_globalSort_L1_L2_1_in_dist0_peek_dout = out_dist_3__dout;
  assign krnl_globalSort_L1_L2_1_in_dist0_peek_empty_n = out_dist_3__empty_n;
  assign krnl_globalSort_L1_L2_1_in_dist0_s_dout = out_dist_3__dout;
  assign krnl_globalSort_L1_L2_1_in_dist0_s_empty_n = out_dist_3__empty_n;
  assign out_dist_3__read = krnl_globalSort_L1_L2_1_in_dist0_s_read;
  assign krnl_globalSort_L1_L2_1_in_dist1_peek_dout = out_dist_4__dout;
  assign krnl_globalSort_L1_L2_1_in_dist1_peek_empty_n = out_dist_4__empty_n;
  assign krnl_globalSort_L1_L2_1_in_dist1_s_dout = out_dist_4__dout;
  assign krnl_globalSort_L1_L2_1_in_dist1_s_empty_n = out_dist_4__empty_n;
  assign out_dist_4__read = krnl_globalSort_L1_L2_1_in_dist1_s_read;
  assign krnl_globalSort_L1_L2_1_in_dist2_peek_dout = out_dist_5__dout;
  assign krnl_globalSort_L1_L2_1_in_dist2_peek_empty_n = out_dist_5__empty_n;
  assign krnl_globalSort_L1_L2_1_in_dist2_s_dout = out_dist_5__dout;
  assign krnl_globalSort_L1_L2_1_in_dist2_s_empty_n = out_dist_5__empty_n;
  assign out_dist_5__read = krnl_globalSort_L1_L2_1_in_dist2_s_read;
  assign krnl_globalSort_L1_L2_1_in_id0_peek_dout = out_id_3__dout;
  assign krnl_globalSort_L1_L2_1_in_id0_peek_empty_n = out_id_3__empty_n;
  assign krnl_globalSort_L1_L2_1_in_id0_s_dout = out_id_3__dout;
  assign krnl_globalSort_L1_L2_1_in_id0_s_empty_n = out_id_3__empty_n;
  assign out_id_3__read = krnl_globalSort_L1_L2_1_in_id0_s_read;
  assign krnl_globalSort_L1_L2_1_in_id1_peek_dout = out_id_4__dout;
  assign krnl_globalSort_L1_L2_1_in_id1_peek_empty_n = out_id_4__empty_n;
  assign krnl_globalSort_L1_L2_1_in_id1_s_dout = out_id_4__dout;
  assign krnl_globalSort_L1_L2_1_in_id1_s_empty_n = out_id_4__empty_n;
  assign out_id_4__read = krnl_globalSort_L1_L2_1_in_id1_s_read;
  assign krnl_globalSort_L1_L2_1_in_id2_peek_dout = out_id_5__dout;
  assign krnl_globalSort_L1_L2_1_in_id2_peek_empty_n = out_id_5__empty_n;
  assign krnl_globalSort_L1_L2_1_in_id2_s_dout = out_id_5__dout;
  assign krnl_globalSort_L1_L2_1_in_id2_s_empty_n = out_id_5__empty_n;
  assign out_id_5__read = krnl_globalSort_L1_L2_1_in_id2_s_read;
  assign L1_out_dist_1__din = krnl_globalSort_L1_L2_1_out_dist_din;
  assign krnl_globalSort_L1_L2_1_out_dist_full_n = L1_out_dist_1__full_n;
  assign L1_out_dist_1__write = krnl_globalSort_L1_L2_1_out_dist_write;
  assign L1_out_id_1__din = krnl_globalSort_L1_L2_1_out_id_din;
  assign krnl_globalSort_L1_L2_1_out_id_full_n = L1_out_id_1__full_n;
  assign L1_out_id_1__write = krnl_globalSort_L1_L2_1_out_id_write;
  assign krnl_globalSort_L1_L2_2_ap_clk = ap_clk;
  assign krnl_globalSort_L1_L2_2__ap_done = krnl_globalSort_L1_L2_2_ap_done;
  assign krnl_globalSort_L1_L2_2__ap_idle = krnl_globalSort_L1_L2_2_ap_idle;
  assign krnl_globalSort_L1_L2_2__ap_ready = krnl_globalSort_L1_L2_2_ap_ready;
  assign krnl_globalSort_L1_L2_2_ap_rst_n = ap_rst_n;
  assign krnl_globalSort_L1_L2_2_ap_start = krnl_globalSort_L1_L2_2__ap_start;
  assign krnl_globalSort_L1_L2_2_in_dist0_peek_dout = out_dist_6__dout;
  assign krnl_globalSort_L1_L2_2_in_dist0_peek_empty_n = out_dist_6__empty_n;
  assign krnl_globalSort_L1_L2_2_in_dist0_s_dout = out_dist_6__dout;
  assign krnl_globalSort_L1_L2_2_in_dist0_s_empty_n = out_dist_6__empty_n;
  assign out_dist_6__read = krnl_globalSort_L1_L2_2_in_dist0_s_read;
  assign krnl_globalSort_L1_L2_2_in_dist1_peek_dout = out_dist_7__dout;
  assign krnl_globalSort_L1_L2_2_in_dist1_peek_empty_n = out_dist_7__empty_n;
  assign krnl_globalSort_L1_L2_2_in_dist1_s_dout = out_dist_7__dout;
  assign krnl_globalSort_L1_L2_2_in_dist1_s_empty_n = out_dist_7__empty_n;
  assign out_dist_7__read = krnl_globalSort_L1_L2_2_in_dist1_s_read;
  assign krnl_globalSort_L1_L2_2_in_dist2_peek_dout = out_dist_8__dout;
  assign krnl_globalSort_L1_L2_2_in_dist2_peek_empty_n = out_dist_8__empty_n;
  assign krnl_globalSort_L1_L2_2_in_dist2_s_dout = out_dist_8__dout;
  assign krnl_globalSort_L1_L2_2_in_dist2_s_empty_n = out_dist_8__empty_n;
  assign out_dist_8__read = krnl_globalSort_L1_L2_2_in_dist2_s_read;
  assign krnl_globalSort_L1_L2_2_in_id0_peek_dout = out_id_6__dout;
  assign krnl_globalSort_L1_L2_2_in_id0_peek_empty_n = out_id_6__empty_n;
  assign krnl_globalSort_L1_L2_2_in_id0_s_dout = out_id_6__dout;
  assign krnl_globalSort_L1_L2_2_in_id0_s_empty_n = out_id_6__empty_n;
  assign out_id_6__read = krnl_globalSort_L1_L2_2_in_id0_s_read;
  assign krnl_globalSort_L1_L2_2_in_id1_peek_dout = out_id_7__dout;
  assign krnl_globalSort_L1_L2_2_in_id1_peek_empty_n = out_id_7__empty_n;
  assign krnl_globalSort_L1_L2_2_in_id1_s_dout = out_id_7__dout;
  assign krnl_globalSort_L1_L2_2_in_id1_s_empty_n = out_id_7__empty_n;
  assign out_id_7__read = krnl_globalSort_L1_L2_2_in_id1_s_read;
  assign krnl_globalSort_L1_L2_2_in_id2_peek_dout = out_id_8__dout;
  assign krnl_globalSort_L1_L2_2_in_id2_peek_empty_n = out_id_8__empty_n;
  assign krnl_globalSort_L1_L2_2_in_id2_s_dout = out_id_8__dout;
  assign krnl_globalSort_L1_L2_2_in_id2_s_empty_n = out_id_8__empty_n;
  assign out_id_8__read = krnl_globalSort_L1_L2_2_in_id2_s_read;
  assign L1_out_dist_2__din = krnl_globalSort_L1_L2_2_out_dist_din;
  assign krnl_globalSort_L1_L2_2_out_dist_full_n = L1_out_dist_2__full_n;
  assign L1_out_dist_2__write = krnl_globalSort_L1_L2_2_out_dist_write;
  assign L1_out_id_2__din = krnl_globalSort_L1_L2_2_out_id_din;
  assign krnl_globalSort_L1_L2_2_out_id_full_n = L1_out_id_2__full_n;
  assign L1_out_id_2__write = krnl_globalSort_L1_L2_2_out_id_write;
  assign krnl_globalSort_L1_L2_3_ap_clk = ap_clk;
  assign krnl_globalSort_L1_L2_3__ap_done = krnl_globalSort_L1_L2_3_ap_done;
  assign krnl_globalSort_L1_L2_3__ap_idle = krnl_globalSort_L1_L2_3_ap_idle;
  assign krnl_globalSort_L1_L2_3__ap_ready = krnl_globalSort_L1_L2_3_ap_ready;
  assign krnl_globalSort_L1_L2_3_ap_rst_n = ap_rst_n;
  assign krnl_globalSort_L1_L2_3_ap_start = krnl_globalSort_L1_L2_3__ap_start;
  assign krnl_globalSort_L1_L2_3_in_dist0_peek_dout = out_dist_9__dout;
  assign krnl_globalSort_L1_L2_3_in_dist0_peek_empty_n = out_dist_9__empty_n;
  assign krnl_globalSort_L1_L2_3_in_dist0_s_dout = out_dist_9__dout;
  assign krnl_globalSort_L1_L2_3_in_dist0_s_empty_n = out_dist_9__empty_n;
  assign out_dist_9__read = krnl_globalSort_L1_L2_3_in_dist0_s_read;
  assign krnl_globalSort_L1_L2_3_in_dist1_peek_dout = out_dist_10__dout;
  assign krnl_globalSort_L1_L2_3_in_dist1_peek_empty_n = out_dist_10__empty_n;
  assign krnl_globalSort_L1_L2_3_in_dist1_s_dout = out_dist_10__dout;
  assign krnl_globalSort_L1_L2_3_in_dist1_s_empty_n = out_dist_10__empty_n;
  assign out_dist_10__read = krnl_globalSort_L1_L2_3_in_dist1_s_read;
  assign krnl_globalSort_L1_L2_3_in_dist2_peek_dout = out_dist_11__dout;
  assign krnl_globalSort_L1_L2_3_in_dist2_peek_empty_n = out_dist_11__empty_n;
  assign krnl_globalSort_L1_L2_3_in_dist2_s_dout = out_dist_11__dout;
  assign krnl_globalSort_L1_L2_3_in_dist2_s_empty_n = out_dist_11__empty_n;
  assign out_dist_11__read = krnl_globalSort_L1_L2_3_in_dist2_s_read;
  assign krnl_globalSort_L1_L2_3_in_id0_peek_dout = out_id_9__dout;
  assign krnl_globalSort_L1_L2_3_in_id0_peek_empty_n = out_id_9__empty_n;
  assign krnl_globalSort_L1_L2_3_in_id0_s_dout = out_id_9__dout;
  assign krnl_globalSort_L1_L2_3_in_id0_s_empty_n = out_id_9__empty_n;
  assign out_id_9__read = krnl_globalSort_L1_L2_3_in_id0_s_read;
  assign krnl_globalSort_L1_L2_3_in_id1_peek_dout = out_id_10__dout;
  assign krnl_globalSort_L1_L2_3_in_id1_peek_empty_n = out_id_10__empty_n;
  assign krnl_globalSort_L1_L2_3_in_id1_s_dout = out_id_10__dout;
  assign krnl_globalSort_L1_L2_3_in_id1_s_empty_n = out_id_10__empty_n;
  assign out_id_10__read = krnl_globalSort_L1_L2_3_in_id1_s_read;
  assign krnl_globalSort_L1_L2_3_in_id2_peek_dout = out_id_11__dout;
  assign krnl_globalSort_L1_L2_3_in_id2_peek_empty_n = out_id_11__empty_n;
  assign krnl_globalSort_L1_L2_3_in_id2_s_dout = out_id_11__dout;
  assign krnl_globalSort_L1_L2_3_in_id2_s_empty_n = out_id_11__empty_n;
  assign out_id_11__read = krnl_globalSort_L1_L2_3_in_id2_s_read;
  assign L1_out_dist_3__din = krnl_globalSort_L1_L2_3_out_dist_din;
  assign krnl_globalSort_L1_L2_3_out_dist_full_n = L1_out_dist_3__full_n;
  assign L1_out_dist_3__write = krnl_globalSort_L1_L2_3_out_dist_write;
  assign L1_out_id_3__din = krnl_globalSort_L1_L2_3_out_id_din;
  assign krnl_globalSort_L1_L2_3_out_id_full_n = L1_out_id_3__full_n;
  assign L1_out_id_3__write = krnl_globalSort_L1_L2_3_out_id_write;
  assign krnl_globalSort_L1_L2_4_ap_clk = ap_clk;
  assign krnl_globalSort_L1_L2_4__ap_done = krnl_globalSort_L1_L2_4_ap_done;
  assign krnl_globalSort_L1_L2_4__ap_idle = krnl_globalSort_L1_L2_4_ap_idle;
  assign krnl_globalSort_L1_L2_4__ap_ready = krnl_globalSort_L1_L2_4_ap_ready;
  assign krnl_globalSort_L1_L2_4_ap_rst_n = ap_rst_n;
  assign krnl_globalSort_L1_L2_4_ap_start = krnl_globalSort_L1_L2_4__ap_start;
  assign krnl_globalSort_L1_L2_4_in_dist0_peek_dout = out_dist_12__dout;
  assign krnl_globalSort_L1_L2_4_in_dist0_peek_empty_n = out_dist_12__empty_n;
  assign krnl_globalSort_L1_L2_4_in_dist0_s_dout = out_dist_12__dout;
  assign krnl_globalSort_L1_L2_4_in_dist0_s_empty_n = out_dist_12__empty_n;
  assign out_dist_12__read = krnl_globalSort_L1_L2_4_in_dist0_s_read;
  assign krnl_globalSort_L1_L2_4_in_dist1_peek_dout = out_dist_13__dout;
  assign krnl_globalSort_L1_L2_4_in_dist1_peek_empty_n = out_dist_13__empty_n;
  assign krnl_globalSort_L1_L2_4_in_dist1_s_dout = out_dist_13__dout;
  assign krnl_globalSort_L1_L2_4_in_dist1_s_empty_n = out_dist_13__empty_n;
  assign out_dist_13__read = krnl_globalSort_L1_L2_4_in_dist1_s_read;
  assign krnl_globalSort_L1_L2_4_in_dist2_peek_dout = out_dist_14__dout;
  assign krnl_globalSort_L1_L2_4_in_dist2_peek_empty_n = out_dist_14__empty_n;
  assign krnl_globalSort_L1_L2_4_in_dist2_s_dout = out_dist_14__dout;
  assign krnl_globalSort_L1_L2_4_in_dist2_s_empty_n = out_dist_14__empty_n;
  assign out_dist_14__read = krnl_globalSort_L1_L2_4_in_dist2_s_read;
  assign krnl_globalSort_L1_L2_4_in_id0_peek_dout = out_id_12__dout;
  assign krnl_globalSort_L1_L2_4_in_id0_peek_empty_n = out_id_12__empty_n;
  assign krnl_globalSort_L1_L2_4_in_id0_s_dout = out_id_12__dout;
  assign krnl_globalSort_L1_L2_4_in_id0_s_empty_n = out_id_12__empty_n;
  assign out_id_12__read = krnl_globalSort_L1_L2_4_in_id0_s_read;
  assign krnl_globalSort_L1_L2_4_in_id1_peek_dout = out_id_13__dout;
  assign krnl_globalSort_L1_L2_4_in_id1_peek_empty_n = out_id_13__empty_n;
  assign krnl_globalSort_L1_L2_4_in_id1_s_dout = out_id_13__dout;
  assign krnl_globalSort_L1_L2_4_in_id1_s_empty_n = out_id_13__empty_n;
  assign out_id_13__read = krnl_globalSort_L1_L2_4_in_id1_s_read;
  assign krnl_globalSort_L1_L2_4_in_id2_peek_dout = out_id_14__dout;
  assign krnl_globalSort_L1_L2_4_in_id2_peek_empty_n = out_id_14__empty_n;
  assign krnl_globalSort_L1_L2_4_in_id2_s_dout = out_id_14__dout;
  assign krnl_globalSort_L1_L2_4_in_id2_s_empty_n = out_id_14__empty_n;
  assign out_id_14__read = krnl_globalSort_L1_L2_4_in_id2_s_read;
  assign L1_out_dist_4__din = krnl_globalSort_L1_L2_4_out_dist_din;
  assign krnl_globalSort_L1_L2_4_out_dist_full_n = L1_out_dist_4__full_n;
  assign L1_out_dist_4__write = krnl_globalSort_L1_L2_4_out_dist_write;
  assign L1_out_id_4__din = krnl_globalSort_L1_L2_4_out_id_din;
  assign krnl_globalSort_L1_L2_4_out_id_full_n = L1_out_id_4__full_n;
  assign L1_out_id_4__write = krnl_globalSort_L1_L2_4_out_id_write;
  assign krnl_globalSort_L1_L2_5_ap_clk = ap_clk;
  assign krnl_globalSort_L1_L2_5__ap_done = krnl_globalSort_L1_L2_5_ap_done;
  assign krnl_globalSort_L1_L2_5__ap_idle = krnl_globalSort_L1_L2_5_ap_idle;
  assign krnl_globalSort_L1_L2_5__ap_ready = krnl_globalSort_L1_L2_5_ap_ready;
  assign krnl_globalSort_L1_L2_5_ap_rst_n = ap_rst_n;
  assign krnl_globalSort_L1_L2_5_ap_start = krnl_globalSort_L1_L2_5__ap_start;
  assign krnl_globalSort_L1_L2_5_in_dist0_peek_dout = out_dist_15__dout;
  assign krnl_globalSort_L1_L2_5_in_dist0_peek_empty_n = out_dist_15__empty_n;
  assign krnl_globalSort_L1_L2_5_in_dist0_s_dout = out_dist_15__dout;
  assign krnl_globalSort_L1_L2_5_in_dist0_s_empty_n = out_dist_15__empty_n;
  assign out_dist_15__read = krnl_globalSort_L1_L2_5_in_dist0_s_read;
  assign krnl_globalSort_L1_L2_5_in_dist1_peek_dout = out_dist_16__dout;
  assign krnl_globalSort_L1_L2_5_in_dist1_peek_empty_n = out_dist_16__empty_n;
  assign krnl_globalSort_L1_L2_5_in_dist1_s_dout = out_dist_16__dout;
  assign krnl_globalSort_L1_L2_5_in_dist1_s_empty_n = out_dist_16__empty_n;
  assign out_dist_16__read = krnl_globalSort_L1_L2_5_in_dist1_s_read;
  assign krnl_globalSort_L1_L2_5_in_dist2_peek_dout = out_dist_17__dout;
  assign krnl_globalSort_L1_L2_5_in_dist2_peek_empty_n = out_dist_17__empty_n;
  assign krnl_globalSort_L1_L2_5_in_dist2_s_dout = out_dist_17__dout;
  assign krnl_globalSort_L1_L2_5_in_dist2_s_empty_n = out_dist_17__empty_n;
  assign out_dist_17__read = krnl_globalSort_L1_L2_5_in_dist2_s_read;
  assign krnl_globalSort_L1_L2_5_in_id0_peek_dout = out_id_15__dout;
  assign krnl_globalSort_L1_L2_5_in_id0_peek_empty_n = out_id_15__empty_n;
  assign krnl_globalSort_L1_L2_5_in_id0_s_dout = out_id_15__dout;
  assign krnl_globalSort_L1_L2_5_in_id0_s_empty_n = out_id_15__empty_n;
  assign out_id_15__read = krnl_globalSort_L1_L2_5_in_id0_s_read;
  assign krnl_globalSort_L1_L2_5_in_id1_peek_dout = out_id_16__dout;
  assign krnl_globalSort_L1_L2_5_in_id1_peek_empty_n = out_id_16__empty_n;
  assign krnl_globalSort_L1_L2_5_in_id1_s_dout = out_id_16__dout;
  assign krnl_globalSort_L1_L2_5_in_id1_s_empty_n = out_id_16__empty_n;
  assign out_id_16__read = krnl_globalSort_L1_L2_5_in_id1_s_read;
  assign krnl_globalSort_L1_L2_5_in_id2_peek_dout = out_id_17__dout;
  assign krnl_globalSort_L1_L2_5_in_id2_peek_empty_n = out_id_17__empty_n;
  assign krnl_globalSort_L1_L2_5_in_id2_s_dout = out_id_17__dout;
  assign krnl_globalSort_L1_L2_5_in_id2_s_empty_n = out_id_17__empty_n;
  assign out_id_17__read = krnl_globalSort_L1_L2_5_in_id2_s_read;
  assign L1_out_dist_5__din = krnl_globalSort_L1_L2_5_out_dist_din;
  assign krnl_globalSort_L1_L2_5_out_dist_full_n = L1_out_dist_5__full_n;
  assign L1_out_dist_5__write = krnl_globalSort_L1_L2_5_out_dist_write;
  assign L1_out_id_5__din = krnl_globalSort_L1_L2_5_out_id_din;
  assign krnl_globalSort_L1_L2_5_out_id_full_n = L1_out_id_5__full_n;
  assign L1_out_id_5__write = krnl_globalSort_L1_L2_5_out_id_write;
  assign krnl_globalSort_L1_L2_6_ap_clk = ap_clk;
  assign krnl_globalSort_L1_L2_6__ap_done = krnl_globalSort_L1_L2_6_ap_done;
  assign krnl_globalSort_L1_L2_6__ap_idle = krnl_globalSort_L1_L2_6_ap_idle;
  assign krnl_globalSort_L1_L2_6__ap_ready = krnl_globalSort_L1_L2_6_ap_ready;
  assign krnl_globalSort_L1_L2_6_ap_rst_n = ap_rst_n;
  assign krnl_globalSort_L1_L2_6_ap_start = krnl_globalSort_L1_L2_6__ap_start;
  assign krnl_globalSort_L1_L2_6_in_dist0_peek_dout = out_dist_18__dout;
  assign krnl_globalSort_L1_L2_6_in_dist0_peek_empty_n = out_dist_18__empty_n;
  assign krnl_globalSort_L1_L2_6_in_dist0_s_dout = out_dist_18__dout;
  assign krnl_globalSort_L1_L2_6_in_dist0_s_empty_n = out_dist_18__empty_n;
  assign out_dist_18__read = krnl_globalSort_L1_L2_6_in_dist0_s_read;
  assign krnl_globalSort_L1_L2_6_in_dist1_peek_dout = out_dist_19__dout;
  assign krnl_globalSort_L1_L2_6_in_dist1_peek_empty_n = out_dist_19__empty_n;
  assign krnl_globalSort_L1_L2_6_in_dist1_s_dout = out_dist_19__dout;
  assign krnl_globalSort_L1_L2_6_in_dist1_s_empty_n = out_dist_19__empty_n;
  assign out_dist_19__read = krnl_globalSort_L1_L2_6_in_dist1_s_read;
  assign krnl_globalSort_L1_L2_6_in_dist2_peek_dout = out_dist_20__dout;
  assign krnl_globalSort_L1_L2_6_in_dist2_peek_empty_n = out_dist_20__empty_n;
  assign krnl_globalSort_L1_L2_6_in_dist2_s_dout = out_dist_20__dout;
  assign krnl_globalSort_L1_L2_6_in_dist2_s_empty_n = out_dist_20__empty_n;
  assign out_dist_20__read = krnl_globalSort_L1_L2_6_in_dist2_s_read;
  assign krnl_globalSort_L1_L2_6_in_id0_peek_dout = out_id_18__dout;
  assign krnl_globalSort_L1_L2_6_in_id0_peek_empty_n = out_id_18__empty_n;
  assign krnl_globalSort_L1_L2_6_in_id0_s_dout = out_id_18__dout;
  assign krnl_globalSort_L1_L2_6_in_id0_s_empty_n = out_id_18__empty_n;
  assign out_id_18__read = krnl_globalSort_L1_L2_6_in_id0_s_read;
  assign krnl_globalSort_L1_L2_6_in_id1_peek_dout = out_id_19__dout;
  assign krnl_globalSort_L1_L2_6_in_id1_peek_empty_n = out_id_19__empty_n;
  assign krnl_globalSort_L1_L2_6_in_id1_s_dout = out_id_19__dout;
  assign krnl_globalSort_L1_L2_6_in_id1_s_empty_n = out_id_19__empty_n;
  assign out_id_19__read = krnl_globalSort_L1_L2_6_in_id1_s_read;
  assign krnl_globalSort_L1_L2_6_in_id2_peek_dout = out_id_20__dout;
  assign krnl_globalSort_L1_L2_6_in_id2_peek_empty_n = out_id_20__empty_n;
  assign krnl_globalSort_L1_L2_6_in_id2_s_dout = out_id_20__dout;
  assign krnl_globalSort_L1_L2_6_in_id2_s_empty_n = out_id_20__empty_n;
  assign out_id_20__read = krnl_globalSort_L1_L2_6_in_id2_s_read;
  assign L1_out_dist_6__din = krnl_globalSort_L1_L2_6_out_dist_din;
  assign krnl_globalSort_L1_L2_6_out_dist_full_n = L1_out_dist_6__full_n;
  assign L1_out_dist_6__write = krnl_globalSort_L1_L2_6_out_dist_write;
  assign L1_out_id_6__din = krnl_globalSort_L1_L2_6_out_id_din;
  assign krnl_globalSort_L1_L2_6_out_id_full_n = L1_out_id_6__full_n;
  assign L1_out_id_6__write = krnl_globalSort_L1_L2_6_out_id_write;
  assign krnl_globalSort_L1_L2_7_ap_clk = ap_clk;
  assign krnl_globalSort_L1_L2_7__ap_done = krnl_globalSort_L1_L2_7_ap_done;
  assign krnl_globalSort_L1_L2_7__ap_idle = krnl_globalSort_L1_L2_7_ap_idle;
  assign krnl_globalSort_L1_L2_7__ap_ready = krnl_globalSort_L1_L2_7_ap_ready;
  assign krnl_globalSort_L1_L2_7_ap_rst_n = ap_rst_n;
  assign krnl_globalSort_L1_L2_7_ap_start = krnl_globalSort_L1_L2_7__ap_start;
  assign krnl_globalSort_L1_L2_7_in_dist0_peek_dout = out_dist_21__dout;
  assign krnl_globalSort_L1_L2_7_in_dist0_peek_empty_n = out_dist_21__empty_n;
  assign krnl_globalSort_L1_L2_7_in_dist0_s_dout = out_dist_21__dout;
  assign krnl_globalSort_L1_L2_7_in_dist0_s_empty_n = out_dist_21__empty_n;
  assign out_dist_21__read = krnl_globalSort_L1_L2_7_in_dist0_s_read;
  assign krnl_globalSort_L1_L2_7_in_dist1_peek_dout = out_dist_22__dout;
  assign krnl_globalSort_L1_L2_7_in_dist1_peek_empty_n = out_dist_22__empty_n;
  assign krnl_globalSort_L1_L2_7_in_dist1_s_dout = out_dist_22__dout;
  assign krnl_globalSort_L1_L2_7_in_dist1_s_empty_n = out_dist_22__empty_n;
  assign out_dist_22__read = krnl_globalSort_L1_L2_7_in_dist1_s_read;
  assign krnl_globalSort_L1_L2_7_in_dist2_peek_dout = out_dist_23__dout;
  assign krnl_globalSort_L1_L2_7_in_dist2_peek_empty_n = out_dist_23__empty_n;
  assign krnl_globalSort_L1_L2_7_in_dist2_s_dout = out_dist_23__dout;
  assign krnl_globalSort_L1_L2_7_in_dist2_s_empty_n = out_dist_23__empty_n;
  assign out_dist_23__read = krnl_globalSort_L1_L2_7_in_dist2_s_read;
  assign krnl_globalSort_L1_L2_7_in_id0_peek_dout = out_id_21__dout;
  assign krnl_globalSort_L1_L2_7_in_id0_peek_empty_n = out_id_21__empty_n;
  assign krnl_globalSort_L1_L2_7_in_id0_s_dout = out_id_21__dout;
  assign krnl_globalSort_L1_L2_7_in_id0_s_empty_n = out_id_21__empty_n;
  assign out_id_21__read = krnl_globalSort_L1_L2_7_in_id0_s_read;
  assign krnl_globalSort_L1_L2_7_in_id1_peek_dout = out_id_22__dout;
  assign krnl_globalSort_L1_L2_7_in_id1_peek_empty_n = out_id_22__empty_n;
  assign krnl_globalSort_L1_L2_7_in_id1_s_dout = out_id_22__dout;
  assign krnl_globalSort_L1_L2_7_in_id1_s_empty_n = out_id_22__empty_n;
  assign out_id_22__read = krnl_globalSort_L1_L2_7_in_id1_s_read;
  assign krnl_globalSort_L1_L2_7_in_id2_peek_dout = out_id_23__dout;
  assign krnl_globalSort_L1_L2_7_in_id2_peek_empty_n = out_id_23__empty_n;
  assign krnl_globalSort_L1_L2_7_in_id2_s_dout = out_id_23__dout;
  assign krnl_globalSort_L1_L2_7_in_id2_s_empty_n = out_id_23__empty_n;
  assign out_id_23__read = krnl_globalSort_L1_L2_7_in_id2_s_read;
  assign L1_out_dist_7__din = krnl_globalSort_L1_L2_7_out_dist_din;
  assign krnl_globalSort_L1_L2_7_out_dist_full_n = L1_out_dist_7__full_n;
  assign L1_out_dist_7__write = krnl_globalSort_L1_L2_7_out_dist_write;
  assign L1_out_id_7__din = krnl_globalSort_L1_L2_7_out_id_din;
  assign krnl_globalSort_L1_L2_7_out_id_full_n = L1_out_id_7__full_n;
  assign L1_out_id_7__write = krnl_globalSort_L1_L2_7_out_id_write;
  assign krnl_globalSort_L1_L2_8_ap_clk = ap_clk;
  assign krnl_globalSort_L1_L2_8__ap_done = krnl_globalSort_L1_L2_8_ap_done;
  assign krnl_globalSort_L1_L2_8__ap_idle = krnl_globalSort_L1_L2_8_ap_idle;
  assign krnl_globalSort_L1_L2_8__ap_ready = krnl_globalSort_L1_L2_8_ap_ready;
  assign krnl_globalSort_L1_L2_8_ap_rst_n = ap_rst_n;
  assign krnl_globalSort_L1_L2_8_ap_start = krnl_globalSort_L1_L2_8__ap_start;
  assign krnl_globalSort_L1_L2_8_in_dist0_peek_dout = out_dist_24__dout;
  assign krnl_globalSort_L1_L2_8_in_dist0_peek_empty_n = out_dist_24__empty_n;
  assign krnl_globalSort_L1_L2_8_in_dist0_s_dout = out_dist_24__dout;
  assign krnl_globalSort_L1_L2_8_in_dist0_s_empty_n = out_dist_24__empty_n;
  assign out_dist_24__read = krnl_globalSort_L1_L2_8_in_dist0_s_read;
  assign krnl_globalSort_L1_L2_8_in_dist1_peek_dout = out_dist_25__dout;
  assign krnl_globalSort_L1_L2_8_in_dist1_peek_empty_n = out_dist_25__empty_n;
  assign krnl_globalSort_L1_L2_8_in_dist1_s_dout = out_dist_25__dout;
  assign krnl_globalSort_L1_L2_8_in_dist1_s_empty_n = out_dist_25__empty_n;
  assign out_dist_25__read = krnl_globalSort_L1_L2_8_in_dist1_s_read;
  assign krnl_globalSort_L1_L2_8_in_dist2_peek_dout = out_dist_26__dout;
  assign krnl_globalSort_L1_L2_8_in_dist2_peek_empty_n = out_dist_26__empty_n;
  assign krnl_globalSort_L1_L2_8_in_dist2_s_dout = out_dist_26__dout;
  assign krnl_globalSort_L1_L2_8_in_dist2_s_empty_n = out_dist_26__empty_n;
  assign out_dist_26__read = krnl_globalSort_L1_L2_8_in_dist2_s_read;
  assign krnl_globalSort_L1_L2_8_in_id0_peek_dout = out_id_24__dout;
  assign krnl_globalSort_L1_L2_8_in_id0_peek_empty_n = out_id_24__empty_n;
  assign krnl_globalSort_L1_L2_8_in_id0_s_dout = out_id_24__dout;
  assign krnl_globalSort_L1_L2_8_in_id0_s_empty_n = out_id_24__empty_n;
  assign out_id_24__read = krnl_globalSort_L1_L2_8_in_id0_s_read;
  assign krnl_globalSort_L1_L2_8_in_id1_peek_dout = out_id_25__dout;
  assign krnl_globalSort_L1_L2_8_in_id1_peek_empty_n = out_id_25__empty_n;
  assign krnl_globalSort_L1_L2_8_in_id1_s_dout = out_id_25__dout;
  assign krnl_globalSort_L1_L2_8_in_id1_s_empty_n = out_id_25__empty_n;
  assign out_id_25__read = krnl_globalSort_L1_L2_8_in_id1_s_read;
  assign krnl_globalSort_L1_L2_8_in_id2_peek_dout = out_id_26__dout;
  assign krnl_globalSort_L1_L2_8_in_id2_peek_empty_n = out_id_26__empty_n;
  assign krnl_globalSort_L1_L2_8_in_id2_s_dout = out_id_26__dout;
  assign krnl_globalSort_L1_L2_8_in_id2_s_empty_n = out_id_26__empty_n;
  assign out_id_26__read = krnl_globalSort_L1_L2_8_in_id2_s_read;
  assign L1_out_dist_8__din = krnl_globalSort_L1_L2_8_out_dist_din;
  assign krnl_globalSort_L1_L2_8_out_dist_full_n = L1_out_dist_8__full_n;
  assign L1_out_dist_8__write = krnl_globalSort_L1_L2_8_out_dist_write;
  assign L1_out_id_8__din = krnl_globalSort_L1_L2_8_out_id_din;
  assign krnl_globalSort_L1_L2_8_out_id_full_n = L1_out_id_8__full_n;
  assign L1_out_id_8__write = krnl_globalSort_L1_L2_8_out_id_write;
  assign krnl_globalSort_L1_L2_9_ap_clk = ap_clk;
  assign krnl_globalSort_L1_L2_9__ap_done = krnl_globalSort_L1_L2_9_ap_done;
  assign krnl_globalSort_L1_L2_9__ap_idle = krnl_globalSort_L1_L2_9_ap_idle;
  assign krnl_globalSort_L1_L2_9__ap_ready = krnl_globalSort_L1_L2_9_ap_ready;
  assign krnl_globalSort_L1_L2_9_ap_rst_n = ap_rst_n;
  assign krnl_globalSort_L1_L2_9_ap_start = krnl_globalSort_L1_L2_9__ap_start;
  assign krnl_globalSort_L1_L2_9_in_dist0_peek_dout = L1_out_dist_0__dout;
  assign krnl_globalSort_L1_L2_9_in_dist0_peek_empty_n = L1_out_dist_0__empty_n;
  assign krnl_globalSort_L1_L2_9_in_dist0_s_dout = L1_out_dist_0__dout;
  assign krnl_globalSort_L1_L2_9_in_dist0_s_empty_n = L1_out_dist_0__empty_n;
  assign L1_out_dist_0__read = krnl_globalSort_L1_L2_9_in_dist0_s_read;
  assign krnl_globalSort_L1_L2_9_in_dist1_peek_dout = L1_out_dist_1__dout;
  assign krnl_globalSort_L1_L2_9_in_dist1_peek_empty_n = L1_out_dist_1__empty_n;
  assign krnl_globalSort_L1_L2_9_in_dist1_s_dout = L1_out_dist_1__dout;
  assign krnl_globalSort_L1_L2_9_in_dist1_s_empty_n = L1_out_dist_1__empty_n;
  assign L1_out_dist_1__read = krnl_globalSort_L1_L2_9_in_dist1_s_read;
  assign krnl_globalSort_L1_L2_9_in_dist2_peek_dout = L1_out_dist_2__dout;
  assign krnl_globalSort_L1_L2_9_in_dist2_peek_empty_n = L1_out_dist_2__empty_n;
  assign krnl_globalSort_L1_L2_9_in_dist2_s_dout = L1_out_dist_2__dout;
  assign krnl_globalSort_L1_L2_9_in_dist2_s_empty_n = L1_out_dist_2__empty_n;
  assign L1_out_dist_2__read = krnl_globalSort_L1_L2_9_in_dist2_s_read;
  assign krnl_globalSort_L1_L2_9_in_id0_peek_dout = L1_out_id_0__dout;
  assign krnl_globalSort_L1_L2_9_in_id0_peek_empty_n = L1_out_id_0__empty_n;
  assign krnl_globalSort_L1_L2_9_in_id0_s_dout = L1_out_id_0__dout;
  assign krnl_globalSort_L1_L2_9_in_id0_s_empty_n = L1_out_id_0__empty_n;
  assign L1_out_id_0__read = krnl_globalSort_L1_L2_9_in_id0_s_read;
  assign krnl_globalSort_L1_L2_9_in_id1_peek_dout = L1_out_id_1__dout;
  assign krnl_globalSort_L1_L2_9_in_id1_peek_empty_n = L1_out_id_1__empty_n;
  assign krnl_globalSort_L1_L2_9_in_id1_s_dout = L1_out_id_1__dout;
  assign krnl_globalSort_L1_L2_9_in_id1_s_empty_n = L1_out_id_1__empty_n;
  assign L1_out_id_1__read = krnl_globalSort_L1_L2_9_in_id1_s_read;
  assign krnl_globalSort_L1_L2_9_in_id2_peek_dout = L1_out_id_2__dout;
  assign krnl_globalSort_L1_L2_9_in_id2_peek_empty_n = L1_out_id_2__empty_n;
  assign krnl_globalSort_L1_L2_9_in_id2_s_dout = L1_out_id_2__dout;
  assign krnl_globalSort_L1_L2_9_in_id2_s_empty_n = L1_out_id_2__empty_n;
  assign L1_out_id_2__read = krnl_globalSort_L1_L2_9_in_id2_s_read;
  assign L2_out_dist0__din = krnl_globalSort_L1_L2_9_out_dist_din;
  assign krnl_globalSort_L1_L2_9_out_dist_full_n = L2_out_dist0__full_n;
  assign L2_out_dist0__write = krnl_globalSort_L1_L2_9_out_dist_write;
  assign L2_out_id0__din = krnl_globalSort_L1_L2_9_out_id_din;
  assign krnl_globalSort_L1_L2_9_out_id_full_n = L2_out_id0__full_n;
  assign L2_out_id0__write = krnl_globalSort_L1_L2_9_out_id_write;
  assign krnl_globalSort_L1_L2_10_ap_clk = ap_clk;
  assign krnl_globalSort_L1_L2_10__ap_done = krnl_globalSort_L1_L2_10_ap_done;
  assign krnl_globalSort_L1_L2_10__ap_idle = krnl_globalSort_L1_L2_10_ap_idle;
  assign krnl_globalSort_L1_L2_10__ap_ready = krnl_globalSort_L1_L2_10_ap_ready;
  assign krnl_globalSort_L1_L2_10_ap_rst_n = ap_rst_n;
  assign krnl_globalSort_L1_L2_10_ap_start = krnl_globalSort_L1_L2_10__ap_start;
  assign krnl_globalSort_L1_L2_10_in_dist0_peek_dout = L1_out_dist_3__dout;
  assign krnl_globalSort_L1_L2_10_in_dist0_peek_empty_n = L1_out_dist_3__empty_n;
  assign krnl_globalSort_L1_L2_10_in_dist0_s_dout = L1_out_dist_3__dout;
  assign krnl_globalSort_L1_L2_10_in_dist0_s_empty_n = L1_out_dist_3__empty_n;
  assign L1_out_dist_3__read = krnl_globalSort_L1_L2_10_in_dist0_s_read;
  assign krnl_globalSort_L1_L2_10_in_dist1_peek_dout = L1_out_dist_4__dout;
  assign krnl_globalSort_L1_L2_10_in_dist1_peek_empty_n = L1_out_dist_4__empty_n;
  assign krnl_globalSort_L1_L2_10_in_dist1_s_dout = L1_out_dist_4__dout;
  assign krnl_globalSort_L1_L2_10_in_dist1_s_empty_n = L1_out_dist_4__empty_n;
  assign L1_out_dist_4__read = krnl_globalSort_L1_L2_10_in_dist1_s_read;
  assign krnl_globalSort_L1_L2_10_in_dist2_peek_dout = L1_out_dist_5__dout;
  assign krnl_globalSort_L1_L2_10_in_dist2_peek_empty_n = L1_out_dist_5__empty_n;
  assign krnl_globalSort_L1_L2_10_in_dist2_s_dout = L1_out_dist_5__dout;
  assign krnl_globalSort_L1_L2_10_in_dist2_s_empty_n = L1_out_dist_5__empty_n;
  assign L1_out_dist_5__read = krnl_globalSort_L1_L2_10_in_dist2_s_read;
  assign krnl_globalSort_L1_L2_10_in_id0_peek_dout = L1_out_id_3__dout;
  assign krnl_globalSort_L1_L2_10_in_id0_peek_empty_n = L1_out_id_3__empty_n;
  assign krnl_globalSort_L1_L2_10_in_id0_s_dout = L1_out_id_3__dout;
  assign krnl_globalSort_L1_L2_10_in_id0_s_empty_n = L1_out_id_3__empty_n;
  assign L1_out_id_3__read = krnl_globalSort_L1_L2_10_in_id0_s_read;
  assign krnl_globalSort_L1_L2_10_in_id1_peek_dout = L1_out_id_4__dout;
  assign krnl_globalSort_L1_L2_10_in_id1_peek_empty_n = L1_out_id_4__empty_n;
  assign krnl_globalSort_L1_L2_10_in_id1_s_dout = L1_out_id_4__dout;
  assign krnl_globalSort_L1_L2_10_in_id1_s_empty_n = L1_out_id_4__empty_n;
  assign L1_out_id_4__read = krnl_globalSort_L1_L2_10_in_id1_s_read;
  assign krnl_globalSort_L1_L2_10_in_id2_peek_dout = L1_out_id_5__dout;
  assign krnl_globalSort_L1_L2_10_in_id2_peek_empty_n = L1_out_id_5__empty_n;
  assign krnl_globalSort_L1_L2_10_in_id2_s_dout = L1_out_id_5__dout;
  assign krnl_globalSort_L1_L2_10_in_id2_s_empty_n = L1_out_id_5__empty_n;
  assign L1_out_id_5__read = krnl_globalSort_L1_L2_10_in_id2_s_read;
  assign L2_out_dist1__din = krnl_globalSort_L1_L2_10_out_dist_din;
  assign krnl_globalSort_L1_L2_10_out_dist_full_n = L2_out_dist1__full_n;
  assign L2_out_dist1__write = krnl_globalSort_L1_L2_10_out_dist_write;
  assign L2_out_id1__din = krnl_globalSort_L1_L2_10_out_id_din;
  assign krnl_globalSort_L1_L2_10_out_id_full_n = L2_out_id1__full_n;
  assign L2_out_id1__write = krnl_globalSort_L1_L2_10_out_id_write;
  assign krnl_globalSort_L1_L2_11_ap_clk = ap_clk;
  assign krnl_globalSort_L1_L2_11__ap_done = krnl_globalSort_L1_L2_11_ap_done;
  assign krnl_globalSort_L1_L2_11__ap_idle = krnl_globalSort_L1_L2_11_ap_idle;
  assign krnl_globalSort_L1_L2_11__ap_ready = krnl_globalSort_L1_L2_11_ap_ready;
  assign krnl_globalSort_L1_L2_11_ap_rst_n = ap_rst_n;
  assign krnl_globalSort_L1_L2_11_ap_start = krnl_globalSort_L1_L2_11__ap_start;
  assign krnl_globalSort_L1_L2_11_in_dist0_peek_dout = L1_out_dist_6__dout;
  assign krnl_globalSort_L1_L2_11_in_dist0_peek_empty_n = L1_out_dist_6__empty_n;
  assign krnl_globalSort_L1_L2_11_in_dist0_s_dout = L1_out_dist_6__dout;
  assign krnl_globalSort_L1_L2_11_in_dist0_s_empty_n = L1_out_dist_6__empty_n;
  assign L1_out_dist_6__read = krnl_globalSort_L1_L2_11_in_dist0_s_read;
  assign krnl_globalSort_L1_L2_11_in_dist1_peek_dout = L1_out_dist_7__dout;
  assign krnl_globalSort_L1_L2_11_in_dist1_peek_empty_n = L1_out_dist_7__empty_n;
  assign krnl_globalSort_L1_L2_11_in_dist1_s_dout = L1_out_dist_7__dout;
  assign krnl_globalSort_L1_L2_11_in_dist1_s_empty_n = L1_out_dist_7__empty_n;
  assign L1_out_dist_7__read = krnl_globalSort_L1_L2_11_in_dist1_s_read;
  assign krnl_globalSort_L1_L2_11_in_dist2_peek_dout = L1_out_dist_8__dout;
  assign krnl_globalSort_L1_L2_11_in_dist2_peek_empty_n = L1_out_dist_8__empty_n;
  assign krnl_globalSort_L1_L2_11_in_dist2_s_dout = L1_out_dist_8__dout;
  assign krnl_globalSort_L1_L2_11_in_dist2_s_empty_n = L1_out_dist_8__empty_n;
  assign L1_out_dist_8__read = krnl_globalSort_L1_L2_11_in_dist2_s_read;
  assign krnl_globalSort_L1_L2_11_in_id0_peek_dout = L1_out_id_6__dout;
  assign krnl_globalSort_L1_L2_11_in_id0_peek_empty_n = L1_out_id_6__empty_n;
  assign krnl_globalSort_L1_L2_11_in_id0_s_dout = L1_out_id_6__dout;
  assign krnl_globalSort_L1_L2_11_in_id0_s_empty_n = L1_out_id_6__empty_n;
  assign L1_out_id_6__read = krnl_globalSort_L1_L2_11_in_id0_s_read;
  assign krnl_globalSort_L1_L2_11_in_id1_peek_dout = L1_out_id_7__dout;
  assign krnl_globalSort_L1_L2_11_in_id1_peek_empty_n = L1_out_id_7__empty_n;
  assign krnl_globalSort_L1_L2_11_in_id1_s_dout = L1_out_id_7__dout;
  assign krnl_globalSort_L1_L2_11_in_id1_s_empty_n = L1_out_id_7__empty_n;
  assign L1_out_id_7__read = krnl_globalSort_L1_L2_11_in_id1_s_read;
  assign krnl_globalSort_L1_L2_11_in_id2_peek_dout = L1_out_id_8__dout;
  assign krnl_globalSort_L1_L2_11_in_id2_peek_empty_n = L1_out_id_8__empty_n;
  assign krnl_globalSort_L1_L2_11_in_id2_s_dout = L1_out_id_8__dout;
  assign krnl_globalSort_L1_L2_11_in_id2_s_empty_n = L1_out_id_8__empty_n;
  assign L1_out_id_8__read = krnl_globalSort_L1_L2_11_in_id2_s_read;
  assign L2_out_dist2__din = krnl_globalSort_L1_L2_11_out_dist_din;
  assign krnl_globalSort_L1_L2_11_out_dist_full_n = L2_out_dist2__full_n;
  assign L2_out_dist2__write = krnl_globalSort_L1_L2_11_out_dist_write;
  assign L2_out_id2__din = krnl_globalSort_L1_L2_11_out_id_din;
  assign krnl_globalSort_L1_L2_11_out_id_full_n = L2_out_id2__full_n;
  assign L2_out_id2__write = krnl_globalSort_L1_L2_11_out_id_write;
  assign krnl_globalSort_L1_L2_12_ap_clk = ap_clk;
  assign krnl_globalSort_L1_L2_12__ap_done = krnl_globalSort_L1_L2_12_ap_done;
  assign krnl_globalSort_L1_L2_12__ap_idle = krnl_globalSort_L1_L2_12_ap_idle;
  assign krnl_globalSort_L1_L2_12__ap_ready = krnl_globalSort_L1_L2_12_ap_ready;
  assign krnl_globalSort_L1_L2_12_ap_rst_n = ap_rst_n;
  assign krnl_globalSort_L1_L2_12_ap_start = krnl_globalSort_L1_L2_12__ap_start;
  assign krnl_globalSort_L1_L2_12_in_dist0_peek_dout = L2_out_dist0__dout;
  assign krnl_globalSort_L1_L2_12_in_dist0_peek_empty_n = L2_out_dist0__empty_n;
  assign krnl_globalSort_L1_L2_12_in_dist0_s_dout = L2_out_dist0__dout;
  assign krnl_globalSort_L1_L2_12_in_dist0_s_empty_n = L2_out_dist0__empty_n;
  assign L2_out_dist0__read = krnl_globalSort_L1_L2_12_in_dist0_s_read;
  assign krnl_globalSort_L1_L2_12_in_dist1_peek_dout = L2_out_dist1__dout;
  assign krnl_globalSort_L1_L2_12_in_dist1_peek_empty_n = L2_out_dist1__empty_n;
  assign krnl_globalSort_L1_L2_12_in_dist1_s_dout = L2_out_dist1__dout;
  assign krnl_globalSort_L1_L2_12_in_dist1_s_empty_n = L2_out_dist1__empty_n;
  assign L2_out_dist1__read = krnl_globalSort_L1_L2_12_in_dist1_s_read;
  assign krnl_globalSort_L1_L2_12_in_dist2_peek_dout = L2_out_dist2__dout;
  assign krnl_globalSort_L1_L2_12_in_dist2_peek_empty_n = L2_out_dist2__empty_n;
  assign krnl_globalSort_L1_L2_12_in_dist2_s_dout = L2_out_dist2__dout;
  assign krnl_globalSort_L1_L2_12_in_dist2_s_empty_n = L2_out_dist2__empty_n;
  assign L2_out_dist2__read = krnl_globalSort_L1_L2_12_in_dist2_s_read;
  assign krnl_globalSort_L1_L2_12_in_id0_peek_dout = L2_out_id0__dout;
  assign krnl_globalSort_L1_L2_12_in_id0_peek_empty_n = L2_out_id0__empty_n;
  assign krnl_globalSort_L1_L2_12_in_id0_s_dout = L2_out_id0__dout;
  assign krnl_globalSort_L1_L2_12_in_id0_s_empty_n = L2_out_id0__empty_n;
  assign L2_out_id0__read = krnl_globalSort_L1_L2_12_in_id0_s_read;
  assign krnl_globalSort_L1_L2_12_in_id1_peek_dout = L2_out_id1__dout;
  assign krnl_globalSort_L1_L2_12_in_id1_peek_empty_n = L2_out_id1__empty_n;
  assign krnl_globalSort_L1_L2_12_in_id1_s_dout = L2_out_id1__dout;
  assign krnl_globalSort_L1_L2_12_in_id1_s_empty_n = L2_out_id1__empty_n;
  assign L2_out_id1__read = krnl_globalSort_L1_L2_12_in_id1_s_read;
  assign krnl_globalSort_L1_L2_12_in_id2_peek_dout = L2_out_id2__dout;
  assign krnl_globalSort_L1_L2_12_in_id2_peek_empty_n = L2_out_id2__empty_n;
  assign krnl_globalSort_L1_L2_12_in_id2_s_dout = L2_out_id2__dout;
  assign krnl_globalSort_L1_L2_12_in_id2_s_empty_n = L2_out_id2__empty_n;
  assign L2_out_id2__read = krnl_globalSort_L1_L2_12_in_id2_s_read;
  assign L3_out_dist_stream__din = krnl_globalSort_L1_L2_12_out_dist_din;
  assign krnl_globalSort_L1_L2_12_out_dist_full_n = L3_out_dist_stream__full_n;
  assign L3_out_dist_stream__write = krnl_globalSort_L1_L2_12_out_dist_write;
  assign L3_out_id_stream__din = krnl_globalSort_L1_L2_12_out_id_din;
  assign krnl_globalSort_L1_L2_12_out_id_full_n = L3_out_id_stream__full_n;
  assign L3_out_id_stream__write = krnl_globalSort_L1_L2_12_out_id_write;
  assign krnl_output_dist_id_0_ap_clk = ap_clk;
  assign krnl_output_dist_id_0__ap_done = krnl_output_dist_id_0_ap_done;
  assign krnl_output_dist_id_0__ap_idle = krnl_output_dist_id_0_ap_idle;
  assign krnl_output_dist_id_0__ap_ready = krnl_output_dist_id_0_ap_ready;
  assign krnl_output_dist_id_0_ap_rst_n = ap_rst_n;
  assign krnl_output_dist_id_0_ap_start = krnl_output_dist_id_0__ap_start;
  assign krnl_output_dist_id_0_in_dist_peek_dout = L3_out_dist_stream__dout;
  assign krnl_output_dist_id_0_in_dist_peek_empty_n = L3_out_dist_stream__empty_n;
  assign krnl_output_dist_id_0_in_dist_s_dout = L3_out_dist_stream__dout;
  assign krnl_output_dist_id_0_in_dist_s_empty_n = L3_out_dist_stream__empty_n;
  assign L3_out_dist_stream__read = krnl_output_dist_id_0_in_dist_s_read;
  assign krnl_output_dist_id_0_in_id_peek_dout = L3_out_id_stream__dout;
  assign krnl_output_dist_id_0_in_id_peek_empty_n = L3_out_id_stream__empty_n;
  assign krnl_output_dist_id_0_in_id_s_dout = L3_out_id_stream__dout;
  assign krnl_output_dist_id_0_in_id_s_empty_n = L3_out_id_stream__empty_n;
  assign L3_out_id_stream__read = krnl_output_dist_id_0_in_id_s_read;
  assign krnl_output_dist_id_0_output_knnDist_read_addr_offset = krnl_output_dist_id_0___L3_out_dist__q0;
  assign L3_out_dist_read_addr__din = krnl_output_dist_id_0_output_knnDist_read_addr_s_din;
  assign krnl_output_dist_id_0_output_knnDist_read_addr_s_full_n = L3_out_dist_read_addr__full_n;
  assign L3_out_dist_read_addr__write = krnl_output_dist_id_0_output_knnDist_read_addr_s_write;
  assign krnl_output_dist_id_0_output_knnDist_read_data_peek_dout = { 1'b0 , L3_out_dist_read_data__dout };
  assign krnl_output_dist_id_0_output_knnDist_read_data_peek_empty_n = L3_out_dist_read_data__empty_n;
  assign krnl_output_dist_id_0_output_knnDist_read_data_s_dout = { 1'b0 , L3_out_dist_read_data__dout };
  assign krnl_output_dist_id_0_output_knnDist_read_data_s_empty_n = L3_out_dist_read_data__empty_n;
  assign L3_out_dist_read_data__read = krnl_output_dist_id_0_output_knnDist_read_data_s_read;
  assign krnl_output_dist_id_0_output_knnDist_write_addr_offset = krnl_output_dist_id_0___L3_out_dist__q0;
  assign L3_out_dist_write_addr__din = krnl_output_dist_id_0_output_knnDist_write_addr_s_din;
  assign krnl_output_dist_id_0_output_knnDist_write_addr_s_full_n = L3_out_dist_write_addr__full_n;
  assign L3_out_dist_write_addr__write = krnl_output_dist_id_0_output_knnDist_write_addr_s_write;
  assign L3_out_dist_write_data__din = krnl_output_dist_id_0_output_knnDist_write_data_din;
  assign krnl_output_dist_id_0_output_knnDist_write_data_full_n = L3_out_dist_write_data__full_n;
  assign L3_out_dist_write_data__write = krnl_output_dist_id_0_output_knnDist_write_data_write;
  assign krnl_output_dist_id_0_output_knnDist_write_resp_peek_dout = { 1'b0 , L3_out_dist_write_resp__dout };
  assign krnl_output_dist_id_0_output_knnDist_write_resp_peek_empty_n = L3_out_dist_write_resp__empty_n;
  assign krnl_output_dist_id_0_output_knnDist_write_resp_s_dout = { 1'b0 , L3_out_dist_write_resp__dout };
  assign krnl_output_dist_id_0_output_knnDist_write_resp_s_empty_n = L3_out_dist_write_resp__empty_n;
  assign L3_out_dist_write_resp__read = krnl_output_dist_id_0_output_knnDist_write_resp_s_read;
  assign krnl_output_dist_id_0_output_knnId_read_addr_offset = krnl_output_dist_id_0___L3_out_id__q0;
  assign L3_out_id_read_addr__din = krnl_output_dist_id_0_output_knnId_read_addr_s_din;
  assign krnl_output_dist_id_0_output_knnId_read_addr_s_full_n = L3_out_id_read_addr__full_n;
  assign L3_out_id_read_addr__write = krnl_output_dist_id_0_output_knnId_read_addr_s_write;
  assign krnl_output_dist_id_0_output_knnId_read_data_peek_dout = { 1'b0 , L3_out_id_read_data__dout };
  assign krnl_output_dist_id_0_output_knnId_read_data_peek_empty_n = L3_out_id_read_data__empty_n;
  assign krnl_output_dist_id_0_output_knnId_read_data_s_dout = { 1'b0 , L3_out_id_read_data__dout };
  assign krnl_output_dist_id_0_output_knnId_read_data_s_empty_n = L3_out_id_read_data__empty_n;
  assign L3_out_id_read_data__read = krnl_output_dist_id_0_output_knnId_read_data_s_read;
  assign krnl_output_dist_id_0_output_knnId_write_addr_offset = krnl_output_dist_id_0___L3_out_id__q0;
  assign L3_out_id_write_addr__din = krnl_output_dist_id_0_output_knnId_write_addr_s_din;
  assign krnl_output_dist_id_0_output_knnId_write_addr_s_full_n = L3_out_id_write_addr__full_n;
  assign L3_out_id_write_addr__write = krnl_output_dist_id_0_output_knnId_write_addr_s_write;
  assign L3_out_id_write_data__din = krnl_output_dist_id_0_output_knnId_write_data_din;
  assign krnl_output_dist_id_0_output_knnId_write_data_full_n = L3_out_id_write_data__full_n;
  assign L3_out_id_write_data__write = krnl_output_dist_id_0_output_knnId_write_data_write;
  assign krnl_output_dist_id_0_output_knnId_write_resp_peek_dout = { 1'b0 , L3_out_id_write_resp__dout };
  assign krnl_output_dist_id_0_output_knnId_write_resp_peek_empty_n = L3_out_id_write_resp__empty_n;
  assign krnl_output_dist_id_0_output_knnId_write_resp_s_dout = { 1'b0 , L3_out_id_write_resp__dout };
  assign krnl_output_dist_id_0_output_knnId_write_resp_s_empty_n = L3_out_id_write_resp__empty_n;
  assign L3_out_id_write_resp__read = krnl_output_dist_id_0_output_knnId_write_resp_s_read;
  assign krnl_partialKnn_wrapper_0_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_0_0__ap_done = krnl_partialKnn_wrapper_0_0_ap_done;
  assign krnl_partialKnn_wrapper_0_0__ap_idle = krnl_partialKnn_wrapper_0_0_ap_idle;
  assign krnl_partialKnn_wrapper_0_0__ap_ready = krnl_partialKnn_wrapper_0_0_ap_ready;
  assign krnl_partialKnn_wrapper_0_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_0_0_ap_start = krnl_partialKnn_wrapper_0_0__ap_start;
  assign out_dist_0__din = krnl_partialKnn_wrapper_0_0_out_dist_din;
  assign krnl_partialKnn_wrapper_0_0_out_dist_full_n = out_dist_0__full_n;
  assign out_dist_0__write = krnl_partialKnn_wrapper_0_0_out_dist_write;
  assign out_id_0__din = krnl_partialKnn_wrapper_0_0_out_id_din;
  assign krnl_partialKnn_wrapper_0_0_out_id_full_n = out_id_0__full_n;
  assign out_id_0__write = krnl_partialKnn_wrapper_0_0_out_id_write;
  assign krnl_partialKnn_wrapper_0_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_0_0___in_0__q0;
  assign in_0_read_addr__din = krnl_partialKnn_wrapper_0_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_0_0_searchSpace_0_read_addr_s_full_n = in_0_read_addr__full_n;
  assign in_0_read_addr__write = krnl_partialKnn_wrapper_0_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_0_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_0_read_data__dout };
  assign krnl_partialKnn_wrapper_0_0_searchSpace_0_read_data_peek_empty_n = in_0_read_data__empty_n;
  assign krnl_partialKnn_wrapper_0_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_0_read_data__dout };
  assign krnl_partialKnn_wrapper_0_0_searchSpace_0_read_data_s_empty_n = in_0_read_data__empty_n;
  assign in_0_read_data__read = krnl_partialKnn_wrapper_0_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_0_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_0_0___in_0__q0;
  assign in_0_write_addr__din = krnl_partialKnn_wrapper_0_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_0_0_searchSpace_0_write_addr_s_full_n = in_0_write_addr__full_n;
  assign in_0_write_addr__write = krnl_partialKnn_wrapper_0_0_searchSpace_0_write_addr_s_write;
  assign in_0_write_data__din = krnl_partialKnn_wrapper_0_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_0_0_searchSpace_0_write_data_full_n = in_0_write_data__full_n;
  assign in_0_write_data__write = krnl_partialKnn_wrapper_0_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_0_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_0_write_resp__dout };
  assign krnl_partialKnn_wrapper_0_0_searchSpace_write_resp_peek_empty_n = in_0_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_0_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_0_write_resp__dout };
  assign krnl_partialKnn_wrapper_0_0_searchSpace_0_write_resp_s_empty_n = in_0_write_resp__empty_n;
  assign in_0_write_resp__read = krnl_partialKnn_wrapper_0_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_0_0_start_id_0 = 64'd0;
  assign krnl_partialKnn_wrapper_1_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_1_0__ap_done = krnl_partialKnn_wrapper_1_0_ap_done;
  assign krnl_partialKnn_wrapper_1_0__ap_idle = krnl_partialKnn_wrapper_1_0_ap_idle;
  assign krnl_partialKnn_wrapper_1_0__ap_ready = krnl_partialKnn_wrapper_1_0_ap_ready;
  assign krnl_partialKnn_wrapper_1_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_1_0_ap_start = krnl_partialKnn_wrapper_1_0__ap_start;
  assign out_dist_1__din = krnl_partialKnn_wrapper_1_0_out_dist_din;
  assign krnl_partialKnn_wrapper_1_0_out_dist_full_n = out_dist_1__full_n;
  assign out_dist_1__write = krnl_partialKnn_wrapper_1_0_out_dist_write;
  assign out_id_1__din = krnl_partialKnn_wrapper_1_0_out_id_din;
  assign krnl_partialKnn_wrapper_1_0_out_id_full_n = out_id_1__full_n;
  assign out_id_1__write = krnl_partialKnn_wrapper_1_0_out_id_write;
  assign krnl_partialKnn_wrapper_1_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_1_0___in_1__q0;
  assign in_1_read_addr__din = krnl_partialKnn_wrapper_1_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_1_0_searchSpace_0_read_addr_s_full_n = in_1_read_addr__full_n;
  assign in_1_read_addr__write = krnl_partialKnn_wrapper_1_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_1_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_1_read_data__dout };
  assign krnl_partialKnn_wrapper_1_0_searchSpace_0_read_data_peek_empty_n = in_1_read_data__empty_n;
  assign krnl_partialKnn_wrapper_1_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_1_read_data__dout };
  assign krnl_partialKnn_wrapper_1_0_searchSpace_0_read_data_s_empty_n = in_1_read_data__empty_n;
  assign in_1_read_data__read = krnl_partialKnn_wrapper_1_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_1_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_1_0___in_1__q0;
  assign in_1_write_addr__din = krnl_partialKnn_wrapper_1_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_1_0_searchSpace_0_write_addr_s_full_n = in_1_write_addr__full_n;
  assign in_1_write_addr__write = krnl_partialKnn_wrapper_1_0_searchSpace_0_write_addr_s_write;
  assign in_1_write_data__din = krnl_partialKnn_wrapper_1_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_1_0_searchSpace_0_write_data_full_n = in_1_write_data__full_n;
  assign in_1_write_data__write = krnl_partialKnn_wrapper_1_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_1_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_1_write_resp__dout };
  assign krnl_partialKnn_wrapper_1_0_searchSpace_write_resp_peek_empty_n = in_1_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_1_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_1_write_resp__dout };
  assign krnl_partialKnn_wrapper_1_0_searchSpace_0_write_resp_s_empty_n = in_1_write_resp__empty_n;
  assign in_1_write_resp__read = krnl_partialKnn_wrapper_1_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_1_0_start_id_0 = 64'd8192;
  assign krnl_partialKnn_wrapper_10_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_10_0__ap_done = krnl_partialKnn_wrapper_10_0_ap_done;
  assign krnl_partialKnn_wrapper_10_0__ap_idle = krnl_partialKnn_wrapper_10_0_ap_idle;
  assign krnl_partialKnn_wrapper_10_0__ap_ready = krnl_partialKnn_wrapper_10_0_ap_ready;
  assign krnl_partialKnn_wrapper_10_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_10_0_ap_start = krnl_partialKnn_wrapper_10_0__ap_start;
  assign out_dist_10__din = krnl_partialKnn_wrapper_10_0_out_dist_din;
  assign krnl_partialKnn_wrapper_10_0_out_dist_full_n = out_dist_10__full_n;
  assign out_dist_10__write = krnl_partialKnn_wrapper_10_0_out_dist_write;
  assign out_id_10__din = krnl_partialKnn_wrapper_10_0_out_id_din;
  assign krnl_partialKnn_wrapper_10_0_out_id_full_n = out_id_10__full_n;
  assign out_id_10__write = krnl_partialKnn_wrapper_10_0_out_id_write;
  assign krnl_partialKnn_wrapper_10_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_10_0___in_10__q0;
  assign in_10_read_addr__din = krnl_partialKnn_wrapper_10_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_10_0_searchSpace_0_read_addr_s_full_n = in_10_read_addr__full_n;
  assign in_10_read_addr__write = krnl_partialKnn_wrapper_10_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_10_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_10_read_data__dout };
  assign krnl_partialKnn_wrapper_10_0_searchSpace_read_data_peek_empty_n = in_10_read_data__empty_n;
  assign krnl_partialKnn_wrapper_10_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_10_read_data__dout };
  assign krnl_partialKnn_wrapper_10_0_searchSpace_0_read_data_s_empty_n = in_10_read_data__empty_n;
  assign in_10_read_data__read = krnl_partialKnn_wrapper_10_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_10_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_10_0___in_10__q0;
  assign in_10_write_addr__din = krnl_partialKnn_wrapper_10_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_10_0_searchSpace_0_write_addr_s_full_n = in_10_write_addr__full_n;
  assign in_10_write_addr__write = krnl_partialKnn_wrapper_10_0_searchSpace_0_write_addr_s_write;
  assign in_10_write_data__din = krnl_partialKnn_wrapper_10_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_10_0_searchSpace_0_write_data_full_n = in_10_write_data__full_n;
  assign in_10_write_data__write = krnl_partialKnn_wrapper_10_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_10_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_10_write_resp__dout };
  assign krnl_partialKnn_wrapper_10_0_searchSpace_write_resp_peek_empty_n = in_10_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_10_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_10_write_resp__dout };
  assign krnl_partialKnn_wrapper_10_0_searchSpace_0_write_resp_s_empty_n = in_10_write_resp__empty_n;
  assign in_10_write_resp__read = krnl_partialKnn_wrapper_10_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_10_0_start_id_0 = 64'd81920;
  assign krnl_partialKnn_wrapper_11_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_11_0__ap_done = krnl_partialKnn_wrapper_11_0_ap_done;
  assign krnl_partialKnn_wrapper_11_0__ap_idle = krnl_partialKnn_wrapper_11_0_ap_idle;
  assign krnl_partialKnn_wrapper_11_0__ap_ready = krnl_partialKnn_wrapper_11_0_ap_ready;
  assign krnl_partialKnn_wrapper_11_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_11_0_ap_start = krnl_partialKnn_wrapper_11_0__ap_start;
  assign out_dist_11__din = krnl_partialKnn_wrapper_11_0_out_dist_din;
  assign krnl_partialKnn_wrapper_11_0_out_dist_full_n = out_dist_11__full_n;
  assign out_dist_11__write = krnl_partialKnn_wrapper_11_0_out_dist_write;
  assign out_id_11__din = krnl_partialKnn_wrapper_11_0_out_id_din;
  assign krnl_partialKnn_wrapper_11_0_out_id_full_n = out_id_11__full_n;
  assign out_id_11__write = krnl_partialKnn_wrapper_11_0_out_id_write;
  assign krnl_partialKnn_wrapper_11_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_11_0___in_11__q0;
  assign in_11_read_addr__din = krnl_partialKnn_wrapper_11_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_11_0_searchSpace_0_read_addr_s_full_n = in_11_read_addr__full_n;
  assign in_11_read_addr__write = krnl_partialKnn_wrapper_11_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_11_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_11_read_data__dout };
  assign krnl_partialKnn_wrapper_11_0_searchSpace_read_data_peek_empty_n = in_11_read_data__empty_n;
  assign krnl_partialKnn_wrapper_11_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_11_read_data__dout };
  assign krnl_partialKnn_wrapper_11_0_searchSpace_0_read_data_s_empty_n = in_11_read_data__empty_n;
  assign in_11_read_data__read = krnl_partialKnn_wrapper_11_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_11_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_11_0___in_11__q0;
  assign in_11_write_addr__din = krnl_partialKnn_wrapper_11_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_11_0_searchSpace_0_write_addr_s_full_n = in_11_write_addr__full_n;
  assign in_11_write_addr__write = krnl_partialKnn_wrapper_11_0_searchSpace_0_write_addr_s_write;
  assign in_11_write_data__din = krnl_partialKnn_wrapper_11_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_11_0_searchSpace_0_write_data_full_n = in_11_write_data__full_n;
  assign in_11_write_data__write = krnl_partialKnn_wrapper_11_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_11_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_11_write_resp__dout };
  assign krnl_partialKnn_wrapper_11_0_searchSpace_write_resp_peek_empty_n = in_11_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_11_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_11_write_resp__dout };
  assign krnl_partialKnn_wrapper_11_0_searchSpace_0_write_resp_s_empty_n = in_11_write_resp__empty_n;
  assign in_11_write_resp__read = krnl_partialKnn_wrapper_11_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_11_0_start_id_0 = 64'd90112;
  assign krnl_partialKnn_wrapper_12_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_12_0__ap_done = krnl_partialKnn_wrapper_12_0_ap_done;
  assign krnl_partialKnn_wrapper_12_0__ap_idle = krnl_partialKnn_wrapper_12_0_ap_idle;
  assign krnl_partialKnn_wrapper_12_0__ap_ready = krnl_partialKnn_wrapper_12_0_ap_ready;
  assign krnl_partialKnn_wrapper_12_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_12_0_ap_start = krnl_partialKnn_wrapper_12_0__ap_start;
  assign out_dist_12__din = krnl_partialKnn_wrapper_12_0_out_dist_din;
  assign krnl_partialKnn_wrapper_12_0_out_dist_full_n = out_dist_12__full_n;
  assign out_dist_12__write = krnl_partialKnn_wrapper_12_0_out_dist_write;
  assign out_id_12__din = krnl_partialKnn_wrapper_12_0_out_id_din;
  assign krnl_partialKnn_wrapper_12_0_out_id_full_n = out_id_12__full_n;
  assign out_id_12__write = krnl_partialKnn_wrapper_12_0_out_id_write;
  assign krnl_partialKnn_wrapper_12_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_12_0___in_12__q0;
  assign in_12_read_addr__din = krnl_partialKnn_wrapper_12_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_12_0_searchSpace_0_read_addr_s_full_n = in_12_read_addr__full_n;
  assign in_12_read_addr__write = krnl_partialKnn_wrapper_12_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_12_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_12_read_data__dout };
  assign krnl_partialKnn_wrapper_12_0_searchSpace_read_data_peek_empty_n = in_12_read_data__empty_n;
  assign krnl_partialKnn_wrapper_12_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_12_read_data__dout };
  assign krnl_partialKnn_wrapper_12_0_searchSpace_0_read_data_s_empty_n = in_12_read_data__empty_n;
  assign in_12_read_data__read = krnl_partialKnn_wrapper_12_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_12_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_12_0___in_12__q0;
  assign in_12_write_addr__din = krnl_partialKnn_wrapper_12_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_12_0_searchSpace_0_write_addr_s_full_n = in_12_write_addr__full_n;
  assign in_12_write_addr__write = krnl_partialKnn_wrapper_12_0_searchSpace_0_write_addr_s_write;
  assign in_12_write_data__din = krnl_partialKnn_wrapper_12_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_12_0_searchSpace_0_write_data_full_n = in_12_write_data__full_n;
  assign in_12_write_data__write = krnl_partialKnn_wrapper_12_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_12_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_12_write_resp__dout };
  assign krnl_partialKnn_wrapper_12_0_searchSpace_write_resp_peek_empty_n = in_12_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_12_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_12_write_resp__dout };
  assign krnl_partialKnn_wrapper_12_0_searchSpace_0_write_resp_s_empty_n = in_12_write_resp__empty_n;
  assign in_12_write_resp__read = krnl_partialKnn_wrapper_12_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_12_0_start_id_0 = 64'd98304;
  assign krnl_partialKnn_wrapper_13_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_13_0__ap_done = krnl_partialKnn_wrapper_13_0_ap_done;
  assign krnl_partialKnn_wrapper_13_0__ap_idle = krnl_partialKnn_wrapper_13_0_ap_idle;
  assign krnl_partialKnn_wrapper_13_0__ap_ready = krnl_partialKnn_wrapper_13_0_ap_ready;
  assign krnl_partialKnn_wrapper_13_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_13_0_ap_start = krnl_partialKnn_wrapper_13_0__ap_start;
  assign out_dist_13__din = krnl_partialKnn_wrapper_13_0_out_dist_din;
  assign krnl_partialKnn_wrapper_13_0_out_dist_full_n = out_dist_13__full_n;
  assign out_dist_13__write = krnl_partialKnn_wrapper_13_0_out_dist_write;
  assign out_id_13__din = krnl_partialKnn_wrapper_13_0_out_id_din;
  assign krnl_partialKnn_wrapper_13_0_out_id_full_n = out_id_13__full_n;
  assign out_id_13__write = krnl_partialKnn_wrapper_13_0_out_id_write;
  assign krnl_partialKnn_wrapper_13_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_13_0___in_13__q0;
  assign in_13_read_addr__din = krnl_partialKnn_wrapper_13_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_13_0_searchSpace_0_read_addr_s_full_n = in_13_read_addr__full_n;
  assign in_13_read_addr__write = krnl_partialKnn_wrapper_13_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_13_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_13_read_data__dout };
  assign krnl_partialKnn_wrapper_13_0_searchSpace_read_data_peek_empty_n = in_13_read_data__empty_n;
  assign krnl_partialKnn_wrapper_13_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_13_read_data__dout };
  assign krnl_partialKnn_wrapper_13_0_searchSpace_0_read_data_s_empty_n = in_13_read_data__empty_n;
  assign in_13_read_data__read = krnl_partialKnn_wrapper_13_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_13_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_13_0___in_13__q0;
  assign in_13_write_addr__din = krnl_partialKnn_wrapper_13_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_13_0_searchSpace_0_write_addr_s_full_n = in_13_write_addr__full_n;
  assign in_13_write_addr__write = krnl_partialKnn_wrapper_13_0_searchSpace_0_write_addr_s_write;
  assign in_13_write_data__din = krnl_partialKnn_wrapper_13_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_13_0_searchSpace_0_write_data_full_n = in_13_write_data__full_n;
  assign in_13_write_data__write = krnl_partialKnn_wrapper_13_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_13_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_13_write_resp__dout };
  assign krnl_partialKnn_wrapper_13_0_searchSpace_write_resp_peek_empty_n = in_13_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_13_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_13_write_resp__dout };
  assign krnl_partialKnn_wrapper_13_0_searchSpace_0_write_resp_s_empty_n = in_13_write_resp__empty_n;
  assign in_13_write_resp__read = krnl_partialKnn_wrapper_13_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_13_0_start_id_0 = 64'd106496;
  assign krnl_partialKnn_wrapper_14_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_14_0__ap_done = krnl_partialKnn_wrapper_14_0_ap_done;
  assign krnl_partialKnn_wrapper_14_0__ap_idle = krnl_partialKnn_wrapper_14_0_ap_idle;
  assign krnl_partialKnn_wrapper_14_0__ap_ready = krnl_partialKnn_wrapper_14_0_ap_ready;
  assign krnl_partialKnn_wrapper_14_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_14_0_ap_start = krnl_partialKnn_wrapper_14_0__ap_start;
  assign out_dist_14__din = krnl_partialKnn_wrapper_14_0_out_dist_din;
  assign krnl_partialKnn_wrapper_14_0_out_dist_full_n = out_dist_14__full_n;
  assign out_dist_14__write = krnl_partialKnn_wrapper_14_0_out_dist_write;
  assign out_id_14__din = krnl_partialKnn_wrapper_14_0_out_id_din;
  assign krnl_partialKnn_wrapper_14_0_out_id_full_n = out_id_14__full_n;
  assign out_id_14__write = krnl_partialKnn_wrapper_14_0_out_id_write;
  assign krnl_partialKnn_wrapper_14_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_14_0___in_14__q0;
  assign in_14_read_addr__din = krnl_partialKnn_wrapper_14_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_14_0_searchSpace_0_read_addr_s_full_n = in_14_read_addr__full_n;
  assign in_14_read_addr__write = krnl_partialKnn_wrapper_14_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_14_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_14_read_data__dout };
  assign krnl_partialKnn_wrapper_14_0_searchSpace_read_data_peek_empty_n = in_14_read_data__empty_n;
  assign krnl_partialKnn_wrapper_14_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_14_read_data__dout };
  assign krnl_partialKnn_wrapper_14_0_searchSpace_0_read_data_s_empty_n = in_14_read_data__empty_n;
  assign in_14_read_data__read = krnl_partialKnn_wrapper_14_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_14_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_14_0___in_14__q0;
  assign in_14_write_addr__din = krnl_partialKnn_wrapper_14_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_14_0_searchSpace_0_write_addr_s_full_n = in_14_write_addr__full_n;
  assign in_14_write_addr__write = krnl_partialKnn_wrapper_14_0_searchSpace_0_write_addr_s_write;
  assign in_14_write_data__din = krnl_partialKnn_wrapper_14_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_14_0_searchSpace_0_write_data_full_n = in_14_write_data__full_n;
  assign in_14_write_data__write = krnl_partialKnn_wrapper_14_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_14_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_14_write_resp__dout };
  assign krnl_partialKnn_wrapper_14_0_searchSpace_write_resp_peek_empty_n = in_14_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_14_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_14_write_resp__dout };
  assign krnl_partialKnn_wrapper_14_0_searchSpace_0_write_resp_s_empty_n = in_14_write_resp__empty_n;
  assign in_14_write_resp__read = krnl_partialKnn_wrapper_14_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_14_0_start_id_0 = 64'd114688;
  assign krnl_partialKnn_wrapper_15_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_15_0__ap_done = krnl_partialKnn_wrapper_15_0_ap_done;
  assign krnl_partialKnn_wrapper_15_0__ap_idle = krnl_partialKnn_wrapper_15_0_ap_idle;
  assign krnl_partialKnn_wrapper_15_0__ap_ready = krnl_partialKnn_wrapper_15_0_ap_ready;
  assign krnl_partialKnn_wrapper_15_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_15_0_ap_start = krnl_partialKnn_wrapper_15_0__ap_start;
  assign out_dist_15__din = krnl_partialKnn_wrapper_15_0_out_dist_din;
  assign krnl_partialKnn_wrapper_15_0_out_dist_full_n = out_dist_15__full_n;
  assign out_dist_15__write = krnl_partialKnn_wrapper_15_0_out_dist_write;
  assign out_id_15__din = krnl_partialKnn_wrapper_15_0_out_id_din;
  assign krnl_partialKnn_wrapper_15_0_out_id_full_n = out_id_15__full_n;
  assign out_id_15__write = krnl_partialKnn_wrapper_15_0_out_id_write;
  assign krnl_partialKnn_wrapper_15_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_15_0___in_15__q0;
  assign in_15_read_addr__din = krnl_partialKnn_wrapper_15_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_15_0_searchSpace_0_read_addr_s_full_n = in_15_read_addr__full_n;
  assign in_15_read_addr__write = krnl_partialKnn_wrapper_15_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_15_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_15_read_data__dout };
  assign krnl_partialKnn_wrapper_15_0_searchSpace_read_data_peek_empty_n = in_15_read_data__empty_n;
  assign krnl_partialKnn_wrapper_15_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_15_read_data__dout };
  assign krnl_partialKnn_wrapper_15_0_searchSpace_0_read_data_s_empty_n = in_15_read_data__empty_n;
  assign in_15_read_data__read = krnl_partialKnn_wrapper_15_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_15_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_15_0___in_15__q0;
  assign in_15_write_addr__din = krnl_partialKnn_wrapper_15_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_15_0_searchSpace_0_write_addr_s_full_n = in_15_write_addr__full_n;
  assign in_15_write_addr__write = krnl_partialKnn_wrapper_15_0_searchSpace_0_write_addr_s_write;
  assign in_15_write_data__din = krnl_partialKnn_wrapper_15_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_15_0_searchSpace_0_write_data_full_n = in_15_write_data__full_n;
  assign in_15_write_data__write = krnl_partialKnn_wrapper_15_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_15_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_15_write_resp__dout };
  assign krnl_partialKnn_wrapper_15_0_searchSpace_write_resp_peek_empty_n = in_15_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_15_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_15_write_resp__dout };
  assign krnl_partialKnn_wrapper_15_0_searchSpace_0_write_resp_s_empty_n = in_15_write_resp__empty_n;
  assign in_15_write_resp__read = krnl_partialKnn_wrapper_15_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_15_0_start_id_0 = 64'd122880;
  assign krnl_partialKnn_wrapper_16_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_16_0__ap_done = krnl_partialKnn_wrapper_16_0_ap_done;
  assign krnl_partialKnn_wrapper_16_0__ap_idle = krnl_partialKnn_wrapper_16_0_ap_idle;
  assign krnl_partialKnn_wrapper_16_0__ap_ready = krnl_partialKnn_wrapper_16_0_ap_ready;
  assign krnl_partialKnn_wrapper_16_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_16_0_ap_start = krnl_partialKnn_wrapper_16_0__ap_start;
  assign out_dist_16__din = krnl_partialKnn_wrapper_16_0_out_dist_din;
  assign krnl_partialKnn_wrapper_16_0_out_dist_full_n = out_dist_16__full_n;
  assign out_dist_16__write = krnl_partialKnn_wrapper_16_0_out_dist_write;
  assign out_id_16__din = krnl_partialKnn_wrapper_16_0_out_id_din;
  assign krnl_partialKnn_wrapper_16_0_out_id_full_n = out_id_16__full_n;
  assign out_id_16__write = krnl_partialKnn_wrapper_16_0_out_id_write;
  assign krnl_partialKnn_wrapper_16_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_16_0___in_16__q0;
  assign in_16_read_addr__din = krnl_partialKnn_wrapper_16_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_16_0_searchSpace_0_read_addr_s_full_n = in_16_read_addr__full_n;
  assign in_16_read_addr__write = krnl_partialKnn_wrapper_16_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_16_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_16_read_data__dout };
  assign krnl_partialKnn_wrapper_16_0_searchSpace_read_data_peek_empty_n = in_16_read_data__empty_n;
  assign krnl_partialKnn_wrapper_16_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_16_read_data__dout };
  assign krnl_partialKnn_wrapper_16_0_searchSpace_0_read_data_s_empty_n = in_16_read_data__empty_n;
  assign in_16_read_data__read = krnl_partialKnn_wrapper_16_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_16_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_16_0___in_16__q0;
  assign in_16_write_addr__din = krnl_partialKnn_wrapper_16_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_16_0_searchSpace_0_write_addr_s_full_n = in_16_write_addr__full_n;
  assign in_16_write_addr__write = krnl_partialKnn_wrapper_16_0_searchSpace_0_write_addr_s_write;
  assign in_16_write_data__din = krnl_partialKnn_wrapper_16_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_16_0_searchSpace_0_write_data_full_n = in_16_write_data__full_n;
  assign in_16_write_data__write = krnl_partialKnn_wrapper_16_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_16_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_16_write_resp__dout };
  assign krnl_partialKnn_wrapper_16_0_searchSpace_write_resp_peek_empty_n = in_16_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_16_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_16_write_resp__dout };
  assign krnl_partialKnn_wrapper_16_0_searchSpace_0_write_resp_s_empty_n = in_16_write_resp__empty_n;
  assign in_16_write_resp__read = krnl_partialKnn_wrapper_16_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_16_0_start_id_0 = 64'd131072;
  assign krnl_partialKnn_wrapper_17_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_17_0__ap_done = krnl_partialKnn_wrapper_17_0_ap_done;
  assign krnl_partialKnn_wrapper_17_0__ap_idle = krnl_partialKnn_wrapper_17_0_ap_idle;
  assign krnl_partialKnn_wrapper_17_0__ap_ready = krnl_partialKnn_wrapper_17_0_ap_ready;
  assign krnl_partialKnn_wrapper_17_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_17_0_ap_start = krnl_partialKnn_wrapper_17_0__ap_start;
  assign out_dist_17__din = krnl_partialKnn_wrapper_17_0_out_dist_din;
  assign krnl_partialKnn_wrapper_17_0_out_dist_full_n = out_dist_17__full_n;
  assign out_dist_17__write = krnl_partialKnn_wrapper_17_0_out_dist_write;
  assign out_id_17__din = krnl_partialKnn_wrapper_17_0_out_id_din;
  assign krnl_partialKnn_wrapper_17_0_out_id_full_n = out_id_17__full_n;
  assign out_id_17__write = krnl_partialKnn_wrapper_17_0_out_id_write;
  assign krnl_partialKnn_wrapper_17_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_17_0___in_17__q0;
  assign in_17_read_addr__din = krnl_partialKnn_wrapper_17_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_17_0_searchSpace_0_read_addr_s_full_n = in_17_read_addr__full_n;
  assign in_17_read_addr__write = krnl_partialKnn_wrapper_17_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_17_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_17_read_data__dout };
  assign krnl_partialKnn_wrapper_17_0_searchSpace_read_data_peek_empty_n = in_17_read_data__empty_n;
  assign krnl_partialKnn_wrapper_17_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_17_read_data__dout };
  assign krnl_partialKnn_wrapper_17_0_searchSpace_0_read_data_s_empty_n = in_17_read_data__empty_n;
  assign in_17_read_data__read = krnl_partialKnn_wrapper_17_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_17_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_17_0___in_17__q0;
  assign in_17_write_addr__din = krnl_partialKnn_wrapper_17_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_17_0_searchSpace_0_write_addr_s_full_n = in_17_write_addr__full_n;
  assign in_17_write_addr__write = krnl_partialKnn_wrapper_17_0_searchSpace_0_write_addr_s_write;
  assign in_17_write_data__din = krnl_partialKnn_wrapper_17_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_17_0_searchSpace_0_write_data_full_n = in_17_write_data__full_n;
  assign in_17_write_data__write = krnl_partialKnn_wrapper_17_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_17_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_17_write_resp__dout };
  assign krnl_partialKnn_wrapper_17_0_searchSpace_write_resp_peek_empty_n = in_17_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_17_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_17_write_resp__dout };
  assign krnl_partialKnn_wrapper_17_0_searchSpace_0_write_resp_s_empty_n = in_17_write_resp__empty_n;
  assign in_17_write_resp__read = krnl_partialKnn_wrapper_17_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_17_0_start_id_0 = 64'd139264;
  assign krnl_partialKnn_wrapper_18_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_18_0__ap_done = krnl_partialKnn_wrapper_18_0_ap_done;
  assign krnl_partialKnn_wrapper_18_0__ap_idle = krnl_partialKnn_wrapper_18_0_ap_idle;
  assign krnl_partialKnn_wrapper_18_0__ap_ready = krnl_partialKnn_wrapper_18_0_ap_ready;
  assign krnl_partialKnn_wrapper_18_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_18_0_ap_start = krnl_partialKnn_wrapper_18_0__ap_start;
  assign out_dist_18__din = krnl_partialKnn_wrapper_18_0_out_dist_din;
  assign krnl_partialKnn_wrapper_18_0_out_dist_full_n = out_dist_18__full_n;
  assign out_dist_18__write = krnl_partialKnn_wrapper_18_0_out_dist_write;
  assign out_id_18__din = krnl_partialKnn_wrapper_18_0_out_id_din;
  assign krnl_partialKnn_wrapper_18_0_out_id_full_n = out_id_18__full_n;
  assign out_id_18__write = krnl_partialKnn_wrapper_18_0_out_id_write;
  assign krnl_partialKnn_wrapper_18_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_18_0___in_18__q0;
  assign in_18_read_addr__din = krnl_partialKnn_wrapper_18_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_18_0_searchSpace_0_read_addr_s_full_n = in_18_read_addr__full_n;
  assign in_18_read_addr__write = krnl_partialKnn_wrapper_18_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_18_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_18_read_data__dout };
  assign krnl_partialKnn_wrapper_18_0_searchSpace_read_data_peek_empty_n = in_18_read_data__empty_n;
  assign krnl_partialKnn_wrapper_18_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_18_read_data__dout };
  assign krnl_partialKnn_wrapper_18_0_searchSpace_0_read_data_s_empty_n = in_18_read_data__empty_n;
  assign in_18_read_data__read = krnl_partialKnn_wrapper_18_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_18_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_18_0___in_18__q0;
  assign in_18_write_addr__din = krnl_partialKnn_wrapper_18_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_18_0_searchSpace_0_write_addr_s_full_n = in_18_write_addr__full_n;
  assign in_18_write_addr__write = krnl_partialKnn_wrapper_18_0_searchSpace_0_write_addr_s_write;
  assign in_18_write_data__din = krnl_partialKnn_wrapper_18_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_18_0_searchSpace_0_write_data_full_n = in_18_write_data__full_n;
  assign in_18_write_data__write = krnl_partialKnn_wrapper_18_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_18_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_18_write_resp__dout };
  assign krnl_partialKnn_wrapper_18_0_searchSpace_write_resp_peek_empty_n = in_18_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_18_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_18_write_resp__dout };
  assign krnl_partialKnn_wrapper_18_0_searchSpace_0_write_resp_s_empty_n = in_18_write_resp__empty_n;
  assign in_18_write_resp__read = krnl_partialKnn_wrapper_18_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_18_0_start_id_0 = 64'd147456;
  assign krnl_partialKnn_wrapper_19_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_19_0__ap_done = krnl_partialKnn_wrapper_19_0_ap_done;
  assign krnl_partialKnn_wrapper_19_0__ap_idle = krnl_partialKnn_wrapper_19_0_ap_idle;
  assign krnl_partialKnn_wrapper_19_0__ap_ready = krnl_partialKnn_wrapper_19_0_ap_ready;
  assign krnl_partialKnn_wrapper_19_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_19_0_ap_start = krnl_partialKnn_wrapper_19_0__ap_start;
  assign out_dist_19__din = krnl_partialKnn_wrapper_19_0_out_dist_din;
  assign krnl_partialKnn_wrapper_19_0_out_dist_full_n = out_dist_19__full_n;
  assign out_dist_19__write = krnl_partialKnn_wrapper_19_0_out_dist_write;
  assign out_id_19__din = krnl_partialKnn_wrapper_19_0_out_id_din;
  assign krnl_partialKnn_wrapper_19_0_out_id_full_n = out_id_19__full_n;
  assign out_id_19__write = krnl_partialKnn_wrapper_19_0_out_id_write;
  assign krnl_partialKnn_wrapper_19_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_19_0___in_19__q0;
  assign in_19_read_addr__din = krnl_partialKnn_wrapper_19_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_19_0_searchSpace_0_read_addr_s_full_n = in_19_read_addr__full_n;
  assign in_19_read_addr__write = krnl_partialKnn_wrapper_19_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_19_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_19_read_data__dout };
  assign krnl_partialKnn_wrapper_19_0_searchSpace_read_data_peek_empty_n = in_19_read_data__empty_n;
  assign krnl_partialKnn_wrapper_19_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_19_read_data__dout };
  assign krnl_partialKnn_wrapper_19_0_searchSpace_0_read_data_s_empty_n = in_19_read_data__empty_n;
  assign in_19_read_data__read = krnl_partialKnn_wrapper_19_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_19_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_19_0___in_19__q0;
  assign in_19_write_addr__din = krnl_partialKnn_wrapper_19_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_19_0_searchSpace_0_write_addr_s_full_n = in_19_write_addr__full_n;
  assign in_19_write_addr__write = krnl_partialKnn_wrapper_19_0_searchSpace_0_write_addr_s_write;
  assign in_19_write_data__din = krnl_partialKnn_wrapper_19_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_19_0_searchSpace_0_write_data_full_n = in_19_write_data__full_n;
  assign in_19_write_data__write = krnl_partialKnn_wrapper_19_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_19_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_19_write_resp__dout };
  assign krnl_partialKnn_wrapper_19_0_searchSpace_write_resp_peek_empty_n = in_19_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_19_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_19_write_resp__dout };
  assign krnl_partialKnn_wrapper_19_0_searchSpace_0_write_resp_s_empty_n = in_19_write_resp__empty_n;
  assign in_19_write_resp__read = krnl_partialKnn_wrapper_19_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_19_0_start_id_0 = 64'd155648;
  assign krnl_partialKnn_wrapper_2_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_2_0__ap_done = krnl_partialKnn_wrapper_2_0_ap_done;
  assign krnl_partialKnn_wrapper_2_0__ap_idle = krnl_partialKnn_wrapper_2_0_ap_idle;
  assign krnl_partialKnn_wrapper_2_0__ap_ready = krnl_partialKnn_wrapper_2_0_ap_ready;
  assign krnl_partialKnn_wrapper_2_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_2_0_ap_start = krnl_partialKnn_wrapper_2_0__ap_start;
  assign out_dist_2__din = krnl_partialKnn_wrapper_2_0_out_dist_din;
  assign krnl_partialKnn_wrapper_2_0_out_dist_full_n = out_dist_2__full_n;
  assign out_dist_2__write = krnl_partialKnn_wrapper_2_0_out_dist_write;
  assign out_id_2__din = krnl_partialKnn_wrapper_2_0_out_id_din;
  assign krnl_partialKnn_wrapper_2_0_out_id_full_n = out_id_2__full_n;
  assign out_id_2__write = krnl_partialKnn_wrapper_2_0_out_id_write;
  assign krnl_partialKnn_wrapper_2_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_2_0___in_2__q0;
  assign in_2_read_addr__din = krnl_partialKnn_wrapper_2_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_2_0_searchSpace_0_read_addr_s_full_n = in_2_read_addr__full_n;
  assign in_2_read_addr__write = krnl_partialKnn_wrapper_2_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_2_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_2_read_data__dout };
  assign krnl_partialKnn_wrapper_2_0_searchSpace_0_read_data_peek_empty_n = in_2_read_data__empty_n;
  assign krnl_partialKnn_wrapper_2_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_2_read_data__dout };
  assign krnl_partialKnn_wrapper_2_0_searchSpace_0_read_data_s_empty_n = in_2_read_data__empty_n;
  assign in_2_read_data__read = krnl_partialKnn_wrapper_2_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_2_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_2_0___in_2__q0;
  assign in_2_write_addr__din = krnl_partialKnn_wrapper_2_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_2_0_searchSpace_0_write_addr_s_full_n = in_2_write_addr__full_n;
  assign in_2_write_addr__write = krnl_partialKnn_wrapper_2_0_searchSpace_0_write_addr_s_write;
  assign in_2_write_data__din = krnl_partialKnn_wrapper_2_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_2_0_searchSpace_0_write_data_full_n = in_2_write_data__full_n;
  assign in_2_write_data__write = krnl_partialKnn_wrapper_2_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_2_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_2_write_resp__dout };
  assign krnl_partialKnn_wrapper_2_0_searchSpace_write_resp_peek_empty_n = in_2_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_2_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_2_write_resp__dout };
  assign krnl_partialKnn_wrapper_2_0_searchSpace_0_write_resp_s_empty_n = in_2_write_resp__empty_n;
  assign in_2_write_resp__read = krnl_partialKnn_wrapper_2_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_2_0_start_id_0 = 64'd16384;
  assign krnl_partialKnn_wrapper_20_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_20_0__ap_done = krnl_partialKnn_wrapper_20_0_ap_done;
  assign krnl_partialKnn_wrapper_20_0__ap_idle = krnl_partialKnn_wrapper_20_0_ap_idle;
  assign krnl_partialKnn_wrapper_20_0__ap_ready = krnl_partialKnn_wrapper_20_0_ap_ready;
  assign krnl_partialKnn_wrapper_20_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_20_0_ap_start = krnl_partialKnn_wrapper_20_0__ap_start;
  assign out_dist_20__din = krnl_partialKnn_wrapper_20_0_out_dist_din;
  assign krnl_partialKnn_wrapper_20_0_out_dist_full_n = out_dist_20__full_n;
  assign out_dist_20__write = krnl_partialKnn_wrapper_20_0_out_dist_write;
  assign out_id_20__din = krnl_partialKnn_wrapper_20_0_out_id_din;
  assign krnl_partialKnn_wrapper_20_0_out_id_full_n = out_id_20__full_n;
  assign out_id_20__write = krnl_partialKnn_wrapper_20_0_out_id_write;
  assign krnl_partialKnn_wrapper_20_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_20_0___in_20__q0;
  assign in_20_read_addr__din = krnl_partialKnn_wrapper_20_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_20_0_searchSpace_0_read_addr_s_full_n = in_20_read_addr__full_n;
  assign in_20_read_addr__write = krnl_partialKnn_wrapper_20_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_20_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_20_read_data__dout };
  assign krnl_partialKnn_wrapper_20_0_searchSpace_read_data_peek_empty_n = in_20_read_data__empty_n;
  assign krnl_partialKnn_wrapper_20_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_20_read_data__dout };
  assign krnl_partialKnn_wrapper_20_0_searchSpace_0_read_data_s_empty_n = in_20_read_data__empty_n;
  assign in_20_read_data__read = krnl_partialKnn_wrapper_20_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_20_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_20_0___in_20__q0;
  assign in_20_write_addr__din = krnl_partialKnn_wrapper_20_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_20_0_searchSpace_0_write_addr_s_full_n = in_20_write_addr__full_n;
  assign in_20_write_addr__write = krnl_partialKnn_wrapper_20_0_searchSpace_0_write_addr_s_write;
  assign in_20_write_data__din = krnl_partialKnn_wrapper_20_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_20_0_searchSpace_0_write_data_full_n = in_20_write_data__full_n;
  assign in_20_write_data__write = krnl_partialKnn_wrapper_20_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_20_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_20_write_resp__dout };
  assign krnl_partialKnn_wrapper_20_0_searchSpace_write_resp_peek_empty_n = in_20_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_20_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_20_write_resp__dout };
  assign krnl_partialKnn_wrapper_20_0_searchSpace_0_write_resp_s_empty_n = in_20_write_resp__empty_n;
  assign in_20_write_resp__read = krnl_partialKnn_wrapper_20_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_20_0_start_id_0 = 64'd163840;
  assign krnl_partialKnn_wrapper_21_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_21_0__ap_done = krnl_partialKnn_wrapper_21_0_ap_done;
  assign krnl_partialKnn_wrapper_21_0__ap_idle = krnl_partialKnn_wrapper_21_0_ap_idle;
  assign krnl_partialKnn_wrapper_21_0__ap_ready = krnl_partialKnn_wrapper_21_0_ap_ready;
  assign krnl_partialKnn_wrapper_21_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_21_0_ap_start = krnl_partialKnn_wrapper_21_0__ap_start;
  assign out_dist_21__din = krnl_partialKnn_wrapper_21_0_out_dist_din;
  assign krnl_partialKnn_wrapper_21_0_out_dist_full_n = out_dist_21__full_n;
  assign out_dist_21__write = krnl_partialKnn_wrapper_21_0_out_dist_write;
  assign out_id_21__din = krnl_partialKnn_wrapper_21_0_out_id_din;
  assign krnl_partialKnn_wrapper_21_0_out_id_full_n = out_id_21__full_n;
  assign out_id_21__write = krnl_partialKnn_wrapper_21_0_out_id_write;
  assign krnl_partialKnn_wrapper_21_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_21_0___in_21__q0;
  assign in_21_read_addr__din = krnl_partialKnn_wrapper_21_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_21_0_searchSpace_0_read_addr_s_full_n = in_21_read_addr__full_n;
  assign in_21_read_addr__write = krnl_partialKnn_wrapper_21_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_21_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_21_read_data__dout };
  assign krnl_partialKnn_wrapper_21_0_searchSpace_read_data_peek_empty_n = in_21_read_data__empty_n;
  assign krnl_partialKnn_wrapper_21_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_21_read_data__dout };
  assign krnl_partialKnn_wrapper_21_0_searchSpace_0_read_data_s_empty_n = in_21_read_data__empty_n;
  assign in_21_read_data__read = krnl_partialKnn_wrapper_21_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_21_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_21_0___in_21__q0;
  assign in_21_write_addr__din = krnl_partialKnn_wrapper_21_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_21_0_searchSpace_0_write_addr_s_full_n = in_21_write_addr__full_n;
  assign in_21_write_addr__write = krnl_partialKnn_wrapper_21_0_searchSpace_0_write_addr_s_write;
  assign in_21_write_data__din = krnl_partialKnn_wrapper_21_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_21_0_searchSpace_0_write_data_full_n = in_21_write_data__full_n;
  assign in_21_write_data__write = krnl_partialKnn_wrapper_21_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_21_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_21_write_resp__dout };
  assign krnl_partialKnn_wrapper_21_0_searchSpace_write_resp_peek_empty_n = in_21_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_21_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_21_write_resp__dout };
  assign krnl_partialKnn_wrapper_21_0_searchSpace_0_write_resp_s_empty_n = in_21_write_resp__empty_n;
  assign in_21_write_resp__read = krnl_partialKnn_wrapper_21_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_21_0_start_id_0 = 64'd172032;
  assign krnl_partialKnn_wrapper_22_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_22_0__ap_done = krnl_partialKnn_wrapper_22_0_ap_done;
  assign krnl_partialKnn_wrapper_22_0__ap_idle = krnl_partialKnn_wrapper_22_0_ap_idle;
  assign krnl_partialKnn_wrapper_22_0__ap_ready = krnl_partialKnn_wrapper_22_0_ap_ready;
  assign krnl_partialKnn_wrapper_22_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_22_0_ap_start = krnl_partialKnn_wrapper_22_0__ap_start;
  assign out_dist_22__din = krnl_partialKnn_wrapper_22_0_out_dist_din;
  assign krnl_partialKnn_wrapper_22_0_out_dist_full_n = out_dist_22__full_n;
  assign out_dist_22__write = krnl_partialKnn_wrapper_22_0_out_dist_write;
  assign out_id_22__din = krnl_partialKnn_wrapper_22_0_out_id_din;
  assign krnl_partialKnn_wrapper_22_0_out_id_full_n = out_id_22__full_n;
  assign out_id_22__write = krnl_partialKnn_wrapper_22_0_out_id_write;
  assign krnl_partialKnn_wrapper_22_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_22_0___in_22__q0;
  assign in_22_read_addr__din = krnl_partialKnn_wrapper_22_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_22_0_searchSpace_0_read_addr_s_full_n = in_22_read_addr__full_n;
  assign in_22_read_addr__write = krnl_partialKnn_wrapper_22_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_22_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_22_read_data__dout };
  assign krnl_partialKnn_wrapper_22_0_searchSpace_read_data_peek_empty_n = in_22_read_data__empty_n;
  assign krnl_partialKnn_wrapper_22_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_22_read_data__dout };
  assign krnl_partialKnn_wrapper_22_0_searchSpace_0_read_data_s_empty_n = in_22_read_data__empty_n;
  assign in_22_read_data__read = krnl_partialKnn_wrapper_22_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_22_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_22_0___in_22__q0;
  assign in_22_write_addr__din = krnl_partialKnn_wrapper_22_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_22_0_searchSpace_0_write_addr_s_full_n = in_22_write_addr__full_n;
  assign in_22_write_addr__write = krnl_partialKnn_wrapper_22_0_searchSpace_0_write_addr_s_write;
  assign in_22_write_data__din = krnl_partialKnn_wrapper_22_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_22_0_searchSpace_0_write_data_full_n = in_22_write_data__full_n;
  assign in_22_write_data__write = krnl_partialKnn_wrapper_22_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_22_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_22_write_resp__dout };
  assign krnl_partialKnn_wrapper_22_0_searchSpace_write_resp_peek_empty_n = in_22_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_22_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_22_write_resp__dout };
  assign krnl_partialKnn_wrapper_22_0_searchSpace_0_write_resp_s_empty_n = in_22_write_resp__empty_n;
  assign in_22_write_resp__read = krnl_partialKnn_wrapper_22_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_22_0_start_id_0 = 64'd180224;
  assign krnl_partialKnn_wrapper_23_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_23_0__ap_done = krnl_partialKnn_wrapper_23_0_ap_done;
  assign krnl_partialKnn_wrapper_23_0__ap_idle = krnl_partialKnn_wrapper_23_0_ap_idle;
  assign krnl_partialKnn_wrapper_23_0__ap_ready = krnl_partialKnn_wrapper_23_0_ap_ready;
  assign krnl_partialKnn_wrapper_23_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_23_0_ap_start = krnl_partialKnn_wrapper_23_0__ap_start;
  assign out_dist_23__din = krnl_partialKnn_wrapper_23_0_out_dist_din;
  assign krnl_partialKnn_wrapper_23_0_out_dist_full_n = out_dist_23__full_n;
  assign out_dist_23__write = krnl_partialKnn_wrapper_23_0_out_dist_write;
  assign out_id_23__din = krnl_partialKnn_wrapper_23_0_out_id_din;
  assign krnl_partialKnn_wrapper_23_0_out_id_full_n = out_id_23__full_n;
  assign out_id_23__write = krnl_partialKnn_wrapper_23_0_out_id_write;
  assign krnl_partialKnn_wrapper_23_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_23_0___in_23__q0;
  assign in_23_read_addr__din = krnl_partialKnn_wrapper_23_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_23_0_searchSpace_0_read_addr_s_full_n = in_23_read_addr__full_n;
  assign in_23_read_addr__write = krnl_partialKnn_wrapper_23_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_23_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_23_read_data__dout };
  assign krnl_partialKnn_wrapper_23_0_searchSpace_read_data_peek_empty_n = in_23_read_data__empty_n;
  assign krnl_partialKnn_wrapper_23_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_23_read_data__dout };
  assign krnl_partialKnn_wrapper_23_0_searchSpace_0_read_data_s_empty_n = in_23_read_data__empty_n;
  assign in_23_read_data__read = krnl_partialKnn_wrapper_23_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_23_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_23_0___in_23__q0;
  assign in_23_write_addr__din = krnl_partialKnn_wrapper_23_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_23_0_searchSpace_0_write_addr_s_full_n = in_23_write_addr__full_n;
  assign in_23_write_addr__write = krnl_partialKnn_wrapper_23_0_searchSpace_0_write_addr_s_write;
  assign in_23_write_data__din = krnl_partialKnn_wrapper_23_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_23_0_searchSpace_0_write_data_full_n = in_23_write_data__full_n;
  assign in_23_write_data__write = krnl_partialKnn_wrapper_23_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_23_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_23_write_resp__dout };
  assign krnl_partialKnn_wrapper_23_0_searchSpace_write_resp_peek_empty_n = in_23_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_23_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_23_write_resp__dout };
  assign krnl_partialKnn_wrapper_23_0_searchSpace_0_write_resp_s_empty_n = in_23_write_resp__empty_n;
  assign in_23_write_resp__read = krnl_partialKnn_wrapper_23_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_23_0_start_id_0 = 64'd188416;
  assign krnl_partialKnn_wrapper_24_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_24_0__ap_done = krnl_partialKnn_wrapper_24_0_ap_done;
  assign krnl_partialKnn_wrapper_24_0__ap_idle = krnl_partialKnn_wrapper_24_0_ap_idle;
  assign krnl_partialKnn_wrapper_24_0__ap_ready = krnl_partialKnn_wrapper_24_0_ap_ready;
  assign krnl_partialKnn_wrapper_24_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_24_0_ap_start = krnl_partialKnn_wrapper_24_0__ap_start;
  assign out_dist_24__din = krnl_partialKnn_wrapper_24_0_out_dist_din;
  assign krnl_partialKnn_wrapper_24_0_out_dist_full_n = out_dist_24__full_n;
  assign out_dist_24__write = krnl_partialKnn_wrapper_24_0_out_dist_write;
  assign out_id_24__din = krnl_partialKnn_wrapper_24_0_out_id_din;
  assign krnl_partialKnn_wrapper_24_0_out_id_full_n = out_id_24__full_n;
  assign out_id_24__write = krnl_partialKnn_wrapper_24_0_out_id_write;
  assign krnl_partialKnn_wrapper_24_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_24_0___in_24__q0;
  assign in_24_read_addr__din = krnl_partialKnn_wrapper_24_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_24_0_searchSpace_0_read_addr_s_full_n = in_24_read_addr__full_n;
  assign in_24_read_addr__write = krnl_partialKnn_wrapper_24_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_24_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_24_read_data__dout };
  assign krnl_partialKnn_wrapper_24_0_searchSpace_read_data_peek_empty_n = in_24_read_data__empty_n;
  assign krnl_partialKnn_wrapper_24_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_24_read_data__dout };
  assign krnl_partialKnn_wrapper_24_0_searchSpace_0_read_data_s_empty_n = in_24_read_data__empty_n;
  assign in_24_read_data__read = krnl_partialKnn_wrapper_24_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_24_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_24_0___in_24__q0;
  assign in_24_write_addr__din = krnl_partialKnn_wrapper_24_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_24_0_searchSpace_0_write_addr_s_full_n = in_24_write_addr__full_n;
  assign in_24_write_addr__write = krnl_partialKnn_wrapper_24_0_searchSpace_0_write_addr_s_write;
  assign in_24_write_data__din = krnl_partialKnn_wrapper_24_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_24_0_searchSpace_0_write_data_full_n = in_24_write_data__full_n;
  assign in_24_write_data__write = krnl_partialKnn_wrapper_24_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_24_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_24_write_resp__dout };
  assign krnl_partialKnn_wrapper_24_0_searchSpace_write_resp_peek_empty_n = in_24_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_24_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_24_write_resp__dout };
  assign krnl_partialKnn_wrapper_24_0_searchSpace_0_write_resp_s_empty_n = in_24_write_resp__empty_n;
  assign in_24_write_resp__read = krnl_partialKnn_wrapper_24_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_24_0_start_id_0 = 64'd196608;
  assign krnl_partialKnn_wrapper_25_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_25_0__ap_done = krnl_partialKnn_wrapper_25_0_ap_done;
  assign krnl_partialKnn_wrapper_25_0__ap_idle = krnl_partialKnn_wrapper_25_0_ap_idle;
  assign krnl_partialKnn_wrapper_25_0__ap_ready = krnl_partialKnn_wrapper_25_0_ap_ready;
  assign krnl_partialKnn_wrapper_25_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_25_0_ap_start = krnl_partialKnn_wrapper_25_0__ap_start;
  assign out_dist_25__din = krnl_partialKnn_wrapper_25_0_out_dist_din;
  assign krnl_partialKnn_wrapper_25_0_out_dist_full_n = out_dist_25__full_n;
  assign out_dist_25__write = krnl_partialKnn_wrapper_25_0_out_dist_write;
  assign out_id_25__din = krnl_partialKnn_wrapper_25_0_out_id_din;
  assign krnl_partialKnn_wrapper_25_0_out_id_full_n = out_id_25__full_n;
  assign out_id_25__write = krnl_partialKnn_wrapper_25_0_out_id_write;
  assign krnl_partialKnn_wrapper_25_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_25_0___in_25__q0;
  assign in_25_read_addr__din = krnl_partialKnn_wrapper_25_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_25_0_searchSpace_0_read_addr_s_full_n = in_25_read_addr__full_n;
  assign in_25_read_addr__write = krnl_partialKnn_wrapper_25_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_25_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_25_read_data__dout };
  assign krnl_partialKnn_wrapper_25_0_searchSpace_read_data_peek_empty_n = in_25_read_data__empty_n;
  assign krnl_partialKnn_wrapper_25_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_25_read_data__dout };
  assign krnl_partialKnn_wrapper_25_0_searchSpace_0_read_data_s_empty_n = in_25_read_data__empty_n;
  assign in_25_read_data__read = krnl_partialKnn_wrapper_25_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_25_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_25_0___in_25__q0;
  assign in_25_write_addr__din = krnl_partialKnn_wrapper_25_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_25_0_searchSpace_0_write_addr_s_full_n = in_25_write_addr__full_n;
  assign in_25_write_addr__write = krnl_partialKnn_wrapper_25_0_searchSpace_0_write_addr_s_write;
  assign in_25_write_data__din = krnl_partialKnn_wrapper_25_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_25_0_searchSpace_0_write_data_full_n = in_25_write_data__full_n;
  assign in_25_write_data__write = krnl_partialKnn_wrapper_25_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_25_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_25_write_resp__dout };
  assign krnl_partialKnn_wrapper_25_0_searchSpace_write_resp_peek_empty_n = in_25_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_25_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_25_write_resp__dout };
  assign krnl_partialKnn_wrapper_25_0_searchSpace_0_write_resp_s_empty_n = in_25_write_resp__empty_n;
  assign in_25_write_resp__read = krnl_partialKnn_wrapper_25_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_25_0_start_id_0 = 64'd204800;
  assign krnl_partialKnn_wrapper_26_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_26_0__ap_done = krnl_partialKnn_wrapper_26_0_ap_done;
  assign krnl_partialKnn_wrapper_26_0__ap_idle = krnl_partialKnn_wrapper_26_0_ap_idle;
  assign krnl_partialKnn_wrapper_26_0__ap_ready = krnl_partialKnn_wrapper_26_0_ap_ready;
  assign krnl_partialKnn_wrapper_26_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_26_0_ap_start = krnl_partialKnn_wrapper_26_0__ap_start;
  assign out_dist_26__din = krnl_partialKnn_wrapper_26_0_out_dist_din;
  assign krnl_partialKnn_wrapper_26_0_out_dist_full_n = out_dist_26__full_n;
  assign out_dist_26__write = krnl_partialKnn_wrapper_26_0_out_dist_write;
  assign out_id_26__din = krnl_partialKnn_wrapper_26_0_out_id_din;
  assign krnl_partialKnn_wrapper_26_0_out_id_full_n = out_id_26__full_n;
  assign out_id_26__write = krnl_partialKnn_wrapper_26_0_out_id_write;
  assign krnl_partialKnn_wrapper_26_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_26_0___in_26__q0;
  assign in_26_read_addr__din = krnl_partialKnn_wrapper_26_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_26_0_searchSpace_0_read_addr_s_full_n = in_26_read_addr__full_n;
  assign in_26_read_addr__write = krnl_partialKnn_wrapper_26_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_26_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_26_read_data__dout };
  assign krnl_partialKnn_wrapper_26_0_searchSpace_read_data_peek_empty_n = in_26_read_data__empty_n;
  assign krnl_partialKnn_wrapper_26_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_26_read_data__dout };
  assign krnl_partialKnn_wrapper_26_0_searchSpace_0_read_data_s_empty_n = in_26_read_data__empty_n;
  assign in_26_read_data__read = krnl_partialKnn_wrapper_26_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_26_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_26_0___in_26__q0;
  assign in_26_write_addr__din = krnl_partialKnn_wrapper_26_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_26_0_searchSpace_0_write_addr_s_full_n = in_26_write_addr__full_n;
  assign in_26_write_addr__write = krnl_partialKnn_wrapper_26_0_searchSpace_0_write_addr_s_write;
  assign in_26_write_data__din = krnl_partialKnn_wrapper_26_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_26_0_searchSpace_0_write_data_full_n = in_26_write_data__full_n;
  assign in_26_write_data__write = krnl_partialKnn_wrapper_26_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_26_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_26_write_resp__dout };
  assign krnl_partialKnn_wrapper_26_0_searchSpace_write_resp_peek_empty_n = in_26_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_26_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_26_write_resp__dout };
  assign krnl_partialKnn_wrapper_26_0_searchSpace_0_write_resp_s_empty_n = in_26_write_resp__empty_n;
  assign in_26_write_resp__read = krnl_partialKnn_wrapper_26_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_26_0_start_id_0 = 64'd212992;
  assign krnl_partialKnn_wrapper_3_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_3_0__ap_done = krnl_partialKnn_wrapper_3_0_ap_done;
  assign krnl_partialKnn_wrapper_3_0__ap_idle = krnl_partialKnn_wrapper_3_0_ap_idle;
  assign krnl_partialKnn_wrapper_3_0__ap_ready = krnl_partialKnn_wrapper_3_0_ap_ready;
  assign krnl_partialKnn_wrapper_3_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_3_0_ap_start = krnl_partialKnn_wrapper_3_0__ap_start;
  assign out_dist_3__din = krnl_partialKnn_wrapper_3_0_out_dist_din;
  assign krnl_partialKnn_wrapper_3_0_out_dist_full_n = out_dist_3__full_n;
  assign out_dist_3__write = krnl_partialKnn_wrapper_3_0_out_dist_write;
  assign out_id_3__din = krnl_partialKnn_wrapper_3_0_out_id_din;
  assign krnl_partialKnn_wrapper_3_0_out_id_full_n = out_id_3__full_n;
  assign out_id_3__write = krnl_partialKnn_wrapper_3_0_out_id_write;
  assign krnl_partialKnn_wrapper_3_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_3_0___in_3__q0;
  assign in_3_read_addr__din = krnl_partialKnn_wrapper_3_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_3_0_searchSpace_0_read_addr_s_full_n = in_3_read_addr__full_n;
  assign in_3_read_addr__write = krnl_partialKnn_wrapper_3_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_3_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_3_read_data__dout };
  assign krnl_partialKnn_wrapper_3_0_searchSpace_0_read_data_peek_empty_n = in_3_read_data__empty_n;
  assign krnl_partialKnn_wrapper_3_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_3_read_data__dout };
  assign krnl_partialKnn_wrapper_3_0_searchSpace_0_read_data_s_empty_n = in_3_read_data__empty_n;
  assign in_3_read_data__read = krnl_partialKnn_wrapper_3_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_3_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_3_0___in_3__q0;
  assign in_3_write_addr__din = krnl_partialKnn_wrapper_3_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_3_0_searchSpace_0_write_addr_s_full_n = in_3_write_addr__full_n;
  assign in_3_write_addr__write = krnl_partialKnn_wrapper_3_0_searchSpace_0_write_addr_s_write;
  assign in_3_write_data__din = krnl_partialKnn_wrapper_3_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_3_0_searchSpace_0_write_data_full_n = in_3_write_data__full_n;
  assign in_3_write_data__write = krnl_partialKnn_wrapper_3_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_3_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_3_write_resp__dout };
  assign krnl_partialKnn_wrapper_3_0_searchSpace_write_resp_peek_empty_n = in_3_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_3_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_3_write_resp__dout };
  assign krnl_partialKnn_wrapper_3_0_searchSpace_0_write_resp_s_empty_n = in_3_write_resp__empty_n;
  assign in_3_write_resp__read = krnl_partialKnn_wrapper_3_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_3_0_start_id_0 = 64'd24576;
  assign krnl_partialKnn_wrapper_4_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_4_0__ap_done = krnl_partialKnn_wrapper_4_0_ap_done;
  assign krnl_partialKnn_wrapper_4_0__ap_idle = krnl_partialKnn_wrapper_4_0_ap_idle;
  assign krnl_partialKnn_wrapper_4_0__ap_ready = krnl_partialKnn_wrapper_4_0_ap_ready;
  assign krnl_partialKnn_wrapper_4_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_4_0_ap_start = krnl_partialKnn_wrapper_4_0__ap_start;
  assign out_dist_4__din = krnl_partialKnn_wrapper_4_0_out_dist_din;
  assign krnl_partialKnn_wrapper_4_0_out_dist_full_n = out_dist_4__full_n;
  assign out_dist_4__write = krnl_partialKnn_wrapper_4_0_out_dist_write;
  assign out_id_4__din = krnl_partialKnn_wrapper_4_0_out_id_din;
  assign krnl_partialKnn_wrapper_4_0_out_id_full_n = out_id_4__full_n;
  assign out_id_4__write = krnl_partialKnn_wrapper_4_0_out_id_write;
  assign krnl_partialKnn_wrapper_4_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_4_0___in_4__q0;
  assign in_4_read_addr__din = krnl_partialKnn_wrapper_4_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_4_0_searchSpace_0_read_addr_s_full_n = in_4_read_addr__full_n;
  assign in_4_read_addr__write = krnl_partialKnn_wrapper_4_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_4_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_4_read_data__dout };
  assign krnl_partialKnn_wrapper_4_0_searchSpace_0_read_data_peek_empty_n = in_4_read_data__empty_n;
  assign krnl_partialKnn_wrapper_4_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_4_read_data__dout };
  assign krnl_partialKnn_wrapper_4_0_searchSpace_0_read_data_s_empty_n = in_4_read_data__empty_n;
  assign in_4_read_data__read = krnl_partialKnn_wrapper_4_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_4_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_4_0___in_4__q0;
  assign in_4_write_addr__din = krnl_partialKnn_wrapper_4_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_4_0_searchSpace_0_write_addr_s_full_n = in_4_write_addr__full_n;
  assign in_4_write_addr__write = krnl_partialKnn_wrapper_4_0_searchSpace_0_write_addr_s_write;
  assign in_4_write_data__din = krnl_partialKnn_wrapper_4_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_4_0_searchSpace_0_write_data_full_n = in_4_write_data__full_n;
  assign in_4_write_data__write = krnl_partialKnn_wrapper_4_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_4_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_4_write_resp__dout };
  assign krnl_partialKnn_wrapper_4_0_searchSpace_write_resp_peek_empty_n = in_4_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_4_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_4_write_resp__dout };
  assign krnl_partialKnn_wrapper_4_0_searchSpace_0_write_resp_s_empty_n = in_4_write_resp__empty_n;
  assign in_4_write_resp__read = krnl_partialKnn_wrapper_4_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_4_0_start_id_0 = 64'd32768;
  assign krnl_partialKnn_wrapper_5_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_5_0__ap_done = krnl_partialKnn_wrapper_5_0_ap_done;
  assign krnl_partialKnn_wrapper_5_0__ap_idle = krnl_partialKnn_wrapper_5_0_ap_idle;
  assign krnl_partialKnn_wrapper_5_0__ap_ready = krnl_partialKnn_wrapper_5_0_ap_ready;
  assign krnl_partialKnn_wrapper_5_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_5_0_ap_start = krnl_partialKnn_wrapper_5_0__ap_start;
  assign out_dist_5__din = krnl_partialKnn_wrapper_5_0_out_dist_din;
  assign krnl_partialKnn_wrapper_5_0_out_dist_full_n = out_dist_5__full_n;
  assign out_dist_5__write = krnl_partialKnn_wrapper_5_0_out_dist_write;
  assign out_id_5__din = krnl_partialKnn_wrapper_5_0_out_id_din;
  assign krnl_partialKnn_wrapper_5_0_out_id_full_n = out_id_5__full_n;
  assign out_id_5__write = krnl_partialKnn_wrapper_5_0_out_id_write;
  assign krnl_partialKnn_wrapper_5_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_5_0___in_5__q0;
  assign in_5_read_addr__din = krnl_partialKnn_wrapper_5_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_5_0_searchSpace_0_read_addr_s_full_n = in_5_read_addr__full_n;
  assign in_5_read_addr__write = krnl_partialKnn_wrapper_5_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_5_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_5_read_data__dout };
  assign krnl_partialKnn_wrapper_5_0_searchSpace_0_read_data_peek_empty_n = in_5_read_data__empty_n;
  assign krnl_partialKnn_wrapper_5_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_5_read_data__dout };
  assign krnl_partialKnn_wrapper_5_0_searchSpace_0_read_data_s_empty_n = in_5_read_data__empty_n;
  assign in_5_read_data__read = krnl_partialKnn_wrapper_5_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_5_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_5_0___in_5__q0;
  assign in_5_write_addr__din = krnl_partialKnn_wrapper_5_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_5_0_searchSpace_0_write_addr_s_full_n = in_5_write_addr__full_n;
  assign in_5_write_addr__write = krnl_partialKnn_wrapper_5_0_searchSpace_0_write_addr_s_write;
  assign in_5_write_data__din = krnl_partialKnn_wrapper_5_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_5_0_searchSpace_0_write_data_full_n = in_5_write_data__full_n;
  assign in_5_write_data__write = krnl_partialKnn_wrapper_5_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_5_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_5_write_resp__dout };
  assign krnl_partialKnn_wrapper_5_0_searchSpace_write_resp_peek_empty_n = in_5_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_5_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_5_write_resp__dout };
  assign krnl_partialKnn_wrapper_5_0_searchSpace_0_write_resp_s_empty_n = in_5_write_resp__empty_n;
  assign in_5_write_resp__read = krnl_partialKnn_wrapper_5_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_5_0_start_id_0 = 64'd40960;
  assign krnl_partialKnn_wrapper_6_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_6_0__ap_done = krnl_partialKnn_wrapper_6_0_ap_done;
  assign krnl_partialKnn_wrapper_6_0__ap_idle = krnl_partialKnn_wrapper_6_0_ap_idle;
  assign krnl_partialKnn_wrapper_6_0__ap_ready = krnl_partialKnn_wrapper_6_0_ap_ready;
  assign krnl_partialKnn_wrapper_6_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_6_0_ap_start = krnl_partialKnn_wrapper_6_0__ap_start;
  assign out_dist_6__din = krnl_partialKnn_wrapper_6_0_out_dist_din;
  assign krnl_partialKnn_wrapper_6_0_out_dist_full_n = out_dist_6__full_n;
  assign out_dist_6__write = krnl_partialKnn_wrapper_6_0_out_dist_write;
  assign out_id_6__din = krnl_partialKnn_wrapper_6_0_out_id_din;
  assign krnl_partialKnn_wrapper_6_0_out_id_full_n = out_id_6__full_n;
  assign out_id_6__write = krnl_partialKnn_wrapper_6_0_out_id_write;
  assign krnl_partialKnn_wrapper_6_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_6_0___in_6__q0;
  assign in_6_read_addr__din = krnl_partialKnn_wrapper_6_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_6_0_searchSpace_0_read_addr_s_full_n = in_6_read_addr__full_n;
  assign in_6_read_addr__write = krnl_partialKnn_wrapper_6_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_6_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_6_read_data__dout };
  assign krnl_partialKnn_wrapper_6_0_searchSpace_0_read_data_peek_empty_n = in_6_read_data__empty_n;
  assign krnl_partialKnn_wrapper_6_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_6_read_data__dout };
  assign krnl_partialKnn_wrapper_6_0_searchSpace_0_read_data_s_empty_n = in_6_read_data__empty_n;
  assign in_6_read_data__read = krnl_partialKnn_wrapper_6_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_6_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_6_0___in_6__q0;
  assign in_6_write_addr__din = krnl_partialKnn_wrapper_6_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_6_0_searchSpace_0_write_addr_s_full_n = in_6_write_addr__full_n;
  assign in_6_write_addr__write = krnl_partialKnn_wrapper_6_0_searchSpace_0_write_addr_s_write;
  assign in_6_write_data__din = krnl_partialKnn_wrapper_6_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_6_0_searchSpace_0_write_data_full_n = in_6_write_data__full_n;
  assign in_6_write_data__write = krnl_partialKnn_wrapper_6_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_6_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_6_write_resp__dout };
  assign krnl_partialKnn_wrapper_6_0_searchSpace_write_resp_peek_empty_n = in_6_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_6_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_6_write_resp__dout };
  assign krnl_partialKnn_wrapper_6_0_searchSpace_0_write_resp_s_empty_n = in_6_write_resp__empty_n;
  assign in_6_write_resp__read = krnl_partialKnn_wrapper_6_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_6_0_start_id_0 = 64'd49152;
  assign krnl_partialKnn_wrapper_7_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_7_0__ap_done = krnl_partialKnn_wrapper_7_0_ap_done;
  assign krnl_partialKnn_wrapper_7_0__ap_idle = krnl_partialKnn_wrapper_7_0_ap_idle;
  assign krnl_partialKnn_wrapper_7_0__ap_ready = krnl_partialKnn_wrapper_7_0_ap_ready;
  assign krnl_partialKnn_wrapper_7_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_7_0_ap_start = krnl_partialKnn_wrapper_7_0__ap_start;
  assign out_dist_7__din = krnl_partialKnn_wrapper_7_0_out_dist_din;
  assign krnl_partialKnn_wrapper_7_0_out_dist_full_n = out_dist_7__full_n;
  assign out_dist_7__write = krnl_partialKnn_wrapper_7_0_out_dist_write;
  assign out_id_7__din = krnl_partialKnn_wrapper_7_0_out_id_din;
  assign krnl_partialKnn_wrapper_7_0_out_id_full_n = out_id_7__full_n;
  assign out_id_7__write = krnl_partialKnn_wrapper_7_0_out_id_write;
  assign krnl_partialKnn_wrapper_7_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_7_0___in_7__q0;
  assign in_7_read_addr__din = krnl_partialKnn_wrapper_7_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_7_0_searchSpace_0_read_addr_s_full_n = in_7_read_addr__full_n;
  assign in_7_read_addr__write = krnl_partialKnn_wrapper_7_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_7_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_7_read_data__dout };
  assign krnl_partialKnn_wrapper_7_0_searchSpace_0_read_data_peek_empty_n = in_7_read_data__empty_n;
  assign krnl_partialKnn_wrapper_7_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_7_read_data__dout };
  assign krnl_partialKnn_wrapper_7_0_searchSpace_0_read_data_s_empty_n = in_7_read_data__empty_n;
  assign in_7_read_data__read = krnl_partialKnn_wrapper_7_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_7_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_7_0___in_7__q0;
  assign in_7_write_addr__din = krnl_partialKnn_wrapper_7_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_7_0_searchSpace_0_write_addr_s_full_n = in_7_write_addr__full_n;
  assign in_7_write_addr__write = krnl_partialKnn_wrapper_7_0_searchSpace_0_write_addr_s_write;
  assign in_7_write_data__din = krnl_partialKnn_wrapper_7_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_7_0_searchSpace_0_write_data_full_n = in_7_write_data__full_n;
  assign in_7_write_data__write = krnl_partialKnn_wrapper_7_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_7_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_7_write_resp__dout };
  assign krnl_partialKnn_wrapper_7_0_searchSpace_write_resp_peek_empty_n = in_7_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_7_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_7_write_resp__dout };
  assign krnl_partialKnn_wrapper_7_0_searchSpace_0_write_resp_s_empty_n = in_7_write_resp__empty_n;
  assign in_7_write_resp__read = krnl_partialKnn_wrapper_7_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_7_0_start_id_0 = 64'd57344;
  assign krnl_partialKnn_wrapper_8_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_8_0__ap_done = krnl_partialKnn_wrapper_8_0_ap_done;
  assign krnl_partialKnn_wrapper_8_0__ap_idle = krnl_partialKnn_wrapper_8_0_ap_idle;
  assign krnl_partialKnn_wrapper_8_0__ap_ready = krnl_partialKnn_wrapper_8_0_ap_ready;
  assign krnl_partialKnn_wrapper_8_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_8_0_ap_start = krnl_partialKnn_wrapper_8_0__ap_start;
  assign out_dist_8__din = krnl_partialKnn_wrapper_8_0_out_dist_din;
  assign krnl_partialKnn_wrapper_8_0_out_dist_full_n = out_dist_8__full_n;
  assign out_dist_8__write = krnl_partialKnn_wrapper_8_0_out_dist_write;
  assign out_id_8__din = krnl_partialKnn_wrapper_8_0_out_id_din;
  assign krnl_partialKnn_wrapper_8_0_out_id_full_n = out_id_8__full_n;
  assign out_id_8__write = krnl_partialKnn_wrapper_8_0_out_id_write;
  assign krnl_partialKnn_wrapper_8_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_8_0___in_8__q0;
  assign in_8_read_addr__din = krnl_partialKnn_wrapper_8_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_8_0_searchSpace_0_read_addr_s_full_n = in_8_read_addr__full_n;
  assign in_8_read_addr__write = krnl_partialKnn_wrapper_8_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_8_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_8_read_data__dout };
  assign krnl_partialKnn_wrapper_8_0_searchSpace_0_read_data_peek_empty_n = in_8_read_data__empty_n;
  assign krnl_partialKnn_wrapper_8_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_8_read_data__dout };
  assign krnl_partialKnn_wrapper_8_0_searchSpace_0_read_data_s_empty_n = in_8_read_data__empty_n;
  assign in_8_read_data__read = krnl_partialKnn_wrapper_8_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_8_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_8_0___in_8__q0;
  assign in_8_write_addr__din = krnl_partialKnn_wrapper_8_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_8_0_searchSpace_0_write_addr_s_full_n = in_8_write_addr__full_n;
  assign in_8_write_addr__write = krnl_partialKnn_wrapper_8_0_searchSpace_0_write_addr_s_write;
  assign in_8_write_data__din = krnl_partialKnn_wrapper_8_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_8_0_searchSpace_0_write_data_full_n = in_8_write_data__full_n;
  assign in_8_write_data__write = krnl_partialKnn_wrapper_8_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_8_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_8_write_resp__dout };
  assign krnl_partialKnn_wrapper_8_0_searchSpace_write_resp_peek_empty_n = in_8_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_8_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_8_write_resp__dout };
  assign krnl_partialKnn_wrapper_8_0_searchSpace_0_write_resp_s_empty_n = in_8_write_resp__empty_n;
  assign in_8_write_resp__read = krnl_partialKnn_wrapper_8_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_8_0_start_id_0 = 64'd65536;
  assign krnl_partialKnn_wrapper_9_0_ap_clk = ap_clk;
  assign krnl_partialKnn_wrapper_9_0__ap_done = krnl_partialKnn_wrapper_9_0_ap_done;
  assign krnl_partialKnn_wrapper_9_0__ap_idle = krnl_partialKnn_wrapper_9_0_ap_idle;
  assign krnl_partialKnn_wrapper_9_0__ap_ready = krnl_partialKnn_wrapper_9_0_ap_ready;
  assign krnl_partialKnn_wrapper_9_0_ap_rst_n = ap_rst_n;
  assign krnl_partialKnn_wrapper_9_0_ap_start = krnl_partialKnn_wrapper_9_0__ap_start;
  assign out_dist_9__din = krnl_partialKnn_wrapper_9_0_out_dist_din;
  assign krnl_partialKnn_wrapper_9_0_out_dist_full_n = out_dist_9__full_n;
  assign out_dist_9__write = krnl_partialKnn_wrapper_9_0_out_dist_write;
  assign out_id_9__din = krnl_partialKnn_wrapper_9_0_out_id_din;
  assign krnl_partialKnn_wrapper_9_0_out_id_full_n = out_id_9__full_n;
  assign out_id_9__write = krnl_partialKnn_wrapper_9_0_out_id_write;
  assign krnl_partialKnn_wrapper_9_0_searchSpace_0_read_addr_offset = krnl_partialKnn_wrapper_9_0___in_9__q0;
  assign in_9_read_addr__din = krnl_partialKnn_wrapper_9_0_searchSpace_0_read_addr_s_din;
  assign krnl_partialKnn_wrapper_9_0_searchSpace_0_read_addr_s_full_n = in_9_read_addr__full_n;
  assign in_9_read_addr__write = krnl_partialKnn_wrapper_9_0_searchSpace_0_read_addr_s_write;
  assign krnl_partialKnn_wrapper_9_0_searchSpace_0_read_data_peek_dout = { 1'b0 , in_9_read_data__dout };
  assign krnl_partialKnn_wrapper_9_0_searchSpace_0_read_data_peek_empty_n = in_9_read_data__empty_n;
  assign krnl_partialKnn_wrapper_9_0_searchSpace_0_read_data_s_dout = { 1'b0 , in_9_read_data__dout };
  assign krnl_partialKnn_wrapper_9_0_searchSpace_0_read_data_s_empty_n = in_9_read_data__empty_n;
  assign in_9_read_data__read = krnl_partialKnn_wrapper_9_0_searchSpace_0_read_data_s_read;
  assign krnl_partialKnn_wrapper_9_0_searchSpace_0_write_addr_offset = krnl_partialKnn_wrapper_9_0___in_9__q0;
  assign in_9_write_addr__din = krnl_partialKnn_wrapper_9_0_searchSpace_0_write_addr_s_din;
  assign krnl_partialKnn_wrapper_9_0_searchSpace_0_write_addr_s_full_n = in_9_write_addr__full_n;
  assign in_9_write_addr__write = krnl_partialKnn_wrapper_9_0_searchSpace_0_write_addr_s_write;
  assign in_9_write_data__din = krnl_partialKnn_wrapper_9_0_searchSpace_0_write_data_din;
  assign krnl_partialKnn_wrapper_9_0_searchSpace_0_write_data_full_n = in_9_write_data__full_n;
  assign in_9_write_data__write = krnl_partialKnn_wrapper_9_0_searchSpace_0_write_data_write;
  assign krnl_partialKnn_wrapper_9_0_searchSpace_0_write_resp_peek_dout = { 1'b0 , in_9_write_resp__dout };
  assign krnl_partialKnn_wrapper_9_0_searchSpace_write_resp_peek_empty_n = in_9_write_resp__empty_n;
  assign krnl_partialKnn_wrapper_9_0_searchSpace_0_write_resp_s_dout = { 1'b0 , in_9_write_resp__dout };
  assign krnl_partialKnn_wrapper_9_0_searchSpace_0_write_resp_s_empty_n = in_9_write_resp__empty_n;
  assign in_9_write_resp__read = krnl_partialKnn_wrapper_9_0_searchSpace_0_write_resp_s_read;
  assign krnl_partialKnn_wrapper_9_0_start_id_0 = 64'd73728;
  assign L3_out_dist__m_axi_clk = ap_clk;
  assign m_axi_L3_out_dist_ARADDR = L3_out_dist__m_axi_m_axi_ARADDR;
  assign m_axi_L3_out_dist_ARBURST = L3_out_dist__m_axi_m_axi_ARBURST;
  assign m_axi_L3_out_dist_ARCACHE = L3_out_dist__m_axi_m_axi_ARCACHE;
  assign m_axi_L3_out_dist_ARID = L3_out_dist__m_axi_m_axi_ARID;
  assign m_axi_L3_out_dist_ARLEN = L3_out_dist__m_axi_m_axi_ARLEN;
  assign m_axi_L3_out_dist_ARLOCK = L3_out_dist__m_axi_m_axi_ARLOCK;
  assign m_axi_L3_out_dist_ARPROT = L3_out_dist__m_axi_m_axi_ARPROT;
  assign m_axi_L3_out_dist_ARQOS = L3_out_dist__m_axi_m_axi_ARQOS;
  assign L3_out_dist__m_axi_m_axi_ARREADY = m_axi_L3_out_dist_ARREADY;
  assign m_axi_L3_out_dist_ARSIZE = L3_out_dist__m_axi_m_axi_ARSIZE;
  assign m_axi_L3_out_dist_ARVALID = L3_out_dist__m_axi_m_axi_ARVALID;
  assign m_axi_L3_out_dist_AWADDR = L3_out_dist__m_axi_m_axi_AWADDR;
  assign m_axi_L3_out_dist_AWBURST = L3_out_dist__m_axi_m_axi_AWBURST;
  assign m_axi_L3_out_dist_AWCACHE = L3_out_dist__m_axi_m_axi_AWCACHE;
  assign m_axi_L3_out_dist_AWID = L3_out_dist__m_axi_m_axi_AWID;
  assign m_axi_L3_out_dist_AWLEN = L3_out_dist__m_axi_m_axi_AWLEN;
  assign m_axi_L3_out_dist_AWLOCK = L3_out_dist__m_axi_m_axi_AWLOCK;
  assign m_axi_L3_out_dist_AWPROT = L3_out_dist__m_axi_m_axi_AWPROT;
  assign m_axi_L3_out_dist_AWQOS = L3_out_dist__m_axi_m_axi_AWQOS;
  assign L3_out_dist__m_axi_m_axi_AWREADY = m_axi_L3_out_dist_AWREADY;
  assign m_axi_L3_out_dist_AWSIZE = L3_out_dist__m_axi_m_axi_AWSIZE;
  assign m_axi_L3_out_dist_AWVALID = L3_out_dist__m_axi_m_axi_AWVALID;
  assign L3_out_dist__m_axi_m_axi_BID = m_axi_L3_out_dist_BID;
  assign m_axi_L3_out_dist_BREADY = L3_out_dist__m_axi_m_axi_BREADY;
  assign L3_out_dist__m_axi_m_axi_BRESP = m_axi_L3_out_dist_BRESP;
  assign L3_out_dist__m_axi_m_axi_BVALID = m_axi_L3_out_dist_BVALID;
  assign L3_out_dist__m_axi_m_axi_RDATA = m_axi_L3_out_dist_RDATA;
  assign L3_out_dist__m_axi_m_axi_RID = m_axi_L3_out_dist_RID;
  assign L3_out_dist__m_axi_m_axi_RLAST = m_axi_L3_out_dist_RLAST;
  assign m_axi_L3_out_dist_RREADY = L3_out_dist__m_axi_m_axi_RREADY;
  assign L3_out_dist__m_axi_m_axi_RRESP = m_axi_L3_out_dist_RRESP;
  assign L3_out_dist__m_axi_m_axi_RVALID = m_axi_L3_out_dist_RVALID;
  assign m_axi_L3_out_dist_WDATA = L3_out_dist__m_axi_m_axi_WDATA;
  assign m_axi_L3_out_dist_WLAST = L3_out_dist__m_axi_m_axi_WLAST;
  assign L3_out_dist__m_axi_m_axi_WREADY = m_axi_L3_out_dist_WREADY;
  assign m_axi_L3_out_dist_WSTRB = L3_out_dist__m_axi_m_axi_WSTRB;
  assign m_axi_L3_out_dist_WVALID = L3_out_dist__m_axi_m_axi_WVALID;
  assign L3_out_dist__m_axi_read_addr_din = L3_out_dist_read_addr__din;
  assign L3_out_dist_read_addr__full_n = L3_out_dist__m_axi_read_addr_full_n;
  assign L3_out_dist__m_axi_read_addr_write = L3_out_dist_read_addr__write;
  assign L3_out_dist_read_data__dout = L3_out_dist__m_axi_read_data_dout;
  assign L3_out_dist_read_data__empty_n = L3_out_dist__m_axi_read_data_empty_n;
  assign L3_out_dist__m_axi_read_data_read = L3_out_dist_read_data__read;
  assign L3_out_dist__m_axi_rst = ~ ap_rst_n;
  assign L3_out_dist__m_axi_write_addr_din = L3_out_dist_write_addr__din;
  assign L3_out_dist_write_addr__full_n = L3_out_dist__m_axi_write_addr_full_n;
  assign L3_out_dist__m_axi_write_addr_write = L3_out_dist_write_addr__write;
  assign L3_out_dist__m_axi_write_data_din = L3_out_dist_write_data__din;
  assign L3_out_dist_write_data__full_n = L3_out_dist__m_axi_write_data_full_n;
  assign L3_out_dist__m_axi_write_data_write = L3_out_dist_write_data__write;
  assign L3_out_dist_write_resp__dout = L3_out_dist__m_axi_write_resp_dout;
  assign L3_out_dist_write_resp__empty_n = L3_out_dist__m_axi_write_resp_empty_n;
  assign L3_out_dist__m_axi_write_resp_read = L3_out_dist_write_resp__read;
  assign L3_out_id__m_axi_clk = ap_clk;
  assign m_axi_L3_out_id_ARADDR = L3_out_id__m_axi_m_axi_ARADDR;
  assign m_axi_L3_out_id_ARBURST = L3_out_id__m_axi_m_axi_ARBURST;
  assign m_axi_L3_out_id_ARCACHE = L3_out_id__m_axi_m_axi_ARCACHE;
  assign m_axi_L3_out_id_ARID = L3_out_id__m_axi_m_axi_ARID;
  assign m_axi_L3_out_id_ARLEN = L3_out_id__m_axi_m_axi_ARLEN;
  assign m_axi_L3_out_id_ARLOCK = L3_out_id__m_axi_m_axi_ARLOCK;
  assign m_axi_L3_out_id_ARPROT = L3_out_id__m_axi_m_axi_ARPROT;
  assign m_axi_L3_out_id_ARQOS = L3_out_id__m_axi_m_axi_ARQOS;
  assign L3_out_id__m_axi_m_axi_ARREADY = m_axi_L3_out_id_ARREADY;
  assign m_axi_L3_out_id_ARSIZE = L3_out_id__m_axi_m_axi_ARSIZE;
  assign m_axi_L3_out_id_ARVALID = L3_out_id__m_axi_m_axi_ARVALID;
  assign m_axi_L3_out_id_AWADDR = L3_out_id__m_axi_m_axi_AWADDR;
  assign m_axi_L3_out_id_AWBURST = L3_out_id__m_axi_m_axi_AWBURST;
  assign m_axi_L3_out_id_AWCACHE = L3_out_id__m_axi_m_axi_AWCACHE;
  assign m_axi_L3_out_id_AWID = L3_out_id__m_axi_m_axi_AWID;
  assign m_axi_L3_out_id_AWLEN = L3_out_id__m_axi_m_axi_AWLEN;
  assign m_axi_L3_out_id_AWLOCK = L3_out_id__m_axi_m_axi_AWLOCK;
  assign m_axi_L3_out_id_AWPROT = L3_out_id__m_axi_m_axi_AWPROT;
  assign m_axi_L3_out_id_AWQOS = L3_out_id__m_axi_m_axi_AWQOS;
  assign L3_out_id__m_axi_m_axi_AWREADY = m_axi_L3_out_id_AWREADY;
  assign m_axi_L3_out_id_AWSIZE = L3_out_id__m_axi_m_axi_AWSIZE;
  assign m_axi_L3_out_id_AWVALID = L3_out_id__m_axi_m_axi_AWVALID;
  assign L3_out_id__m_axi_m_axi_BID = m_axi_L3_out_id_BID;
  assign m_axi_L3_out_id_BREADY = L3_out_id__m_axi_m_axi_BREADY;
  assign L3_out_id__m_axi_m_axi_BRESP = m_axi_L3_out_id_BRESP;
  assign L3_out_id__m_axi_m_axi_BVALID = m_axi_L3_out_id_BVALID;
  assign L3_out_id__m_axi_m_axi_RDATA = m_axi_L3_out_id_RDATA;
  assign L3_out_id__m_axi_m_axi_RID = m_axi_L3_out_id_RID;
  assign L3_out_id__m_axi_m_axi_RLAST = m_axi_L3_out_id_RLAST;
  assign m_axi_L3_out_id_RREADY = L3_out_id__m_axi_m_axi_RREADY;
  assign L3_out_id__m_axi_m_axi_RRESP = m_axi_L3_out_id_RRESP;
  assign L3_out_id__m_axi_m_axi_RVALID = m_axi_L3_out_id_RVALID;
  assign m_axi_L3_out_id_WDATA = L3_out_id__m_axi_m_axi_WDATA;
  assign m_axi_L3_out_id_WLAST = L3_out_id__m_axi_m_axi_WLAST;
  assign L3_out_id__m_axi_m_axi_WREADY = m_axi_L3_out_id_WREADY;
  assign m_axi_L3_out_id_WSTRB = L3_out_id__m_axi_m_axi_WSTRB;
  assign m_axi_L3_out_id_WVALID = L3_out_id__m_axi_m_axi_WVALID;
  assign L3_out_id__m_axi_read_addr_din = L3_out_id_read_addr__din;
  assign L3_out_id_read_addr__full_n = L3_out_id__m_axi_read_addr_full_n;
  assign L3_out_id__m_axi_read_addr_write = L3_out_id_read_addr__write;
  assign L3_out_id_read_data__dout = L3_out_id__m_axi_read_data_dout;
  assign L3_out_id_read_data__empty_n = L3_out_id__m_axi_read_data_empty_n;
  assign L3_out_id__m_axi_read_data_read = L3_out_id_read_data__read;
  assign L3_out_id__m_axi_rst = ~ ap_rst_n;
  assign L3_out_id__m_axi_write_addr_din = L3_out_id_write_addr__din;
  assign L3_out_id_write_addr__full_n = L3_out_id__m_axi_write_addr_full_n;
  assign L3_out_id__m_axi_write_addr_write = L3_out_id_write_addr__write;
  assign L3_out_id__m_axi_write_data_din = L3_out_id_write_data__din;
  assign L3_out_id_write_data__full_n = L3_out_id__m_axi_write_data_full_n;
  assign L3_out_id__m_axi_write_data_write = L3_out_id_write_data__write;
  assign L3_out_id_write_resp__dout = L3_out_id__m_axi_write_resp_dout;
  assign L3_out_id_write_resp__empty_n = L3_out_id__m_axi_write_resp_empty_n;
  assign L3_out_id__m_axi_write_resp_read = L3_out_id_write_resp__read;
  assign in_0__m_axi_clk = ap_clk;
  assign m_axi_in_0_ARADDR = in_0__m_axi_m_axi_ARADDR;
  assign m_axi_in_0_ARBURST = in_0__m_axi_m_axi_ARBURST;
  assign m_axi_in_0_ARCACHE = in_0__m_axi_m_axi_ARCACHE;
  assign m_axi_in_0_ARID = in_0__m_axi_m_axi_ARID;
  assign m_axi_in_0_ARLEN = in_0__m_axi_m_axi_ARLEN;
  assign m_axi_in_0_ARLOCK = in_0__m_axi_m_axi_ARLOCK;
  assign m_axi_in_0_ARPROT = in_0__m_axi_m_axi_ARPROT;
  assign m_axi_in_0_ARQOS = in_0__m_axi_m_axi_ARQOS;
  assign in_0__m_axi_m_axi_ARREADY = m_axi_in_0_ARREADY;
  assign m_axi_in_0_ARSIZE = in_0__m_axi_m_axi_ARSIZE;
  assign m_axi_in_0_ARVALID = in_0__m_axi_m_axi_ARVALID;
  assign m_axi_in_0_AWADDR = in_0__m_axi_m_axi_AWADDR;
  assign m_axi_in_0_AWBURST = in_0__m_axi_m_axi_AWBURST;
  assign m_axi_in_0_AWCACHE = in_0__m_axi_m_axi_AWCACHE;
  assign m_axi_in_0_AWID = in_0__m_axi_m_axi_AWID;
  assign m_axi_in_0_AWLEN = in_0__m_axi_m_axi_AWLEN;
  assign m_axi_in_0_AWLOCK = in_0__m_axi_m_axi_AWLOCK;
  assign m_axi_in_0_AWPROT = in_0__m_axi_m_axi_AWPROT;
  assign m_axi_in_0_AWQOS = in_0__m_axi_m_axi_AWQOS;
  assign in_0__m_axi_m_axi_AWREADY = m_axi_in_0_AWREADY;
  assign m_axi_in_0_AWSIZE = in_0__m_axi_m_axi_AWSIZE;
  assign m_axi_in_0_AWVALID = in_0__m_axi_m_axi_AWVALID;
  assign in_0__m_axi_m_axi_BID = m_axi_in_0_BID;
  assign m_axi_in_0_BREADY = in_0__m_axi_m_axi_BREADY;
  assign in_0__m_axi_m_axi_BRESP = m_axi_in_0_BRESP;
  assign in_0__m_axi_m_axi_BVALID = m_axi_in_0_BVALID;
  assign in_0__m_axi_m_axi_RDATA = m_axi_in_0_RDATA;
  assign in_0__m_axi_m_axi_RID = m_axi_in_0_RID;
  assign in_0__m_axi_m_axi_RLAST = m_axi_in_0_RLAST;
  assign m_axi_in_0_RREADY = in_0__m_axi_m_axi_RREADY;
  assign in_0__m_axi_m_axi_RRESP = m_axi_in_0_RRESP;
  assign in_0__m_axi_m_axi_RVALID = m_axi_in_0_RVALID;
  assign m_axi_in_0_WDATA = in_0__m_axi_m_axi_WDATA;
  assign m_axi_in_0_WLAST = in_0__m_axi_m_axi_WLAST;
  assign in_0__m_axi_m_axi_WREADY = m_axi_in_0_WREADY;
  assign m_axi_in_0_WSTRB = in_0__m_axi_m_axi_WSTRB;
  assign m_axi_in_0_WVALID = in_0__m_axi_m_axi_WVALID;
  assign in_0__m_axi_read_addr_din = in_0_read_addr__din;
  assign in_0_read_addr__full_n = in_0__m_axi_read_addr_full_n;
  assign in_0__m_axi_read_addr_write = in_0_read_addr__write;
  assign in_0_read_data__dout = in_0__m_axi_read_data_dout;
  assign in_0_read_data__empty_n = in_0__m_axi_read_data_empty_n;
  assign in_0__m_axi_read_data_read = in_0_read_data__read;
  assign in_0__m_axi_rst = ~ ap_rst_n;
  assign in_0__m_axi_write_addr_din = in_0_write_addr__din;
  assign in_0_write_addr__full_n = in_0__m_axi_write_addr_full_n;
  assign in_0__m_axi_write_addr_write = in_0_write_addr__write;
  assign in_0__m_axi_write_data_din = in_0_write_data__din;
  assign in_0_write_data__full_n = in_0__m_axi_write_data_full_n;
  assign in_0__m_axi_write_data_write = in_0_write_data__write;
  assign in_0_write_resp__dout = in_0__m_axi_write_resp_dout;
  assign in_0_write_resp__empty_n = in_0__m_axi_write_resp_empty_n;
  assign in_0__m_axi_write_resp_read = in_0_write_resp__read;
  assign in_1__m_axi_clk = ap_clk;
  assign m_axi_in_1_ARADDR = in_1__m_axi_m_axi_ARADDR;
  assign m_axi_in_1_ARBURST = in_1__m_axi_m_axi_ARBURST;
  assign m_axi_in_1_ARCACHE = in_1__m_axi_m_axi_ARCACHE;
  assign m_axi_in_1_ARID = in_1__m_axi_m_axi_ARID;
  assign m_axi_in_1_ARLEN = in_1__m_axi_m_axi_ARLEN;
  assign m_axi_in_1_ARLOCK = in_1__m_axi_m_axi_ARLOCK;
  assign m_axi_in_1_ARPROT = in_1__m_axi_m_axi_ARPROT;
  assign m_axi_in_1_ARQOS = in_1__m_axi_m_axi_ARQOS;
  assign in_1__m_axi_m_axi_ARREADY = m_axi_in_1_ARREADY;
  assign m_axi_in_1_ARSIZE = in_1__m_axi_m_axi_ARSIZE;
  assign m_axi_in_1_ARVALID = in_1__m_axi_m_axi_ARVALID;
  assign m_axi_in_1_AWADDR = in_1__m_axi_m_axi_AWADDR;
  assign m_axi_in_1_AWBURST = in_1__m_axi_m_axi_AWBURST;
  assign m_axi_in_1_AWCACHE = in_1__m_axi_m_axi_AWCACHE;
  assign m_axi_in_1_AWID = in_1__m_axi_m_axi_AWID;
  assign m_axi_in_1_AWLEN = in_1__m_axi_m_axi_AWLEN;
  assign m_axi_in_1_AWLOCK = in_1__m_axi_m_axi_AWLOCK;
  assign m_axi_in_1_AWPROT = in_1__m_axi_m_axi_AWPROT;
  assign m_axi_in_1_AWQOS = in_1__m_axi_m_axi_AWQOS;
  assign in_1__m_axi_m_axi_AWREADY = m_axi_in_1_AWREADY;
  assign m_axi_in_1_AWSIZE = in_1__m_axi_m_axi_AWSIZE;
  assign m_axi_in_1_AWVALID = in_1__m_axi_m_axi_AWVALID;
  assign in_1__m_axi_m_axi_BID = m_axi_in_1_BID;
  assign m_axi_in_1_BREADY = in_1__m_axi_m_axi_BREADY;
  assign in_1__m_axi_m_axi_BRESP = m_axi_in_1_BRESP;
  assign in_1__m_axi_m_axi_BVALID = m_axi_in_1_BVALID;
  assign in_1__m_axi_m_axi_RDATA = m_axi_in_1_RDATA;
  assign in_1__m_axi_m_axi_RID = m_axi_in_1_RID;
  assign in_1__m_axi_m_axi_RLAST = m_axi_in_1_RLAST;
  assign m_axi_in_1_RREADY = in_1__m_axi_m_axi_RREADY;
  assign in_1__m_axi_m_axi_RRESP = m_axi_in_1_RRESP;
  assign in_1__m_axi_m_axi_RVALID = m_axi_in_1_RVALID;
  assign m_axi_in_1_WDATA = in_1__m_axi_m_axi_WDATA;
  assign m_axi_in_1_WLAST = in_1__m_axi_m_axi_WLAST;
  assign in_1__m_axi_m_axi_WREADY = m_axi_in_1_WREADY;
  assign m_axi_in_1_WSTRB = in_1__m_axi_m_axi_WSTRB;
  assign m_axi_in_1_WVALID = in_1__m_axi_m_axi_WVALID;
  assign in_1__m_axi_read_addr_din = in_1_read_addr__din;
  assign in_1_read_addr__full_n = in_1__m_axi_read_addr_full_n;
  assign in_1__m_axi_read_addr_write = in_1_read_addr__write;
  assign in_1_read_data__dout = in_1__m_axi_read_data_dout;
  assign in_1_read_data__empty_n = in_1__m_axi_read_data_empty_n;
  assign in_1__m_axi_read_data_read = in_1_read_data__read;
  assign in_1__m_axi_rst = ~ ap_rst_n;
  assign in_1__m_axi_write_addr_din = in_1_write_addr__din;
  assign in_1_write_addr__full_n = in_1__m_axi_write_addr_full_n;
  assign in_1__m_axi_write_addr_write = in_1_write_addr__write;
  assign in_1__m_axi_write_data_din = in_1_write_data__din;
  assign in_1_write_data__full_n = in_1__m_axi_write_data_full_n;
  assign in_1__m_axi_write_data_write = in_1_write_data__write;
  assign in_1_write_resp__dout = in_1__m_axi_write_resp_dout;
  assign in_1_write_resp__empty_n = in_1__m_axi_write_resp_empty_n;
  assign in_1__m_axi_write_resp_read = in_1_write_resp__read;
  assign in_10__m_axi_clk = ap_clk;
  assign m_axi_in_10_ARADDR = in_10__m_axi_m_axi_ARADDR;
  assign m_axi_in_10_ARBURST = in_10__m_axi_m_axi_ARBURST;
  assign m_axi_in_10_ARCACHE = in_10__m_axi_m_axi_ARCACHE;
  assign m_axi_in_10_ARID = in_10__m_axi_m_axi_ARID;
  assign m_axi_in_10_ARLEN = in_10__m_axi_m_axi_ARLEN;
  assign m_axi_in_10_ARLOCK = in_10__m_axi_m_axi_ARLOCK;
  assign m_axi_in_10_ARPROT = in_10__m_axi_m_axi_ARPROT;
  assign m_axi_in_10_ARQOS = in_10__m_axi_m_axi_ARQOS;
  assign in_10__m_axi_m_axi_ARREADY = m_axi_in_10_ARREADY;
  assign m_axi_in_10_ARSIZE = in_10__m_axi_m_axi_ARSIZE;
  assign m_axi_in_10_ARVALID = in_10__m_axi_m_axi_ARVALID;
  assign m_axi_in_10_AWADDR = in_10__m_axi_m_axi_AWADDR;
  assign m_axi_in_10_AWBURST = in_10__m_axi_m_axi_AWBURST;
  assign m_axi_in_10_AWCACHE = in_10__m_axi_m_axi_AWCACHE;
  assign m_axi_in_10_AWID = in_10__m_axi_m_axi_AWID;
  assign m_axi_in_10_AWLEN = in_10__m_axi_m_axi_AWLEN;
  assign m_axi_in_10_AWLOCK = in_10__m_axi_m_axi_AWLOCK;
  assign m_axi_in_10_AWPROT = in_10__m_axi_m_axi_AWPROT;
  assign m_axi_in_10_AWQOS = in_10__m_axi_m_axi_AWQOS;
  assign in_10__m_axi_m_axi_AWREADY = m_axi_in_10_AWREADY;
  assign m_axi_in_10_AWSIZE = in_10__m_axi_m_axi_AWSIZE;
  assign m_axi_in_10_AWVALID = in_10__m_axi_m_axi_AWVALID;
  assign in_10__m_axi_m_axi_BID = m_axi_in_10_BID;
  assign m_axi_in_10_BREADY = in_10__m_axi_m_axi_BREADY;
  assign in_10__m_axi_m_axi_BRESP = m_axi_in_10_BRESP;
  assign in_10__m_axi_m_axi_BVALID = m_axi_in_10_BVALID;
  assign in_10__m_axi_m_axi_RDATA = m_axi_in_10_RDATA;
  assign in_10__m_axi_m_axi_RID = m_axi_in_10_RID;
  assign in_10__m_axi_m_axi_RLAST = m_axi_in_10_RLAST;
  assign m_axi_in_10_RREADY = in_10__m_axi_m_axi_RREADY;
  assign in_10__m_axi_m_axi_RRESP = m_axi_in_10_RRESP;
  assign in_10__m_axi_m_axi_RVALID = m_axi_in_10_RVALID;
  assign m_axi_in_10_WDATA = in_10__m_axi_m_axi_WDATA;
  assign m_axi_in_10_WLAST = in_10__m_axi_m_axi_WLAST;
  assign in_10__m_axi_m_axi_WREADY = m_axi_in_10_WREADY;
  assign m_axi_in_10_WSTRB = in_10__m_axi_m_axi_WSTRB;
  assign m_axi_in_10_WVALID = in_10__m_axi_m_axi_WVALID;
  assign in_10__m_axi_read_addr_din = in_10_read_addr__din;
  assign in_10_read_addr__full_n = in_10__m_axi_read_addr_full_n;
  assign in_10__m_axi_read_addr_write = in_10_read_addr__write;
  assign in_10_read_data__dout = in_10__m_axi_read_data_dout;
  assign in_10_read_data__empty_n = in_10__m_axi_read_data_empty_n;
  assign in_10__m_axi_read_data_read = in_10_read_data__read;
  assign in_10__m_axi_rst = ~ ap_rst_n;
  assign in_10__m_axi_write_addr_din = in_10_write_addr__din;
  assign in_10_write_addr__full_n = in_10__m_axi_write_addr_full_n;
  assign in_10__m_axi_write_addr_write = in_10_write_addr__write;
  assign in_10__m_axi_write_data_din = in_10_write_data__din;
  assign in_10_write_data__full_n = in_10__m_axi_write_data_full_n;
  assign in_10__m_axi_write_data_write = in_10_write_data__write;
  assign in_10_write_resp__dout = in_10__m_axi_write_resp_dout;
  assign in_10_write_resp__empty_n = in_10__m_axi_write_resp_empty_n;
  assign in_10__m_axi_write_resp_read = in_10_write_resp__read;
  assign in_11__m_axi_clk = ap_clk;
  assign m_axi_in_11_ARADDR = in_11__m_axi_m_axi_ARADDR;
  assign m_axi_in_11_ARBURST = in_11__m_axi_m_axi_ARBURST;
  assign m_axi_in_11_ARCACHE = in_11__m_axi_m_axi_ARCACHE;
  assign m_axi_in_11_ARID = in_11__m_axi_m_axi_ARID;
  assign m_axi_in_11_ARLEN = in_11__m_axi_m_axi_ARLEN;
  assign m_axi_in_11_ARLOCK = in_11__m_axi_m_axi_ARLOCK;
  assign m_axi_in_11_ARPROT = in_11__m_axi_m_axi_ARPROT;
  assign m_axi_in_11_ARQOS = in_11__m_axi_m_axi_ARQOS;
  assign in_11__m_axi_m_axi_ARREADY = m_axi_in_11_ARREADY;
  assign m_axi_in_11_ARSIZE = in_11__m_axi_m_axi_ARSIZE;
  assign m_axi_in_11_ARVALID = in_11__m_axi_m_axi_ARVALID;
  assign m_axi_in_11_AWADDR = in_11__m_axi_m_axi_AWADDR;
  assign m_axi_in_11_AWBURST = in_11__m_axi_m_axi_AWBURST;
  assign m_axi_in_11_AWCACHE = in_11__m_axi_m_axi_AWCACHE;
  assign m_axi_in_11_AWID = in_11__m_axi_m_axi_AWID;
  assign m_axi_in_11_AWLEN = in_11__m_axi_m_axi_AWLEN;
  assign m_axi_in_11_AWLOCK = in_11__m_axi_m_axi_AWLOCK;
  assign m_axi_in_11_AWPROT = in_11__m_axi_m_axi_AWPROT;
  assign m_axi_in_11_AWQOS = in_11__m_axi_m_axi_AWQOS;
  assign in_11__m_axi_m_axi_AWREADY = m_axi_in_11_AWREADY;
  assign m_axi_in_11_AWSIZE = in_11__m_axi_m_axi_AWSIZE;
  assign m_axi_in_11_AWVALID = in_11__m_axi_m_axi_AWVALID;
  assign in_11__m_axi_m_axi_BID = m_axi_in_11_BID;
  assign m_axi_in_11_BREADY = in_11__m_axi_m_axi_BREADY;
  assign in_11__m_axi_m_axi_BRESP = m_axi_in_11_BRESP;
  assign in_11__m_axi_m_axi_BVALID = m_axi_in_11_BVALID;
  assign in_11__m_axi_m_axi_RDATA = m_axi_in_11_RDATA;
  assign in_11__m_axi_m_axi_RID = m_axi_in_11_RID;
  assign in_11__m_axi_m_axi_RLAST = m_axi_in_11_RLAST;
  assign m_axi_in_11_RREADY = in_11__m_axi_m_axi_RREADY;
  assign in_11__m_axi_m_axi_RRESP = m_axi_in_11_RRESP;
  assign in_11__m_axi_m_axi_RVALID = m_axi_in_11_RVALID;
  assign m_axi_in_11_WDATA = in_11__m_axi_m_axi_WDATA;
  assign m_axi_in_11_WLAST = in_11__m_axi_m_axi_WLAST;
  assign in_11__m_axi_m_axi_WREADY = m_axi_in_11_WREADY;
  assign m_axi_in_11_WSTRB = in_11__m_axi_m_axi_WSTRB;
  assign m_axi_in_11_WVALID = in_11__m_axi_m_axi_WVALID;
  assign in_11__m_axi_read_addr_din = in_11_read_addr__din;
  assign in_11_read_addr__full_n = in_11__m_axi_read_addr_full_n;
  assign in_11__m_axi_read_addr_write = in_11_read_addr__write;
  assign in_11_read_data__dout = in_11__m_axi_read_data_dout;
  assign in_11_read_data__empty_n = in_11__m_axi_read_data_empty_n;
  assign in_11__m_axi_read_data_read = in_11_read_data__read;
  assign in_11__m_axi_rst = ~ ap_rst_n;
  assign in_11__m_axi_write_addr_din = in_11_write_addr__din;
  assign in_11_write_addr__full_n = in_11__m_axi_write_addr_full_n;
  assign in_11__m_axi_write_addr_write = in_11_write_addr__write;
  assign in_11__m_axi_write_data_din = in_11_write_data__din;
  assign in_11_write_data__full_n = in_11__m_axi_write_data_full_n;
  assign in_11__m_axi_write_data_write = in_11_write_data__write;
  assign in_11_write_resp__dout = in_11__m_axi_write_resp_dout;
  assign in_11_write_resp__empty_n = in_11__m_axi_write_resp_empty_n;
  assign in_11__m_axi_write_resp_read = in_11_write_resp__read;
  assign in_12__m_axi_clk = ap_clk;
  assign m_axi_in_12_ARADDR = in_12__m_axi_m_axi_ARADDR;
  assign m_axi_in_12_ARBURST = in_12__m_axi_m_axi_ARBURST;
  assign m_axi_in_12_ARCACHE = in_12__m_axi_m_axi_ARCACHE;
  assign m_axi_in_12_ARID = in_12__m_axi_m_axi_ARID;
  assign m_axi_in_12_ARLEN = in_12__m_axi_m_axi_ARLEN;
  assign m_axi_in_12_ARLOCK = in_12__m_axi_m_axi_ARLOCK;
  assign m_axi_in_12_ARPROT = in_12__m_axi_m_axi_ARPROT;
  assign m_axi_in_12_ARQOS = in_12__m_axi_m_axi_ARQOS;
  assign in_12__m_axi_m_axi_ARREADY = m_axi_in_12_ARREADY;
  assign m_axi_in_12_ARSIZE = in_12__m_axi_m_axi_ARSIZE;
  assign m_axi_in_12_ARVALID = in_12__m_axi_m_axi_ARVALID;
  assign m_axi_in_12_AWADDR = in_12__m_axi_m_axi_AWADDR;
  assign m_axi_in_12_AWBURST = in_12__m_axi_m_axi_AWBURST;
  assign m_axi_in_12_AWCACHE = in_12__m_axi_m_axi_AWCACHE;
  assign m_axi_in_12_AWID = in_12__m_axi_m_axi_AWID;
  assign m_axi_in_12_AWLEN = in_12__m_axi_m_axi_AWLEN;
  assign m_axi_in_12_AWLOCK = in_12__m_axi_m_axi_AWLOCK;
  assign m_axi_in_12_AWPROT = in_12__m_axi_m_axi_AWPROT;
  assign m_axi_in_12_AWQOS = in_12__m_axi_m_axi_AWQOS;
  assign in_12__m_axi_m_axi_AWREADY = m_axi_in_12_AWREADY;
  assign m_axi_in_12_AWSIZE = in_12__m_axi_m_axi_AWSIZE;
  assign m_axi_in_12_AWVALID = in_12__m_axi_m_axi_AWVALID;
  assign in_12__m_axi_m_axi_BID = m_axi_in_12_BID;
  assign m_axi_in_12_BREADY = in_12__m_axi_m_axi_BREADY;
  assign in_12__m_axi_m_axi_BRESP = m_axi_in_12_BRESP;
  assign in_12__m_axi_m_axi_BVALID = m_axi_in_12_BVALID;
  assign in_12__m_axi_m_axi_RDATA = m_axi_in_12_RDATA;
  assign in_12__m_axi_m_axi_RID = m_axi_in_12_RID;
  assign in_12__m_axi_m_axi_RLAST = m_axi_in_12_RLAST;
  assign m_axi_in_12_RREADY = in_12__m_axi_m_axi_RREADY;
  assign in_12__m_axi_m_axi_RRESP = m_axi_in_12_RRESP;
  assign in_12__m_axi_m_axi_RVALID = m_axi_in_12_RVALID;
  assign m_axi_in_12_WDATA = in_12__m_axi_m_axi_WDATA;
  assign m_axi_in_12_WLAST = in_12__m_axi_m_axi_WLAST;
  assign in_12__m_axi_m_axi_WREADY = m_axi_in_12_WREADY;
  assign m_axi_in_12_WSTRB = in_12__m_axi_m_axi_WSTRB;
  assign m_axi_in_12_WVALID = in_12__m_axi_m_axi_WVALID;
  assign in_12__m_axi_read_addr_din = in_12_read_addr__din;
  assign in_12_read_addr__full_n = in_12__m_axi_read_addr_full_n;
  assign in_12__m_axi_read_addr_write = in_12_read_addr__write;
  assign in_12_read_data__dout = in_12__m_axi_read_data_dout;
  assign in_12_read_data__empty_n = in_12__m_axi_read_data_empty_n;
  assign in_12__m_axi_read_data_read = in_12_read_data__read;
  assign in_12__m_axi_rst = ~ ap_rst_n;
  assign in_12__m_axi_write_addr_din = in_12_write_addr__din;
  assign in_12_write_addr__full_n = in_12__m_axi_write_addr_full_n;
  assign in_12__m_axi_write_addr_write = in_12_write_addr__write;
  assign in_12__m_axi_write_data_din = in_12_write_data__din;
  assign in_12_write_data__full_n = in_12__m_axi_write_data_full_n;
  assign in_12__m_axi_write_data_write = in_12_write_data__write;
  assign in_12_write_resp__dout = in_12__m_axi_write_resp_dout;
  assign in_12_write_resp__empty_n = in_12__m_axi_write_resp_empty_n;
  assign in_12__m_axi_write_resp_read = in_12_write_resp__read;
  assign in_13__m_axi_clk = ap_clk;
  assign m_axi_in_13_ARADDR = in_13__m_axi_m_axi_ARADDR;
  assign m_axi_in_13_ARBURST = in_13__m_axi_m_axi_ARBURST;
  assign m_axi_in_13_ARCACHE = in_13__m_axi_m_axi_ARCACHE;
  assign m_axi_in_13_ARID = in_13__m_axi_m_axi_ARID;
  assign m_axi_in_13_ARLEN = in_13__m_axi_m_axi_ARLEN;
  assign m_axi_in_13_ARLOCK = in_13__m_axi_m_axi_ARLOCK;
  assign m_axi_in_13_ARPROT = in_13__m_axi_m_axi_ARPROT;
  assign m_axi_in_13_ARQOS = in_13__m_axi_m_axi_ARQOS;
  assign in_13__m_axi_m_axi_ARREADY = m_axi_in_13_ARREADY;
  assign m_axi_in_13_ARSIZE = in_13__m_axi_m_axi_ARSIZE;
  assign m_axi_in_13_ARVALID = in_13__m_axi_m_axi_ARVALID;
  assign m_axi_in_13_AWADDR = in_13__m_axi_m_axi_AWADDR;
  assign m_axi_in_13_AWBURST = in_13__m_axi_m_axi_AWBURST;
  assign m_axi_in_13_AWCACHE = in_13__m_axi_m_axi_AWCACHE;
  assign m_axi_in_13_AWID = in_13__m_axi_m_axi_AWID;
  assign m_axi_in_13_AWLEN = in_13__m_axi_m_axi_AWLEN;
  assign m_axi_in_13_AWLOCK = in_13__m_axi_m_axi_AWLOCK;
  assign m_axi_in_13_AWPROT = in_13__m_axi_m_axi_AWPROT;
  assign m_axi_in_13_AWQOS = in_13__m_axi_m_axi_AWQOS;
  assign in_13__m_axi_m_axi_AWREADY = m_axi_in_13_AWREADY;
  assign m_axi_in_13_AWSIZE = in_13__m_axi_m_axi_AWSIZE;
  assign m_axi_in_13_AWVALID = in_13__m_axi_m_axi_AWVALID;
  assign in_13__m_axi_m_axi_BID = m_axi_in_13_BID;
  assign m_axi_in_13_BREADY = in_13__m_axi_m_axi_BREADY;
  assign in_13__m_axi_m_axi_BRESP = m_axi_in_13_BRESP;
  assign in_13__m_axi_m_axi_BVALID = m_axi_in_13_BVALID;
  assign in_13__m_axi_m_axi_RDATA = m_axi_in_13_RDATA;
  assign in_13__m_axi_m_axi_RID = m_axi_in_13_RID;
  assign in_13__m_axi_m_axi_RLAST = m_axi_in_13_RLAST;
  assign m_axi_in_13_RREADY = in_13__m_axi_m_axi_RREADY;
  assign in_13__m_axi_m_axi_RRESP = m_axi_in_13_RRESP;
  assign in_13__m_axi_m_axi_RVALID = m_axi_in_13_RVALID;
  assign m_axi_in_13_WDATA = in_13__m_axi_m_axi_WDATA;
  assign m_axi_in_13_WLAST = in_13__m_axi_m_axi_WLAST;
  assign in_13__m_axi_m_axi_WREADY = m_axi_in_13_WREADY;
  assign m_axi_in_13_WSTRB = in_13__m_axi_m_axi_WSTRB;
  assign m_axi_in_13_WVALID = in_13__m_axi_m_axi_WVALID;
  assign in_13__m_axi_read_addr_din = in_13_read_addr__din;
  assign in_13_read_addr__full_n = in_13__m_axi_read_addr_full_n;
  assign in_13__m_axi_read_addr_write = in_13_read_addr__write;
  assign in_13_read_data__dout = in_13__m_axi_read_data_dout;
  assign in_13_read_data__empty_n = in_13__m_axi_read_data_empty_n;
  assign in_13__m_axi_read_data_read = in_13_read_data__read;
  assign in_13__m_axi_rst = ~ ap_rst_n;
  assign in_13__m_axi_write_addr_din = in_13_write_addr__din;
  assign in_13_write_addr__full_n = in_13__m_axi_write_addr_full_n;
  assign in_13__m_axi_write_addr_write = in_13_write_addr__write;
  assign in_13__m_axi_write_data_din = in_13_write_data__din;
  assign in_13_write_data__full_n = in_13__m_axi_write_data_full_n;
  assign in_13__m_axi_write_data_write = in_13_write_data__write;
  assign in_13_write_resp__dout = in_13__m_axi_write_resp_dout;
  assign in_13_write_resp__empty_n = in_13__m_axi_write_resp_empty_n;
  assign in_13__m_axi_write_resp_read = in_13_write_resp__read;
  assign in_14__m_axi_clk = ap_clk;
  assign m_axi_in_14_ARADDR = in_14__m_axi_m_axi_ARADDR;
  assign m_axi_in_14_ARBURST = in_14__m_axi_m_axi_ARBURST;
  assign m_axi_in_14_ARCACHE = in_14__m_axi_m_axi_ARCACHE;
  assign m_axi_in_14_ARID = in_14__m_axi_m_axi_ARID;
  assign m_axi_in_14_ARLEN = in_14__m_axi_m_axi_ARLEN;
  assign m_axi_in_14_ARLOCK = in_14__m_axi_m_axi_ARLOCK;
  assign m_axi_in_14_ARPROT = in_14__m_axi_m_axi_ARPROT;
  assign m_axi_in_14_ARQOS = in_14__m_axi_m_axi_ARQOS;
  assign in_14__m_axi_m_axi_ARREADY = m_axi_in_14_ARREADY;
  assign m_axi_in_14_ARSIZE = in_14__m_axi_m_axi_ARSIZE;
  assign m_axi_in_14_ARVALID = in_14__m_axi_m_axi_ARVALID;
  assign m_axi_in_14_AWADDR = in_14__m_axi_m_axi_AWADDR;
  assign m_axi_in_14_AWBURST = in_14__m_axi_m_axi_AWBURST;
  assign m_axi_in_14_AWCACHE = in_14__m_axi_m_axi_AWCACHE;
  assign m_axi_in_14_AWID = in_14__m_axi_m_axi_AWID;
  assign m_axi_in_14_AWLEN = in_14__m_axi_m_axi_AWLEN;
  assign m_axi_in_14_AWLOCK = in_14__m_axi_m_axi_AWLOCK;
  assign m_axi_in_14_AWPROT = in_14__m_axi_m_axi_AWPROT;
  assign m_axi_in_14_AWQOS = in_14__m_axi_m_axi_AWQOS;
  assign in_14__m_axi_m_axi_AWREADY = m_axi_in_14_AWREADY;
  assign m_axi_in_14_AWSIZE = in_14__m_axi_m_axi_AWSIZE;
  assign m_axi_in_14_AWVALID = in_14__m_axi_m_axi_AWVALID;
  assign in_14__m_axi_m_axi_BID = m_axi_in_14_BID;
  assign m_axi_in_14_BREADY = in_14__m_axi_m_axi_BREADY;
  assign in_14__m_axi_m_axi_BRESP = m_axi_in_14_BRESP;
  assign in_14__m_axi_m_axi_BVALID = m_axi_in_14_BVALID;
  assign in_14__m_axi_m_axi_RDATA = m_axi_in_14_RDATA;
  assign in_14__m_axi_m_axi_RID = m_axi_in_14_RID;
  assign in_14__m_axi_m_axi_RLAST = m_axi_in_14_RLAST;
  assign m_axi_in_14_RREADY = in_14__m_axi_m_axi_RREADY;
  assign in_14__m_axi_m_axi_RRESP = m_axi_in_14_RRESP;
  assign in_14__m_axi_m_axi_RVALID = m_axi_in_14_RVALID;
  assign m_axi_in_14_WDATA = in_14__m_axi_m_axi_WDATA;
  assign m_axi_in_14_WLAST = in_14__m_axi_m_axi_WLAST;
  assign in_14__m_axi_m_axi_WREADY = m_axi_in_14_WREADY;
  assign m_axi_in_14_WSTRB = in_14__m_axi_m_axi_WSTRB;
  assign m_axi_in_14_WVALID = in_14__m_axi_m_axi_WVALID;
  assign in_14__m_axi_read_addr_din = in_14_read_addr__din;
  assign in_14_read_addr__full_n = in_14__m_axi_read_addr_full_n;
  assign in_14__m_axi_read_addr_write = in_14_read_addr__write;
  assign in_14_read_data__dout = in_14__m_axi_read_data_dout;
  assign in_14_read_data__empty_n = in_14__m_axi_read_data_empty_n;
  assign in_14__m_axi_read_data_read = in_14_read_data__read;
  assign in_14__m_axi_rst = ~ ap_rst_n;
  assign in_14__m_axi_write_addr_din = in_14_write_addr__din;
  assign in_14_write_addr__full_n = in_14__m_axi_write_addr_full_n;
  assign in_14__m_axi_write_addr_write = in_14_write_addr__write;
  assign in_14__m_axi_write_data_din = in_14_write_data__din;
  assign in_14_write_data__full_n = in_14__m_axi_write_data_full_n;
  assign in_14__m_axi_write_data_write = in_14_write_data__write;
  assign in_14_write_resp__dout = in_14__m_axi_write_resp_dout;
  assign in_14_write_resp__empty_n = in_14__m_axi_write_resp_empty_n;
  assign in_14__m_axi_write_resp_read = in_14_write_resp__read;
  assign in_15__m_axi_clk = ap_clk;
  assign m_axi_in_15_ARADDR = in_15__m_axi_m_axi_ARADDR;
  assign m_axi_in_15_ARBURST = in_15__m_axi_m_axi_ARBURST;
  assign m_axi_in_15_ARCACHE = in_15__m_axi_m_axi_ARCACHE;
  assign m_axi_in_15_ARID = in_15__m_axi_m_axi_ARID;
  assign m_axi_in_15_ARLEN = in_15__m_axi_m_axi_ARLEN;
  assign m_axi_in_15_ARLOCK = in_15__m_axi_m_axi_ARLOCK;
  assign m_axi_in_15_ARPROT = in_15__m_axi_m_axi_ARPROT;
  assign m_axi_in_15_ARQOS = in_15__m_axi_m_axi_ARQOS;
  assign in_15__m_axi_m_axi_ARREADY = m_axi_in_15_ARREADY;
  assign m_axi_in_15_ARSIZE = in_15__m_axi_m_axi_ARSIZE;
  assign m_axi_in_15_ARVALID = in_15__m_axi_m_axi_ARVALID;
  assign m_axi_in_15_AWADDR = in_15__m_axi_m_axi_AWADDR;
  assign m_axi_in_15_AWBURST = in_15__m_axi_m_axi_AWBURST;
  assign m_axi_in_15_AWCACHE = in_15__m_axi_m_axi_AWCACHE;
  assign m_axi_in_15_AWID = in_15__m_axi_m_axi_AWID;
  assign m_axi_in_15_AWLEN = in_15__m_axi_m_axi_AWLEN;
  assign m_axi_in_15_AWLOCK = in_15__m_axi_m_axi_AWLOCK;
  assign m_axi_in_15_AWPROT = in_15__m_axi_m_axi_AWPROT;
  assign m_axi_in_15_AWQOS = in_15__m_axi_m_axi_AWQOS;
  assign in_15__m_axi_m_axi_AWREADY = m_axi_in_15_AWREADY;
  assign m_axi_in_15_AWSIZE = in_15__m_axi_m_axi_AWSIZE;
  assign m_axi_in_15_AWVALID = in_15__m_axi_m_axi_AWVALID;
  assign in_15__m_axi_m_axi_BID = m_axi_in_15_BID;
  assign m_axi_in_15_BREADY = in_15__m_axi_m_axi_BREADY;
  assign in_15__m_axi_m_axi_BRESP = m_axi_in_15_BRESP;
  assign in_15__m_axi_m_axi_BVALID = m_axi_in_15_BVALID;
  assign in_15__m_axi_m_axi_RDATA = m_axi_in_15_RDATA;
  assign in_15__m_axi_m_axi_RID = m_axi_in_15_RID;
  assign in_15__m_axi_m_axi_RLAST = m_axi_in_15_RLAST;
  assign m_axi_in_15_RREADY = in_15__m_axi_m_axi_RREADY;
  assign in_15__m_axi_m_axi_RRESP = m_axi_in_15_RRESP;
  assign in_15__m_axi_m_axi_RVALID = m_axi_in_15_RVALID;
  assign m_axi_in_15_WDATA = in_15__m_axi_m_axi_WDATA;
  assign m_axi_in_15_WLAST = in_15__m_axi_m_axi_WLAST;
  assign in_15__m_axi_m_axi_WREADY = m_axi_in_15_WREADY;
  assign m_axi_in_15_WSTRB = in_15__m_axi_m_axi_WSTRB;
  assign m_axi_in_15_WVALID = in_15__m_axi_m_axi_WVALID;
  assign in_15__m_axi_read_addr_din = in_15_read_addr__din;
  assign in_15_read_addr__full_n = in_15__m_axi_read_addr_full_n;
  assign in_15__m_axi_read_addr_write = in_15_read_addr__write;
  assign in_15_read_data__dout = in_15__m_axi_read_data_dout;
  assign in_15_read_data__empty_n = in_15__m_axi_read_data_empty_n;
  assign in_15__m_axi_read_data_read = in_15_read_data__read;
  assign in_15__m_axi_rst = ~ ap_rst_n;
  assign in_15__m_axi_write_addr_din = in_15_write_addr__din;
  assign in_15_write_addr__full_n = in_15__m_axi_write_addr_full_n;
  assign in_15__m_axi_write_addr_write = in_15_write_addr__write;
  assign in_15__m_axi_write_data_din = in_15_write_data__din;
  assign in_15_write_data__full_n = in_15__m_axi_write_data_full_n;
  assign in_15__m_axi_write_data_write = in_15_write_data__write;
  assign in_15_write_resp__dout = in_15__m_axi_write_resp_dout;
  assign in_15_write_resp__empty_n = in_15__m_axi_write_resp_empty_n;
  assign in_15__m_axi_write_resp_read = in_15_write_resp__read;
  assign in_16__m_axi_clk = ap_clk;
  assign m_axi_in_16_ARADDR = in_16__m_axi_m_axi_ARADDR;
  assign m_axi_in_16_ARBURST = in_16__m_axi_m_axi_ARBURST;
  assign m_axi_in_16_ARCACHE = in_16__m_axi_m_axi_ARCACHE;
  assign m_axi_in_16_ARID = in_16__m_axi_m_axi_ARID;
  assign m_axi_in_16_ARLEN = in_16__m_axi_m_axi_ARLEN;
  assign m_axi_in_16_ARLOCK = in_16__m_axi_m_axi_ARLOCK;
  assign m_axi_in_16_ARPROT = in_16__m_axi_m_axi_ARPROT;
  assign m_axi_in_16_ARQOS = in_16__m_axi_m_axi_ARQOS;
  assign in_16__m_axi_m_axi_ARREADY = m_axi_in_16_ARREADY;
  assign m_axi_in_16_ARSIZE = in_16__m_axi_m_axi_ARSIZE;
  assign m_axi_in_16_ARVALID = in_16__m_axi_m_axi_ARVALID;
  assign m_axi_in_16_AWADDR = in_16__m_axi_m_axi_AWADDR;
  assign m_axi_in_16_AWBURST = in_16__m_axi_m_axi_AWBURST;
  assign m_axi_in_16_AWCACHE = in_16__m_axi_m_axi_AWCACHE;
  assign m_axi_in_16_AWID = in_16__m_axi_m_axi_AWID;
  assign m_axi_in_16_AWLEN = in_16__m_axi_m_axi_AWLEN;
  assign m_axi_in_16_AWLOCK = in_16__m_axi_m_axi_AWLOCK;
  assign m_axi_in_16_AWPROT = in_16__m_axi_m_axi_AWPROT;
  assign m_axi_in_16_AWQOS = in_16__m_axi_m_axi_AWQOS;
  assign in_16__m_axi_m_axi_AWREADY = m_axi_in_16_AWREADY;
  assign m_axi_in_16_AWSIZE = in_16__m_axi_m_axi_AWSIZE;
  assign m_axi_in_16_AWVALID = in_16__m_axi_m_axi_AWVALID;
  assign in_16__m_axi_m_axi_BID = m_axi_in_16_BID;
  assign m_axi_in_16_BREADY = in_16__m_axi_m_axi_BREADY;
  assign in_16__m_axi_m_axi_BRESP = m_axi_in_16_BRESP;
  assign in_16__m_axi_m_axi_BVALID = m_axi_in_16_BVALID;
  assign in_16__m_axi_m_axi_RDATA = m_axi_in_16_RDATA;
  assign in_16__m_axi_m_axi_RID = m_axi_in_16_RID;
  assign in_16__m_axi_m_axi_RLAST = m_axi_in_16_RLAST;
  assign m_axi_in_16_RREADY = in_16__m_axi_m_axi_RREADY;
  assign in_16__m_axi_m_axi_RRESP = m_axi_in_16_RRESP;
  assign in_16__m_axi_m_axi_RVALID = m_axi_in_16_RVALID;
  assign m_axi_in_16_WDATA = in_16__m_axi_m_axi_WDATA;
  assign m_axi_in_16_WLAST = in_16__m_axi_m_axi_WLAST;
  assign in_16__m_axi_m_axi_WREADY = m_axi_in_16_WREADY;
  assign m_axi_in_16_WSTRB = in_16__m_axi_m_axi_WSTRB;
  assign m_axi_in_16_WVALID = in_16__m_axi_m_axi_WVALID;
  assign in_16__m_axi_read_addr_din = in_16_read_addr__din;
  assign in_16_read_addr__full_n = in_16__m_axi_read_addr_full_n;
  assign in_16__m_axi_read_addr_write = in_16_read_addr__write;
  assign in_16_read_data__dout = in_16__m_axi_read_data_dout;
  assign in_16_read_data__empty_n = in_16__m_axi_read_data_empty_n;
  assign in_16__m_axi_read_data_read = in_16_read_data__read;
  assign in_16__m_axi_rst = ~ ap_rst_n;
  assign in_16__m_axi_write_addr_din = in_16_write_addr__din;
  assign in_16_write_addr__full_n = in_16__m_axi_write_addr_full_n;
  assign in_16__m_axi_write_addr_write = in_16_write_addr__write;
  assign in_16__m_axi_write_data_din = in_16_write_data__din;
  assign in_16_write_data__full_n = in_16__m_axi_write_data_full_n;
  assign in_16__m_axi_write_data_write = in_16_write_data__write;
  assign in_16_write_resp__dout = in_16__m_axi_write_resp_dout;
  assign in_16_write_resp__empty_n = in_16__m_axi_write_resp_empty_n;
  assign in_16__m_axi_write_resp_read = in_16_write_resp__read;
  assign in_17__m_axi_clk = ap_clk;
  assign m_axi_in_17_ARADDR = in_17__m_axi_m_axi_ARADDR;
  assign m_axi_in_17_ARBURST = in_17__m_axi_m_axi_ARBURST;
  assign m_axi_in_17_ARCACHE = in_17__m_axi_m_axi_ARCACHE;
  assign m_axi_in_17_ARID = in_17__m_axi_m_axi_ARID;
  assign m_axi_in_17_ARLEN = in_17__m_axi_m_axi_ARLEN;
  assign m_axi_in_17_ARLOCK = in_17__m_axi_m_axi_ARLOCK;
  assign m_axi_in_17_ARPROT = in_17__m_axi_m_axi_ARPROT;
  assign m_axi_in_17_ARQOS = in_17__m_axi_m_axi_ARQOS;
  assign in_17__m_axi_m_axi_ARREADY = m_axi_in_17_ARREADY;
  assign m_axi_in_17_ARSIZE = in_17__m_axi_m_axi_ARSIZE;
  assign m_axi_in_17_ARVALID = in_17__m_axi_m_axi_ARVALID;
  assign m_axi_in_17_AWADDR = in_17__m_axi_m_axi_AWADDR;
  assign m_axi_in_17_AWBURST = in_17__m_axi_m_axi_AWBURST;
  assign m_axi_in_17_AWCACHE = in_17__m_axi_m_axi_AWCACHE;
  assign m_axi_in_17_AWID = in_17__m_axi_m_axi_AWID;
  assign m_axi_in_17_AWLEN = in_17__m_axi_m_axi_AWLEN;
  assign m_axi_in_17_AWLOCK = in_17__m_axi_m_axi_AWLOCK;
  assign m_axi_in_17_AWPROT = in_17__m_axi_m_axi_AWPROT;
  assign m_axi_in_17_AWQOS = in_17__m_axi_m_axi_AWQOS;
  assign in_17__m_axi_m_axi_AWREADY = m_axi_in_17_AWREADY;
  assign m_axi_in_17_AWSIZE = in_17__m_axi_m_axi_AWSIZE;
  assign m_axi_in_17_AWVALID = in_17__m_axi_m_axi_AWVALID;
  assign in_17__m_axi_m_axi_BID = m_axi_in_17_BID;
  assign m_axi_in_17_BREADY = in_17__m_axi_m_axi_BREADY;
  assign in_17__m_axi_m_axi_BRESP = m_axi_in_17_BRESP;
  assign in_17__m_axi_m_axi_BVALID = m_axi_in_17_BVALID;
  assign in_17__m_axi_m_axi_RDATA = m_axi_in_17_RDATA;
  assign in_17__m_axi_m_axi_RID = m_axi_in_17_RID;
  assign in_17__m_axi_m_axi_RLAST = m_axi_in_17_RLAST;
  assign m_axi_in_17_RREADY = in_17__m_axi_m_axi_RREADY;
  assign in_17__m_axi_m_axi_RRESP = m_axi_in_17_RRESP;
  assign in_17__m_axi_m_axi_RVALID = m_axi_in_17_RVALID;
  assign m_axi_in_17_WDATA = in_17__m_axi_m_axi_WDATA;
  assign m_axi_in_17_WLAST = in_17__m_axi_m_axi_WLAST;
  assign in_17__m_axi_m_axi_WREADY = m_axi_in_17_WREADY;
  assign m_axi_in_17_WSTRB = in_17__m_axi_m_axi_WSTRB;
  assign m_axi_in_17_WVALID = in_17__m_axi_m_axi_WVALID;
  assign in_17__m_axi_read_addr_din = in_17_read_addr__din;
  assign in_17_read_addr__full_n = in_17__m_axi_read_addr_full_n;
  assign in_17__m_axi_read_addr_write = in_17_read_addr__write;
  assign in_17_read_data__dout = in_17__m_axi_read_data_dout;
  assign in_17_read_data__empty_n = in_17__m_axi_read_data_empty_n;
  assign in_17__m_axi_read_data_read = in_17_read_data__read;
  assign in_17__m_axi_rst = ~ ap_rst_n;
  assign in_17__m_axi_write_addr_din = in_17_write_addr__din;
  assign in_17_write_addr__full_n = in_17__m_axi_write_addr_full_n;
  assign in_17__m_axi_write_addr_write = in_17_write_addr__write;
  assign in_17__m_axi_write_data_din = in_17_write_data__din;
  assign in_17_write_data__full_n = in_17__m_axi_write_data_full_n;
  assign in_17__m_axi_write_data_write = in_17_write_data__write;
  assign in_17_write_resp__dout = in_17__m_axi_write_resp_dout;
  assign in_17_write_resp__empty_n = in_17__m_axi_write_resp_empty_n;
  assign in_17__m_axi_write_resp_read = in_17_write_resp__read;
  assign in_18__m_axi_clk = ap_clk;
  assign m_axi_in_18_ARADDR = in_18__m_axi_m_axi_ARADDR;
  assign m_axi_in_18_ARBURST = in_18__m_axi_m_axi_ARBURST;
  assign m_axi_in_18_ARCACHE = in_18__m_axi_m_axi_ARCACHE;
  assign m_axi_in_18_ARID = in_18__m_axi_m_axi_ARID;
  assign m_axi_in_18_ARLEN = in_18__m_axi_m_axi_ARLEN;
  assign m_axi_in_18_ARLOCK = in_18__m_axi_m_axi_ARLOCK;
  assign m_axi_in_18_ARPROT = in_18__m_axi_m_axi_ARPROT;
  assign m_axi_in_18_ARQOS = in_18__m_axi_m_axi_ARQOS;
  assign in_18__m_axi_m_axi_ARREADY = m_axi_in_18_ARREADY;
  assign m_axi_in_18_ARSIZE = in_18__m_axi_m_axi_ARSIZE;
  assign m_axi_in_18_ARVALID = in_18__m_axi_m_axi_ARVALID;
  assign m_axi_in_18_AWADDR = in_18__m_axi_m_axi_AWADDR;
  assign m_axi_in_18_AWBURST = in_18__m_axi_m_axi_AWBURST;
  assign m_axi_in_18_AWCACHE = in_18__m_axi_m_axi_AWCACHE;
  assign m_axi_in_18_AWID = in_18__m_axi_m_axi_AWID;
  assign m_axi_in_18_AWLEN = in_18__m_axi_m_axi_AWLEN;
  assign m_axi_in_18_AWLOCK = in_18__m_axi_m_axi_AWLOCK;
  assign m_axi_in_18_AWPROT = in_18__m_axi_m_axi_AWPROT;
  assign m_axi_in_18_AWQOS = in_18__m_axi_m_axi_AWQOS;
  assign in_18__m_axi_m_axi_AWREADY = m_axi_in_18_AWREADY;
  assign m_axi_in_18_AWSIZE = in_18__m_axi_m_axi_AWSIZE;
  assign m_axi_in_18_AWVALID = in_18__m_axi_m_axi_AWVALID;
  assign in_18__m_axi_m_axi_BID = m_axi_in_18_BID;
  assign m_axi_in_18_BREADY = in_18__m_axi_m_axi_BREADY;
  assign in_18__m_axi_m_axi_BRESP = m_axi_in_18_BRESP;
  assign in_18__m_axi_m_axi_BVALID = m_axi_in_18_BVALID;
  assign in_18__m_axi_m_axi_RDATA = m_axi_in_18_RDATA;
  assign in_18__m_axi_m_axi_RID = m_axi_in_18_RID;
  assign in_18__m_axi_m_axi_RLAST = m_axi_in_18_RLAST;
  assign m_axi_in_18_RREADY = in_18__m_axi_m_axi_RREADY;
  assign in_18__m_axi_m_axi_RRESP = m_axi_in_18_RRESP;
  assign in_18__m_axi_m_axi_RVALID = m_axi_in_18_RVALID;
  assign m_axi_in_18_WDATA = in_18__m_axi_m_axi_WDATA;
  assign m_axi_in_18_WLAST = in_18__m_axi_m_axi_WLAST;
  assign in_18__m_axi_m_axi_WREADY = m_axi_in_18_WREADY;
  assign m_axi_in_18_WSTRB = in_18__m_axi_m_axi_WSTRB;
  assign m_axi_in_18_WVALID = in_18__m_axi_m_axi_WVALID;
  assign in_18__m_axi_read_addr_din = in_18_read_addr__din;
  assign in_18_read_addr__full_n = in_18__m_axi_read_addr_full_n;
  assign in_18__m_axi_read_addr_write = in_18_read_addr__write;
  assign in_18_read_data__dout = in_18__m_axi_read_data_dout;
  assign in_18_read_data__empty_n = in_18__m_axi_read_data_empty_n;
  assign in_18__m_axi_read_data_read = in_18_read_data__read;
  assign in_18__m_axi_rst = ~ ap_rst_n;
  assign in_18__m_axi_write_addr_din = in_18_write_addr__din;
  assign in_18_write_addr__full_n = in_18__m_axi_write_addr_full_n;
  assign in_18__m_axi_write_addr_write = in_18_write_addr__write;
  assign in_18__m_axi_write_data_din = in_18_write_data__din;
  assign in_18_write_data__full_n = in_18__m_axi_write_data_full_n;
  assign in_18__m_axi_write_data_write = in_18_write_data__write;
  assign in_18_write_resp__dout = in_18__m_axi_write_resp_dout;
  assign in_18_write_resp__empty_n = in_18__m_axi_write_resp_empty_n;
  assign in_18__m_axi_write_resp_read = in_18_write_resp__read;
  assign in_19__m_axi_clk = ap_clk;
  assign m_axi_in_19_ARADDR = in_19__m_axi_m_axi_ARADDR;
  assign m_axi_in_19_ARBURST = in_19__m_axi_m_axi_ARBURST;
  assign m_axi_in_19_ARCACHE = in_19__m_axi_m_axi_ARCACHE;
  assign m_axi_in_19_ARID = in_19__m_axi_m_axi_ARID;
  assign m_axi_in_19_ARLEN = in_19__m_axi_m_axi_ARLEN;
  assign m_axi_in_19_ARLOCK = in_19__m_axi_m_axi_ARLOCK;
  assign m_axi_in_19_ARPROT = in_19__m_axi_m_axi_ARPROT;
  assign m_axi_in_19_ARQOS = in_19__m_axi_m_axi_ARQOS;
  assign in_19__m_axi_m_axi_ARREADY = m_axi_in_19_ARREADY;
  assign m_axi_in_19_ARSIZE = in_19__m_axi_m_axi_ARSIZE;
  assign m_axi_in_19_ARVALID = in_19__m_axi_m_axi_ARVALID;
  assign m_axi_in_19_AWADDR = in_19__m_axi_m_axi_AWADDR;
  assign m_axi_in_19_AWBURST = in_19__m_axi_m_axi_AWBURST;
  assign m_axi_in_19_AWCACHE = in_19__m_axi_m_axi_AWCACHE;
  assign m_axi_in_19_AWID = in_19__m_axi_m_axi_AWID;
  assign m_axi_in_19_AWLEN = in_19__m_axi_m_axi_AWLEN;
  assign m_axi_in_19_AWLOCK = in_19__m_axi_m_axi_AWLOCK;
  assign m_axi_in_19_AWPROT = in_19__m_axi_m_axi_AWPROT;
  assign m_axi_in_19_AWQOS = in_19__m_axi_m_axi_AWQOS;
  assign in_19__m_axi_m_axi_AWREADY = m_axi_in_19_AWREADY;
  assign m_axi_in_19_AWSIZE = in_19__m_axi_m_axi_AWSIZE;
  assign m_axi_in_19_AWVALID = in_19__m_axi_m_axi_AWVALID;
  assign in_19__m_axi_m_axi_BID = m_axi_in_19_BID;
  assign m_axi_in_19_BREADY = in_19__m_axi_m_axi_BREADY;
  assign in_19__m_axi_m_axi_BRESP = m_axi_in_19_BRESP;
  assign in_19__m_axi_m_axi_BVALID = m_axi_in_19_BVALID;
  assign in_19__m_axi_m_axi_RDATA = m_axi_in_19_RDATA;
  assign in_19__m_axi_m_axi_RID = m_axi_in_19_RID;
  assign in_19__m_axi_m_axi_RLAST = m_axi_in_19_RLAST;
  assign m_axi_in_19_RREADY = in_19__m_axi_m_axi_RREADY;
  assign in_19__m_axi_m_axi_RRESP = m_axi_in_19_RRESP;
  assign in_19__m_axi_m_axi_RVALID = m_axi_in_19_RVALID;
  assign m_axi_in_19_WDATA = in_19__m_axi_m_axi_WDATA;
  assign m_axi_in_19_WLAST = in_19__m_axi_m_axi_WLAST;
  assign in_19__m_axi_m_axi_WREADY = m_axi_in_19_WREADY;
  assign m_axi_in_19_WSTRB = in_19__m_axi_m_axi_WSTRB;
  assign m_axi_in_19_WVALID = in_19__m_axi_m_axi_WVALID;
  assign in_19__m_axi_read_addr_din = in_19_read_addr__din;
  assign in_19_read_addr__full_n = in_19__m_axi_read_addr_full_n;
  assign in_19__m_axi_read_addr_write = in_19_read_addr__write;
  assign in_19_read_data__dout = in_19__m_axi_read_data_dout;
  assign in_19_read_data__empty_n = in_19__m_axi_read_data_empty_n;
  assign in_19__m_axi_read_data_read = in_19_read_data__read;
  assign in_19__m_axi_rst = ~ ap_rst_n;
  assign in_19__m_axi_write_addr_din = in_19_write_addr__din;
  assign in_19_write_addr__full_n = in_19__m_axi_write_addr_full_n;
  assign in_19__m_axi_write_addr_write = in_19_write_addr__write;
  assign in_19__m_axi_write_data_din = in_19_write_data__din;
  assign in_19_write_data__full_n = in_19__m_axi_write_data_full_n;
  assign in_19__m_axi_write_data_write = in_19_write_data__write;
  assign in_19_write_resp__dout = in_19__m_axi_write_resp_dout;
  assign in_19_write_resp__empty_n = in_19__m_axi_write_resp_empty_n;
  assign in_19__m_axi_write_resp_read = in_19_write_resp__read;
  assign in_2__m_axi_clk = ap_clk;
  assign m_axi_in_2_ARADDR = in_2__m_axi_m_axi_ARADDR;
  assign m_axi_in_2_ARBURST = in_2__m_axi_m_axi_ARBURST;
  assign m_axi_in_2_ARCACHE = in_2__m_axi_m_axi_ARCACHE;
  assign m_axi_in_2_ARID = in_2__m_axi_m_axi_ARID;
  assign m_axi_in_2_ARLEN = in_2__m_axi_m_axi_ARLEN;
  assign m_axi_in_2_ARLOCK = in_2__m_axi_m_axi_ARLOCK;
  assign m_axi_in_2_ARPROT = in_2__m_axi_m_axi_ARPROT;
  assign m_axi_in_2_ARQOS = in_2__m_axi_m_axi_ARQOS;
  assign in_2__m_axi_m_axi_ARREADY = m_axi_in_2_ARREADY;
  assign m_axi_in_2_ARSIZE = in_2__m_axi_m_axi_ARSIZE;
  assign m_axi_in_2_ARVALID = in_2__m_axi_m_axi_ARVALID;
  assign m_axi_in_2_AWADDR = in_2__m_axi_m_axi_AWADDR;
  assign m_axi_in_2_AWBURST = in_2__m_axi_m_axi_AWBURST;
  assign m_axi_in_2_AWCACHE = in_2__m_axi_m_axi_AWCACHE;
  assign m_axi_in_2_AWID = in_2__m_axi_m_axi_AWID;
  assign m_axi_in_2_AWLEN = in_2__m_axi_m_axi_AWLEN;
  assign m_axi_in_2_AWLOCK = in_2__m_axi_m_axi_AWLOCK;
  assign m_axi_in_2_AWPROT = in_2__m_axi_m_axi_AWPROT;
  assign m_axi_in_2_AWQOS = in_2__m_axi_m_axi_AWQOS;
  assign in_2__m_axi_m_axi_AWREADY = m_axi_in_2_AWREADY;
  assign m_axi_in_2_AWSIZE = in_2__m_axi_m_axi_AWSIZE;
  assign m_axi_in_2_AWVALID = in_2__m_axi_m_axi_AWVALID;
  assign in_2__m_axi_m_axi_BID = m_axi_in_2_BID;
  assign m_axi_in_2_BREADY = in_2__m_axi_m_axi_BREADY;
  assign in_2__m_axi_m_axi_BRESP = m_axi_in_2_BRESP;
  assign in_2__m_axi_m_axi_BVALID = m_axi_in_2_BVALID;
  assign in_2__m_axi_m_axi_RDATA = m_axi_in_2_RDATA;
  assign in_2__m_axi_m_axi_RID = m_axi_in_2_RID;
  assign in_2__m_axi_m_axi_RLAST = m_axi_in_2_RLAST;
  assign m_axi_in_2_RREADY = in_2__m_axi_m_axi_RREADY;
  assign in_2__m_axi_m_axi_RRESP = m_axi_in_2_RRESP;
  assign in_2__m_axi_m_axi_RVALID = m_axi_in_2_RVALID;
  assign m_axi_in_2_WDATA = in_2__m_axi_m_axi_WDATA;
  assign m_axi_in_2_WLAST = in_2__m_axi_m_axi_WLAST;
  assign in_2__m_axi_m_axi_WREADY = m_axi_in_2_WREADY;
  assign m_axi_in_2_WSTRB = in_2__m_axi_m_axi_WSTRB;
  assign m_axi_in_2_WVALID = in_2__m_axi_m_axi_WVALID;
  assign in_2__m_axi_read_addr_din = in_2_read_addr__din;
  assign in_2_read_addr__full_n = in_2__m_axi_read_addr_full_n;
  assign in_2__m_axi_read_addr_write = in_2_read_addr__write;
  assign in_2_read_data__dout = in_2__m_axi_read_data_dout;
  assign in_2_read_data__empty_n = in_2__m_axi_read_data_empty_n;
  assign in_2__m_axi_read_data_read = in_2_read_data__read;
  assign in_2__m_axi_rst = ~ ap_rst_n;
  assign in_2__m_axi_write_addr_din = in_2_write_addr__din;
  assign in_2_write_addr__full_n = in_2__m_axi_write_addr_full_n;
  assign in_2__m_axi_write_addr_write = in_2_write_addr__write;
  assign in_2__m_axi_write_data_din = in_2_write_data__din;
  assign in_2_write_data__full_n = in_2__m_axi_write_data_full_n;
  assign in_2__m_axi_write_data_write = in_2_write_data__write;
  assign in_2_write_resp__dout = in_2__m_axi_write_resp_dout;
  assign in_2_write_resp__empty_n = in_2__m_axi_write_resp_empty_n;
  assign in_2__m_axi_write_resp_read = in_2_write_resp__read;
  assign in_20__m_axi_clk = ap_clk;
  assign m_axi_in_20_ARADDR = in_20__m_axi_m_axi_ARADDR;
  assign m_axi_in_20_ARBURST = in_20__m_axi_m_axi_ARBURST;
  assign m_axi_in_20_ARCACHE = in_20__m_axi_m_axi_ARCACHE;
  assign m_axi_in_20_ARID = in_20__m_axi_m_axi_ARID;
  assign m_axi_in_20_ARLEN = in_20__m_axi_m_axi_ARLEN;
  assign m_axi_in_20_ARLOCK = in_20__m_axi_m_axi_ARLOCK;
  assign m_axi_in_20_ARPROT = in_20__m_axi_m_axi_ARPROT;
  assign m_axi_in_20_ARQOS = in_20__m_axi_m_axi_ARQOS;
  assign in_20__m_axi_m_axi_ARREADY = m_axi_in_20_ARREADY;
  assign m_axi_in_20_ARSIZE = in_20__m_axi_m_axi_ARSIZE;
  assign m_axi_in_20_ARVALID = in_20__m_axi_m_axi_ARVALID;
  assign m_axi_in_20_AWADDR = in_20__m_axi_m_axi_AWADDR;
  assign m_axi_in_20_AWBURST = in_20__m_axi_m_axi_AWBURST;
  assign m_axi_in_20_AWCACHE = in_20__m_axi_m_axi_AWCACHE;
  assign m_axi_in_20_AWID = in_20__m_axi_m_axi_AWID;
  assign m_axi_in_20_AWLEN = in_20__m_axi_m_axi_AWLEN;
  assign m_axi_in_20_AWLOCK = in_20__m_axi_m_axi_AWLOCK;
  assign m_axi_in_20_AWPROT = in_20__m_axi_m_axi_AWPROT;
  assign m_axi_in_20_AWQOS = in_20__m_axi_m_axi_AWQOS;
  assign in_20__m_axi_m_axi_AWREADY = m_axi_in_20_AWREADY;
  assign m_axi_in_20_AWSIZE = in_20__m_axi_m_axi_AWSIZE;
  assign m_axi_in_20_AWVALID = in_20__m_axi_m_axi_AWVALID;
  assign in_20__m_axi_m_axi_BID = m_axi_in_20_BID;
  assign m_axi_in_20_BREADY = in_20__m_axi_m_axi_BREADY;
  assign in_20__m_axi_m_axi_BRESP = m_axi_in_20_BRESP;
  assign in_20__m_axi_m_axi_BVALID = m_axi_in_20_BVALID;
  assign in_20__m_axi_m_axi_RDATA = m_axi_in_20_RDATA;
  assign in_20__m_axi_m_axi_RID = m_axi_in_20_RID;
  assign in_20__m_axi_m_axi_RLAST = m_axi_in_20_RLAST;
  assign m_axi_in_20_RREADY = in_20__m_axi_m_axi_RREADY;
  assign in_20__m_axi_m_axi_RRESP = m_axi_in_20_RRESP;
  assign in_20__m_axi_m_axi_RVALID = m_axi_in_20_RVALID;
  assign m_axi_in_20_WDATA = in_20__m_axi_m_axi_WDATA;
  assign m_axi_in_20_WLAST = in_20__m_axi_m_axi_WLAST;
  assign in_20__m_axi_m_axi_WREADY = m_axi_in_20_WREADY;
  assign m_axi_in_20_WSTRB = in_20__m_axi_m_axi_WSTRB;
  assign m_axi_in_20_WVALID = in_20__m_axi_m_axi_WVALID;
  assign in_20__m_axi_read_addr_din = in_20_read_addr__din;
  assign in_20_read_addr__full_n = in_20__m_axi_read_addr_full_n;
  assign in_20__m_axi_read_addr_write = in_20_read_addr__write;
  assign in_20_read_data__dout = in_20__m_axi_read_data_dout;
  assign in_20_read_data__empty_n = in_20__m_axi_read_data_empty_n;
  assign in_20__m_axi_read_data_read = in_20_read_data__read;
  assign in_20__m_axi_rst = ~ ap_rst_n;
  assign in_20__m_axi_write_addr_din = in_20_write_addr__din;
  assign in_20_write_addr__full_n = in_20__m_axi_write_addr_full_n;
  assign in_20__m_axi_write_addr_write = in_20_write_addr__write;
  assign in_20__m_axi_write_data_din = in_20_write_data__din;
  assign in_20_write_data__full_n = in_20__m_axi_write_data_full_n;
  assign in_20__m_axi_write_data_write = in_20_write_data__write;
  assign in_20_write_resp__dout = in_20__m_axi_write_resp_dout;
  assign in_20_write_resp__empty_n = in_20__m_axi_write_resp_empty_n;
  assign in_20__m_axi_write_resp_read = in_20_write_resp__read;
  assign in_21__m_axi_clk = ap_clk;
  assign m_axi_in_21_ARADDR = in_21__m_axi_m_axi_ARADDR;
  assign m_axi_in_21_ARBURST = in_21__m_axi_m_axi_ARBURST;
  assign m_axi_in_21_ARCACHE = in_21__m_axi_m_axi_ARCACHE;
  assign m_axi_in_21_ARID = in_21__m_axi_m_axi_ARID;
  assign m_axi_in_21_ARLEN = in_21__m_axi_m_axi_ARLEN;
  assign m_axi_in_21_ARLOCK = in_21__m_axi_m_axi_ARLOCK;
  assign m_axi_in_21_ARPROT = in_21__m_axi_m_axi_ARPROT;
  assign m_axi_in_21_ARQOS = in_21__m_axi_m_axi_ARQOS;
  assign in_21__m_axi_m_axi_ARREADY = m_axi_in_21_ARREADY;
  assign m_axi_in_21_ARSIZE = in_21__m_axi_m_axi_ARSIZE;
  assign m_axi_in_21_ARVALID = in_21__m_axi_m_axi_ARVALID;
  assign m_axi_in_21_AWADDR = in_21__m_axi_m_axi_AWADDR;
  assign m_axi_in_21_AWBURST = in_21__m_axi_m_axi_AWBURST;
  assign m_axi_in_21_AWCACHE = in_21__m_axi_m_axi_AWCACHE;
  assign m_axi_in_21_AWID = in_21__m_axi_m_axi_AWID;
  assign m_axi_in_21_AWLEN = in_21__m_axi_m_axi_AWLEN;
  assign m_axi_in_21_AWLOCK = in_21__m_axi_m_axi_AWLOCK;
  assign m_axi_in_21_AWPROT = in_21__m_axi_m_axi_AWPROT;
  assign m_axi_in_21_AWQOS = in_21__m_axi_m_axi_AWQOS;
  assign in_21__m_axi_m_axi_AWREADY = m_axi_in_21_AWREADY;
  assign m_axi_in_21_AWSIZE = in_21__m_axi_m_axi_AWSIZE;
  assign m_axi_in_21_AWVALID = in_21__m_axi_m_axi_AWVALID;
  assign in_21__m_axi_m_axi_BID = m_axi_in_21_BID;
  assign m_axi_in_21_BREADY = in_21__m_axi_m_axi_BREADY;
  assign in_21__m_axi_m_axi_BRESP = m_axi_in_21_BRESP;
  assign in_21__m_axi_m_axi_BVALID = m_axi_in_21_BVALID;
  assign in_21__m_axi_m_axi_RDATA = m_axi_in_21_RDATA;
  assign in_21__m_axi_m_axi_RID = m_axi_in_21_RID;
  assign in_21__m_axi_m_axi_RLAST = m_axi_in_21_RLAST;
  assign m_axi_in_21_RREADY = in_21__m_axi_m_axi_RREADY;
  assign in_21__m_axi_m_axi_RRESP = m_axi_in_21_RRESP;
  assign in_21__m_axi_m_axi_RVALID = m_axi_in_21_RVALID;
  assign m_axi_in_21_WDATA = in_21__m_axi_m_axi_WDATA;
  assign m_axi_in_21_WLAST = in_21__m_axi_m_axi_WLAST;
  assign in_21__m_axi_m_axi_WREADY = m_axi_in_21_WREADY;
  assign m_axi_in_21_WSTRB = in_21__m_axi_m_axi_WSTRB;
  assign m_axi_in_21_WVALID = in_21__m_axi_m_axi_WVALID;
  assign in_21__m_axi_read_addr_din = in_21_read_addr__din;
  assign in_21_read_addr__full_n = in_21__m_axi_read_addr_full_n;
  assign in_21__m_axi_read_addr_write = in_21_read_addr__write;
  assign in_21_read_data__dout = in_21__m_axi_read_data_dout;
  assign in_21_read_data__empty_n = in_21__m_axi_read_data_empty_n;
  assign in_21__m_axi_read_data_read = in_21_read_data__read;
  assign in_21__m_axi_rst = ~ ap_rst_n;
  assign in_21__m_axi_write_addr_din = in_21_write_addr__din;
  assign in_21_write_addr__full_n = in_21__m_axi_write_addr_full_n;
  assign in_21__m_axi_write_addr_write = in_21_write_addr__write;
  assign in_21__m_axi_write_data_din = in_21_write_data__din;
  assign in_21_write_data__full_n = in_21__m_axi_write_data_full_n;
  assign in_21__m_axi_write_data_write = in_21_write_data__write;
  assign in_21_write_resp__dout = in_21__m_axi_write_resp_dout;
  assign in_21_write_resp__empty_n = in_21__m_axi_write_resp_empty_n;
  assign in_21__m_axi_write_resp_read = in_21_write_resp__read;
  assign in_22__m_axi_clk = ap_clk;
  assign m_axi_in_22_ARADDR = in_22__m_axi_m_axi_ARADDR;
  assign m_axi_in_22_ARBURST = in_22__m_axi_m_axi_ARBURST;
  assign m_axi_in_22_ARCACHE = in_22__m_axi_m_axi_ARCACHE;
  assign m_axi_in_22_ARID = in_22__m_axi_m_axi_ARID;
  assign m_axi_in_22_ARLEN = in_22__m_axi_m_axi_ARLEN;
  assign m_axi_in_22_ARLOCK = in_22__m_axi_m_axi_ARLOCK;
  assign m_axi_in_22_ARPROT = in_22__m_axi_m_axi_ARPROT;
  assign m_axi_in_22_ARQOS = in_22__m_axi_m_axi_ARQOS;
  assign in_22__m_axi_m_axi_ARREADY = m_axi_in_22_ARREADY;
  assign m_axi_in_22_ARSIZE = in_22__m_axi_m_axi_ARSIZE;
  assign m_axi_in_22_ARVALID = in_22__m_axi_m_axi_ARVALID;
  assign m_axi_in_22_AWADDR = in_22__m_axi_m_axi_AWADDR;
  assign m_axi_in_22_AWBURST = in_22__m_axi_m_axi_AWBURST;
  assign m_axi_in_22_AWCACHE = in_22__m_axi_m_axi_AWCACHE;
  assign m_axi_in_22_AWID = in_22__m_axi_m_axi_AWID;
  assign m_axi_in_22_AWLEN = in_22__m_axi_m_axi_AWLEN;
  assign m_axi_in_22_AWLOCK = in_22__m_axi_m_axi_AWLOCK;
  assign m_axi_in_22_AWPROT = in_22__m_axi_m_axi_AWPROT;
  assign m_axi_in_22_AWQOS = in_22__m_axi_m_axi_AWQOS;
  assign in_22__m_axi_m_axi_AWREADY = m_axi_in_22_AWREADY;
  assign m_axi_in_22_AWSIZE = in_22__m_axi_m_axi_AWSIZE;
  assign m_axi_in_22_AWVALID = in_22__m_axi_m_axi_AWVALID;
  assign in_22__m_axi_m_axi_BID = m_axi_in_22_BID;
  assign m_axi_in_22_BREADY = in_22__m_axi_m_axi_BREADY;
  assign in_22__m_axi_m_axi_BRESP = m_axi_in_22_BRESP;
  assign in_22__m_axi_m_axi_BVALID = m_axi_in_22_BVALID;
  assign in_22__m_axi_m_axi_RDATA = m_axi_in_22_RDATA;
  assign in_22__m_axi_m_axi_RID = m_axi_in_22_RID;
  assign in_22__m_axi_m_axi_RLAST = m_axi_in_22_RLAST;
  assign m_axi_in_22_RREADY = in_22__m_axi_m_axi_RREADY;
  assign in_22__m_axi_m_axi_RRESP = m_axi_in_22_RRESP;
  assign in_22__m_axi_m_axi_RVALID = m_axi_in_22_RVALID;
  assign m_axi_in_22_WDATA = in_22__m_axi_m_axi_WDATA;
  assign m_axi_in_22_WLAST = in_22__m_axi_m_axi_WLAST;
  assign in_22__m_axi_m_axi_WREADY = m_axi_in_22_WREADY;
  assign m_axi_in_22_WSTRB = in_22__m_axi_m_axi_WSTRB;
  assign m_axi_in_22_WVALID = in_22__m_axi_m_axi_WVALID;
  assign in_22__m_axi_read_addr_din = in_22_read_addr__din;
  assign in_22_read_addr__full_n = in_22__m_axi_read_addr_full_n;
  assign in_22__m_axi_read_addr_write = in_22_read_addr__write;
  assign in_22_read_data__dout = in_22__m_axi_read_data_dout;
  assign in_22_read_data__empty_n = in_22__m_axi_read_data_empty_n;
  assign in_22__m_axi_read_data_read = in_22_read_data__read;
  assign in_22__m_axi_rst = ~ ap_rst_n;
  assign in_22__m_axi_write_addr_din = in_22_write_addr__din;
  assign in_22_write_addr__full_n = in_22__m_axi_write_addr_full_n;
  assign in_22__m_axi_write_addr_write = in_22_write_addr__write;
  assign in_22__m_axi_write_data_din = in_22_write_data__din;
  assign in_22_write_data__full_n = in_22__m_axi_write_data_full_n;
  assign in_22__m_axi_write_data_write = in_22_write_data__write;
  assign in_22_write_resp__dout = in_22__m_axi_write_resp_dout;
  assign in_22_write_resp__empty_n = in_22__m_axi_write_resp_empty_n;
  assign in_22__m_axi_write_resp_read = in_22_write_resp__read;
  assign in_23__m_axi_clk = ap_clk;
  assign m_axi_in_23_ARADDR = in_23__m_axi_m_axi_ARADDR;
  assign m_axi_in_23_ARBURST = in_23__m_axi_m_axi_ARBURST;
  assign m_axi_in_23_ARCACHE = in_23__m_axi_m_axi_ARCACHE;
  assign m_axi_in_23_ARID = in_23__m_axi_m_axi_ARID;
  assign m_axi_in_23_ARLEN = in_23__m_axi_m_axi_ARLEN;
  assign m_axi_in_23_ARLOCK = in_23__m_axi_m_axi_ARLOCK;
  assign m_axi_in_23_ARPROT = in_23__m_axi_m_axi_ARPROT;
  assign m_axi_in_23_ARQOS = in_23__m_axi_m_axi_ARQOS;
  assign in_23__m_axi_m_axi_ARREADY = m_axi_in_23_ARREADY;
  assign m_axi_in_23_ARSIZE = in_23__m_axi_m_axi_ARSIZE;
  assign m_axi_in_23_ARVALID = in_23__m_axi_m_axi_ARVALID;
  assign m_axi_in_23_AWADDR = in_23__m_axi_m_axi_AWADDR;
  assign m_axi_in_23_AWBURST = in_23__m_axi_m_axi_AWBURST;
  assign m_axi_in_23_AWCACHE = in_23__m_axi_m_axi_AWCACHE;
  assign m_axi_in_23_AWID = in_23__m_axi_m_axi_AWID;
  assign m_axi_in_23_AWLEN = in_23__m_axi_m_axi_AWLEN;
  assign m_axi_in_23_AWLOCK = in_23__m_axi_m_axi_AWLOCK;
  assign m_axi_in_23_AWPROT = in_23__m_axi_m_axi_AWPROT;
  assign m_axi_in_23_AWQOS = in_23__m_axi_m_axi_AWQOS;
  assign in_23__m_axi_m_axi_AWREADY = m_axi_in_23_AWREADY;
  assign m_axi_in_23_AWSIZE = in_23__m_axi_m_axi_AWSIZE;
  assign m_axi_in_23_AWVALID = in_23__m_axi_m_axi_AWVALID;
  assign in_23__m_axi_m_axi_BID = m_axi_in_23_BID;
  assign m_axi_in_23_BREADY = in_23__m_axi_m_axi_BREADY;
  assign in_23__m_axi_m_axi_BRESP = m_axi_in_23_BRESP;
  assign in_23__m_axi_m_axi_BVALID = m_axi_in_23_BVALID;
  assign in_23__m_axi_m_axi_RDATA = m_axi_in_23_RDATA;
  assign in_23__m_axi_m_axi_RID = m_axi_in_23_RID;
  assign in_23__m_axi_m_axi_RLAST = m_axi_in_23_RLAST;
  assign m_axi_in_23_RREADY = in_23__m_axi_m_axi_RREADY;
  assign in_23__m_axi_m_axi_RRESP = m_axi_in_23_RRESP;
  assign in_23__m_axi_m_axi_RVALID = m_axi_in_23_RVALID;
  assign m_axi_in_23_WDATA = in_23__m_axi_m_axi_WDATA;
  assign m_axi_in_23_WLAST = in_23__m_axi_m_axi_WLAST;
  assign in_23__m_axi_m_axi_WREADY = m_axi_in_23_WREADY;
  assign m_axi_in_23_WSTRB = in_23__m_axi_m_axi_WSTRB;
  assign m_axi_in_23_WVALID = in_23__m_axi_m_axi_WVALID;
  assign in_23__m_axi_read_addr_din = in_23_read_addr__din;
  assign in_23_read_addr__full_n = in_23__m_axi_read_addr_full_n;
  assign in_23__m_axi_read_addr_write = in_23_read_addr__write;
  assign in_23_read_data__dout = in_23__m_axi_read_data_dout;
  assign in_23_read_data__empty_n = in_23__m_axi_read_data_empty_n;
  assign in_23__m_axi_read_data_read = in_23_read_data__read;
  assign in_23__m_axi_rst = ~ ap_rst_n;
  assign in_23__m_axi_write_addr_din = in_23_write_addr__din;
  assign in_23_write_addr__full_n = in_23__m_axi_write_addr_full_n;
  assign in_23__m_axi_write_addr_write = in_23_write_addr__write;
  assign in_23__m_axi_write_data_din = in_23_write_data__din;
  assign in_23_write_data__full_n = in_23__m_axi_write_data_full_n;
  assign in_23__m_axi_write_data_write = in_23_write_data__write;
  assign in_23_write_resp__dout = in_23__m_axi_write_resp_dout;
  assign in_23_write_resp__empty_n = in_23__m_axi_write_resp_empty_n;
  assign in_23__m_axi_write_resp_read = in_23_write_resp__read;
  assign in_24__m_axi_clk = ap_clk;
  assign m_axi_in_24_ARADDR = in_24__m_axi_m_axi_ARADDR;
  assign m_axi_in_24_ARBURST = in_24__m_axi_m_axi_ARBURST;
  assign m_axi_in_24_ARCACHE = in_24__m_axi_m_axi_ARCACHE;
  assign m_axi_in_24_ARID = in_24__m_axi_m_axi_ARID;
  assign m_axi_in_24_ARLEN = in_24__m_axi_m_axi_ARLEN;
  assign m_axi_in_24_ARLOCK = in_24__m_axi_m_axi_ARLOCK;
  assign m_axi_in_24_ARPROT = in_24__m_axi_m_axi_ARPROT;
  assign m_axi_in_24_ARQOS = in_24__m_axi_m_axi_ARQOS;
  assign in_24__m_axi_m_axi_ARREADY = m_axi_in_24_ARREADY;
  assign m_axi_in_24_ARSIZE = in_24__m_axi_m_axi_ARSIZE;
  assign m_axi_in_24_ARVALID = in_24__m_axi_m_axi_ARVALID;
  assign m_axi_in_24_AWADDR = in_24__m_axi_m_axi_AWADDR;
  assign m_axi_in_24_AWBURST = in_24__m_axi_m_axi_AWBURST;
  assign m_axi_in_24_AWCACHE = in_24__m_axi_m_axi_AWCACHE;
  assign m_axi_in_24_AWID = in_24__m_axi_m_axi_AWID;
  assign m_axi_in_24_AWLEN = in_24__m_axi_m_axi_AWLEN;
  assign m_axi_in_24_AWLOCK = in_24__m_axi_m_axi_AWLOCK;
  assign m_axi_in_24_AWPROT = in_24__m_axi_m_axi_AWPROT;
  assign m_axi_in_24_AWQOS = in_24__m_axi_m_axi_AWQOS;
  assign in_24__m_axi_m_axi_AWREADY = m_axi_in_24_AWREADY;
  assign m_axi_in_24_AWSIZE = in_24__m_axi_m_axi_AWSIZE;
  assign m_axi_in_24_AWVALID = in_24__m_axi_m_axi_AWVALID;
  assign in_24__m_axi_m_axi_BID = m_axi_in_24_BID;
  assign m_axi_in_24_BREADY = in_24__m_axi_m_axi_BREADY;
  assign in_24__m_axi_m_axi_BRESP = m_axi_in_24_BRESP;
  assign in_24__m_axi_m_axi_BVALID = m_axi_in_24_BVALID;
  assign in_24__m_axi_m_axi_RDATA = m_axi_in_24_RDATA;
  assign in_24__m_axi_m_axi_RID = m_axi_in_24_RID;
  assign in_24__m_axi_m_axi_RLAST = m_axi_in_24_RLAST;
  assign m_axi_in_24_RREADY = in_24__m_axi_m_axi_RREADY;
  assign in_24__m_axi_m_axi_RRESP = m_axi_in_24_RRESP;
  assign in_24__m_axi_m_axi_RVALID = m_axi_in_24_RVALID;
  assign m_axi_in_24_WDATA = in_24__m_axi_m_axi_WDATA;
  assign m_axi_in_24_WLAST = in_24__m_axi_m_axi_WLAST;
  assign in_24__m_axi_m_axi_WREADY = m_axi_in_24_WREADY;
  assign m_axi_in_24_WSTRB = in_24__m_axi_m_axi_WSTRB;
  assign m_axi_in_24_WVALID = in_24__m_axi_m_axi_WVALID;
  assign in_24__m_axi_read_addr_din = in_24_read_addr__din;
  assign in_24_read_addr__full_n = in_24__m_axi_read_addr_full_n;
  assign in_24__m_axi_read_addr_write = in_24_read_addr__write;
  assign in_24_read_data__dout = in_24__m_axi_read_data_dout;
  assign in_24_read_data__empty_n = in_24__m_axi_read_data_empty_n;
  assign in_24__m_axi_read_data_read = in_24_read_data__read;
  assign in_24__m_axi_rst = ~ ap_rst_n;
  assign in_24__m_axi_write_addr_din = in_24_write_addr__din;
  assign in_24_write_addr__full_n = in_24__m_axi_write_addr_full_n;
  assign in_24__m_axi_write_addr_write = in_24_write_addr__write;
  assign in_24__m_axi_write_data_din = in_24_write_data__din;
  assign in_24_write_data__full_n = in_24__m_axi_write_data_full_n;
  assign in_24__m_axi_write_data_write = in_24_write_data__write;
  assign in_24_write_resp__dout = in_24__m_axi_write_resp_dout;
  assign in_24_write_resp__empty_n = in_24__m_axi_write_resp_empty_n;
  assign in_24__m_axi_write_resp_read = in_24_write_resp__read;
  assign in_25__m_axi_clk = ap_clk;
  assign m_axi_in_25_ARADDR = in_25__m_axi_m_axi_ARADDR;
  assign m_axi_in_25_ARBURST = in_25__m_axi_m_axi_ARBURST;
  assign m_axi_in_25_ARCACHE = in_25__m_axi_m_axi_ARCACHE;
  assign m_axi_in_25_ARID = in_25__m_axi_m_axi_ARID;
  assign m_axi_in_25_ARLEN = in_25__m_axi_m_axi_ARLEN;
  assign m_axi_in_25_ARLOCK = in_25__m_axi_m_axi_ARLOCK;
  assign m_axi_in_25_ARPROT = in_25__m_axi_m_axi_ARPROT;
  assign m_axi_in_25_ARQOS = in_25__m_axi_m_axi_ARQOS;
  assign in_25__m_axi_m_axi_ARREADY = m_axi_in_25_ARREADY;
  assign m_axi_in_25_ARSIZE = in_25__m_axi_m_axi_ARSIZE;
  assign m_axi_in_25_ARVALID = in_25__m_axi_m_axi_ARVALID;
  assign m_axi_in_25_AWADDR = in_25__m_axi_m_axi_AWADDR;
  assign m_axi_in_25_AWBURST = in_25__m_axi_m_axi_AWBURST;
  assign m_axi_in_25_AWCACHE = in_25__m_axi_m_axi_AWCACHE;
  assign m_axi_in_25_AWID = in_25__m_axi_m_axi_AWID;
  assign m_axi_in_25_AWLEN = in_25__m_axi_m_axi_AWLEN;
  assign m_axi_in_25_AWLOCK = in_25__m_axi_m_axi_AWLOCK;
  assign m_axi_in_25_AWPROT = in_25__m_axi_m_axi_AWPROT;
  assign m_axi_in_25_AWQOS = in_25__m_axi_m_axi_AWQOS;
  assign in_25__m_axi_m_axi_AWREADY = m_axi_in_25_AWREADY;
  assign m_axi_in_25_AWSIZE = in_25__m_axi_m_axi_AWSIZE;
  assign m_axi_in_25_AWVALID = in_25__m_axi_m_axi_AWVALID;
  assign in_25__m_axi_m_axi_BID = m_axi_in_25_BID;
  assign m_axi_in_25_BREADY = in_25__m_axi_m_axi_BREADY;
  assign in_25__m_axi_m_axi_BRESP = m_axi_in_25_BRESP;
  assign in_25__m_axi_m_axi_BVALID = m_axi_in_25_BVALID;
  assign in_25__m_axi_m_axi_RDATA = m_axi_in_25_RDATA;
  assign in_25__m_axi_m_axi_RID = m_axi_in_25_RID;
  assign in_25__m_axi_m_axi_RLAST = m_axi_in_25_RLAST;
  assign m_axi_in_25_RREADY = in_25__m_axi_m_axi_RREADY;
  assign in_25__m_axi_m_axi_RRESP = m_axi_in_25_RRESP;
  assign in_25__m_axi_m_axi_RVALID = m_axi_in_25_RVALID;
  assign m_axi_in_25_WDATA = in_25__m_axi_m_axi_WDATA;
  assign m_axi_in_25_WLAST = in_25__m_axi_m_axi_WLAST;
  assign in_25__m_axi_m_axi_WREADY = m_axi_in_25_WREADY;
  assign m_axi_in_25_WSTRB = in_25__m_axi_m_axi_WSTRB;
  assign m_axi_in_25_WVALID = in_25__m_axi_m_axi_WVALID;
  assign in_25__m_axi_read_addr_din = in_25_read_addr__din;
  assign in_25_read_addr__full_n = in_25__m_axi_read_addr_full_n;
  assign in_25__m_axi_read_addr_write = in_25_read_addr__write;
  assign in_25_read_data__dout = in_25__m_axi_read_data_dout;
  assign in_25_read_data__empty_n = in_25__m_axi_read_data_empty_n;
  assign in_25__m_axi_read_data_read = in_25_read_data__read;
  assign in_25__m_axi_rst = ~ ap_rst_n;
  assign in_25__m_axi_write_addr_din = in_25_write_addr__din;
  assign in_25_write_addr__full_n = in_25__m_axi_write_addr_full_n;
  assign in_25__m_axi_write_addr_write = in_25_write_addr__write;
  assign in_25__m_axi_write_data_din = in_25_write_data__din;
  assign in_25_write_data__full_n = in_25__m_axi_write_data_full_n;
  assign in_25__m_axi_write_data_write = in_25_write_data__write;
  assign in_25_write_resp__dout = in_25__m_axi_write_resp_dout;
  assign in_25_write_resp__empty_n = in_25__m_axi_write_resp_empty_n;
  assign in_25__m_axi_write_resp_read = in_25_write_resp__read;
  assign in_26__m_axi_clk = ap_clk;
  assign m_axi_in_26_ARADDR = in_26__m_axi_m_axi_ARADDR;
  assign m_axi_in_26_ARBURST = in_26__m_axi_m_axi_ARBURST;
  assign m_axi_in_26_ARCACHE = in_26__m_axi_m_axi_ARCACHE;
  assign m_axi_in_26_ARID = in_26__m_axi_m_axi_ARID;
  assign m_axi_in_26_ARLEN = in_26__m_axi_m_axi_ARLEN;
  assign m_axi_in_26_ARLOCK = in_26__m_axi_m_axi_ARLOCK;
  assign m_axi_in_26_ARPROT = in_26__m_axi_m_axi_ARPROT;
  assign m_axi_in_26_ARQOS = in_26__m_axi_m_axi_ARQOS;
  assign in_26__m_axi_m_axi_ARREADY = m_axi_in_26_ARREADY;
  assign m_axi_in_26_ARSIZE = in_26__m_axi_m_axi_ARSIZE;
  assign m_axi_in_26_ARVALID = in_26__m_axi_m_axi_ARVALID;
  assign m_axi_in_26_AWADDR = in_26__m_axi_m_axi_AWADDR;
  assign m_axi_in_26_AWBURST = in_26__m_axi_m_axi_AWBURST;
  assign m_axi_in_26_AWCACHE = in_26__m_axi_m_axi_AWCACHE;
  assign m_axi_in_26_AWID = in_26__m_axi_m_axi_AWID;
  assign m_axi_in_26_AWLEN = in_26__m_axi_m_axi_AWLEN;
  assign m_axi_in_26_AWLOCK = in_26__m_axi_m_axi_AWLOCK;
  assign m_axi_in_26_AWPROT = in_26__m_axi_m_axi_AWPROT;
  assign m_axi_in_26_AWQOS = in_26__m_axi_m_axi_AWQOS;
  assign in_26__m_axi_m_axi_AWREADY = m_axi_in_26_AWREADY;
  assign m_axi_in_26_AWSIZE = in_26__m_axi_m_axi_AWSIZE;
  assign m_axi_in_26_AWVALID = in_26__m_axi_m_axi_AWVALID;
  assign in_26__m_axi_m_axi_BID = m_axi_in_26_BID;
  assign m_axi_in_26_BREADY = in_26__m_axi_m_axi_BREADY;
  assign in_26__m_axi_m_axi_BRESP = m_axi_in_26_BRESP;
  assign in_26__m_axi_m_axi_BVALID = m_axi_in_26_BVALID;
  assign in_26__m_axi_m_axi_RDATA = m_axi_in_26_RDATA;
  assign in_26__m_axi_m_axi_RID = m_axi_in_26_RID;
  assign in_26__m_axi_m_axi_RLAST = m_axi_in_26_RLAST;
  assign m_axi_in_26_RREADY = in_26__m_axi_m_axi_RREADY;
  assign in_26__m_axi_m_axi_RRESP = m_axi_in_26_RRESP;
  assign in_26__m_axi_m_axi_RVALID = m_axi_in_26_RVALID;
  assign m_axi_in_26_WDATA = in_26__m_axi_m_axi_WDATA;
  assign m_axi_in_26_WLAST = in_26__m_axi_m_axi_WLAST;
  assign in_26__m_axi_m_axi_WREADY = m_axi_in_26_WREADY;
  assign m_axi_in_26_WSTRB = in_26__m_axi_m_axi_WSTRB;
  assign m_axi_in_26_WVALID = in_26__m_axi_m_axi_WVALID;
  assign in_26__m_axi_read_addr_din = in_26_read_addr__din;
  assign in_26_read_addr__full_n = in_26__m_axi_read_addr_full_n;
  assign in_26__m_axi_read_addr_write = in_26_read_addr__write;
  assign in_26_read_data__dout = in_26__m_axi_read_data_dout;
  assign in_26_read_data__empty_n = in_26__m_axi_read_data_empty_n;
  assign in_26__m_axi_read_data_read = in_26_read_data__read;
  assign in_26__m_axi_rst = ~ ap_rst_n;
  assign in_26__m_axi_write_addr_din = in_26_write_addr__din;
  assign in_26_write_addr__full_n = in_26__m_axi_write_addr_full_n;
  assign in_26__m_axi_write_addr_write = in_26_write_addr__write;
  assign in_26__m_axi_write_data_din = in_26_write_data__din;
  assign in_26_write_data__full_n = in_26__m_axi_write_data_full_n;
  assign in_26__m_axi_write_data_write = in_26_write_data__write;
  assign in_26_write_resp__dout = in_26__m_axi_write_resp_dout;
  assign in_26_write_resp__empty_n = in_26__m_axi_write_resp_empty_n;
  assign in_26__m_axi_write_resp_read = in_26_write_resp__read;
  assign in_3__m_axi_clk = ap_clk;
  assign m_axi_in_3_ARADDR = in_3__m_axi_m_axi_ARADDR;
  assign m_axi_in_3_ARBURST = in_3__m_axi_m_axi_ARBURST;
  assign m_axi_in_3_ARCACHE = in_3__m_axi_m_axi_ARCACHE;
  assign m_axi_in_3_ARID = in_3__m_axi_m_axi_ARID;
  assign m_axi_in_3_ARLEN = in_3__m_axi_m_axi_ARLEN;
  assign m_axi_in_3_ARLOCK = in_3__m_axi_m_axi_ARLOCK;
  assign m_axi_in_3_ARPROT = in_3__m_axi_m_axi_ARPROT;
  assign m_axi_in_3_ARQOS = in_3__m_axi_m_axi_ARQOS;
  assign in_3__m_axi_m_axi_ARREADY = m_axi_in_3_ARREADY;
  assign m_axi_in_3_ARSIZE = in_3__m_axi_m_axi_ARSIZE;
  assign m_axi_in_3_ARVALID = in_3__m_axi_m_axi_ARVALID;
  assign m_axi_in_3_AWADDR = in_3__m_axi_m_axi_AWADDR;
  assign m_axi_in_3_AWBURST = in_3__m_axi_m_axi_AWBURST;
  assign m_axi_in_3_AWCACHE = in_3__m_axi_m_axi_AWCACHE;
  assign m_axi_in_3_AWID = in_3__m_axi_m_axi_AWID;
  assign m_axi_in_3_AWLEN = in_3__m_axi_m_axi_AWLEN;
  assign m_axi_in_3_AWLOCK = in_3__m_axi_m_axi_AWLOCK;
  assign m_axi_in_3_AWPROT = in_3__m_axi_m_axi_AWPROT;
  assign m_axi_in_3_AWQOS = in_3__m_axi_m_axi_AWQOS;
  assign in_3__m_axi_m_axi_AWREADY = m_axi_in_3_AWREADY;
  assign m_axi_in_3_AWSIZE = in_3__m_axi_m_axi_AWSIZE;
  assign m_axi_in_3_AWVALID = in_3__m_axi_m_axi_AWVALID;
  assign in_3__m_axi_m_axi_BID = m_axi_in_3_BID;
  assign m_axi_in_3_BREADY = in_3__m_axi_m_axi_BREADY;
  assign in_3__m_axi_m_axi_BRESP = m_axi_in_3_BRESP;
  assign in_3__m_axi_m_axi_BVALID = m_axi_in_3_BVALID;
  assign in_3__m_axi_m_axi_RDATA = m_axi_in_3_RDATA;
  assign in_3__m_axi_m_axi_RID = m_axi_in_3_RID;
  assign in_3__m_axi_m_axi_RLAST = m_axi_in_3_RLAST;
  assign m_axi_in_3_RREADY = in_3__m_axi_m_axi_RREADY;
  assign in_3__m_axi_m_axi_RRESP = m_axi_in_3_RRESP;
  assign in_3__m_axi_m_axi_RVALID = m_axi_in_3_RVALID;
  assign m_axi_in_3_WDATA = in_3__m_axi_m_axi_WDATA;
  assign m_axi_in_3_WLAST = in_3__m_axi_m_axi_WLAST;
  assign in_3__m_axi_m_axi_WREADY = m_axi_in_3_WREADY;
  assign m_axi_in_3_WSTRB = in_3__m_axi_m_axi_WSTRB;
  assign m_axi_in_3_WVALID = in_3__m_axi_m_axi_WVALID;
  assign in_3__m_axi_read_addr_din = in_3_read_addr__din;
  assign in_3_read_addr__full_n = in_3__m_axi_read_addr_full_n;
  assign in_3__m_axi_read_addr_write = in_3_read_addr__write;
  assign in_3_read_data__dout = in_3__m_axi_read_data_dout;
  assign in_3_read_data__empty_n = in_3__m_axi_read_data_empty_n;
  assign in_3__m_axi_read_data_read = in_3_read_data__read;
  assign in_3__m_axi_rst = ~ ap_rst_n;
  assign in_3__m_axi_write_addr_din = in_3_write_addr__din;
  assign in_3_write_addr__full_n = in_3__m_axi_write_addr_full_n;
  assign in_3__m_axi_write_addr_write = in_3_write_addr__write;
  assign in_3__m_axi_write_data_din = in_3_write_data__din;
  assign in_3_write_data__full_n = in_3__m_axi_write_data_full_n;
  assign in_3__m_axi_write_data_write = in_3_write_data__write;
  assign in_3_write_resp__dout = in_3__m_axi_write_resp_dout;
  assign in_3_write_resp__empty_n = in_3__m_axi_write_resp_empty_n;
  assign in_3__m_axi_write_resp_read = in_3_write_resp__read;
  assign in_4__m_axi_clk = ap_clk;
  assign m_axi_in_4_ARADDR = in_4__m_axi_m_axi_ARADDR;
  assign m_axi_in_4_ARBURST = in_4__m_axi_m_axi_ARBURST;
  assign m_axi_in_4_ARCACHE = in_4__m_axi_m_axi_ARCACHE;
  assign m_axi_in_4_ARID = in_4__m_axi_m_axi_ARID;
  assign m_axi_in_4_ARLEN = in_4__m_axi_m_axi_ARLEN;
  assign m_axi_in_4_ARLOCK = in_4__m_axi_m_axi_ARLOCK;
  assign m_axi_in_4_ARPROT = in_4__m_axi_m_axi_ARPROT;
  assign m_axi_in_4_ARQOS = in_4__m_axi_m_axi_ARQOS;
  assign in_4__m_axi_m_axi_ARREADY = m_axi_in_4_ARREADY;
  assign m_axi_in_4_ARSIZE = in_4__m_axi_m_axi_ARSIZE;
  assign m_axi_in_4_ARVALID = in_4__m_axi_m_axi_ARVALID;
  assign m_axi_in_4_AWADDR = in_4__m_axi_m_axi_AWADDR;
  assign m_axi_in_4_AWBURST = in_4__m_axi_m_axi_AWBURST;
  assign m_axi_in_4_AWCACHE = in_4__m_axi_m_axi_AWCACHE;
  assign m_axi_in_4_AWID = in_4__m_axi_m_axi_AWID;
  assign m_axi_in_4_AWLEN = in_4__m_axi_m_axi_AWLEN;
  assign m_axi_in_4_AWLOCK = in_4__m_axi_m_axi_AWLOCK;
  assign m_axi_in_4_AWPROT = in_4__m_axi_m_axi_AWPROT;
  assign m_axi_in_4_AWQOS = in_4__m_axi_m_axi_AWQOS;
  assign in_4__m_axi_m_axi_AWREADY = m_axi_in_4_AWREADY;
  assign m_axi_in_4_AWSIZE = in_4__m_axi_m_axi_AWSIZE;
  assign m_axi_in_4_AWVALID = in_4__m_axi_m_axi_AWVALID;
  assign in_4__m_axi_m_axi_BID = m_axi_in_4_BID;
  assign m_axi_in_4_BREADY = in_4__m_axi_m_axi_BREADY;
  assign in_4__m_axi_m_axi_BRESP = m_axi_in_4_BRESP;
  assign in_4__m_axi_m_axi_BVALID = m_axi_in_4_BVALID;
  assign in_4__m_axi_m_axi_RDATA = m_axi_in_4_RDATA;
  assign in_4__m_axi_m_axi_RID = m_axi_in_4_RID;
  assign in_4__m_axi_m_axi_RLAST = m_axi_in_4_RLAST;
  assign m_axi_in_4_RREADY = in_4__m_axi_m_axi_RREADY;
  assign in_4__m_axi_m_axi_RRESP = m_axi_in_4_RRESP;
  assign in_4__m_axi_m_axi_RVALID = m_axi_in_4_RVALID;
  assign m_axi_in_4_WDATA = in_4__m_axi_m_axi_WDATA;
  assign m_axi_in_4_WLAST = in_4__m_axi_m_axi_WLAST;
  assign in_4__m_axi_m_axi_WREADY = m_axi_in_4_WREADY;
  assign m_axi_in_4_WSTRB = in_4__m_axi_m_axi_WSTRB;
  assign m_axi_in_4_WVALID = in_4__m_axi_m_axi_WVALID;
  assign in_4__m_axi_read_addr_din = in_4_read_addr__din;
  assign in_4_read_addr__full_n = in_4__m_axi_read_addr_full_n;
  assign in_4__m_axi_read_addr_write = in_4_read_addr__write;
  assign in_4_read_data__dout = in_4__m_axi_read_data_dout;
  assign in_4_read_data__empty_n = in_4__m_axi_read_data_empty_n;
  assign in_4__m_axi_read_data_read = in_4_read_data__read;
  assign in_4__m_axi_rst = ~ ap_rst_n;
  assign in_4__m_axi_write_addr_din = in_4_write_addr__din;
  assign in_4_write_addr__full_n = in_4__m_axi_write_addr_full_n;
  assign in_4__m_axi_write_addr_write = in_4_write_addr__write;
  assign in_4__m_axi_write_data_din = in_4_write_data__din;
  assign in_4_write_data__full_n = in_4__m_axi_write_data_full_n;
  assign in_4__m_axi_write_data_write = in_4_write_data__write;
  assign in_4_write_resp__dout = in_4__m_axi_write_resp_dout;
  assign in_4_write_resp__empty_n = in_4__m_axi_write_resp_empty_n;
  assign in_4__m_axi_write_resp_read = in_4_write_resp__read;
  assign in_5__m_axi_clk = ap_clk;
  assign m_axi_in_5_ARADDR = in_5__m_axi_m_axi_ARADDR;
  assign m_axi_in_5_ARBURST = in_5__m_axi_m_axi_ARBURST;
  assign m_axi_in_5_ARCACHE = in_5__m_axi_m_axi_ARCACHE;
  assign m_axi_in_5_ARID = in_5__m_axi_m_axi_ARID;
  assign m_axi_in_5_ARLEN = in_5__m_axi_m_axi_ARLEN;
  assign m_axi_in_5_ARLOCK = in_5__m_axi_m_axi_ARLOCK;
  assign m_axi_in_5_ARPROT = in_5__m_axi_m_axi_ARPROT;
  assign m_axi_in_5_ARQOS = in_5__m_axi_m_axi_ARQOS;
  assign in_5__m_axi_m_axi_ARREADY = m_axi_in_5_ARREADY;
  assign m_axi_in_5_ARSIZE = in_5__m_axi_m_axi_ARSIZE;
  assign m_axi_in_5_ARVALID = in_5__m_axi_m_axi_ARVALID;
  assign m_axi_in_5_AWADDR = in_5__m_axi_m_axi_AWADDR;
  assign m_axi_in_5_AWBURST = in_5__m_axi_m_axi_AWBURST;
  assign m_axi_in_5_AWCACHE = in_5__m_axi_m_axi_AWCACHE;
  assign m_axi_in_5_AWID = in_5__m_axi_m_axi_AWID;
  assign m_axi_in_5_AWLEN = in_5__m_axi_m_axi_AWLEN;
  assign m_axi_in_5_AWLOCK = in_5__m_axi_m_axi_AWLOCK;
  assign m_axi_in_5_AWPROT = in_5__m_axi_m_axi_AWPROT;
  assign m_axi_in_5_AWQOS = in_5__m_axi_m_axi_AWQOS;
  assign in_5__m_axi_m_axi_AWREADY = m_axi_in_5_AWREADY;
  assign m_axi_in_5_AWSIZE = in_5__m_axi_m_axi_AWSIZE;
  assign m_axi_in_5_AWVALID = in_5__m_axi_m_axi_AWVALID;
  assign in_5__m_axi_m_axi_BID = m_axi_in_5_BID;
  assign m_axi_in_5_BREADY = in_5__m_axi_m_axi_BREADY;
  assign in_5__m_axi_m_axi_BRESP = m_axi_in_5_BRESP;
  assign in_5__m_axi_m_axi_BVALID = m_axi_in_5_BVALID;
  assign in_5__m_axi_m_axi_RDATA = m_axi_in_5_RDATA;
  assign in_5__m_axi_m_axi_RID = m_axi_in_5_RID;
  assign in_5__m_axi_m_axi_RLAST = m_axi_in_5_RLAST;
  assign m_axi_in_5_RREADY = in_5__m_axi_m_axi_RREADY;
  assign in_5__m_axi_m_axi_RRESP = m_axi_in_5_RRESP;
  assign in_5__m_axi_m_axi_RVALID = m_axi_in_5_RVALID;
  assign m_axi_in_5_WDATA = in_5__m_axi_m_axi_WDATA;
  assign m_axi_in_5_WLAST = in_5__m_axi_m_axi_WLAST;
  assign in_5__m_axi_m_axi_WREADY = m_axi_in_5_WREADY;
  assign m_axi_in_5_WSTRB = in_5__m_axi_m_axi_WSTRB;
  assign m_axi_in_5_WVALID = in_5__m_axi_m_axi_WVALID;
  assign in_5__m_axi_read_addr_din = in_5_read_addr__din;
  assign in_5_read_addr__full_n = in_5__m_axi_read_addr_full_n;
  assign in_5__m_axi_read_addr_write = in_5_read_addr__write;
  assign in_5_read_data__dout = in_5__m_axi_read_data_dout;
  assign in_5_read_data__empty_n = in_5__m_axi_read_data_empty_n;
  assign in_5__m_axi_read_data_read = in_5_read_data__read;
  assign in_5__m_axi_rst = ~ ap_rst_n;
  assign in_5__m_axi_write_addr_din = in_5_write_addr__din;
  assign in_5_write_addr__full_n = in_5__m_axi_write_addr_full_n;
  assign in_5__m_axi_write_addr_write = in_5_write_addr__write;
  assign in_5__m_axi_write_data_din = in_5_write_data__din;
  assign in_5_write_data__full_n = in_5__m_axi_write_data_full_n;
  assign in_5__m_axi_write_data_write = in_5_write_data__write;
  assign in_5_write_resp__dout = in_5__m_axi_write_resp_dout;
  assign in_5_write_resp__empty_n = in_5__m_axi_write_resp_empty_n;
  assign in_5__m_axi_write_resp_read = in_5_write_resp__read;
  assign in_6__m_axi_clk = ap_clk;
  assign m_axi_in_6_ARADDR = in_6__m_axi_m_axi_ARADDR;
  assign m_axi_in_6_ARBURST = in_6__m_axi_m_axi_ARBURST;
  assign m_axi_in_6_ARCACHE = in_6__m_axi_m_axi_ARCACHE;
  assign m_axi_in_6_ARID = in_6__m_axi_m_axi_ARID;
  assign m_axi_in_6_ARLEN = in_6__m_axi_m_axi_ARLEN;
  assign m_axi_in_6_ARLOCK = in_6__m_axi_m_axi_ARLOCK;
  assign m_axi_in_6_ARPROT = in_6__m_axi_m_axi_ARPROT;
  assign m_axi_in_6_ARQOS = in_6__m_axi_m_axi_ARQOS;
  assign in_6__m_axi_m_axi_ARREADY = m_axi_in_6_ARREADY;
  assign m_axi_in_6_ARSIZE = in_6__m_axi_m_axi_ARSIZE;
  assign m_axi_in_6_ARVALID = in_6__m_axi_m_axi_ARVALID;
  assign m_axi_in_6_AWADDR = in_6__m_axi_m_axi_AWADDR;
  assign m_axi_in_6_AWBURST = in_6__m_axi_m_axi_AWBURST;
  assign m_axi_in_6_AWCACHE = in_6__m_axi_m_axi_AWCACHE;
  assign m_axi_in_6_AWID = in_6__m_axi_m_axi_AWID;
  assign m_axi_in_6_AWLEN = in_6__m_axi_m_axi_AWLEN;
  assign m_axi_in_6_AWLOCK = in_6__m_axi_m_axi_AWLOCK;
  assign m_axi_in_6_AWPROT = in_6__m_axi_m_axi_AWPROT;
  assign m_axi_in_6_AWQOS = in_6__m_axi_m_axi_AWQOS;
  assign in_6__m_axi_m_axi_AWREADY = m_axi_in_6_AWREADY;
  assign m_axi_in_6_AWSIZE = in_6__m_axi_m_axi_AWSIZE;
  assign m_axi_in_6_AWVALID = in_6__m_axi_m_axi_AWVALID;
  assign in_6__m_axi_m_axi_BID = m_axi_in_6_BID;
  assign m_axi_in_6_BREADY = in_6__m_axi_m_axi_BREADY;
  assign in_6__m_axi_m_axi_BRESP = m_axi_in_6_BRESP;
  assign in_6__m_axi_m_axi_BVALID = m_axi_in_6_BVALID;
  assign in_6__m_axi_m_axi_RDATA = m_axi_in_6_RDATA;
  assign in_6__m_axi_m_axi_RID = m_axi_in_6_RID;
  assign in_6__m_axi_m_axi_RLAST = m_axi_in_6_RLAST;
  assign m_axi_in_6_RREADY = in_6__m_axi_m_axi_RREADY;
  assign in_6__m_axi_m_axi_RRESP = m_axi_in_6_RRESP;
  assign in_6__m_axi_m_axi_RVALID = m_axi_in_6_RVALID;
  assign m_axi_in_6_WDATA = in_6__m_axi_m_axi_WDATA;
  assign m_axi_in_6_WLAST = in_6__m_axi_m_axi_WLAST;
  assign in_6__m_axi_m_axi_WREADY = m_axi_in_6_WREADY;
  assign m_axi_in_6_WSTRB = in_6__m_axi_m_axi_WSTRB;
  assign m_axi_in_6_WVALID = in_6__m_axi_m_axi_WVALID;
  assign in_6__m_axi_read_addr_din = in_6_read_addr__din;
  assign in_6_read_addr__full_n = in_6__m_axi_read_addr_full_n;
  assign in_6__m_axi_read_addr_write = in_6_read_addr__write;
  assign in_6_read_data__dout = in_6__m_axi_read_data_dout;
  assign in_6_read_data__empty_n = in_6__m_axi_read_data_empty_n;
  assign in_6__m_axi_read_data_read = in_6_read_data__read;
  assign in_6__m_axi_rst = ~ ap_rst_n;
  assign in_6__m_axi_write_addr_din = in_6_write_addr__din;
  assign in_6_write_addr__full_n = in_6__m_axi_write_addr_full_n;
  assign in_6__m_axi_write_addr_write = in_6_write_addr__write;
  assign in_6__m_axi_write_data_din = in_6_write_data__din;
  assign in_6_write_data__full_n = in_6__m_axi_write_data_full_n;
  assign in_6__m_axi_write_data_write = in_6_write_data__write;
  assign in_6_write_resp__dout = in_6__m_axi_write_resp_dout;
  assign in_6_write_resp__empty_n = in_6__m_axi_write_resp_empty_n;
  assign in_6__m_axi_write_resp_read = in_6_write_resp__read;
  assign in_7__m_axi_clk = ap_clk;
  assign m_axi_in_7_ARADDR = in_7__m_axi_m_axi_ARADDR;
  assign m_axi_in_7_ARBURST = in_7__m_axi_m_axi_ARBURST;
  assign m_axi_in_7_ARCACHE = in_7__m_axi_m_axi_ARCACHE;
  assign m_axi_in_7_ARID = in_7__m_axi_m_axi_ARID;
  assign m_axi_in_7_ARLEN = in_7__m_axi_m_axi_ARLEN;
  assign m_axi_in_7_ARLOCK = in_7__m_axi_m_axi_ARLOCK;
  assign m_axi_in_7_ARPROT = in_7__m_axi_m_axi_ARPROT;
  assign m_axi_in_7_ARQOS = in_7__m_axi_m_axi_ARQOS;
  assign in_7__m_axi_m_axi_ARREADY = m_axi_in_7_ARREADY;
  assign m_axi_in_7_ARSIZE = in_7__m_axi_m_axi_ARSIZE;
  assign m_axi_in_7_ARVALID = in_7__m_axi_m_axi_ARVALID;
  assign m_axi_in_7_AWADDR = in_7__m_axi_m_axi_AWADDR;
  assign m_axi_in_7_AWBURST = in_7__m_axi_m_axi_AWBURST;
  assign m_axi_in_7_AWCACHE = in_7__m_axi_m_axi_AWCACHE;
  assign m_axi_in_7_AWID = in_7__m_axi_m_axi_AWID;
  assign m_axi_in_7_AWLEN = in_7__m_axi_m_axi_AWLEN;
  assign m_axi_in_7_AWLOCK = in_7__m_axi_m_axi_AWLOCK;
  assign m_axi_in_7_AWPROT = in_7__m_axi_m_axi_AWPROT;
  assign m_axi_in_7_AWQOS = in_7__m_axi_m_axi_AWQOS;
  assign in_7__m_axi_m_axi_AWREADY = m_axi_in_7_AWREADY;
  assign m_axi_in_7_AWSIZE = in_7__m_axi_m_axi_AWSIZE;
  assign m_axi_in_7_AWVALID = in_7__m_axi_m_axi_AWVALID;
  assign in_7__m_axi_m_axi_BID = m_axi_in_7_BID;
  assign m_axi_in_7_BREADY = in_7__m_axi_m_axi_BREADY;
  assign in_7__m_axi_m_axi_BRESP = m_axi_in_7_BRESP;
  assign in_7__m_axi_m_axi_BVALID = m_axi_in_7_BVALID;
  assign in_7__m_axi_m_axi_RDATA = m_axi_in_7_RDATA;
  assign in_7__m_axi_m_axi_RID = m_axi_in_7_RID;
  assign in_7__m_axi_m_axi_RLAST = m_axi_in_7_RLAST;
  assign m_axi_in_7_RREADY = in_7__m_axi_m_axi_RREADY;
  assign in_7__m_axi_m_axi_RRESP = m_axi_in_7_RRESP;
  assign in_7__m_axi_m_axi_RVALID = m_axi_in_7_RVALID;
  assign m_axi_in_7_WDATA = in_7__m_axi_m_axi_WDATA;
  assign m_axi_in_7_WLAST = in_7__m_axi_m_axi_WLAST;
  assign in_7__m_axi_m_axi_WREADY = m_axi_in_7_WREADY;
  assign m_axi_in_7_WSTRB = in_7__m_axi_m_axi_WSTRB;
  assign m_axi_in_7_WVALID = in_7__m_axi_m_axi_WVALID;
  assign in_7__m_axi_read_addr_din = in_7_read_addr__din;
  assign in_7_read_addr__full_n = in_7__m_axi_read_addr_full_n;
  assign in_7__m_axi_read_addr_write = in_7_read_addr__write;
  assign in_7_read_data__dout = in_7__m_axi_read_data_dout;
  assign in_7_read_data__empty_n = in_7__m_axi_read_data_empty_n;
  assign in_7__m_axi_read_data_read = in_7_read_data__read;
  assign in_7__m_axi_rst = ~ ap_rst_n;
  assign in_7__m_axi_write_addr_din = in_7_write_addr__din;
  assign in_7_write_addr__full_n = in_7__m_axi_write_addr_full_n;
  assign in_7__m_axi_write_addr_write = in_7_write_addr__write;
  assign in_7__m_axi_write_data_din = in_7_write_data__din;
  assign in_7_write_data__full_n = in_7__m_axi_write_data_full_n;
  assign in_7__m_axi_write_data_write = in_7_write_data__write;
  assign in_7_write_resp__dout = in_7__m_axi_write_resp_dout;
  assign in_7_write_resp__empty_n = in_7__m_axi_write_resp_empty_n;
  assign in_7__m_axi_write_resp_read = in_7_write_resp__read;
  assign in_8__m_axi_clk = ap_clk;
  assign m_axi_in_8_ARADDR = in_8__m_axi_m_axi_ARADDR;
  assign m_axi_in_8_ARBURST = in_8__m_axi_m_axi_ARBURST;
  assign m_axi_in_8_ARCACHE = in_8__m_axi_m_axi_ARCACHE;
  assign m_axi_in_8_ARID = in_8__m_axi_m_axi_ARID;
  assign m_axi_in_8_ARLEN = in_8__m_axi_m_axi_ARLEN;
  assign m_axi_in_8_ARLOCK = in_8__m_axi_m_axi_ARLOCK;
  assign m_axi_in_8_ARPROT = in_8__m_axi_m_axi_ARPROT;
  assign m_axi_in_8_ARQOS = in_8__m_axi_m_axi_ARQOS;
  assign in_8__m_axi_m_axi_ARREADY = m_axi_in_8_ARREADY;
  assign m_axi_in_8_ARSIZE = in_8__m_axi_m_axi_ARSIZE;
  assign m_axi_in_8_ARVALID = in_8__m_axi_m_axi_ARVALID;
  assign m_axi_in_8_AWADDR = in_8__m_axi_m_axi_AWADDR;
  assign m_axi_in_8_AWBURST = in_8__m_axi_m_axi_AWBURST;
  assign m_axi_in_8_AWCACHE = in_8__m_axi_m_axi_AWCACHE;
  assign m_axi_in_8_AWID = in_8__m_axi_m_axi_AWID;
  assign m_axi_in_8_AWLEN = in_8__m_axi_m_axi_AWLEN;
  assign m_axi_in_8_AWLOCK = in_8__m_axi_m_axi_AWLOCK;
  assign m_axi_in_8_AWPROT = in_8__m_axi_m_axi_AWPROT;
  assign m_axi_in_8_AWQOS = in_8__m_axi_m_axi_AWQOS;
  assign in_8__m_axi_m_axi_AWREADY = m_axi_in_8_AWREADY;
  assign m_axi_in_8_AWSIZE = in_8__m_axi_m_axi_AWSIZE;
  assign m_axi_in_8_AWVALID = in_8__m_axi_m_axi_AWVALID;
  assign in_8__m_axi_m_axi_BID = m_axi_in_8_BID;
  assign m_axi_in_8_BREADY = in_8__m_axi_m_axi_BREADY;
  assign in_8__m_axi_m_axi_BRESP = m_axi_in_8_BRESP;
  assign in_8__m_axi_m_axi_BVALID = m_axi_in_8_BVALID;
  assign in_8__m_axi_m_axi_RDATA = m_axi_in_8_RDATA;
  assign in_8__m_axi_m_axi_RID = m_axi_in_8_RID;
  assign in_8__m_axi_m_axi_RLAST = m_axi_in_8_RLAST;
  assign m_axi_in_8_RREADY = in_8__m_axi_m_axi_RREADY;
  assign in_8__m_axi_m_axi_RRESP = m_axi_in_8_RRESP;
  assign in_8__m_axi_m_axi_RVALID = m_axi_in_8_RVALID;
  assign m_axi_in_8_WDATA = in_8__m_axi_m_axi_WDATA;
  assign m_axi_in_8_WLAST = in_8__m_axi_m_axi_WLAST;
  assign in_8__m_axi_m_axi_WREADY = m_axi_in_8_WREADY;
  assign m_axi_in_8_WSTRB = in_8__m_axi_m_axi_WSTRB;
  assign m_axi_in_8_WVALID = in_8__m_axi_m_axi_WVALID;
  assign in_8__m_axi_read_addr_din = in_8_read_addr__din;
  assign in_8_read_addr__full_n = in_8__m_axi_read_addr_full_n;
  assign in_8__m_axi_read_addr_write = in_8_read_addr__write;
  assign in_8_read_data__dout = in_8__m_axi_read_data_dout;
  assign in_8_read_data__empty_n = in_8__m_axi_read_data_empty_n;
  assign in_8__m_axi_read_data_read = in_8_read_data__read;
  assign in_8__m_axi_rst = ~ ap_rst_n;
  assign in_8__m_axi_write_addr_din = in_8_write_addr__din;
  assign in_8_write_addr__full_n = in_8__m_axi_write_addr_full_n;
  assign in_8__m_axi_write_addr_write = in_8_write_addr__write;
  assign in_8__m_axi_write_data_din = in_8_write_data__din;
  assign in_8_write_data__full_n = in_8__m_axi_write_data_full_n;
  assign in_8__m_axi_write_data_write = in_8_write_data__write;
  assign in_8_write_resp__dout = in_8__m_axi_write_resp_dout;
  assign in_8_write_resp__empty_n = in_8__m_axi_write_resp_empty_n;
  assign in_8__m_axi_write_resp_read = in_8_write_resp__read;
  assign in_9__m_axi_clk = ap_clk;
  assign m_axi_in_9_ARADDR = in_9__m_axi_m_axi_ARADDR;
  assign m_axi_in_9_ARBURST = in_9__m_axi_m_axi_ARBURST;
  assign m_axi_in_9_ARCACHE = in_9__m_axi_m_axi_ARCACHE;
  assign m_axi_in_9_ARID = in_9__m_axi_m_axi_ARID;
  assign m_axi_in_9_ARLEN = in_9__m_axi_m_axi_ARLEN;
  assign m_axi_in_9_ARLOCK = in_9__m_axi_m_axi_ARLOCK;
  assign m_axi_in_9_ARPROT = in_9__m_axi_m_axi_ARPROT;
  assign m_axi_in_9_ARQOS = in_9__m_axi_m_axi_ARQOS;
  assign in_9__m_axi_m_axi_ARREADY = m_axi_in_9_ARREADY;
  assign m_axi_in_9_ARSIZE = in_9__m_axi_m_axi_ARSIZE;
  assign m_axi_in_9_ARVALID = in_9__m_axi_m_axi_ARVALID;
  assign m_axi_in_9_AWADDR = in_9__m_axi_m_axi_AWADDR;
  assign m_axi_in_9_AWBURST = in_9__m_axi_m_axi_AWBURST;
  assign m_axi_in_9_AWCACHE = in_9__m_axi_m_axi_AWCACHE;
  assign m_axi_in_9_AWID = in_9__m_axi_m_axi_AWID;
  assign m_axi_in_9_AWLEN = in_9__m_axi_m_axi_AWLEN;
  assign m_axi_in_9_AWLOCK = in_9__m_axi_m_axi_AWLOCK;
  assign m_axi_in_9_AWPROT = in_9__m_axi_m_axi_AWPROT;
  assign m_axi_in_9_AWQOS = in_9__m_axi_m_axi_AWQOS;
  assign in_9__m_axi_m_axi_AWREADY = m_axi_in_9_AWREADY;
  assign m_axi_in_9_AWSIZE = in_9__m_axi_m_axi_AWSIZE;
  assign m_axi_in_9_AWVALID = in_9__m_axi_m_axi_AWVALID;
  assign in_9__m_axi_m_axi_BID = m_axi_in_9_BID;
  assign m_axi_in_9_BREADY = in_9__m_axi_m_axi_BREADY;
  assign in_9__m_axi_m_axi_BRESP = m_axi_in_9_BRESP;
  assign in_9__m_axi_m_axi_BVALID = m_axi_in_9_BVALID;
  assign in_9__m_axi_m_axi_RDATA = m_axi_in_9_RDATA;
  assign in_9__m_axi_m_axi_RID = m_axi_in_9_RID;
  assign in_9__m_axi_m_axi_RLAST = m_axi_in_9_RLAST;
  assign m_axi_in_9_RREADY = in_9__m_axi_m_axi_RREADY;
  assign in_9__m_axi_m_axi_RRESP = m_axi_in_9_RRESP;
  assign in_9__m_axi_m_axi_RVALID = m_axi_in_9_RVALID;
  assign m_axi_in_9_WDATA = in_9__m_axi_m_axi_WDATA;
  assign m_axi_in_9_WLAST = in_9__m_axi_m_axi_WLAST;
  assign in_9__m_axi_m_axi_WREADY = m_axi_in_9_WREADY;
  assign m_axi_in_9_WSTRB = in_9__m_axi_m_axi_WSTRB;
  assign m_axi_in_9_WVALID = in_9__m_axi_m_axi_WVALID;
  assign in_9__m_axi_read_addr_din = in_9_read_addr__din;
  assign in_9_read_addr__full_n = in_9__m_axi_read_addr_full_n;
  assign in_9__m_axi_read_addr_write = in_9_read_addr__write;
  assign in_9_read_data__dout = in_9__m_axi_read_data_dout;
  assign in_9_read_data__empty_n = in_9__m_axi_read_data_empty_n;
  assign in_9__m_axi_read_data_read = in_9_read_data__read;
  assign in_9__m_axi_rst = ~ ap_rst_n;
  assign in_9__m_axi_write_addr_din = in_9_write_addr__din;
  assign in_9_write_addr__full_n = in_9__m_axi_write_addr_full_n;
  assign in_9__m_axi_write_addr_write = in_9_write_addr__write;
  assign in_9__m_axi_write_data_din = in_9_write_data__din;
  assign in_9_write_data__full_n = in_9__m_axi_write_data_full_n;
  assign in_9__m_axi_write_data_write = in_9_write_data__write;
  assign in_9_write_resp__dout = in_9__m_axi_write_resp_dout;
  assign in_9_write_resp__empty_n = in_9__m_axi_write_resp_empty_n;
  assign in_9__m_axi_write_resp_read = in_9_write_resp__read;
  assign __tapa_fsm_unit_L3_out_dist = L3_out_dist;
  assign __tapa_fsm_unit_L3_out_id = L3_out_id;
  assign __tapa_fsm_unit_ap_clk = ap_clk;
  assign ap_done = __tapa_fsm_unit_ap_done;
  assign ap_idle = __tapa_fsm_unit_ap_idle;
  assign ap_ready = __tapa_fsm_unit_ap_ready;
  assign __tapa_fsm_unit_ap_rst_n = ap_rst_n;
  assign __tapa_fsm_unit_ap_start = ap_start;
  assign __tapa_fsm_unit_in_0 = in_0;
  assign __tapa_fsm_unit_in_1 = in_1;
  assign __tapa_fsm_unit_in_10 = in_10;
  assign __tapa_fsm_unit_in_11 = in_11;
  assign __tapa_fsm_unit_in_12 = in_12;
  assign __tapa_fsm_unit_in_13 = in_13;
  assign __tapa_fsm_unit_in_14 = in_14;
  assign __tapa_fsm_unit_in_15 = in_15;
  assign __tapa_fsm_unit_in_16 = in_16;
  assign __tapa_fsm_unit_in_17 = in_17;
  assign __tapa_fsm_unit_in_18 = in_18;
  assign __tapa_fsm_unit_in_19 = in_19;
  assign __tapa_fsm_unit_in_2 = in_2;
  assign __tapa_fsm_unit_in_20 = in_20;
  assign __tapa_fsm_unit_in_21 = in_21;
  assign __tapa_fsm_unit_in_22 = in_22;
  assign __tapa_fsm_unit_in_23 = in_23;
  assign __tapa_fsm_unit_in_24 = in_24;
  assign __tapa_fsm_unit_in_25 = in_25;
  assign __tapa_fsm_unit_in_26 = in_26;
  assign __tapa_fsm_unit_in_3 = in_3;
  assign __tapa_fsm_unit_in_4 = in_4;
  assign __tapa_fsm_unit_in_5 = in_5;
  assign __tapa_fsm_unit_in_6 = in_6;
  assign __tapa_fsm_unit_in_7 = in_7;
  assign __tapa_fsm_unit_in_8 = in_8;
  assign __tapa_fsm_unit_in_9 = in_9;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_0__ap_done = krnl_globalSort_L1_L2_0__ap_done;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_0__ap_idle = krnl_globalSort_L1_L2_0__ap_idle;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_0__ap_ready = krnl_globalSort_L1_L2_0__ap_ready;
  assign krnl_globalSort_L1_L2_0__ap_start = __tapa_fsm_unit_krnl_globalSort_L1_L2_0__ap_start;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_10__ap_done = krnl_globalSort_L1_L2_10__ap_done;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_10__ap_idle = krnl_globalSort_L1_L2_10__ap_idle;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_10__ap_ready = krnl_globalSort_L1_L2_10__ap_ready;
  assign krnl_globalSort_L1_L2_10__ap_start = __tapa_fsm_unit_krnl_globalSort_L1_L2_10__ap_start;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_11__ap_done = krnl_globalSort_L1_L2_11__ap_done;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_11__ap_idle = krnl_globalSort_L1_L2_11__ap_idle;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_11__ap_ready = krnl_globalSort_L1_L2_11__ap_ready;
  assign krnl_globalSort_L1_L2_11__ap_start = __tapa_fsm_unit_krnl_globalSort_L1_L2_11__ap_start;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_12__ap_done = krnl_globalSort_L1_L2_12__ap_done;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_12__ap_idle = krnl_globalSort_L1_L2_12__ap_idle;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_12__ap_ready = krnl_globalSort_L1_L2_12__ap_ready;
  assign krnl_globalSort_L1_L2_12__ap_start = __tapa_fsm_unit_krnl_globalSort_L1_L2_12__ap_start;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_1__ap_done = krnl_globalSort_L1_L2_1__ap_done;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_1__ap_idle = krnl_globalSort_L1_L2_1__ap_idle;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_1__ap_ready = krnl_globalSort_L1_L2_1__ap_ready;
  assign krnl_globalSort_L1_L2_1__ap_start = __tapa_fsm_unit_krnl_globalSort_L1_L2_1__ap_start;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_2__ap_done = krnl_globalSort_L1_L2_2__ap_done;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_2__ap_idle = krnl_globalSort_L1_L2_2__ap_idle;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_2__ap_ready = krnl_globalSort_L1_L2_2__ap_ready;
  assign krnl_globalSort_L1_L2_2__ap_start = __tapa_fsm_unit_krnl_globalSort_L1_L2_2__ap_start;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_3__ap_done = krnl_globalSort_L1_L2_3__ap_done;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_3__ap_idle = krnl_globalSort_L1_L2_3__ap_idle;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_3__ap_ready = krnl_globalSort_L1_L2_3__ap_ready;
  assign krnl_globalSort_L1_L2_3__ap_start = __tapa_fsm_unit_krnl_globalSort_L1_L2_3__ap_start;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_4__ap_done = krnl_globalSort_L1_L2_4__ap_done;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_4__ap_idle = krnl_globalSort_L1_L2_4__ap_idle;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_4__ap_ready = krnl_globalSort_L1_L2_4__ap_ready;
  assign krnl_globalSort_L1_L2_4__ap_start = __tapa_fsm_unit_krnl_globalSort_L1_L2_4__ap_start;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_5__ap_done = krnl_globalSort_L1_L2_5__ap_done;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_5__ap_idle = krnl_globalSort_L1_L2_5__ap_idle;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_5__ap_ready = krnl_globalSort_L1_L2_5__ap_ready;
  assign krnl_globalSort_L1_L2_5__ap_start = __tapa_fsm_unit_krnl_globalSort_L1_L2_5__ap_start;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_6__ap_done = krnl_globalSort_L1_L2_6__ap_done;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_6__ap_idle = krnl_globalSort_L1_L2_6__ap_idle;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_6__ap_ready = krnl_globalSort_L1_L2_6__ap_ready;
  assign krnl_globalSort_L1_L2_6__ap_start = __tapa_fsm_unit_krnl_globalSort_L1_L2_6__ap_start;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_7__ap_done = krnl_globalSort_L1_L2_7__ap_done;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_7__ap_idle = krnl_globalSort_L1_L2_7__ap_idle;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_7__ap_ready = krnl_globalSort_L1_L2_7__ap_ready;
  assign krnl_globalSort_L1_L2_7__ap_start = __tapa_fsm_unit_krnl_globalSort_L1_L2_7__ap_start;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_8__ap_done = krnl_globalSort_L1_L2_8__ap_done;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_8__ap_idle = krnl_globalSort_L1_L2_8__ap_idle;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_8__ap_ready = krnl_globalSort_L1_L2_8__ap_ready;
  assign krnl_globalSort_L1_L2_8__ap_start = __tapa_fsm_unit_krnl_globalSort_L1_L2_8__ap_start;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_9__ap_done = krnl_globalSort_L1_L2_9__ap_done;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_9__ap_idle = krnl_globalSort_L1_L2_9__ap_idle;
  assign __tapa_fsm_unit_krnl_globalSort_L1_L2_9__ap_ready = krnl_globalSort_L1_L2_9__ap_ready;
  assign krnl_globalSort_L1_L2_9__ap_start = __tapa_fsm_unit_krnl_globalSort_L1_L2_9__ap_start;
  assign krnl_output_dist_id_0___L3_out_dist__q0 = __tapa_fsm_unit_krnl_output_dist_id_0___L3_out_dist__q0;
  assign krnl_output_dist_id_0___L3_out_id__q0 = __tapa_fsm_unit_krnl_output_dist_id_0___L3_out_id__q0;
  assign __tapa_fsm_unit_krnl_output_dist_id_0__ap_done = krnl_output_dist_id_0__ap_done;
  assign __tapa_fsm_unit_krnl_output_dist_id_0__ap_idle = krnl_output_dist_id_0__ap_idle;
  assign __tapa_fsm_unit_krnl_output_dist_id_0__ap_ready = krnl_output_dist_id_0__ap_ready;
  assign krnl_output_dist_id_0__ap_start = __tapa_fsm_unit_krnl_output_dist_id_0__ap_start;
  assign krnl_partialKnn_wrapper_0_0___in_0__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_0_0___in_0__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_0_0__ap_done = krnl_partialKnn_wrapper_0_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_0_0__ap_idle = krnl_partialKnn_wrapper_0_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_0_0__ap_ready = krnl_partialKnn_wrapper_0_0__ap_ready;
  assign krnl_partialKnn_wrapper_0_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_0_0__ap_start;
  assign krnl_partialKnn_wrapper_10_0___in_10__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_10_0___in_10__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_10_0__ap_done = krnl_partialKnn_wrapper_10_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_10_0__ap_idle = krnl_partialKnn_wrapper_10_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_10_0__ap_ready = krnl_partialKnn_wrapper_10_0__ap_ready;
  assign krnl_partialKnn_wrapper_10_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_10_0__ap_start;
  assign krnl_partialKnn_wrapper_11_0___in_11__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_11_0___in_11__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_11_0__ap_done = krnl_partialKnn_wrapper_11_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_11_0__ap_idle = krnl_partialKnn_wrapper_11_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_11_0__ap_ready = krnl_partialKnn_wrapper_11_0__ap_ready;
  assign krnl_partialKnn_wrapper_11_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_11_0__ap_start;
  assign krnl_partialKnn_wrapper_12_0___in_12__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_12_0___in_12__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_12_0__ap_done = krnl_partialKnn_wrapper_12_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_12_0__ap_idle = krnl_partialKnn_wrapper_12_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_12_0__ap_ready = krnl_partialKnn_wrapper_12_0__ap_ready;
  assign krnl_partialKnn_wrapper_12_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_12_0__ap_start;
  assign krnl_partialKnn_wrapper_13_0___in_13__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_13_0___in_13__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_13_0__ap_done = krnl_partialKnn_wrapper_13_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_13_0__ap_idle = krnl_partialKnn_wrapper_13_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_13_0__ap_ready = krnl_partialKnn_wrapper_13_0__ap_ready;
  assign krnl_partialKnn_wrapper_13_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_13_0__ap_start;
  assign krnl_partialKnn_wrapper_14_0___in_14__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_14_0___in_14__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_14_0__ap_done = krnl_partialKnn_wrapper_14_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_14_0__ap_idle = krnl_partialKnn_wrapper_14_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_14_0__ap_ready = krnl_partialKnn_wrapper_14_0__ap_ready;
  assign krnl_partialKnn_wrapper_14_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_14_0__ap_start;
  assign krnl_partialKnn_wrapper_15_0___in_15__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_15_0___in_15__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_15_0__ap_done = krnl_partialKnn_wrapper_15_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_15_0__ap_idle = krnl_partialKnn_wrapper_15_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_15_0__ap_ready = krnl_partialKnn_wrapper_15_0__ap_ready;
  assign krnl_partialKnn_wrapper_15_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_15_0__ap_start;
  assign krnl_partialKnn_wrapper_16_0___in_16__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_16_0___in_16__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_16_0__ap_done = krnl_partialKnn_wrapper_16_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_16_0__ap_idle = krnl_partialKnn_wrapper_16_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_16_0__ap_ready = krnl_partialKnn_wrapper_16_0__ap_ready;
  assign krnl_partialKnn_wrapper_16_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_16_0__ap_start;
  assign krnl_partialKnn_wrapper_17_0___in_17__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_17_0___in_17__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_17_0__ap_done = krnl_partialKnn_wrapper_17_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_17_0__ap_idle = krnl_partialKnn_wrapper_17_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_17_0__ap_ready = krnl_partialKnn_wrapper_17_0__ap_ready;
  assign krnl_partialKnn_wrapper_17_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_17_0__ap_start;
  assign krnl_partialKnn_wrapper_18_0___in_18__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_18_0___in_18__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_18_0__ap_done = krnl_partialKnn_wrapper_18_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_18_0__ap_idle = krnl_partialKnn_wrapper_18_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_18_0__ap_ready = krnl_partialKnn_wrapper_18_0__ap_ready;
  assign krnl_partialKnn_wrapper_18_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_18_0__ap_start;
  assign krnl_partialKnn_wrapper_19_0___in_19__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_19_0___in_19__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_19_0__ap_done = krnl_partialKnn_wrapper_19_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_19_0__ap_idle = krnl_partialKnn_wrapper_19_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_19_0__ap_ready = krnl_partialKnn_wrapper_19_0__ap_ready;
  assign krnl_partialKnn_wrapper_19_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_19_0__ap_start;
  assign krnl_partialKnn_wrapper_1_0___in_1__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_1_0___in_1__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_1_0__ap_done = krnl_partialKnn_wrapper_1_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_1_0__ap_idle = krnl_partialKnn_wrapper_1_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_1_0__ap_ready = krnl_partialKnn_wrapper_1_0__ap_ready;
  assign krnl_partialKnn_wrapper_1_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_1_0__ap_start;
  assign krnl_partialKnn_wrapper_20_0___in_20__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_20_0___in_20__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_20_0__ap_done = krnl_partialKnn_wrapper_20_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_20_0__ap_idle = krnl_partialKnn_wrapper_20_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_20_0__ap_ready = krnl_partialKnn_wrapper_20_0__ap_ready;
  assign krnl_partialKnn_wrapper_20_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_20_0__ap_start;
  assign krnl_partialKnn_wrapper_21_0___in_21__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_21_0___in_21__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_21_0__ap_done = krnl_partialKnn_wrapper_21_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_21_0__ap_idle = krnl_partialKnn_wrapper_21_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_21_0__ap_ready = krnl_partialKnn_wrapper_21_0__ap_ready;
  assign krnl_partialKnn_wrapper_21_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_21_0__ap_start;
  assign krnl_partialKnn_wrapper_22_0___in_22__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_22_0___in_22__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_22_0__ap_done = krnl_partialKnn_wrapper_22_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_22_0__ap_idle = krnl_partialKnn_wrapper_22_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_22_0__ap_ready = krnl_partialKnn_wrapper_22_0__ap_ready;
  assign krnl_partialKnn_wrapper_22_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_22_0__ap_start;
  assign krnl_partialKnn_wrapper_23_0___in_23__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_23_0___in_23__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_23_0__ap_done = krnl_partialKnn_wrapper_23_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_23_0__ap_idle = krnl_partialKnn_wrapper_23_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_23_0__ap_ready = krnl_partialKnn_wrapper_23_0__ap_ready;
  assign krnl_partialKnn_wrapper_23_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_23_0__ap_start;
  assign krnl_partialKnn_wrapper_24_0___in_24__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_24_0___in_24__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_24_0__ap_done = krnl_partialKnn_wrapper_24_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_24_0__ap_idle = krnl_partialKnn_wrapper_24_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_24_0__ap_ready = krnl_partialKnn_wrapper_24_0__ap_ready;
  assign krnl_partialKnn_wrapper_24_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_24_0__ap_start;
  assign krnl_partialKnn_wrapper_25_0___in_25__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_25_0___in_25__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_25_0__ap_done = krnl_partialKnn_wrapper_25_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_25_0__ap_idle = krnl_partialKnn_wrapper_25_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_25_0__ap_ready = krnl_partialKnn_wrapper_25_0__ap_ready;
  assign krnl_partialKnn_wrapper_25_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_25_0__ap_start;
  assign krnl_partialKnn_wrapper_26_0___in_26__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_26_0___in_26__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_26_0__ap_done = krnl_partialKnn_wrapper_26_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_26_0__ap_idle = krnl_partialKnn_wrapper_26_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_26_0__ap_ready = krnl_partialKnn_wrapper_26_0__ap_ready;
  assign krnl_partialKnn_wrapper_26_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_26_0__ap_start;
  assign krnl_partialKnn_wrapper_2_0___in_2__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_2_0___in_2__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_2_0__ap_done = krnl_partialKnn_wrapper_2_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_2_0__ap_idle = krnl_partialKnn_wrapper_2_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_2_0__ap_ready = krnl_partialKnn_wrapper_2_0__ap_ready;
  assign krnl_partialKnn_wrapper_2_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_2_0__ap_start;
  assign krnl_partialKnn_wrapper_3_0___in_3__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_3_0___in_3__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_3_0__ap_done = krnl_partialKnn_wrapper_3_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_3_0__ap_idle = krnl_partialKnn_wrapper_3_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_3_0__ap_ready = krnl_partialKnn_wrapper_3_0__ap_ready;
  assign krnl_partialKnn_wrapper_3_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_3_0__ap_start;
  assign krnl_partialKnn_wrapper_4_0___in_4__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_4_0___in_4__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_4_0__ap_done = krnl_partialKnn_wrapper_4_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_4_0__ap_idle = krnl_partialKnn_wrapper_4_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_4_0__ap_ready = krnl_partialKnn_wrapper_4_0__ap_ready;
  assign krnl_partialKnn_wrapper_4_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_4_0__ap_start;
  assign krnl_partialKnn_wrapper_5_0___in_5__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_5_0___in_5__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_5_0__ap_done = krnl_partialKnn_wrapper_5_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_5_0__ap_idle = krnl_partialKnn_wrapper_5_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_5_0__ap_ready = krnl_partialKnn_wrapper_5_0__ap_ready;
  assign krnl_partialKnn_wrapper_5_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_5_0__ap_start;
  assign krnl_partialKnn_wrapper_6_0___in_6__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_6_0___in_6__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_6_0__ap_done = krnl_partialKnn_wrapper_6_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_6_0__ap_idle = krnl_partialKnn_wrapper_6_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_6_0__ap_ready = krnl_partialKnn_wrapper_6_0__ap_ready;
  assign krnl_partialKnn_wrapper_6_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_6_0__ap_start;
  assign krnl_partialKnn_wrapper_7_0___in_7__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_7_0___in_7__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_7_0__ap_done = krnl_partialKnn_wrapper_7_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_7_0__ap_idle = krnl_partialKnn_wrapper_7_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_7_0__ap_ready = krnl_partialKnn_wrapper_7_0__ap_ready;
  assign krnl_partialKnn_wrapper_7_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_7_0__ap_start;
  assign krnl_partialKnn_wrapper_8_0___in_8__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_8_0___in_8__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_8_0__ap_done = krnl_partialKnn_wrapper_8_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_8_0__ap_idle = krnl_partialKnn_wrapper_8_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_8_0__ap_ready = krnl_partialKnn_wrapper_8_0__ap_ready;
  assign krnl_partialKnn_wrapper_8_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_8_0__ap_start;
  assign krnl_partialKnn_wrapper_9_0___in_9__q0 = __tapa_fsm_unit_krnl_partialKnn_wrapper_9_0___in_9__q0;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_9_0__ap_done = krnl_partialKnn_wrapper_9_0__ap_done;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_9_0__ap_idle = krnl_partialKnn_wrapper_9_0__ap_idle;
  assign __tapa_fsm_unit_krnl_partialKnn_wrapper_9_0__ap_ready = krnl_partialKnn_wrapper_9_0__ap_ready;
  assign krnl_partialKnn_wrapper_9_0__ap_start = __tapa_fsm_unit_krnl_partialKnn_wrapper_9_0__ap_start;
endmodule