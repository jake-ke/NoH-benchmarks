

module Serpens_fsm
(
  ap_clk,
  ap_rst_n,
  ap_start,
  ap_ready,
  ap_done,
  ap_idle,
  M,
  P_N,
  alpha_u,
  beta_u,
  NUM_A_LEN,
  edge_list_ch_0,
  edge_list_ch_1,
  edge_list_ch_2,
  edge_list_ch_3,
  edge_list_ch_4,
  edge_list_ch_5,
  edge_list_ch_6,
  edge_list_ch_7,
  edge_list_ch_8,
  edge_list_ch_9,
  edge_list_ch_10,
  edge_list_ch_11,
  edge_list_ch_12,
  edge_list_ch_13,
  edge_list_ch_14,
  edge_list_ch_15,
  edge_list_ch_16,
  edge_list_ch_17,
  edge_list_ch_18,
  edge_list_ch_19,
  edge_list_ch_20,
  edge_list_ch_21,
  edge_list_ch_22,
  edge_list_ch_23,
  edge_list_ch_24,
  edge_list_ch_25,
  edge_list_ch_26,
  edge_list_ch_27,
  edge_list_ch_28,
  edge_list_ch_29,
  edge_list_ch_30,
  edge_list_ch_31,
  edge_list_ch_32,
  edge_list_ch_33,
  edge_list_ch_34,
  edge_list_ch_35,
  edge_list_ch_36,
  edge_list_ch_37,
  edge_list_ch_38,
  edge_list_ch_39,
  edge_list_ch_40,
  edge_list_ch_41,
  edge_list_ch_42,
  edge_list_ch_43,
  edge_list_ch_44,
  edge_list_ch_45,
  edge_list_ch_46,
  edge_list_ch_47,
  K,
  vec_X,
  vec_Y,
  NUM_ITE,
  edge_list_ptr,
  vec_Y_out,
  Arbiter_Y_0___M__q0,
  Arbiter_Y_0___P_N__q0,
  Arbiter_Y_0__ap_start,
  Arbiter_Y_0__ap_ready,
  Arbiter_Y_0__ap_done,
  Arbiter_Y_0__ap_idle,
  Arbiter_Y_1___M__q0,
  Arbiter_Y_1___P_N__q0,
  Arbiter_Y_1__ap_start,
  Arbiter_Y_1__ap_ready,
  Arbiter_Y_1__ap_done,
  Arbiter_Y_1__ap_idle,
  Arbiter_Y_2___M__q0,
  Arbiter_Y_2___P_N__q0,
  Arbiter_Y_2__ap_start,
  Arbiter_Y_2__ap_ready,
  Arbiter_Y_2__ap_done,
  Arbiter_Y_2__ap_idle,
  Arbiter_Y_3___M__q0,
  Arbiter_Y_3___P_N__q0,
  Arbiter_Y_3__ap_start,
  Arbiter_Y_3__ap_ready,
  Arbiter_Y_3__ap_done,
  Arbiter_Y_3__ap_idle,
  Arbiter_Y_4___M__q0,
  Arbiter_Y_4___P_N__q0,
  Arbiter_Y_4__ap_start,
  Arbiter_Y_4__ap_ready,
  Arbiter_Y_4__ap_done,
  Arbiter_Y_4__ap_idle,
  Arbiter_Y_5___M__q0,
  Arbiter_Y_5___P_N__q0,
  Arbiter_Y_5__ap_start,
  Arbiter_Y_5__ap_ready,
  Arbiter_Y_5__ap_done,
  Arbiter_Y_5__ap_idle,
  Arbiter_Y_6___M__q0,
  Arbiter_Y_6___P_N__q0,
  Arbiter_Y_6__ap_start,
  Arbiter_Y_6__ap_ready,
  Arbiter_Y_6__ap_done,
  Arbiter_Y_6__ap_idle,
  Arbiter_Y_7___M__q0,
  Arbiter_Y_7___P_N__q0,
  Arbiter_Y_7__ap_start,
  Arbiter_Y_7__ap_ready,
  Arbiter_Y_7__ap_done,
  Arbiter_Y_7__ap_idle,
  FloatvAddFloatv_0__ap_start,
  FloatvMultConst_0___M__q0,
  FloatvMultConst_0___P_N__q0,
  FloatvMultConst_0___alpha_u__q0,
  FloatvMultConst_0__ap_start,
  FloatvMultConst_0__ap_ready,
  FloatvMultConst_0__ap_done,
  FloatvMultConst_0__ap_idle,
  FloatvMultConst_1___M__q0,
  FloatvMultConst_1___P_N__q0,
  FloatvMultConst_1___beta_u__q0,
  FloatvMultConst_1__ap_start,
  FloatvMultConst_1__ap_ready,
  FloatvMultConst_1__ap_done,
  FloatvMultConst_1__ap_idle,
  Merger_Y_0__ap_start,
  PEG_Xvec_0__ap_start,
  PEG_Xvec_0__ap_ready,
  PEG_Xvec_0__ap_done,
  PEG_Xvec_0__ap_idle,
  PEG_Xvec_1__ap_start,
  PEG_Xvec_1__ap_ready,
  PEG_Xvec_1__ap_done,
  PEG_Xvec_1__ap_idle,
  PEG_Xvec_2__ap_start,
  PEG_Xvec_2__ap_ready,
  PEG_Xvec_2__ap_done,
  PEG_Xvec_2__ap_idle,
  PEG_Xvec_3__ap_start,
  PEG_Xvec_3__ap_ready,
  PEG_Xvec_3__ap_done,
  PEG_Xvec_3__ap_idle,
  PEG_Xvec_4__ap_start,
  PEG_Xvec_4__ap_ready,
  PEG_Xvec_4__ap_done,
  PEG_Xvec_4__ap_idle,
  PEG_Xvec_5__ap_start,
  PEG_Xvec_5__ap_ready,
  PEG_Xvec_5__ap_done,
  PEG_Xvec_5__ap_idle,
  PEG_Xvec_6__ap_start,
  PEG_Xvec_6__ap_ready,
  PEG_Xvec_6__ap_done,
  PEG_Xvec_6__ap_idle,
  PEG_Xvec_7__ap_start,
  PEG_Xvec_7__ap_ready,
  PEG_Xvec_7__ap_done,
  PEG_Xvec_7__ap_idle,
  PEG_Xvec_8__ap_start,
  PEG_Xvec_8__ap_ready,
  PEG_Xvec_8__ap_done,
  PEG_Xvec_8__ap_idle,
  PEG_Xvec_9__ap_start,
  PEG_Xvec_9__ap_ready,
  PEG_Xvec_9__ap_done,
  PEG_Xvec_9__ap_idle,
  PEG_Xvec_10__ap_start,
  PEG_Xvec_10__ap_ready,
  PEG_Xvec_10__ap_done,
  PEG_Xvec_10__ap_idle,
  PEG_Xvec_11__ap_start,
  PEG_Xvec_11__ap_ready,
  PEG_Xvec_11__ap_done,
  PEG_Xvec_11__ap_idle,
  PEG_Xvec_12__ap_start,
  PEG_Xvec_12__ap_ready,
  PEG_Xvec_12__ap_done,
  PEG_Xvec_12__ap_idle,
  PEG_Xvec_13__ap_start,
  PEG_Xvec_13__ap_ready,
  PEG_Xvec_13__ap_done,
  PEG_Xvec_13__ap_idle,
  PEG_Xvec_14__ap_start,
  PEG_Xvec_14__ap_ready,
  PEG_Xvec_14__ap_done,
  PEG_Xvec_14__ap_idle,
  PEG_Xvec_15__ap_start,
  PEG_Xvec_15__ap_ready,
  PEG_Xvec_15__ap_done,
  PEG_Xvec_15__ap_idle,
  PEG_Xvec_16__ap_start,
  PEG_Xvec_16__ap_ready,
  PEG_Xvec_16__ap_done,
  PEG_Xvec_16__ap_idle,
  PEG_Xvec_17__ap_start,
  PEG_Xvec_17__ap_ready,
  PEG_Xvec_17__ap_done,
  PEG_Xvec_17__ap_idle,
  PEG_Xvec_18__ap_start,
  PEG_Xvec_18__ap_ready,
  PEG_Xvec_18__ap_done,
  PEG_Xvec_18__ap_idle,
  PEG_Xvec_19__ap_start,
  PEG_Xvec_19__ap_ready,
  PEG_Xvec_19__ap_done,
  PEG_Xvec_19__ap_idle,
  PEG_Xvec_20__ap_start,
  PEG_Xvec_20__ap_ready,
  PEG_Xvec_20__ap_done,
  PEG_Xvec_20__ap_idle,
  PEG_Xvec_21__ap_start,
  PEG_Xvec_21__ap_ready,
  PEG_Xvec_21__ap_done,
  PEG_Xvec_21__ap_idle,
  PEG_Xvec_22__ap_start,
  PEG_Xvec_22__ap_ready,
  PEG_Xvec_22__ap_done,
  PEG_Xvec_22__ap_idle,
  PEG_Xvec_23__ap_start,
  PEG_Xvec_23__ap_ready,
  PEG_Xvec_23__ap_done,
  PEG_Xvec_23__ap_idle,
  PEG_Xvec_24__ap_start,
  PEG_Xvec_24__ap_ready,
  PEG_Xvec_24__ap_done,
  PEG_Xvec_24__ap_idle,
  PEG_Xvec_25__ap_start,
  PEG_Xvec_25__ap_ready,
  PEG_Xvec_25__ap_done,
  PEG_Xvec_25__ap_idle,
  PEG_Xvec_26__ap_start,
  PEG_Xvec_26__ap_ready,
  PEG_Xvec_26__ap_done,
  PEG_Xvec_26__ap_idle,
  PEG_Xvec_27__ap_start,
  PEG_Xvec_27__ap_ready,
  PEG_Xvec_27__ap_done,
  PEG_Xvec_27__ap_idle,
  PEG_Xvec_28__ap_start,
  PEG_Xvec_28__ap_ready,
  PEG_Xvec_28__ap_done,
  PEG_Xvec_28__ap_idle,
  PEG_Xvec_29__ap_start,
  PEG_Xvec_29__ap_ready,
  PEG_Xvec_29__ap_done,
  PEG_Xvec_29__ap_idle,
  PEG_Xvec_30__ap_start,
  PEG_Xvec_30__ap_ready,
  PEG_Xvec_30__ap_done,
  PEG_Xvec_30__ap_idle,
  PEG_Xvec_31__ap_start,
  PEG_Xvec_31__ap_ready,
  PEG_Xvec_31__ap_done,
  PEG_Xvec_31__ap_idle,
  PEG_Xvec_32__ap_start,
  PEG_Xvec_32__ap_ready,
  PEG_Xvec_32__ap_done,
  PEG_Xvec_32__ap_idle,
  PEG_Xvec_33__ap_start,
  PEG_Xvec_33__ap_ready,
  PEG_Xvec_33__ap_done,
  PEG_Xvec_33__ap_idle,
  PEG_Xvec_34__ap_start,
  PEG_Xvec_34__ap_ready,
  PEG_Xvec_34__ap_done,
  PEG_Xvec_34__ap_idle,
  PEG_Xvec_35__ap_start,
  PEG_Xvec_35__ap_ready,
  PEG_Xvec_35__ap_done,
  PEG_Xvec_35__ap_idle,
  PEG_Xvec_36__ap_start,
  PEG_Xvec_36__ap_ready,
  PEG_Xvec_36__ap_done,
  PEG_Xvec_36__ap_idle,
  PEG_Xvec_37__ap_start,
  PEG_Xvec_37__ap_ready,
  PEG_Xvec_37__ap_done,
  PEG_Xvec_37__ap_idle,
  PEG_Xvec_38__ap_start,
  PEG_Xvec_38__ap_ready,
  PEG_Xvec_38__ap_done,
  PEG_Xvec_38__ap_idle,
  PEG_Xvec_39__ap_start,
  PEG_Xvec_39__ap_ready,
  PEG_Xvec_39__ap_done,
  PEG_Xvec_39__ap_idle,
  PEG_Xvec_40__ap_start,
  PEG_Xvec_40__ap_ready,
  PEG_Xvec_40__ap_done,
  PEG_Xvec_40__ap_idle,
  PEG_Xvec_41__ap_start,
  PEG_Xvec_41__ap_ready,
  PEG_Xvec_41__ap_done,
  PEG_Xvec_41__ap_idle,
  PEG_Xvec_42__ap_start,
  PEG_Xvec_42__ap_ready,
  PEG_Xvec_42__ap_done,
  PEG_Xvec_42__ap_idle,
  PEG_Xvec_43__ap_start,
  PEG_Xvec_43__ap_ready,
  PEG_Xvec_43__ap_done,
  PEG_Xvec_43__ap_idle,
  PEG_Xvec_44__ap_start,
  PEG_Xvec_44__ap_ready,
  PEG_Xvec_44__ap_done,
  PEG_Xvec_44__ap_idle,
  PEG_Xvec_45__ap_start,
  PEG_Xvec_45__ap_ready,
  PEG_Xvec_45__ap_done,
  PEG_Xvec_45__ap_idle,
  PEG_Xvec_46__ap_start,
  PEG_Xvec_46__ap_ready,
  PEG_Xvec_46__ap_done,
  PEG_Xvec_46__ap_idle,
  PEG_Xvec_47__ap_start,
  PEG_Xvec_47__ap_ready,
  PEG_Xvec_47__ap_done,
  PEG_Xvec_47__ap_idle,
  PEG_Yvec_0__ap_start,
  PEG_Yvec_0__ap_ready,
  PEG_Yvec_0__ap_done,
  PEG_Yvec_0__ap_idle,
  PEG_Yvec_1__ap_start,
  PEG_Yvec_1__ap_ready,
  PEG_Yvec_1__ap_done,
  PEG_Yvec_1__ap_idle,
  PEG_Yvec_2__ap_start,
  PEG_Yvec_2__ap_ready,
  PEG_Yvec_2__ap_done,
  PEG_Yvec_2__ap_idle,
  PEG_Yvec_3__ap_start,
  PEG_Yvec_3__ap_ready,
  PEG_Yvec_3__ap_done,
  PEG_Yvec_3__ap_idle,
  PEG_Yvec_4__ap_start,
  PEG_Yvec_4__ap_ready,
  PEG_Yvec_4__ap_done,
  PEG_Yvec_4__ap_idle,
  PEG_Yvec_5__ap_start,
  PEG_Yvec_5__ap_ready,
  PEG_Yvec_5__ap_done,
  PEG_Yvec_5__ap_idle,
  PEG_Yvec_6__ap_start,
  PEG_Yvec_6__ap_ready,
  PEG_Yvec_6__ap_done,
  PEG_Yvec_6__ap_idle,
  PEG_Yvec_7__ap_start,
  PEG_Yvec_7__ap_ready,
  PEG_Yvec_7__ap_done,
  PEG_Yvec_7__ap_idle,
  PEG_Yvec_8__ap_start,
  PEG_Yvec_8__ap_ready,
  PEG_Yvec_8__ap_done,
  PEG_Yvec_8__ap_idle,
  PEG_Yvec_9__ap_start,
  PEG_Yvec_9__ap_ready,
  PEG_Yvec_9__ap_done,
  PEG_Yvec_9__ap_idle,
  PEG_Yvec_10__ap_start,
  PEG_Yvec_10__ap_ready,
  PEG_Yvec_10__ap_done,
  PEG_Yvec_10__ap_idle,
  PEG_Yvec_11__ap_start,
  PEG_Yvec_11__ap_ready,
  PEG_Yvec_11__ap_done,
  PEG_Yvec_11__ap_idle,
  PEG_Yvec_12__ap_start,
  PEG_Yvec_12__ap_ready,
  PEG_Yvec_12__ap_done,
  PEG_Yvec_12__ap_idle,
  PEG_Yvec_13__ap_start,
  PEG_Yvec_13__ap_ready,
  PEG_Yvec_13__ap_done,
  PEG_Yvec_13__ap_idle,
  PEG_Yvec_14__ap_start,
  PEG_Yvec_14__ap_ready,
  PEG_Yvec_14__ap_done,
  PEG_Yvec_14__ap_idle,
  PEG_Yvec_15__ap_start,
  PEG_Yvec_15__ap_ready,
  PEG_Yvec_15__ap_done,
  PEG_Yvec_15__ap_idle,
  PEG_Yvec_16__ap_start,
  PEG_Yvec_16__ap_ready,
  PEG_Yvec_16__ap_done,
  PEG_Yvec_16__ap_idle,
  PEG_Yvec_17__ap_start,
  PEG_Yvec_17__ap_ready,
  PEG_Yvec_17__ap_done,
  PEG_Yvec_17__ap_idle,
  PEG_Yvec_18__ap_start,
  PEG_Yvec_18__ap_ready,
  PEG_Yvec_18__ap_done,
  PEG_Yvec_18__ap_idle,
  PEG_Yvec_19__ap_start,
  PEG_Yvec_19__ap_ready,
  PEG_Yvec_19__ap_done,
  PEG_Yvec_19__ap_idle,
  PEG_Yvec_20__ap_start,
  PEG_Yvec_20__ap_ready,
  PEG_Yvec_20__ap_done,
  PEG_Yvec_20__ap_idle,
  PEG_Yvec_21__ap_start,
  PEG_Yvec_21__ap_ready,
  PEG_Yvec_21__ap_done,
  PEG_Yvec_21__ap_idle,
  PEG_Yvec_22__ap_start,
  PEG_Yvec_22__ap_ready,
  PEG_Yvec_22__ap_done,
  PEG_Yvec_22__ap_idle,
  PEG_Yvec_23__ap_start,
  PEG_Yvec_23__ap_ready,
  PEG_Yvec_23__ap_done,
  PEG_Yvec_23__ap_idle,
  PEG_Yvec_24__ap_start,
  PEG_Yvec_24__ap_ready,
  PEG_Yvec_24__ap_done,
  PEG_Yvec_24__ap_idle,
  PEG_Yvec_25__ap_start,
  PEG_Yvec_25__ap_ready,
  PEG_Yvec_25__ap_done,
  PEG_Yvec_25__ap_idle,
  PEG_Yvec_26__ap_start,
  PEG_Yvec_26__ap_ready,
  PEG_Yvec_26__ap_done,
  PEG_Yvec_26__ap_idle,
  PEG_Yvec_27__ap_start,
  PEG_Yvec_27__ap_ready,
  PEG_Yvec_27__ap_done,
  PEG_Yvec_27__ap_idle,
  PEG_Yvec_28__ap_start,
  PEG_Yvec_28__ap_ready,
  PEG_Yvec_28__ap_done,
  PEG_Yvec_28__ap_idle,
  PEG_Yvec_29__ap_start,
  PEG_Yvec_29__ap_ready,
  PEG_Yvec_29__ap_done,
  PEG_Yvec_29__ap_idle,
  PEG_Yvec_30__ap_start,
  PEG_Yvec_30__ap_ready,
  PEG_Yvec_30__ap_done,
  PEG_Yvec_30__ap_idle,
  PEG_Yvec_31__ap_start,
  PEG_Yvec_31__ap_ready,
  PEG_Yvec_31__ap_done,
  PEG_Yvec_31__ap_idle,
  PEG_Yvec_32__ap_start,
  PEG_Yvec_32__ap_ready,
  PEG_Yvec_32__ap_done,
  PEG_Yvec_32__ap_idle,
  PEG_Yvec_33__ap_start,
  PEG_Yvec_33__ap_ready,
  PEG_Yvec_33__ap_done,
  PEG_Yvec_33__ap_idle,
  PEG_Yvec_34__ap_start,
  PEG_Yvec_34__ap_ready,
  PEG_Yvec_34__ap_done,
  PEG_Yvec_34__ap_idle,
  PEG_Yvec_35__ap_start,
  PEG_Yvec_35__ap_ready,
  PEG_Yvec_35__ap_done,
  PEG_Yvec_35__ap_idle,
  PEG_Yvec_36__ap_start,
  PEG_Yvec_36__ap_ready,
  PEG_Yvec_36__ap_done,
  PEG_Yvec_36__ap_idle,
  PEG_Yvec_37__ap_start,
  PEG_Yvec_37__ap_ready,
  PEG_Yvec_37__ap_done,
  PEG_Yvec_37__ap_idle,
  PEG_Yvec_38__ap_start,
  PEG_Yvec_38__ap_ready,
  PEG_Yvec_38__ap_done,
  PEG_Yvec_38__ap_idle,
  PEG_Yvec_39__ap_start,
  PEG_Yvec_39__ap_ready,
  PEG_Yvec_39__ap_done,
  PEG_Yvec_39__ap_idle,
  PEG_Yvec_40__ap_start,
  PEG_Yvec_40__ap_ready,
  PEG_Yvec_40__ap_done,
  PEG_Yvec_40__ap_idle,
  PEG_Yvec_41__ap_start,
  PEG_Yvec_41__ap_ready,
  PEG_Yvec_41__ap_done,
  PEG_Yvec_41__ap_idle,
  PEG_Yvec_42__ap_start,
  PEG_Yvec_42__ap_ready,
  PEG_Yvec_42__ap_done,
  PEG_Yvec_42__ap_idle,
  PEG_Yvec_43__ap_start,
  PEG_Yvec_43__ap_ready,
  PEG_Yvec_43__ap_done,
  PEG_Yvec_43__ap_idle,
  PEG_Yvec_44__ap_start,
  PEG_Yvec_44__ap_ready,
  PEG_Yvec_44__ap_done,
  PEG_Yvec_44__ap_idle,
  PEG_Yvec_45__ap_start,
  PEG_Yvec_45__ap_ready,
  PEG_Yvec_45__ap_done,
  PEG_Yvec_45__ap_idle,
  PEG_Yvec_46__ap_start,
  PEG_Yvec_46__ap_ready,
  PEG_Yvec_46__ap_done,
  PEG_Yvec_46__ap_idle,
  PEG_Yvec_47__ap_start,
  PEG_Yvec_47__ap_ready,
  PEG_Yvec_47__ap_done,
  PEG_Yvec_47__ap_idle,
  black_hole_float_v16_0__ap_start,
  black_hole_int_0__ap_start,
  read_A_0___NUM_A_LEN__q0,
  read_A_0___P_N__q0,
  read_A_0___edge_list_ch_0__q0,
  read_A_0__ap_start,
  read_A_0__ap_ready,
  read_A_0__ap_done,
  read_A_0__ap_idle,
  read_A_1___NUM_A_LEN__q0,
  read_A_1___P_N__q0,
  read_A_1___edge_list_ch_1__q0,
  read_A_1__ap_start,
  read_A_1__ap_ready,
  read_A_1__ap_done,
  read_A_1__ap_idle,
  read_A_2___NUM_A_LEN__q0,
  read_A_2___P_N__q0,
  read_A_2___edge_list_ch_2__q0,
  read_A_2__ap_start,
  read_A_2__ap_ready,
  read_A_2__ap_done,
  read_A_2__ap_idle,
  read_A_3___NUM_A_LEN__q0,
  read_A_3___P_N__q0,
  read_A_3___edge_list_ch_3__q0,
  read_A_3__ap_start,
  read_A_3__ap_ready,
  read_A_3__ap_done,
  read_A_3__ap_idle,
  read_A_4___NUM_A_LEN__q0,
  read_A_4___P_N__q0,
  read_A_4___edge_list_ch_4__q0,
  read_A_4__ap_start,
  read_A_4__ap_ready,
  read_A_4__ap_done,
  read_A_4__ap_idle,
  read_A_5___NUM_A_LEN__q0,
  read_A_5___P_N__q0,
  read_A_5___edge_list_ch_5__q0,
  read_A_5__ap_start,
  read_A_5__ap_ready,
  read_A_5__ap_done,
  read_A_5__ap_idle,
  read_A_6___NUM_A_LEN__q0,
  read_A_6___P_N__q0,
  read_A_6___edge_list_ch_6__q0,
  read_A_6__ap_start,
  read_A_6__ap_ready,
  read_A_6__ap_done,
  read_A_6__ap_idle,
  read_A_7___NUM_A_LEN__q0,
  read_A_7___P_N__q0,
  read_A_7___edge_list_ch_7__q0,
  read_A_7__ap_start,
  read_A_7__ap_ready,
  read_A_7__ap_done,
  read_A_7__ap_idle,
  read_A_8___NUM_A_LEN__q0,
  read_A_8___P_N__q0,
  read_A_8___edge_list_ch_8__q0,
  read_A_8__ap_start,
  read_A_8__ap_ready,
  read_A_8__ap_done,
  read_A_8__ap_idle,
  read_A_9___NUM_A_LEN__q0,
  read_A_9___P_N__q0,
  read_A_9___edge_list_ch_9__q0,
  read_A_9__ap_start,
  read_A_9__ap_ready,
  read_A_9__ap_done,
  read_A_9__ap_idle,
  read_A_10___NUM_A_LEN__q0,
  read_A_10___P_N__q0,
  read_A_10___edge_list_ch_10__q0,
  read_A_10__ap_start,
  read_A_10__ap_ready,
  read_A_10__ap_done,
  read_A_10__ap_idle,
  read_A_11___NUM_A_LEN__q0,
  read_A_11___P_N__q0,
  read_A_11___edge_list_ch_11__q0,
  read_A_11__ap_start,
  read_A_11__ap_ready,
  read_A_11__ap_done,
  read_A_11__ap_idle,
  read_A_12___NUM_A_LEN__q0,
  read_A_12___P_N__q0,
  read_A_12___edge_list_ch_12__q0,
  read_A_12__ap_start,
  read_A_12__ap_ready,
  read_A_12__ap_done,
  read_A_12__ap_idle,
  read_A_13___NUM_A_LEN__q0,
  read_A_13___P_N__q0,
  read_A_13___edge_list_ch_13__q0,
  read_A_13__ap_start,
  read_A_13__ap_ready,
  read_A_13__ap_done,
  read_A_13__ap_idle,
  read_A_14___NUM_A_LEN__q0,
  read_A_14___P_N__q0,
  read_A_14___edge_list_ch_14__q0,
  read_A_14__ap_start,
  read_A_14__ap_ready,
  read_A_14__ap_done,
  read_A_14__ap_idle,
  read_A_15___NUM_A_LEN__q0,
  read_A_15___P_N__q0,
  read_A_15___edge_list_ch_15__q0,
  read_A_15__ap_start,
  read_A_15__ap_ready,
  read_A_15__ap_done,
  read_A_15__ap_idle,
  read_A_16___NUM_A_LEN__q0,
  read_A_16___P_N__q0,
  read_A_16___edge_list_ch_16__q0,
  read_A_16__ap_start,
  read_A_16__ap_ready,
  read_A_16__ap_done,
  read_A_16__ap_idle,
  read_A_17___NUM_A_LEN__q0,
  read_A_17___P_N__q0,
  read_A_17___edge_list_ch_17__q0,
  read_A_17__ap_start,
  read_A_17__ap_ready,
  read_A_17__ap_done,
  read_A_17__ap_idle,
  read_A_18___NUM_A_LEN__q0,
  read_A_18___P_N__q0,
  read_A_18___edge_list_ch_18__q0,
  read_A_18__ap_start,
  read_A_18__ap_ready,
  read_A_18__ap_done,
  read_A_18__ap_idle,
  read_A_19___NUM_A_LEN__q0,
  read_A_19___P_N__q0,
  read_A_19___edge_list_ch_19__q0,
  read_A_19__ap_start,
  read_A_19__ap_ready,
  read_A_19__ap_done,
  read_A_19__ap_idle,
  read_A_20___NUM_A_LEN__q0,
  read_A_20___P_N__q0,
  read_A_20___edge_list_ch_20__q0,
  read_A_20__ap_start,
  read_A_20__ap_ready,
  read_A_20__ap_done,
  read_A_20__ap_idle,
  read_A_21___NUM_A_LEN__q0,
  read_A_21___P_N__q0,
  read_A_21___edge_list_ch_21__q0,
  read_A_21__ap_start,
  read_A_21__ap_ready,
  read_A_21__ap_done,
  read_A_21__ap_idle,
  read_A_22___NUM_A_LEN__q0,
  read_A_22___P_N__q0,
  read_A_22___edge_list_ch_22__q0,
  read_A_22__ap_start,
  read_A_22__ap_ready,
  read_A_22__ap_done,
  read_A_22__ap_idle,
  read_A_23___NUM_A_LEN__q0,
  read_A_23___P_N__q0,
  read_A_23___edge_list_ch_23__q0,
  read_A_23__ap_start,
  read_A_23__ap_ready,
  read_A_23__ap_done,
  read_A_23__ap_idle,
  read_A_24___NUM_A_LEN__q0,
  read_A_24___P_N__q0,
  read_A_24___edge_list_ch_24__q0,
  read_A_24__ap_start,
  read_A_24__ap_ready,
  read_A_24__ap_done,
  read_A_24__ap_idle,
  read_A_25___NUM_A_LEN__q0,
  read_A_25___P_N__q0,
  read_A_25___edge_list_ch_25__q0,
  read_A_25__ap_start,
  read_A_25__ap_ready,
  read_A_25__ap_done,
  read_A_25__ap_idle,
  read_A_26___NUM_A_LEN__q0,
  read_A_26___P_N__q0,
  read_A_26___edge_list_ch_26__q0,
  read_A_26__ap_start,
  read_A_26__ap_ready,
  read_A_26__ap_done,
  read_A_26__ap_idle,
  read_A_27___NUM_A_LEN__q0,
  read_A_27___P_N__q0,
  read_A_27___edge_list_ch_27__q0,
  read_A_27__ap_start,
  read_A_27__ap_ready,
  read_A_27__ap_done,
  read_A_27__ap_idle,
  read_A_28___NUM_A_LEN__q0,
  read_A_28___P_N__q0,
  read_A_28___edge_list_ch_28__q0,
  read_A_28__ap_start,
  read_A_28__ap_ready,
  read_A_28__ap_done,
  read_A_28__ap_idle,
  read_A_29___NUM_A_LEN__q0,
  read_A_29___P_N__q0,
  read_A_29___edge_list_ch_29__q0,
  read_A_29__ap_start,
  read_A_29__ap_ready,
  read_A_29__ap_done,
  read_A_29__ap_idle,
  read_A_30___NUM_A_LEN__q0,
  read_A_30___P_N__q0,
  read_A_30___edge_list_ch_30__q0,
  read_A_30__ap_start,
  read_A_30__ap_ready,
  read_A_30__ap_done,
  read_A_30__ap_idle,
  read_A_31___NUM_A_LEN__q0,
  read_A_31___P_N__q0,
  read_A_31___edge_list_ch_31__q0,
  read_A_31__ap_start,
  read_A_31__ap_ready,
  read_A_31__ap_done,
  read_A_31__ap_idle,
  read_A_32___NUM_A_LEN__q0,
  read_A_32___P_N__q0,
  read_A_32___edge_list_ch_32__q0,
  read_A_32__ap_start,
  read_A_32__ap_ready,
  read_A_32__ap_done,
  read_A_32__ap_idle,
  read_A_33___NUM_A_LEN__q0,
  read_A_33___P_N__q0,
  read_A_33___edge_list_ch_33__q0,
  read_A_33__ap_start,
  read_A_33__ap_ready,
  read_A_33__ap_done,
  read_A_33__ap_idle,
  read_A_34___NUM_A_LEN__q0,
  read_A_34___P_N__q0,
  read_A_34___edge_list_ch_34__q0,
  read_A_34__ap_start,
  read_A_34__ap_ready,
  read_A_34__ap_done,
  read_A_34__ap_idle,
  read_A_35___NUM_A_LEN__q0,
  read_A_35___P_N__q0,
  read_A_35___edge_list_ch_35__q0,
  read_A_35__ap_start,
  read_A_35__ap_ready,
  read_A_35__ap_done,
  read_A_35__ap_idle,
  read_A_36___NUM_A_LEN__q0,
  read_A_36___P_N__q0,
  read_A_36___edge_list_ch_36__q0,
  read_A_36__ap_start,
  read_A_36__ap_ready,
  read_A_36__ap_done,
  read_A_36__ap_idle,
  read_A_37___NUM_A_LEN__q0,
  read_A_37___P_N__q0,
  read_A_37___edge_list_ch_37__q0,
  read_A_37__ap_start,
  read_A_37__ap_ready,
  read_A_37__ap_done,
  read_A_37__ap_idle,
  read_A_38___NUM_A_LEN__q0,
  read_A_38___P_N__q0,
  read_A_38___edge_list_ch_38__q0,
  read_A_38__ap_start,
  read_A_38__ap_ready,
  read_A_38__ap_done,
  read_A_38__ap_idle,
  read_A_39___NUM_A_LEN__q0,
  read_A_39___P_N__q0,
  read_A_39___edge_list_ch_39__q0,
  read_A_39__ap_start,
  read_A_39__ap_ready,
  read_A_39__ap_done,
  read_A_39__ap_idle,
  read_A_40___NUM_A_LEN__q0,
  read_A_40___P_N__q0,
  read_A_40___edge_list_ch_40__q0,
  read_A_40__ap_start,
  read_A_40__ap_ready,
  read_A_40__ap_done,
  read_A_40__ap_idle,
  read_A_41___NUM_A_LEN__q0,
  read_A_41___P_N__q0,
  read_A_41___edge_list_ch_41__q0,
  read_A_41__ap_start,
  read_A_41__ap_ready,
  read_A_41__ap_done,
  read_A_41__ap_idle,
  read_A_42___NUM_A_LEN__q0,
  read_A_42___P_N__q0,
  read_A_42___edge_list_ch_42__q0,
  read_A_42__ap_start,
  read_A_42__ap_ready,
  read_A_42__ap_done,
  read_A_42__ap_idle,
  read_A_43___NUM_A_LEN__q0,
  read_A_43___P_N__q0,
  read_A_43___edge_list_ch_43__q0,
  read_A_43__ap_start,
  read_A_43__ap_ready,
  read_A_43__ap_done,
  read_A_43__ap_idle,
  read_A_44___NUM_A_LEN__q0,
  read_A_44___P_N__q0,
  read_A_44___edge_list_ch_44__q0,
  read_A_44__ap_start,
  read_A_44__ap_ready,
  read_A_44__ap_done,
  read_A_44__ap_idle,
  read_A_45___NUM_A_LEN__q0,
  read_A_45___P_N__q0,
  read_A_45___edge_list_ch_45__q0,
  read_A_45__ap_start,
  read_A_45__ap_ready,
  read_A_45__ap_done,
  read_A_45__ap_idle,
  read_A_46___NUM_A_LEN__q0,
  read_A_46___P_N__q0,
  read_A_46___edge_list_ch_46__q0,
  read_A_46__ap_start,
  read_A_46__ap_ready,
  read_A_46__ap_done,
  read_A_46__ap_idle,
  read_A_47___NUM_A_LEN__q0,
  read_A_47___P_N__q0,
  read_A_47___edge_list_ch_47__q0,
  read_A_47__ap_start,
  read_A_47__ap_ready,
  read_A_47__ap_done,
  read_A_47__ap_idle,
  read_X_0___K__q0,
  read_X_0___P_N__q0,
  read_X_0___vec_X__q0,
  read_X_0__ap_start,
  read_X_0__ap_ready,
  read_X_0__ap_done,
  read_X_0__ap_idle,
  read_Y_0___M__q0,
  read_Y_0___P_N__q0,
  read_Y_0___vec_Y__q0,
  read_Y_0__ap_start,
  read_Y_0__ap_ready,
  read_Y_0__ap_done,
  read_Y_0__ap_idle,
  read_edge_list_ptr_0___K__q0,
  read_edge_list_ptr_0___M__q0,
  read_edge_list_ptr_0___NUM_ITE__q0,
  read_edge_list_ptr_0___P_N__q0,
  read_edge_list_ptr_0___edge_list_ptr__q0,
  read_edge_list_ptr_0__ap_start,
  read_edge_list_ptr_0__ap_ready,
  read_edge_list_ptr_0__ap_done,
  read_edge_list_ptr_0__ap_idle,
  write_Y_0___M__q0,
  write_Y_0___P_N__q0,
  write_Y_0___vec_Y_out__q0,
  write_Y_0__ap_start,
  write_Y_0__ap_ready,
  write_Y_0__ap_done,
  write_Y_0__ap_idle
);

  // pragma RS clk port=ap_clk
  // pragma RS rst port=ap_rst_n active=low
  // pragma RS ap-ctrl ap_start=ap_start ap_done=ap_done ap_idle=ap_idle ap_ready=ap_ready scalar=(edge_list_ptr|edge_list_ch_0|edge_list_ch_1|edge_list_ch_2|edge_list_ch_3|edge_list_ch_4|edge_list_ch_5|edge_list_ch_6|edge_list_ch_7|edge_list_ch_8|edge_list_ch_9|edge_list_ch_10|edge_list_ch_11|edge_list_ch_12|edge_list_ch_13|edge_list_ch_14|edge_list_ch_15|edge_list_ch_16|edge_list_ch_17|edge_list_ch_18|edge_list_ch_19|edge_list_ch_20|edge_list_ch_21|edge_list_ch_22|edge_list_ch_23|edge_list_ch_24|edge_list_ch_25|edge_list_ch_26|edge_list_ch_27|edge_list_ch_28|edge_list_ch_29|edge_list_ch_30|edge_list_ch_31|edge_list_ch_32|edge_list_ch_33|edge_list_ch_34|edge_list_ch_35|edge_list_ch_36|edge_list_ch_37|edge_list_ch_38|edge_list_ch_39|edge_list_ch_40|edge_list_ch_41|edge_list_ch_42|edge_list_ch_43|edge_list_ch_44|edge_list_ch_45|edge_list_ch_46|edge_list_ch_47|vec_X|vec_Y|vec_Y_out|NUM_ITE|NUM_A_LEN|M|K|P_N|alpha_u|beta_u)
  // pragma RS ap-ctrl ap_start=Arbiter_Y_0__ap_start ap_done=Arbiter_Y_0__ap_done ap_idle=Arbiter_Y_0__ap_idle ap_ready=Arbiter_Y_0__ap_ready scalar=Arbiter_Y_0___.*
  // pragma RS ap-ctrl ap_start=Arbiter_Y_1__ap_start ap_done=Arbiter_Y_1__ap_done ap_idle=Arbiter_Y_1__ap_idle ap_ready=Arbiter_Y_1__ap_ready scalar=Arbiter_Y_1___.*
  // pragma RS ap-ctrl ap_start=Arbiter_Y_2__ap_start ap_done=Arbiter_Y_2__ap_done ap_idle=Arbiter_Y_2__ap_idle ap_ready=Arbiter_Y_2__ap_ready scalar=Arbiter_Y_2___.*
  // pragma RS ap-ctrl ap_start=Arbiter_Y_3__ap_start ap_done=Arbiter_Y_3__ap_done ap_idle=Arbiter_Y_3__ap_idle ap_ready=Arbiter_Y_3__ap_ready scalar=Arbiter_Y_3___.*
  // pragma RS ap-ctrl ap_start=Arbiter_Y_4__ap_start ap_done=Arbiter_Y_4__ap_done ap_idle=Arbiter_Y_4__ap_idle ap_ready=Arbiter_Y_4__ap_ready scalar=Arbiter_Y_4___.*
  // pragma RS ap-ctrl ap_start=Arbiter_Y_5__ap_start ap_done=Arbiter_Y_5__ap_done ap_idle=Arbiter_Y_5__ap_idle ap_ready=Arbiter_Y_5__ap_ready scalar=Arbiter_Y_5___.*
  // pragma RS ap-ctrl ap_start=Arbiter_Y_6__ap_start ap_done=Arbiter_Y_6__ap_done ap_idle=Arbiter_Y_6__ap_idle ap_ready=Arbiter_Y_6__ap_ready scalar=Arbiter_Y_6___.*
  // pragma RS ap-ctrl ap_start=Arbiter_Y_7__ap_start ap_done=Arbiter_Y_7__ap_done ap_idle=Arbiter_Y_7__ap_idle ap_ready=Arbiter_Y_7__ap_ready scalar=Arbiter_Y_7___.*
  // pragma RS ap-ctrl ap_start=FloatvAddFloatv_0__ap_start
  // pragma RS ap-ctrl ap_start=FloatvMultConst_0__ap_start ap_done=FloatvMultConst_0__ap_done ap_idle=FloatvMultConst_0__ap_idle ap_ready=FloatvMultConst_0__ap_ready scalar=FloatvMultConst_0___.*
  // pragma RS ap-ctrl ap_start=FloatvMultConst_1__ap_start ap_done=FloatvMultConst_1__ap_done ap_idle=FloatvMultConst_1__ap_idle ap_ready=FloatvMultConst_1__ap_ready scalar=FloatvMultConst_1___.*
  // pragma RS ap-ctrl ap_start=Merger_Y_0__ap_start
  // pragma RS ap-ctrl ap_start=PEG_Xvec_0__ap_start ap_done=PEG_Xvec_0__ap_done ap_idle=PEG_Xvec_0__ap_idle ap_ready=PEG_Xvec_0__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_1__ap_start ap_done=PEG_Xvec_1__ap_done ap_idle=PEG_Xvec_1__ap_idle ap_ready=PEG_Xvec_1__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_2__ap_start ap_done=PEG_Xvec_2__ap_done ap_idle=PEG_Xvec_2__ap_idle ap_ready=PEG_Xvec_2__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_3__ap_start ap_done=PEG_Xvec_3__ap_done ap_idle=PEG_Xvec_3__ap_idle ap_ready=PEG_Xvec_3__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_4__ap_start ap_done=PEG_Xvec_4__ap_done ap_idle=PEG_Xvec_4__ap_idle ap_ready=PEG_Xvec_4__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_5__ap_start ap_done=PEG_Xvec_5__ap_done ap_idle=PEG_Xvec_5__ap_idle ap_ready=PEG_Xvec_5__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_6__ap_start ap_done=PEG_Xvec_6__ap_done ap_idle=PEG_Xvec_6__ap_idle ap_ready=PEG_Xvec_6__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_7__ap_start ap_done=PEG_Xvec_7__ap_done ap_idle=PEG_Xvec_7__ap_idle ap_ready=PEG_Xvec_7__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_8__ap_start ap_done=PEG_Xvec_8__ap_done ap_idle=PEG_Xvec_8__ap_idle ap_ready=PEG_Xvec_8__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_9__ap_start ap_done=PEG_Xvec_9__ap_done ap_idle=PEG_Xvec_9__ap_idle ap_ready=PEG_Xvec_9__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_10__ap_start ap_done=PEG_Xvec_10__ap_done ap_idle=PEG_Xvec_10__ap_idle ap_ready=PEG_Xvec_10__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_11__ap_start ap_done=PEG_Xvec_11__ap_done ap_idle=PEG_Xvec_11__ap_idle ap_ready=PEG_Xvec_11__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_12__ap_start ap_done=PEG_Xvec_12__ap_done ap_idle=PEG_Xvec_12__ap_idle ap_ready=PEG_Xvec_12__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_13__ap_start ap_done=PEG_Xvec_13__ap_done ap_idle=PEG_Xvec_13__ap_idle ap_ready=PEG_Xvec_13__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_14__ap_start ap_done=PEG_Xvec_14__ap_done ap_idle=PEG_Xvec_14__ap_idle ap_ready=PEG_Xvec_14__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_15__ap_start ap_done=PEG_Xvec_15__ap_done ap_idle=PEG_Xvec_15__ap_idle ap_ready=PEG_Xvec_15__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_16__ap_start ap_done=PEG_Xvec_16__ap_done ap_idle=PEG_Xvec_16__ap_idle ap_ready=PEG_Xvec_16__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_17__ap_start ap_done=PEG_Xvec_17__ap_done ap_idle=PEG_Xvec_17__ap_idle ap_ready=PEG_Xvec_17__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_18__ap_start ap_done=PEG_Xvec_18__ap_done ap_idle=PEG_Xvec_18__ap_idle ap_ready=PEG_Xvec_18__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_19__ap_start ap_done=PEG_Xvec_19__ap_done ap_idle=PEG_Xvec_19__ap_idle ap_ready=PEG_Xvec_19__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_20__ap_start ap_done=PEG_Xvec_20__ap_done ap_idle=PEG_Xvec_20__ap_idle ap_ready=PEG_Xvec_20__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_21__ap_start ap_done=PEG_Xvec_21__ap_done ap_idle=PEG_Xvec_21__ap_idle ap_ready=PEG_Xvec_21__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_22__ap_start ap_done=PEG_Xvec_22__ap_done ap_idle=PEG_Xvec_22__ap_idle ap_ready=PEG_Xvec_22__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_23__ap_start ap_done=PEG_Xvec_23__ap_done ap_idle=PEG_Xvec_23__ap_idle ap_ready=PEG_Xvec_23__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_24__ap_start ap_done=PEG_Xvec_24__ap_done ap_idle=PEG_Xvec_24__ap_idle ap_ready=PEG_Xvec_24__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_25__ap_start ap_done=PEG_Xvec_25__ap_done ap_idle=PEG_Xvec_25__ap_idle ap_ready=PEG_Xvec_25__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_26__ap_start ap_done=PEG_Xvec_26__ap_done ap_idle=PEG_Xvec_26__ap_idle ap_ready=PEG_Xvec_26__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_27__ap_start ap_done=PEG_Xvec_27__ap_done ap_idle=PEG_Xvec_27__ap_idle ap_ready=PEG_Xvec_27__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_28__ap_start ap_done=PEG_Xvec_28__ap_done ap_idle=PEG_Xvec_28__ap_idle ap_ready=PEG_Xvec_28__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_29__ap_start ap_done=PEG_Xvec_29__ap_done ap_idle=PEG_Xvec_29__ap_idle ap_ready=PEG_Xvec_29__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_30__ap_start ap_done=PEG_Xvec_30__ap_done ap_idle=PEG_Xvec_30__ap_idle ap_ready=PEG_Xvec_30__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_31__ap_start ap_done=PEG_Xvec_31__ap_done ap_idle=PEG_Xvec_31__ap_idle ap_ready=PEG_Xvec_31__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_32__ap_start ap_done=PEG_Xvec_32__ap_done ap_idle=PEG_Xvec_32__ap_idle ap_ready=PEG_Xvec_32__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_33__ap_start ap_done=PEG_Xvec_33__ap_done ap_idle=PEG_Xvec_33__ap_idle ap_ready=PEG_Xvec_33__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_34__ap_start ap_done=PEG_Xvec_34__ap_done ap_idle=PEG_Xvec_34__ap_idle ap_ready=PEG_Xvec_34__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_35__ap_start ap_done=PEG_Xvec_35__ap_done ap_idle=PEG_Xvec_35__ap_idle ap_ready=PEG_Xvec_35__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_36__ap_start ap_done=PEG_Xvec_36__ap_done ap_idle=PEG_Xvec_36__ap_idle ap_ready=PEG_Xvec_36__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_37__ap_start ap_done=PEG_Xvec_37__ap_done ap_idle=PEG_Xvec_37__ap_idle ap_ready=PEG_Xvec_37__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_38__ap_start ap_done=PEG_Xvec_38__ap_done ap_idle=PEG_Xvec_38__ap_idle ap_ready=PEG_Xvec_38__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_39__ap_start ap_done=PEG_Xvec_39__ap_done ap_idle=PEG_Xvec_39__ap_idle ap_ready=PEG_Xvec_39__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_40__ap_start ap_done=PEG_Xvec_40__ap_done ap_idle=PEG_Xvec_40__ap_idle ap_ready=PEG_Xvec_40__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_41__ap_start ap_done=PEG_Xvec_41__ap_done ap_idle=PEG_Xvec_41__ap_idle ap_ready=PEG_Xvec_41__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_42__ap_start ap_done=PEG_Xvec_42__ap_done ap_idle=PEG_Xvec_42__ap_idle ap_ready=PEG_Xvec_42__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_43__ap_start ap_done=PEG_Xvec_43__ap_done ap_idle=PEG_Xvec_43__ap_idle ap_ready=PEG_Xvec_43__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_44__ap_start ap_done=PEG_Xvec_44__ap_done ap_idle=PEG_Xvec_44__ap_idle ap_ready=PEG_Xvec_44__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_45__ap_start ap_done=PEG_Xvec_45__ap_done ap_idle=PEG_Xvec_45__ap_idle ap_ready=PEG_Xvec_45__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_46__ap_start ap_done=PEG_Xvec_46__ap_done ap_idle=PEG_Xvec_46__ap_idle ap_ready=PEG_Xvec_46__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Xvec_47__ap_start ap_done=PEG_Xvec_47__ap_done ap_idle=PEG_Xvec_47__ap_idle ap_ready=PEG_Xvec_47__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_0__ap_start ap_done=PEG_Yvec_0__ap_done ap_idle=PEG_Yvec_0__ap_idle ap_ready=PEG_Yvec_0__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_1__ap_start ap_done=PEG_Yvec_1__ap_done ap_idle=PEG_Yvec_1__ap_idle ap_ready=PEG_Yvec_1__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_2__ap_start ap_done=PEG_Yvec_2__ap_done ap_idle=PEG_Yvec_2__ap_idle ap_ready=PEG_Yvec_2__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_3__ap_start ap_done=PEG_Yvec_3__ap_done ap_idle=PEG_Yvec_3__ap_idle ap_ready=PEG_Yvec_3__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_4__ap_start ap_done=PEG_Yvec_4__ap_done ap_idle=PEG_Yvec_4__ap_idle ap_ready=PEG_Yvec_4__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_5__ap_start ap_done=PEG_Yvec_5__ap_done ap_idle=PEG_Yvec_5__ap_idle ap_ready=PEG_Yvec_5__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_6__ap_start ap_done=PEG_Yvec_6__ap_done ap_idle=PEG_Yvec_6__ap_idle ap_ready=PEG_Yvec_6__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_7__ap_start ap_done=PEG_Yvec_7__ap_done ap_idle=PEG_Yvec_7__ap_idle ap_ready=PEG_Yvec_7__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_8__ap_start ap_done=PEG_Yvec_8__ap_done ap_idle=PEG_Yvec_8__ap_idle ap_ready=PEG_Yvec_8__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_9__ap_start ap_done=PEG_Yvec_9__ap_done ap_idle=PEG_Yvec_9__ap_idle ap_ready=PEG_Yvec_9__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_10__ap_start ap_done=PEG_Yvec_10__ap_done ap_idle=PEG_Yvec_10__ap_idle ap_ready=PEG_Yvec_10__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_11__ap_start ap_done=PEG_Yvec_11__ap_done ap_idle=PEG_Yvec_11__ap_idle ap_ready=PEG_Yvec_11__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_12__ap_start ap_done=PEG_Yvec_12__ap_done ap_idle=PEG_Yvec_12__ap_idle ap_ready=PEG_Yvec_12__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_13__ap_start ap_done=PEG_Yvec_13__ap_done ap_idle=PEG_Yvec_13__ap_idle ap_ready=PEG_Yvec_13__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_14__ap_start ap_done=PEG_Yvec_14__ap_done ap_idle=PEG_Yvec_14__ap_idle ap_ready=PEG_Yvec_14__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_15__ap_start ap_done=PEG_Yvec_15__ap_done ap_idle=PEG_Yvec_15__ap_idle ap_ready=PEG_Yvec_15__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_16__ap_start ap_done=PEG_Yvec_16__ap_done ap_idle=PEG_Yvec_16__ap_idle ap_ready=PEG_Yvec_16__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_17__ap_start ap_done=PEG_Yvec_17__ap_done ap_idle=PEG_Yvec_17__ap_idle ap_ready=PEG_Yvec_17__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_18__ap_start ap_done=PEG_Yvec_18__ap_done ap_idle=PEG_Yvec_18__ap_idle ap_ready=PEG_Yvec_18__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_19__ap_start ap_done=PEG_Yvec_19__ap_done ap_idle=PEG_Yvec_19__ap_idle ap_ready=PEG_Yvec_19__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_20__ap_start ap_done=PEG_Yvec_20__ap_done ap_idle=PEG_Yvec_20__ap_idle ap_ready=PEG_Yvec_20__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_21__ap_start ap_done=PEG_Yvec_21__ap_done ap_idle=PEG_Yvec_21__ap_idle ap_ready=PEG_Yvec_21__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_22__ap_start ap_done=PEG_Yvec_22__ap_done ap_idle=PEG_Yvec_22__ap_idle ap_ready=PEG_Yvec_22__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_23__ap_start ap_done=PEG_Yvec_23__ap_done ap_idle=PEG_Yvec_23__ap_idle ap_ready=PEG_Yvec_23__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_24__ap_start ap_done=PEG_Yvec_24__ap_done ap_idle=PEG_Yvec_24__ap_idle ap_ready=PEG_Yvec_24__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_25__ap_start ap_done=PEG_Yvec_25__ap_done ap_idle=PEG_Yvec_25__ap_idle ap_ready=PEG_Yvec_25__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_26__ap_start ap_done=PEG_Yvec_26__ap_done ap_idle=PEG_Yvec_26__ap_idle ap_ready=PEG_Yvec_26__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_27__ap_start ap_done=PEG_Yvec_27__ap_done ap_idle=PEG_Yvec_27__ap_idle ap_ready=PEG_Yvec_27__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_28__ap_start ap_done=PEG_Yvec_28__ap_done ap_idle=PEG_Yvec_28__ap_idle ap_ready=PEG_Yvec_28__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_29__ap_start ap_done=PEG_Yvec_29__ap_done ap_idle=PEG_Yvec_29__ap_idle ap_ready=PEG_Yvec_29__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_30__ap_start ap_done=PEG_Yvec_30__ap_done ap_idle=PEG_Yvec_30__ap_idle ap_ready=PEG_Yvec_30__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_31__ap_start ap_done=PEG_Yvec_31__ap_done ap_idle=PEG_Yvec_31__ap_idle ap_ready=PEG_Yvec_31__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_32__ap_start ap_done=PEG_Yvec_32__ap_done ap_idle=PEG_Yvec_32__ap_idle ap_ready=PEG_Yvec_32__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_33__ap_start ap_done=PEG_Yvec_33__ap_done ap_idle=PEG_Yvec_33__ap_idle ap_ready=PEG_Yvec_33__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_34__ap_start ap_done=PEG_Yvec_34__ap_done ap_idle=PEG_Yvec_34__ap_idle ap_ready=PEG_Yvec_34__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_35__ap_start ap_done=PEG_Yvec_35__ap_done ap_idle=PEG_Yvec_35__ap_idle ap_ready=PEG_Yvec_35__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_36__ap_start ap_done=PEG_Yvec_36__ap_done ap_idle=PEG_Yvec_36__ap_idle ap_ready=PEG_Yvec_36__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_37__ap_start ap_done=PEG_Yvec_37__ap_done ap_idle=PEG_Yvec_37__ap_idle ap_ready=PEG_Yvec_37__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_38__ap_start ap_done=PEG_Yvec_38__ap_done ap_idle=PEG_Yvec_38__ap_idle ap_ready=PEG_Yvec_38__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_39__ap_start ap_done=PEG_Yvec_39__ap_done ap_idle=PEG_Yvec_39__ap_idle ap_ready=PEG_Yvec_39__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_40__ap_start ap_done=PEG_Yvec_40__ap_done ap_idle=PEG_Yvec_40__ap_idle ap_ready=PEG_Yvec_40__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_41__ap_start ap_done=PEG_Yvec_41__ap_done ap_idle=PEG_Yvec_41__ap_idle ap_ready=PEG_Yvec_41__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_42__ap_start ap_done=PEG_Yvec_42__ap_done ap_idle=PEG_Yvec_42__ap_idle ap_ready=PEG_Yvec_42__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_43__ap_start ap_done=PEG_Yvec_43__ap_done ap_idle=PEG_Yvec_43__ap_idle ap_ready=PEG_Yvec_43__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_44__ap_start ap_done=PEG_Yvec_44__ap_done ap_idle=PEG_Yvec_44__ap_idle ap_ready=PEG_Yvec_44__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_45__ap_start ap_done=PEG_Yvec_45__ap_done ap_idle=PEG_Yvec_45__ap_idle ap_ready=PEG_Yvec_45__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_46__ap_start ap_done=PEG_Yvec_46__ap_done ap_idle=PEG_Yvec_46__ap_idle ap_ready=PEG_Yvec_46__ap_ready
  // pragma RS ap-ctrl ap_start=PEG_Yvec_47__ap_start ap_done=PEG_Yvec_47__ap_done ap_idle=PEG_Yvec_47__ap_idle ap_ready=PEG_Yvec_47__ap_ready
  // pragma RS ap-ctrl ap_start=black_hole_float_v16_0__ap_start
  // pragma RS ap-ctrl ap_start=black_hole_int_0__ap_start
  // pragma RS ap-ctrl ap_start=read_A_0__ap_start ap_done=read_A_0__ap_done ap_idle=read_A_0__ap_idle ap_ready=read_A_0__ap_ready scalar=read_A_0___.*
  // pragma RS ap-ctrl ap_start=read_A_1__ap_start ap_done=read_A_1__ap_done ap_idle=read_A_1__ap_idle ap_ready=read_A_1__ap_ready scalar=read_A_1___.*
  // pragma RS ap-ctrl ap_start=read_A_2__ap_start ap_done=read_A_2__ap_done ap_idle=read_A_2__ap_idle ap_ready=read_A_2__ap_ready scalar=read_A_2___.*
  // pragma RS ap-ctrl ap_start=read_A_3__ap_start ap_done=read_A_3__ap_done ap_idle=read_A_3__ap_idle ap_ready=read_A_3__ap_ready scalar=read_A_3___.*
  // pragma RS ap-ctrl ap_start=read_A_4__ap_start ap_done=read_A_4__ap_done ap_idle=read_A_4__ap_idle ap_ready=read_A_4__ap_ready scalar=read_A_4___.*
  // pragma RS ap-ctrl ap_start=read_A_5__ap_start ap_done=read_A_5__ap_done ap_idle=read_A_5__ap_idle ap_ready=read_A_5__ap_ready scalar=read_A_5___.*
  // pragma RS ap-ctrl ap_start=read_A_6__ap_start ap_done=read_A_6__ap_done ap_idle=read_A_6__ap_idle ap_ready=read_A_6__ap_ready scalar=read_A_6___.*
  // pragma RS ap-ctrl ap_start=read_A_7__ap_start ap_done=read_A_7__ap_done ap_idle=read_A_7__ap_idle ap_ready=read_A_7__ap_ready scalar=read_A_7___.*
  // pragma RS ap-ctrl ap_start=read_A_8__ap_start ap_done=read_A_8__ap_done ap_idle=read_A_8__ap_idle ap_ready=read_A_8__ap_ready scalar=read_A_8___.*
  // pragma RS ap-ctrl ap_start=read_A_9__ap_start ap_done=read_A_9__ap_done ap_idle=read_A_9__ap_idle ap_ready=read_A_9__ap_ready scalar=read_A_9___.*
  // pragma RS ap-ctrl ap_start=read_A_10__ap_start ap_done=read_A_10__ap_done ap_idle=read_A_10__ap_idle ap_ready=read_A_10__ap_ready scalar=read_A_10___.*
  // pragma RS ap-ctrl ap_start=read_A_11__ap_start ap_done=read_A_11__ap_done ap_idle=read_A_11__ap_idle ap_ready=read_A_11__ap_ready scalar=read_A_11___.*
  // pragma RS ap-ctrl ap_start=read_A_12__ap_start ap_done=read_A_12__ap_done ap_idle=read_A_12__ap_idle ap_ready=read_A_12__ap_ready scalar=read_A_12___.*
  // pragma RS ap-ctrl ap_start=read_A_13__ap_start ap_done=read_A_13__ap_done ap_idle=read_A_13__ap_idle ap_ready=read_A_13__ap_ready scalar=read_A_13___.*
  // pragma RS ap-ctrl ap_start=read_A_14__ap_start ap_done=read_A_14__ap_done ap_idle=read_A_14__ap_idle ap_ready=read_A_14__ap_ready scalar=read_A_14___.*
  // pragma RS ap-ctrl ap_start=read_A_15__ap_start ap_done=read_A_15__ap_done ap_idle=read_A_15__ap_idle ap_ready=read_A_15__ap_ready scalar=read_A_15___.*
  // pragma RS ap-ctrl ap_start=read_A_16__ap_start ap_done=read_A_16__ap_done ap_idle=read_A_16__ap_idle ap_ready=read_A_16__ap_ready scalar=read_A_16___.*
  // pragma RS ap-ctrl ap_start=read_A_17__ap_start ap_done=read_A_17__ap_done ap_idle=read_A_17__ap_idle ap_ready=read_A_17__ap_ready scalar=read_A_17___.*
  // pragma RS ap-ctrl ap_start=read_A_18__ap_start ap_done=read_A_18__ap_done ap_idle=read_A_18__ap_idle ap_ready=read_A_18__ap_ready scalar=read_A_18___.*
  // pragma RS ap-ctrl ap_start=read_A_19__ap_start ap_done=read_A_19__ap_done ap_idle=read_A_19__ap_idle ap_ready=read_A_19__ap_ready scalar=read_A_19___.*
  // pragma RS ap-ctrl ap_start=read_A_20__ap_start ap_done=read_A_20__ap_done ap_idle=read_A_20__ap_idle ap_ready=read_A_20__ap_ready scalar=read_A_20___.*
  // pragma RS ap-ctrl ap_start=read_A_21__ap_start ap_done=read_A_21__ap_done ap_idle=read_A_21__ap_idle ap_ready=read_A_21__ap_ready scalar=read_A_21___.*
  // pragma RS ap-ctrl ap_start=read_A_22__ap_start ap_done=read_A_22__ap_done ap_idle=read_A_22__ap_idle ap_ready=read_A_22__ap_ready scalar=read_A_22___.*
  // pragma RS ap-ctrl ap_start=read_A_23__ap_start ap_done=read_A_23__ap_done ap_idle=read_A_23__ap_idle ap_ready=read_A_23__ap_ready scalar=read_A_23___.*
  // pragma RS ap-ctrl ap_start=read_A_24__ap_start ap_done=read_A_24__ap_done ap_idle=read_A_24__ap_idle ap_ready=read_A_24__ap_ready scalar=read_A_24___.*
  // pragma RS ap-ctrl ap_start=read_A_25__ap_start ap_done=read_A_25__ap_done ap_idle=read_A_25__ap_idle ap_ready=read_A_25__ap_ready scalar=read_A_25___.*
  // pragma RS ap-ctrl ap_start=read_A_26__ap_start ap_done=read_A_26__ap_done ap_idle=read_A_26__ap_idle ap_ready=read_A_26__ap_ready scalar=read_A_26___.*
  // pragma RS ap-ctrl ap_start=read_A_27__ap_start ap_done=read_A_27__ap_done ap_idle=read_A_27__ap_idle ap_ready=read_A_27__ap_ready scalar=read_A_27___.*
  // pragma RS ap-ctrl ap_start=read_A_28__ap_start ap_done=read_A_28__ap_done ap_idle=read_A_28__ap_idle ap_ready=read_A_28__ap_ready scalar=read_A_28___.*
  // pragma RS ap-ctrl ap_start=read_A_29__ap_start ap_done=read_A_29__ap_done ap_idle=read_A_29__ap_idle ap_ready=read_A_29__ap_ready scalar=read_A_29___.*
  // pragma RS ap-ctrl ap_start=read_A_30__ap_start ap_done=read_A_30__ap_done ap_idle=read_A_30__ap_idle ap_ready=read_A_30__ap_ready scalar=read_A_30___.*
  // pragma RS ap-ctrl ap_start=read_A_31__ap_start ap_done=read_A_31__ap_done ap_idle=read_A_31__ap_idle ap_ready=read_A_31__ap_ready scalar=read_A_31___.*
  // pragma RS ap-ctrl ap_start=read_A_32__ap_start ap_done=read_A_32__ap_done ap_idle=read_A_32__ap_idle ap_ready=read_A_32__ap_ready scalar=read_A_32___.*
  // pragma RS ap-ctrl ap_start=read_A_33__ap_start ap_done=read_A_33__ap_done ap_idle=read_A_33__ap_idle ap_ready=read_A_33__ap_ready scalar=read_A_33___.*
  // pragma RS ap-ctrl ap_start=read_A_34__ap_start ap_done=read_A_34__ap_done ap_idle=read_A_34__ap_idle ap_ready=read_A_34__ap_ready scalar=read_A_34___.*
  // pragma RS ap-ctrl ap_start=read_A_35__ap_start ap_done=read_A_35__ap_done ap_idle=read_A_35__ap_idle ap_ready=read_A_35__ap_ready scalar=read_A_35___.*
  // pragma RS ap-ctrl ap_start=read_A_36__ap_start ap_done=read_A_36__ap_done ap_idle=read_A_36__ap_idle ap_ready=read_A_36__ap_ready scalar=read_A_36___.*
  // pragma RS ap-ctrl ap_start=read_A_37__ap_start ap_done=read_A_37__ap_done ap_idle=read_A_37__ap_idle ap_ready=read_A_37__ap_ready scalar=read_A_37___.*
  // pragma RS ap-ctrl ap_start=read_A_38__ap_start ap_done=read_A_38__ap_done ap_idle=read_A_38__ap_idle ap_ready=read_A_38__ap_ready scalar=read_A_38___.*
  // pragma RS ap-ctrl ap_start=read_A_39__ap_start ap_done=read_A_39__ap_done ap_idle=read_A_39__ap_idle ap_ready=read_A_39__ap_ready scalar=read_A_39___.*
  // pragma RS ap-ctrl ap_start=read_A_40__ap_start ap_done=read_A_40__ap_done ap_idle=read_A_40__ap_idle ap_ready=read_A_40__ap_ready scalar=read_A_40___.*
  // pragma RS ap-ctrl ap_start=read_A_41__ap_start ap_done=read_A_41__ap_done ap_idle=read_A_41__ap_idle ap_ready=read_A_41__ap_ready scalar=read_A_41___.*
  // pragma RS ap-ctrl ap_start=read_A_42__ap_start ap_done=read_A_42__ap_done ap_idle=read_A_42__ap_idle ap_ready=read_A_42__ap_ready scalar=read_A_42___.*
  // pragma RS ap-ctrl ap_start=read_A_43__ap_start ap_done=read_A_43__ap_done ap_idle=read_A_43__ap_idle ap_ready=read_A_43__ap_ready scalar=read_A_43___.*
  // pragma RS ap-ctrl ap_start=read_A_44__ap_start ap_done=read_A_44__ap_done ap_idle=read_A_44__ap_idle ap_ready=read_A_44__ap_ready scalar=read_A_44___.*
  // pragma RS ap-ctrl ap_start=read_A_45__ap_start ap_done=read_A_45__ap_done ap_idle=read_A_45__ap_idle ap_ready=read_A_45__ap_ready scalar=read_A_45___.*
  // pragma RS ap-ctrl ap_start=read_A_46__ap_start ap_done=read_A_46__ap_done ap_idle=read_A_46__ap_idle ap_ready=read_A_46__ap_ready scalar=read_A_46___.*
  // pragma RS ap-ctrl ap_start=read_A_47__ap_start ap_done=read_A_47__ap_done ap_idle=read_A_47__ap_idle ap_ready=read_A_47__ap_ready scalar=read_A_47___.*
  // pragma RS ap-ctrl ap_start=read_X_0__ap_start ap_done=read_X_0__ap_done ap_idle=read_X_0__ap_idle ap_ready=read_X_0__ap_ready scalar=read_X_0___.*
  // pragma RS ap-ctrl ap_start=read_Y_0__ap_start ap_done=read_Y_0__ap_done ap_idle=read_Y_0__ap_idle ap_ready=read_Y_0__ap_ready scalar=read_Y_0___.*
  // pragma RS ap-ctrl ap_start=read_edge_list_ptr_0__ap_start ap_done=read_edge_list_ptr_0__ap_done ap_idle=read_edge_list_ptr_0__ap_idle ap_ready=read_edge_list_ptr_0__ap_ready scalar=read_edge_list_ptr_0___.*
  // pragma RS ap-ctrl ap_start=write_Y_0__ap_start ap_done=write_Y_0__ap_done ap_idle=write_Y_0__ap_idle ap_ready=write_Y_0__ap_ready scalar=write_Y_0___.*

  input ap_clk;
  input ap_rst_n;
  input ap_start;
  output ap_ready;
  output ap_done;
  output ap_idle;
  input [31:0] M;
  input [31:0] P_N;
  input [31:0] alpha_u;
  input [31:0] beta_u;
  input [31:0] NUM_A_LEN;
  input [63:0] edge_list_ch_0;
  input [63:0] edge_list_ch_1;
  input [63:0] edge_list_ch_2;
  input [63:0] edge_list_ch_3;
  input [63:0] edge_list_ch_4;
  input [63:0] edge_list_ch_5;
  input [63:0] edge_list_ch_6;
  input [63:0] edge_list_ch_7;
  input [63:0] edge_list_ch_8;
  input [63:0] edge_list_ch_9;
  input [63:0] edge_list_ch_10;
  input [63:0] edge_list_ch_11;
  input [63:0] edge_list_ch_12;
  input [63:0] edge_list_ch_13;
  input [63:0] edge_list_ch_14;
  input [63:0] edge_list_ch_15;
  input [63:0] edge_list_ch_16;
  input [63:0] edge_list_ch_17;
  input [63:0] edge_list_ch_18;
  input [63:0] edge_list_ch_19;
  input [63:0] edge_list_ch_20;
  input [63:0] edge_list_ch_21;
  input [63:0] edge_list_ch_22;
  input [63:0] edge_list_ch_23;
  input [63:0] edge_list_ch_24;
  input [63:0] edge_list_ch_25;
  input [63:0] edge_list_ch_26;
  input [63:0] edge_list_ch_27;
  input [63:0] edge_list_ch_28;
  input [63:0] edge_list_ch_29;
  input [63:0] edge_list_ch_30;
  input [63:0] edge_list_ch_31;
  input [63:0] edge_list_ch_32;
  input [63:0] edge_list_ch_33;
  input [63:0] edge_list_ch_34;
  input [63:0] edge_list_ch_35;
  input [63:0] edge_list_ch_36;
  input [63:0] edge_list_ch_37;
  input [63:0] edge_list_ch_38;
  input [63:0] edge_list_ch_39;
  input [63:0] edge_list_ch_40;
  input [63:0] edge_list_ch_41;
  input [63:0] edge_list_ch_42;
  input [63:0] edge_list_ch_43;
  input [63:0] edge_list_ch_44;
  input [63:0] edge_list_ch_45;
  input [63:0] edge_list_ch_46;
  input [63:0] edge_list_ch_47;
  input [31:0] K;
  input [63:0] vec_X;
  input [63:0] vec_Y;
  input [31:0] NUM_ITE;
  input [63:0] edge_list_ptr;
  input [63:0] vec_Y_out;
  output [31:0] Arbiter_Y_0___M__q0;
  output [31:0] Arbiter_Y_0___P_N__q0;
  output Arbiter_Y_0__ap_start;
  input Arbiter_Y_0__ap_ready;
  input Arbiter_Y_0__ap_done;
  input Arbiter_Y_0__ap_idle;
  output [31:0] Arbiter_Y_1___M__q0;
  output [31:0] Arbiter_Y_1___P_N__q0;
  output Arbiter_Y_1__ap_start;
  input Arbiter_Y_1__ap_ready;
  input Arbiter_Y_1__ap_done;
  input Arbiter_Y_1__ap_idle;
  output [31:0] Arbiter_Y_2___M__q0;
  output [31:0] Arbiter_Y_2___P_N__q0;
  output Arbiter_Y_2__ap_start;
  input Arbiter_Y_2__ap_ready;
  input Arbiter_Y_2__ap_done;
  input Arbiter_Y_2__ap_idle;
  output [31:0] Arbiter_Y_3___M__q0;
  output [31:0] Arbiter_Y_3___P_N__q0;
  output Arbiter_Y_3__ap_start;
  input Arbiter_Y_3__ap_ready;
  input Arbiter_Y_3__ap_done;
  input Arbiter_Y_3__ap_idle;
  output [31:0] Arbiter_Y_4___M__q0;
  output [31:0] Arbiter_Y_4___P_N__q0;
  output Arbiter_Y_4__ap_start;
  input Arbiter_Y_4__ap_ready;
  input Arbiter_Y_4__ap_done;
  input Arbiter_Y_4__ap_idle;
  output [31:0] Arbiter_Y_5___M__q0;
  output [31:0] Arbiter_Y_5___P_N__q0;
  output Arbiter_Y_5__ap_start;
  input Arbiter_Y_5__ap_ready;
  input Arbiter_Y_5__ap_done;
  input Arbiter_Y_5__ap_idle;
  output [31:0] Arbiter_Y_6___M__q0;
  output [31:0] Arbiter_Y_6___P_N__q0;
  output Arbiter_Y_6__ap_start;
  input Arbiter_Y_6__ap_ready;
  input Arbiter_Y_6__ap_done;
  input Arbiter_Y_6__ap_idle;
  output [31:0] Arbiter_Y_7___M__q0;
  output [31:0] Arbiter_Y_7___P_N__q0;
  output Arbiter_Y_7__ap_start;
  input Arbiter_Y_7__ap_ready;
  input Arbiter_Y_7__ap_done;
  input Arbiter_Y_7__ap_idle;
  output FloatvAddFloatv_0__ap_start;
  output [31:0] FloatvMultConst_0___M__q0;
  output [31:0] FloatvMultConst_0___P_N__q0;
  output [31:0] FloatvMultConst_0___alpha_u__q0;
  output FloatvMultConst_0__ap_start;
  input FloatvMultConst_0__ap_ready;
  input FloatvMultConst_0__ap_done;
  input FloatvMultConst_0__ap_idle;
  output [31:0] FloatvMultConst_1___M__q0;
  output [31:0] FloatvMultConst_1___P_N__q0;
  output [31:0] FloatvMultConst_1___beta_u__q0;
  output FloatvMultConst_1__ap_start;
  input FloatvMultConst_1__ap_ready;
  input FloatvMultConst_1__ap_done;
  input FloatvMultConst_1__ap_idle;
  output Merger_Y_0__ap_start;
  output PEG_Xvec_0__ap_start;
  input PEG_Xvec_0__ap_ready;
  input PEG_Xvec_0__ap_done;
  input PEG_Xvec_0__ap_idle;
  output PEG_Xvec_1__ap_start;
  input PEG_Xvec_1__ap_ready;
  input PEG_Xvec_1__ap_done;
  input PEG_Xvec_1__ap_idle;
  output PEG_Xvec_2__ap_start;
  input PEG_Xvec_2__ap_ready;
  input PEG_Xvec_2__ap_done;
  input PEG_Xvec_2__ap_idle;
  output PEG_Xvec_3__ap_start;
  input PEG_Xvec_3__ap_ready;
  input PEG_Xvec_3__ap_done;
  input PEG_Xvec_3__ap_idle;
  output PEG_Xvec_4__ap_start;
  input PEG_Xvec_4__ap_ready;
  input PEG_Xvec_4__ap_done;
  input PEG_Xvec_4__ap_idle;
  output PEG_Xvec_5__ap_start;
  input PEG_Xvec_5__ap_ready;
  input PEG_Xvec_5__ap_done;
  input PEG_Xvec_5__ap_idle;
  output PEG_Xvec_6__ap_start;
  input PEG_Xvec_6__ap_ready;
  input PEG_Xvec_6__ap_done;
  input PEG_Xvec_6__ap_idle;
  output PEG_Xvec_7__ap_start;
  input PEG_Xvec_7__ap_ready;
  input PEG_Xvec_7__ap_done;
  input PEG_Xvec_7__ap_idle;
  output PEG_Xvec_8__ap_start;
  input PEG_Xvec_8__ap_ready;
  input PEG_Xvec_8__ap_done;
  input PEG_Xvec_8__ap_idle;
  output PEG_Xvec_9__ap_start;
  input PEG_Xvec_9__ap_ready;
  input PEG_Xvec_9__ap_done;
  input PEG_Xvec_9__ap_idle;
  output PEG_Xvec_10__ap_start;
  input PEG_Xvec_10__ap_ready;
  input PEG_Xvec_10__ap_done;
  input PEG_Xvec_10__ap_idle;
  output PEG_Xvec_11__ap_start;
  input PEG_Xvec_11__ap_ready;
  input PEG_Xvec_11__ap_done;
  input PEG_Xvec_11__ap_idle;
  output PEG_Xvec_12__ap_start;
  input PEG_Xvec_12__ap_ready;
  input PEG_Xvec_12__ap_done;
  input PEG_Xvec_12__ap_idle;
  output PEG_Xvec_13__ap_start;
  input PEG_Xvec_13__ap_ready;
  input PEG_Xvec_13__ap_done;
  input PEG_Xvec_13__ap_idle;
  output PEG_Xvec_14__ap_start;
  input PEG_Xvec_14__ap_ready;
  input PEG_Xvec_14__ap_done;
  input PEG_Xvec_14__ap_idle;
  output PEG_Xvec_15__ap_start;
  input PEG_Xvec_15__ap_ready;
  input PEG_Xvec_15__ap_done;
  input PEG_Xvec_15__ap_idle;
  output PEG_Xvec_16__ap_start;
  input PEG_Xvec_16__ap_ready;
  input PEG_Xvec_16__ap_done;
  input PEG_Xvec_16__ap_idle;
  output PEG_Xvec_17__ap_start;
  input PEG_Xvec_17__ap_ready;
  input PEG_Xvec_17__ap_done;
  input PEG_Xvec_17__ap_idle;
  output PEG_Xvec_18__ap_start;
  input PEG_Xvec_18__ap_ready;
  input PEG_Xvec_18__ap_done;
  input PEG_Xvec_18__ap_idle;
  output PEG_Xvec_19__ap_start;
  input PEG_Xvec_19__ap_ready;
  input PEG_Xvec_19__ap_done;
  input PEG_Xvec_19__ap_idle;
  output PEG_Xvec_20__ap_start;
  input PEG_Xvec_20__ap_ready;
  input PEG_Xvec_20__ap_done;
  input PEG_Xvec_20__ap_idle;
  output PEG_Xvec_21__ap_start;
  input PEG_Xvec_21__ap_ready;
  input PEG_Xvec_21__ap_done;
  input PEG_Xvec_21__ap_idle;
  output PEG_Xvec_22__ap_start;
  input PEG_Xvec_22__ap_ready;
  input PEG_Xvec_22__ap_done;
  input PEG_Xvec_22__ap_idle;
  output PEG_Xvec_23__ap_start;
  input PEG_Xvec_23__ap_ready;
  input PEG_Xvec_23__ap_done;
  input PEG_Xvec_23__ap_idle;
  output PEG_Xvec_24__ap_start;
  input PEG_Xvec_24__ap_ready;
  input PEG_Xvec_24__ap_done;
  input PEG_Xvec_24__ap_idle;
  output PEG_Xvec_25__ap_start;
  input PEG_Xvec_25__ap_ready;
  input PEG_Xvec_25__ap_done;
  input PEG_Xvec_25__ap_idle;
  output PEG_Xvec_26__ap_start;
  input PEG_Xvec_26__ap_ready;
  input PEG_Xvec_26__ap_done;
  input PEG_Xvec_26__ap_idle;
  output PEG_Xvec_27__ap_start;
  input PEG_Xvec_27__ap_ready;
  input PEG_Xvec_27__ap_done;
  input PEG_Xvec_27__ap_idle;
  output PEG_Xvec_28__ap_start;
  input PEG_Xvec_28__ap_ready;
  input PEG_Xvec_28__ap_done;
  input PEG_Xvec_28__ap_idle;
  output PEG_Xvec_29__ap_start;
  input PEG_Xvec_29__ap_ready;
  input PEG_Xvec_29__ap_done;
  input PEG_Xvec_29__ap_idle;
  output PEG_Xvec_30__ap_start;
  input PEG_Xvec_30__ap_ready;
  input PEG_Xvec_30__ap_done;
  input PEG_Xvec_30__ap_idle;
  output PEG_Xvec_31__ap_start;
  input PEG_Xvec_31__ap_ready;
  input PEG_Xvec_31__ap_done;
  input PEG_Xvec_31__ap_idle;
  output PEG_Xvec_32__ap_start;
  input PEG_Xvec_32__ap_ready;
  input PEG_Xvec_32__ap_done;
  input PEG_Xvec_32__ap_idle;
  output PEG_Xvec_33__ap_start;
  input PEG_Xvec_33__ap_ready;
  input PEG_Xvec_33__ap_done;
  input PEG_Xvec_33__ap_idle;
  output PEG_Xvec_34__ap_start;
  input PEG_Xvec_34__ap_ready;
  input PEG_Xvec_34__ap_done;
  input PEG_Xvec_34__ap_idle;
  output PEG_Xvec_35__ap_start;
  input PEG_Xvec_35__ap_ready;
  input PEG_Xvec_35__ap_done;
  input PEG_Xvec_35__ap_idle;
  output PEG_Xvec_36__ap_start;
  input PEG_Xvec_36__ap_ready;
  input PEG_Xvec_36__ap_done;
  input PEG_Xvec_36__ap_idle;
  output PEG_Xvec_37__ap_start;
  input PEG_Xvec_37__ap_ready;
  input PEG_Xvec_37__ap_done;
  input PEG_Xvec_37__ap_idle;
  output PEG_Xvec_38__ap_start;
  input PEG_Xvec_38__ap_ready;
  input PEG_Xvec_38__ap_done;
  input PEG_Xvec_38__ap_idle;
  output PEG_Xvec_39__ap_start;
  input PEG_Xvec_39__ap_ready;
  input PEG_Xvec_39__ap_done;
  input PEG_Xvec_39__ap_idle;
  output PEG_Xvec_40__ap_start;
  input PEG_Xvec_40__ap_ready;
  input PEG_Xvec_40__ap_done;
  input PEG_Xvec_40__ap_idle;
  output PEG_Xvec_41__ap_start;
  input PEG_Xvec_41__ap_ready;
  input PEG_Xvec_41__ap_done;
  input PEG_Xvec_41__ap_idle;
  output PEG_Xvec_42__ap_start;
  input PEG_Xvec_42__ap_ready;
  input PEG_Xvec_42__ap_done;
  input PEG_Xvec_42__ap_idle;
  output PEG_Xvec_43__ap_start;
  input PEG_Xvec_43__ap_ready;
  input PEG_Xvec_43__ap_done;
  input PEG_Xvec_43__ap_idle;
  output PEG_Xvec_44__ap_start;
  input PEG_Xvec_44__ap_ready;
  input PEG_Xvec_44__ap_done;
  input PEG_Xvec_44__ap_idle;
  output PEG_Xvec_45__ap_start;
  input PEG_Xvec_45__ap_ready;
  input PEG_Xvec_45__ap_done;
  input PEG_Xvec_45__ap_idle;
  output PEG_Xvec_46__ap_start;
  input PEG_Xvec_46__ap_ready;
  input PEG_Xvec_46__ap_done;
  input PEG_Xvec_46__ap_idle;
  output PEG_Xvec_47__ap_start;
  input PEG_Xvec_47__ap_ready;
  input PEG_Xvec_47__ap_done;
  input PEG_Xvec_47__ap_idle;
  output PEG_Yvec_0__ap_start;
  input PEG_Yvec_0__ap_ready;
  input PEG_Yvec_0__ap_done;
  input PEG_Yvec_0__ap_idle;
  output PEG_Yvec_1__ap_start;
  input PEG_Yvec_1__ap_ready;
  input PEG_Yvec_1__ap_done;
  input PEG_Yvec_1__ap_idle;
  output PEG_Yvec_2__ap_start;
  input PEG_Yvec_2__ap_ready;
  input PEG_Yvec_2__ap_done;
  input PEG_Yvec_2__ap_idle;
  output PEG_Yvec_3__ap_start;
  input PEG_Yvec_3__ap_ready;
  input PEG_Yvec_3__ap_done;
  input PEG_Yvec_3__ap_idle;
  output PEG_Yvec_4__ap_start;
  input PEG_Yvec_4__ap_ready;
  input PEG_Yvec_4__ap_done;
  input PEG_Yvec_4__ap_idle;
  output PEG_Yvec_5__ap_start;
  input PEG_Yvec_5__ap_ready;
  input PEG_Yvec_5__ap_done;
  input PEG_Yvec_5__ap_idle;
  output PEG_Yvec_6__ap_start;
  input PEG_Yvec_6__ap_ready;
  input PEG_Yvec_6__ap_done;
  input PEG_Yvec_6__ap_idle;
  output PEG_Yvec_7__ap_start;
  input PEG_Yvec_7__ap_ready;
  input PEG_Yvec_7__ap_done;
  input PEG_Yvec_7__ap_idle;
  output PEG_Yvec_8__ap_start;
  input PEG_Yvec_8__ap_ready;
  input PEG_Yvec_8__ap_done;
  input PEG_Yvec_8__ap_idle;
  output PEG_Yvec_9__ap_start;
  input PEG_Yvec_9__ap_ready;
  input PEG_Yvec_9__ap_done;
  input PEG_Yvec_9__ap_idle;
  output PEG_Yvec_10__ap_start;
  input PEG_Yvec_10__ap_ready;
  input PEG_Yvec_10__ap_done;
  input PEG_Yvec_10__ap_idle;
  output PEG_Yvec_11__ap_start;
  input PEG_Yvec_11__ap_ready;
  input PEG_Yvec_11__ap_done;
  input PEG_Yvec_11__ap_idle;
  output PEG_Yvec_12__ap_start;
  input PEG_Yvec_12__ap_ready;
  input PEG_Yvec_12__ap_done;
  input PEG_Yvec_12__ap_idle;
  output PEG_Yvec_13__ap_start;
  input PEG_Yvec_13__ap_ready;
  input PEG_Yvec_13__ap_done;
  input PEG_Yvec_13__ap_idle;
  output PEG_Yvec_14__ap_start;
  input PEG_Yvec_14__ap_ready;
  input PEG_Yvec_14__ap_done;
  input PEG_Yvec_14__ap_idle;
  output PEG_Yvec_15__ap_start;
  input PEG_Yvec_15__ap_ready;
  input PEG_Yvec_15__ap_done;
  input PEG_Yvec_15__ap_idle;
  output PEG_Yvec_16__ap_start;
  input PEG_Yvec_16__ap_ready;
  input PEG_Yvec_16__ap_done;
  input PEG_Yvec_16__ap_idle;
  output PEG_Yvec_17__ap_start;
  input PEG_Yvec_17__ap_ready;
  input PEG_Yvec_17__ap_done;
  input PEG_Yvec_17__ap_idle;
  output PEG_Yvec_18__ap_start;
  input PEG_Yvec_18__ap_ready;
  input PEG_Yvec_18__ap_done;
  input PEG_Yvec_18__ap_idle;
  output PEG_Yvec_19__ap_start;
  input PEG_Yvec_19__ap_ready;
  input PEG_Yvec_19__ap_done;
  input PEG_Yvec_19__ap_idle;
  output PEG_Yvec_20__ap_start;
  input PEG_Yvec_20__ap_ready;
  input PEG_Yvec_20__ap_done;
  input PEG_Yvec_20__ap_idle;
  output PEG_Yvec_21__ap_start;
  input PEG_Yvec_21__ap_ready;
  input PEG_Yvec_21__ap_done;
  input PEG_Yvec_21__ap_idle;
  output PEG_Yvec_22__ap_start;
  input PEG_Yvec_22__ap_ready;
  input PEG_Yvec_22__ap_done;
  input PEG_Yvec_22__ap_idle;
  output PEG_Yvec_23__ap_start;
  input PEG_Yvec_23__ap_ready;
  input PEG_Yvec_23__ap_done;
  input PEG_Yvec_23__ap_idle;
  output PEG_Yvec_24__ap_start;
  input PEG_Yvec_24__ap_ready;
  input PEG_Yvec_24__ap_done;
  input PEG_Yvec_24__ap_idle;
  output PEG_Yvec_25__ap_start;
  input PEG_Yvec_25__ap_ready;
  input PEG_Yvec_25__ap_done;
  input PEG_Yvec_25__ap_idle;
  output PEG_Yvec_26__ap_start;
  input PEG_Yvec_26__ap_ready;
  input PEG_Yvec_26__ap_done;
  input PEG_Yvec_26__ap_idle;
  output PEG_Yvec_27__ap_start;
  input PEG_Yvec_27__ap_ready;
  input PEG_Yvec_27__ap_done;
  input PEG_Yvec_27__ap_idle;
  output PEG_Yvec_28__ap_start;
  input PEG_Yvec_28__ap_ready;
  input PEG_Yvec_28__ap_done;
  input PEG_Yvec_28__ap_idle;
  output PEG_Yvec_29__ap_start;
  input PEG_Yvec_29__ap_ready;
  input PEG_Yvec_29__ap_done;
  input PEG_Yvec_29__ap_idle;
  output PEG_Yvec_30__ap_start;
  input PEG_Yvec_30__ap_ready;
  input PEG_Yvec_30__ap_done;
  input PEG_Yvec_30__ap_idle;
  output PEG_Yvec_31__ap_start;
  input PEG_Yvec_31__ap_ready;
  input PEG_Yvec_31__ap_done;
  input PEG_Yvec_31__ap_idle;
  output PEG_Yvec_32__ap_start;
  input PEG_Yvec_32__ap_ready;
  input PEG_Yvec_32__ap_done;
  input PEG_Yvec_32__ap_idle;
  output PEG_Yvec_33__ap_start;
  input PEG_Yvec_33__ap_ready;
  input PEG_Yvec_33__ap_done;
  input PEG_Yvec_33__ap_idle;
  output PEG_Yvec_34__ap_start;
  input PEG_Yvec_34__ap_ready;
  input PEG_Yvec_34__ap_done;
  input PEG_Yvec_34__ap_idle;
  output PEG_Yvec_35__ap_start;
  input PEG_Yvec_35__ap_ready;
  input PEG_Yvec_35__ap_done;
  input PEG_Yvec_35__ap_idle;
  output PEG_Yvec_36__ap_start;
  input PEG_Yvec_36__ap_ready;
  input PEG_Yvec_36__ap_done;
  input PEG_Yvec_36__ap_idle;
  output PEG_Yvec_37__ap_start;
  input PEG_Yvec_37__ap_ready;
  input PEG_Yvec_37__ap_done;
  input PEG_Yvec_37__ap_idle;
  output PEG_Yvec_38__ap_start;
  input PEG_Yvec_38__ap_ready;
  input PEG_Yvec_38__ap_done;
  input PEG_Yvec_38__ap_idle;
  output PEG_Yvec_39__ap_start;
  input PEG_Yvec_39__ap_ready;
  input PEG_Yvec_39__ap_done;
  input PEG_Yvec_39__ap_idle;
  output PEG_Yvec_40__ap_start;
  input PEG_Yvec_40__ap_ready;
  input PEG_Yvec_40__ap_done;
  input PEG_Yvec_40__ap_idle;
  output PEG_Yvec_41__ap_start;
  input PEG_Yvec_41__ap_ready;
  input PEG_Yvec_41__ap_done;
  input PEG_Yvec_41__ap_idle;
  output PEG_Yvec_42__ap_start;
  input PEG_Yvec_42__ap_ready;
  input PEG_Yvec_42__ap_done;
  input PEG_Yvec_42__ap_idle;
  output PEG_Yvec_43__ap_start;
  input PEG_Yvec_43__ap_ready;
  input PEG_Yvec_43__ap_done;
  input PEG_Yvec_43__ap_idle;
  output PEG_Yvec_44__ap_start;
  input PEG_Yvec_44__ap_ready;
  input PEG_Yvec_44__ap_done;
  input PEG_Yvec_44__ap_idle;
  output PEG_Yvec_45__ap_start;
  input PEG_Yvec_45__ap_ready;
  input PEG_Yvec_45__ap_done;
  input PEG_Yvec_45__ap_idle;
  output PEG_Yvec_46__ap_start;
  input PEG_Yvec_46__ap_ready;
  input PEG_Yvec_46__ap_done;
  input PEG_Yvec_46__ap_idle;
  output PEG_Yvec_47__ap_start;
  input PEG_Yvec_47__ap_ready;
  input PEG_Yvec_47__ap_done;
  input PEG_Yvec_47__ap_idle;
  output black_hole_float_v16_0__ap_start;
  output black_hole_int_0__ap_start;
  output [31:0] read_A_0___NUM_A_LEN__q0;
  output [31:0] read_A_0___P_N__q0;
  output [63:0] read_A_0___edge_list_ch_0__q0;
  output read_A_0__ap_start;
  input read_A_0__ap_ready;
  input read_A_0__ap_done;
  input read_A_0__ap_idle;
  output [31:0] read_A_1___NUM_A_LEN__q0;
  output [31:0] read_A_1___P_N__q0;
  output [63:0] read_A_1___edge_list_ch_1__q0;
  output read_A_1__ap_start;
  input read_A_1__ap_ready;
  input read_A_1__ap_done;
  input read_A_1__ap_idle;
  output [31:0] read_A_2___NUM_A_LEN__q0;
  output [31:0] read_A_2___P_N__q0;
  output [63:0] read_A_2___edge_list_ch_2__q0;
  output read_A_2__ap_start;
  input read_A_2__ap_ready;
  input read_A_2__ap_done;
  input read_A_2__ap_idle;
  output [31:0] read_A_3___NUM_A_LEN__q0;
  output [31:0] read_A_3___P_N__q0;
  output [63:0] read_A_3___edge_list_ch_3__q0;
  output read_A_3__ap_start;
  input read_A_3__ap_ready;
  input read_A_3__ap_done;
  input read_A_3__ap_idle;
  output [31:0] read_A_4___NUM_A_LEN__q0;
  output [31:0] read_A_4___P_N__q0;
  output [63:0] read_A_4___edge_list_ch_4__q0;
  output read_A_4__ap_start;
  input read_A_4__ap_ready;
  input read_A_4__ap_done;
  input read_A_4__ap_idle;
  output [31:0] read_A_5___NUM_A_LEN__q0;
  output [31:0] read_A_5___P_N__q0;
  output [63:0] read_A_5___edge_list_ch_5__q0;
  output read_A_5__ap_start;
  input read_A_5__ap_ready;
  input read_A_5__ap_done;
  input read_A_5__ap_idle;
  output [31:0] read_A_6___NUM_A_LEN__q0;
  output [31:0] read_A_6___P_N__q0;
  output [63:0] read_A_6___edge_list_ch_6__q0;
  output read_A_6__ap_start;
  input read_A_6__ap_ready;
  input read_A_6__ap_done;
  input read_A_6__ap_idle;
  output [31:0] read_A_7___NUM_A_LEN__q0;
  output [31:0] read_A_7___P_N__q0;
  output [63:0] read_A_7___edge_list_ch_7__q0;
  output read_A_7__ap_start;
  input read_A_7__ap_ready;
  input read_A_7__ap_done;
  input read_A_7__ap_idle;
  output [31:0] read_A_8___NUM_A_LEN__q0;
  output [31:0] read_A_8___P_N__q0;
  output [63:0] read_A_8___edge_list_ch_8__q0;
  output read_A_8__ap_start;
  input read_A_8__ap_ready;
  input read_A_8__ap_done;
  input read_A_8__ap_idle;
  output [31:0] read_A_9___NUM_A_LEN__q0;
  output [31:0] read_A_9___P_N__q0;
  output [63:0] read_A_9___edge_list_ch_9__q0;
  output read_A_9__ap_start;
  input read_A_9__ap_ready;
  input read_A_9__ap_done;
  input read_A_9__ap_idle;
  output [31:0] read_A_10___NUM_A_LEN__q0;
  output [31:0] read_A_10___P_N__q0;
  output [63:0] read_A_10___edge_list_ch_10__q0;
  output read_A_10__ap_start;
  input read_A_10__ap_ready;
  input read_A_10__ap_done;
  input read_A_10__ap_idle;
  output [31:0] read_A_11___NUM_A_LEN__q0;
  output [31:0] read_A_11___P_N__q0;
  output [63:0] read_A_11___edge_list_ch_11__q0;
  output read_A_11__ap_start;
  input read_A_11__ap_ready;
  input read_A_11__ap_done;
  input read_A_11__ap_idle;
  output [31:0] read_A_12___NUM_A_LEN__q0;
  output [31:0] read_A_12___P_N__q0;
  output [63:0] read_A_12___edge_list_ch_12__q0;
  output read_A_12__ap_start;
  input read_A_12__ap_ready;
  input read_A_12__ap_done;
  input read_A_12__ap_idle;
  output [31:0] read_A_13___NUM_A_LEN__q0;
  output [31:0] read_A_13___P_N__q0;
  output [63:0] read_A_13___edge_list_ch_13__q0;
  output read_A_13__ap_start;
  input read_A_13__ap_ready;
  input read_A_13__ap_done;
  input read_A_13__ap_idle;
  output [31:0] read_A_14___NUM_A_LEN__q0;
  output [31:0] read_A_14___P_N__q0;
  output [63:0] read_A_14___edge_list_ch_14__q0;
  output read_A_14__ap_start;
  input read_A_14__ap_ready;
  input read_A_14__ap_done;
  input read_A_14__ap_idle;
  output [31:0] read_A_15___NUM_A_LEN__q0;
  output [31:0] read_A_15___P_N__q0;
  output [63:0] read_A_15___edge_list_ch_15__q0;
  output read_A_15__ap_start;
  input read_A_15__ap_ready;
  input read_A_15__ap_done;
  input read_A_15__ap_idle;
  output [31:0] read_A_16___NUM_A_LEN__q0;
  output [31:0] read_A_16___P_N__q0;
  output [63:0] read_A_16___edge_list_ch_16__q0;
  output read_A_16__ap_start;
  input read_A_16__ap_ready;
  input read_A_16__ap_done;
  input read_A_16__ap_idle;
  output [31:0] read_A_17___NUM_A_LEN__q0;
  output [31:0] read_A_17___P_N__q0;
  output [63:0] read_A_17___edge_list_ch_17__q0;
  output read_A_17__ap_start;
  input read_A_17__ap_ready;
  input read_A_17__ap_done;
  input read_A_17__ap_idle;
  output [31:0] read_A_18___NUM_A_LEN__q0;
  output [31:0] read_A_18___P_N__q0;
  output [63:0] read_A_18___edge_list_ch_18__q0;
  output read_A_18__ap_start;
  input read_A_18__ap_ready;
  input read_A_18__ap_done;
  input read_A_18__ap_idle;
  output [31:0] read_A_19___NUM_A_LEN__q0;
  output [31:0] read_A_19___P_N__q0;
  output [63:0] read_A_19___edge_list_ch_19__q0;
  output read_A_19__ap_start;
  input read_A_19__ap_ready;
  input read_A_19__ap_done;
  input read_A_19__ap_idle;
  output [31:0] read_A_20___NUM_A_LEN__q0;
  output [31:0] read_A_20___P_N__q0;
  output [63:0] read_A_20___edge_list_ch_20__q0;
  output read_A_20__ap_start;
  input read_A_20__ap_ready;
  input read_A_20__ap_done;
  input read_A_20__ap_idle;
  output [31:0] read_A_21___NUM_A_LEN__q0;
  output [31:0] read_A_21___P_N__q0;
  output [63:0] read_A_21___edge_list_ch_21__q0;
  output read_A_21__ap_start;
  input read_A_21__ap_ready;
  input read_A_21__ap_done;
  input read_A_21__ap_idle;
  output [31:0] read_A_22___NUM_A_LEN__q0;
  output [31:0] read_A_22___P_N__q0;
  output [63:0] read_A_22___edge_list_ch_22__q0;
  output read_A_22__ap_start;
  input read_A_22__ap_ready;
  input read_A_22__ap_done;
  input read_A_22__ap_idle;
  output [31:0] read_A_23___NUM_A_LEN__q0;
  output [31:0] read_A_23___P_N__q0;
  output [63:0] read_A_23___edge_list_ch_23__q0;
  output read_A_23__ap_start;
  input read_A_23__ap_ready;
  input read_A_23__ap_done;
  input read_A_23__ap_idle;
  output [31:0] read_A_24___NUM_A_LEN__q0;
  output [31:0] read_A_24___P_N__q0;
  output [63:0] read_A_24___edge_list_ch_24__q0;
  output read_A_24__ap_start;
  input read_A_24__ap_ready;
  input read_A_24__ap_done;
  input read_A_24__ap_idle;
  output [31:0] read_A_25___NUM_A_LEN__q0;
  output [31:0] read_A_25___P_N__q0;
  output [63:0] read_A_25___edge_list_ch_25__q0;
  output read_A_25__ap_start;
  input read_A_25__ap_ready;
  input read_A_25__ap_done;
  input read_A_25__ap_idle;
  output [31:0] read_A_26___NUM_A_LEN__q0;
  output [31:0] read_A_26___P_N__q0;
  output [63:0] read_A_26___edge_list_ch_26__q0;
  output read_A_26__ap_start;
  input read_A_26__ap_ready;
  input read_A_26__ap_done;
  input read_A_26__ap_idle;
  output [31:0] read_A_27___NUM_A_LEN__q0;
  output [31:0] read_A_27___P_N__q0;
  output [63:0] read_A_27___edge_list_ch_27__q0;
  output read_A_27__ap_start;
  input read_A_27__ap_ready;
  input read_A_27__ap_done;
  input read_A_27__ap_idle;
  output [31:0] read_A_28___NUM_A_LEN__q0;
  output [31:0] read_A_28___P_N__q0;
  output [63:0] read_A_28___edge_list_ch_28__q0;
  output read_A_28__ap_start;
  input read_A_28__ap_ready;
  input read_A_28__ap_done;
  input read_A_28__ap_idle;
  output [31:0] read_A_29___NUM_A_LEN__q0;
  output [31:0] read_A_29___P_N__q0;
  output [63:0] read_A_29___edge_list_ch_29__q0;
  output read_A_29__ap_start;
  input read_A_29__ap_ready;
  input read_A_29__ap_done;
  input read_A_29__ap_idle;
  output [31:0] read_A_30___NUM_A_LEN__q0;
  output [31:0] read_A_30___P_N__q0;
  output [63:0] read_A_30___edge_list_ch_30__q0;
  output read_A_30__ap_start;
  input read_A_30__ap_ready;
  input read_A_30__ap_done;
  input read_A_30__ap_idle;
  output [31:0] read_A_31___NUM_A_LEN__q0;
  output [31:0] read_A_31___P_N__q0;
  output [63:0] read_A_31___edge_list_ch_31__q0;
  output read_A_31__ap_start;
  input read_A_31__ap_ready;
  input read_A_31__ap_done;
  input read_A_31__ap_idle;
  output [31:0] read_A_32___NUM_A_LEN__q0;
  output [31:0] read_A_32___P_N__q0;
  output [63:0] read_A_32___edge_list_ch_32__q0;
  output read_A_32__ap_start;
  input read_A_32__ap_ready;
  input read_A_32__ap_done;
  input read_A_32__ap_idle;
  output [31:0] read_A_33___NUM_A_LEN__q0;
  output [31:0] read_A_33___P_N__q0;
  output [63:0] read_A_33___edge_list_ch_33__q0;
  output read_A_33__ap_start;
  input read_A_33__ap_ready;
  input read_A_33__ap_done;
  input read_A_33__ap_idle;
  output [31:0] read_A_34___NUM_A_LEN__q0;
  output [31:0] read_A_34___P_N__q0;
  output [63:0] read_A_34___edge_list_ch_34__q0;
  output read_A_34__ap_start;
  input read_A_34__ap_ready;
  input read_A_34__ap_done;
  input read_A_34__ap_idle;
  output [31:0] read_A_35___NUM_A_LEN__q0;
  output [31:0] read_A_35___P_N__q0;
  output [63:0] read_A_35___edge_list_ch_35__q0;
  output read_A_35__ap_start;
  input read_A_35__ap_ready;
  input read_A_35__ap_done;
  input read_A_35__ap_idle;
  output [31:0] read_A_36___NUM_A_LEN__q0;
  output [31:0] read_A_36___P_N__q0;
  output [63:0] read_A_36___edge_list_ch_36__q0;
  output read_A_36__ap_start;
  input read_A_36__ap_ready;
  input read_A_36__ap_done;
  input read_A_36__ap_idle;
  output [31:0] read_A_37___NUM_A_LEN__q0;
  output [31:0] read_A_37___P_N__q0;
  output [63:0] read_A_37___edge_list_ch_37__q0;
  output read_A_37__ap_start;
  input read_A_37__ap_ready;
  input read_A_37__ap_done;
  input read_A_37__ap_idle;
  output [31:0] read_A_38___NUM_A_LEN__q0;
  output [31:0] read_A_38___P_N__q0;
  output [63:0] read_A_38___edge_list_ch_38__q0;
  output read_A_38__ap_start;
  input read_A_38__ap_ready;
  input read_A_38__ap_done;
  input read_A_38__ap_idle;
  output [31:0] read_A_39___NUM_A_LEN__q0;
  output [31:0] read_A_39___P_N__q0;
  output [63:0] read_A_39___edge_list_ch_39__q0;
  output read_A_39__ap_start;
  input read_A_39__ap_ready;
  input read_A_39__ap_done;
  input read_A_39__ap_idle;
  output [31:0] read_A_40___NUM_A_LEN__q0;
  output [31:0] read_A_40___P_N__q0;
  output [63:0] read_A_40___edge_list_ch_40__q0;
  output read_A_40__ap_start;
  input read_A_40__ap_ready;
  input read_A_40__ap_done;
  input read_A_40__ap_idle;
  output [31:0] read_A_41___NUM_A_LEN__q0;
  output [31:0] read_A_41___P_N__q0;
  output [63:0] read_A_41___edge_list_ch_41__q0;
  output read_A_41__ap_start;
  input read_A_41__ap_ready;
  input read_A_41__ap_done;
  input read_A_41__ap_idle;
  output [31:0] read_A_42___NUM_A_LEN__q0;
  output [31:0] read_A_42___P_N__q0;
  output [63:0] read_A_42___edge_list_ch_42__q0;
  output read_A_42__ap_start;
  input read_A_42__ap_ready;
  input read_A_42__ap_done;
  input read_A_42__ap_idle;
  output [31:0] read_A_43___NUM_A_LEN__q0;
  output [31:0] read_A_43___P_N__q0;
  output [63:0] read_A_43___edge_list_ch_43__q0;
  output read_A_43__ap_start;
  input read_A_43__ap_ready;
  input read_A_43__ap_done;
  input read_A_43__ap_idle;
  output [31:0] read_A_44___NUM_A_LEN__q0;
  output [31:0] read_A_44___P_N__q0;
  output [63:0] read_A_44___edge_list_ch_44__q0;
  output read_A_44__ap_start;
  input read_A_44__ap_ready;
  input read_A_44__ap_done;
  input read_A_44__ap_idle;
  output [31:0] read_A_45___NUM_A_LEN__q0;
  output [31:0] read_A_45___P_N__q0;
  output [63:0] read_A_45___edge_list_ch_45__q0;
  output read_A_45__ap_start;
  input read_A_45__ap_ready;
  input read_A_45__ap_done;
  input read_A_45__ap_idle;
  output [31:0] read_A_46___NUM_A_LEN__q0;
  output [31:0] read_A_46___P_N__q0;
  output [63:0] read_A_46___edge_list_ch_46__q0;
  output read_A_46__ap_start;
  input read_A_46__ap_ready;
  input read_A_46__ap_done;
  input read_A_46__ap_idle;
  output [31:0] read_A_47___NUM_A_LEN__q0;
  output [31:0] read_A_47___P_N__q0;
  output [63:0] read_A_47___edge_list_ch_47__q0;
  output read_A_47__ap_start;
  input read_A_47__ap_ready;
  input read_A_47__ap_done;
  input read_A_47__ap_idle;
  output [31:0] read_X_0___K__q0;
  output [31:0] read_X_0___P_N__q0;
  output [63:0] read_X_0___vec_X__q0;
  output read_X_0__ap_start;
  input read_X_0__ap_ready;
  input read_X_0__ap_done;
  input read_X_0__ap_idle;
  output [31:0] read_Y_0___M__q0;
  output [31:0] read_Y_0___P_N__q0;
  output [63:0] read_Y_0___vec_Y__q0;
  output read_Y_0__ap_start;
  input read_Y_0__ap_ready;
  input read_Y_0__ap_done;
  input read_Y_0__ap_idle;
  output [31:0] read_edge_list_ptr_0___K__q0;
  output [31:0] read_edge_list_ptr_0___M__q0;
  output [31:0] read_edge_list_ptr_0___NUM_ITE__q0;
  output [31:0] read_edge_list_ptr_0___P_N__q0;
  output [63:0] read_edge_list_ptr_0___edge_list_ptr__q0;
  output read_edge_list_ptr_0__ap_start;
  input read_edge_list_ptr_0__ap_ready;
  input read_edge_list_ptr_0__ap_done;
  input read_edge_list_ptr_0__ap_idle;
  output [31:0] write_Y_0___M__q0;
  output [31:0] write_Y_0___P_N__q0;
  output [63:0] write_Y_0___vec_Y_out__q0;
  output write_Y_0__ap_start;
  input write_Y_0__ap_ready;
  input write_Y_0__ap_done;
  input write_Y_0__ap_idle;
  wire [31:0] Arbiter_Y_0___M__q0;
  wire [31:0] Arbiter_Y_0___P_N__q0;
  wire Arbiter_Y_0__ap_start_global__q0;
  wire Arbiter_Y_0__is_done__q0;
  wire Arbiter_Y_0__ap_done_global__q0;
  wire Arbiter_Y_0__ap_start;
  wire Arbiter_Y_0__ap_ready;
  wire Arbiter_Y_0__ap_done;
  wire Arbiter_Y_0__ap_idle;
  reg [1:0] Arbiter_Y_0__state;
  wire [31:0] Arbiter_Y_1___M__q0;
  wire [31:0] Arbiter_Y_1___P_N__q0;
  wire Arbiter_Y_1__ap_start_global__q0;
  wire Arbiter_Y_1__is_done__q0;
  wire Arbiter_Y_1__ap_done_global__q0;
  wire Arbiter_Y_1__ap_start;
  wire Arbiter_Y_1__ap_ready;
  wire Arbiter_Y_1__ap_done;
  wire Arbiter_Y_1__ap_idle;
  reg [1:0] Arbiter_Y_1__state;
  wire [31:0] Arbiter_Y_2___M__q0;
  wire [31:0] Arbiter_Y_2___P_N__q0;
  wire Arbiter_Y_2__ap_start_global__q0;
  wire Arbiter_Y_2__is_done__q0;
  wire Arbiter_Y_2__ap_done_global__q0;
  wire Arbiter_Y_2__ap_start;
  wire Arbiter_Y_2__ap_ready;
  wire Arbiter_Y_2__ap_done;
  wire Arbiter_Y_2__ap_idle;
  reg [1:0] Arbiter_Y_2__state;
  wire [31:0] Arbiter_Y_3___M__q0;
  wire [31:0] Arbiter_Y_3___P_N__q0;
  wire Arbiter_Y_3__ap_start_global__q0;
  wire Arbiter_Y_3__is_done__q0;
  wire Arbiter_Y_3__ap_done_global__q0;
  wire Arbiter_Y_3__ap_start;
  wire Arbiter_Y_3__ap_ready;
  wire Arbiter_Y_3__ap_done;
  wire Arbiter_Y_3__ap_idle;
  reg [1:0] Arbiter_Y_3__state;
  wire [31:0] Arbiter_Y_4___M__q0;
  wire [31:0] Arbiter_Y_4___P_N__q0;
  wire Arbiter_Y_4__ap_start_global__q0;
  wire Arbiter_Y_4__is_done__q0;
  wire Arbiter_Y_4__ap_done_global__q0;
  wire Arbiter_Y_4__ap_start;
  wire Arbiter_Y_4__ap_ready;
  wire Arbiter_Y_4__ap_done;
  wire Arbiter_Y_4__ap_idle;
  reg [1:0] Arbiter_Y_4__state;
  wire [31:0] Arbiter_Y_5___M__q0;
  wire [31:0] Arbiter_Y_5___P_N__q0;
  wire Arbiter_Y_5__ap_start_global__q0;
  wire Arbiter_Y_5__is_done__q0;
  wire Arbiter_Y_5__ap_done_global__q0;
  wire Arbiter_Y_5__ap_start;
  wire Arbiter_Y_5__ap_ready;
  wire Arbiter_Y_5__ap_done;
  wire Arbiter_Y_5__ap_idle;
  reg [1:0] Arbiter_Y_5__state;
  wire [31:0] Arbiter_Y_6___M__q0;
  wire [31:0] Arbiter_Y_6___P_N__q0;
  wire Arbiter_Y_6__ap_start_global__q0;
  wire Arbiter_Y_6__is_done__q0;
  wire Arbiter_Y_6__ap_done_global__q0;
  wire Arbiter_Y_6__ap_start;
  wire Arbiter_Y_6__ap_ready;
  wire Arbiter_Y_6__ap_done;
  wire Arbiter_Y_6__ap_idle;
  reg [1:0] Arbiter_Y_6__state;
  wire [31:0] Arbiter_Y_7___M__q0;
  wire [31:0] Arbiter_Y_7___P_N__q0;
  wire Arbiter_Y_7__ap_start_global__q0;
  wire Arbiter_Y_7__is_done__q0;
  wire Arbiter_Y_7__ap_done_global__q0;
  wire Arbiter_Y_7__ap_start;
  wire Arbiter_Y_7__ap_ready;
  wire Arbiter_Y_7__ap_done;
  wire Arbiter_Y_7__ap_idle;
  reg [1:0] Arbiter_Y_7__state;
  wire FloatvAddFloatv_0__ap_start_global__q0;
  reg FloatvAddFloatv_0__ap_start;
  wire [31:0] FloatvMultConst_0___M__q0;
  wire [31:0] FloatvMultConst_0___P_N__q0;
  wire [31:0] FloatvMultConst_0___alpha_u__q0;
  wire FloatvMultConst_0__ap_start_global__q0;
  wire FloatvMultConst_0__is_done__q0;
  wire FloatvMultConst_0__ap_done_global__q0;
  wire FloatvMultConst_0__ap_start;
  wire FloatvMultConst_0__ap_ready;
  wire FloatvMultConst_0__ap_done;
  wire FloatvMultConst_0__ap_idle;
  reg [1:0] FloatvMultConst_0__state;
  wire [31:0] FloatvMultConst_1___M__q0;
  wire [31:0] FloatvMultConst_1___P_N__q0;
  wire [31:0] FloatvMultConst_1___beta_u__q0;
  wire FloatvMultConst_1__ap_start_global__q0;
  wire FloatvMultConst_1__is_done__q0;
  wire FloatvMultConst_1__ap_done_global__q0;
  wire FloatvMultConst_1__ap_start;
  wire FloatvMultConst_1__ap_ready;
  wire FloatvMultConst_1__ap_done;
  wire FloatvMultConst_1__ap_idle;
  reg [1:0] FloatvMultConst_1__state;
  wire Merger_Y_0__ap_start_global__q0;
  reg Merger_Y_0__ap_start;
  wire PEG_Xvec_0__ap_start_global__q0;
  wire PEG_Xvec_0__is_done__q0;
  wire PEG_Xvec_0__ap_done_global__q0;
  wire PEG_Xvec_0__ap_start;
  wire PEG_Xvec_0__ap_ready;
  wire PEG_Xvec_0__ap_done;
  wire PEG_Xvec_0__ap_idle;
  reg [1:0] PEG_Xvec_0__state;
  wire PEG_Xvec_1__ap_start_global__q0;
  wire PEG_Xvec_1__is_done__q0;
  wire PEG_Xvec_1__ap_done_global__q0;
  wire PEG_Xvec_1__ap_start;
  wire PEG_Xvec_1__ap_ready;
  wire PEG_Xvec_1__ap_done;
  wire PEG_Xvec_1__ap_idle;
  reg [1:0] PEG_Xvec_1__state;
  wire PEG_Xvec_2__ap_start_global__q0;
  wire PEG_Xvec_2__is_done__q0;
  wire PEG_Xvec_2__ap_done_global__q0;
  wire PEG_Xvec_2__ap_start;
  wire PEG_Xvec_2__ap_ready;
  wire PEG_Xvec_2__ap_done;
  wire PEG_Xvec_2__ap_idle;
  reg [1:0] PEG_Xvec_2__state;
  wire PEG_Xvec_3__ap_start_global__q0;
  wire PEG_Xvec_3__is_done__q0;
  wire PEG_Xvec_3__ap_done_global__q0;
  wire PEG_Xvec_3__ap_start;
  wire PEG_Xvec_3__ap_ready;
  wire PEG_Xvec_3__ap_done;
  wire PEG_Xvec_3__ap_idle;
  reg [1:0] PEG_Xvec_3__state;
  wire PEG_Xvec_4__ap_start_global__q0;
  wire PEG_Xvec_4__is_done__q0;
  wire PEG_Xvec_4__ap_done_global__q0;
  wire PEG_Xvec_4__ap_start;
  wire PEG_Xvec_4__ap_ready;
  wire PEG_Xvec_4__ap_done;
  wire PEG_Xvec_4__ap_idle;
  reg [1:0] PEG_Xvec_4__state;
  wire PEG_Xvec_5__ap_start_global__q0;
  wire PEG_Xvec_5__is_done__q0;
  wire PEG_Xvec_5__ap_done_global__q0;
  wire PEG_Xvec_5__ap_start;
  wire PEG_Xvec_5__ap_ready;
  wire PEG_Xvec_5__ap_done;
  wire PEG_Xvec_5__ap_idle;
  reg [1:0] PEG_Xvec_5__state;
  wire PEG_Xvec_6__ap_start_global__q0;
  wire PEG_Xvec_6__is_done__q0;
  wire PEG_Xvec_6__ap_done_global__q0;
  wire PEG_Xvec_6__ap_start;
  wire PEG_Xvec_6__ap_ready;
  wire PEG_Xvec_6__ap_done;
  wire PEG_Xvec_6__ap_idle;
  reg [1:0] PEG_Xvec_6__state;
  wire PEG_Xvec_7__ap_start_global__q0;
  wire PEG_Xvec_7__is_done__q0;
  wire PEG_Xvec_7__ap_done_global__q0;
  wire PEG_Xvec_7__ap_start;
  wire PEG_Xvec_7__ap_ready;
  wire PEG_Xvec_7__ap_done;
  wire PEG_Xvec_7__ap_idle;
  reg [1:0] PEG_Xvec_7__state;
  wire PEG_Xvec_8__ap_start_global__q0;
  wire PEG_Xvec_8__is_done__q0;
  wire PEG_Xvec_8__ap_done_global__q0;
  wire PEG_Xvec_8__ap_start;
  wire PEG_Xvec_8__ap_ready;
  wire PEG_Xvec_8__ap_done;
  wire PEG_Xvec_8__ap_idle;
  reg [1:0] PEG_Xvec_8__state;
  wire PEG_Xvec_9__ap_start_global__q0;
  wire PEG_Xvec_9__is_done__q0;
  wire PEG_Xvec_9__ap_done_global__q0;
  wire PEG_Xvec_9__ap_start;
  wire PEG_Xvec_9__ap_ready;
  wire PEG_Xvec_9__ap_done;
  wire PEG_Xvec_9__ap_idle;
  reg [1:0] PEG_Xvec_9__state;
  wire PEG_Xvec_10__ap_start_global__q0;
  wire PEG_Xvec_10__is_done__q0;
  wire PEG_Xvec_10__ap_done_global__q0;
  wire PEG_Xvec_10__ap_start;
  wire PEG_Xvec_10__ap_ready;
  wire PEG_Xvec_10__ap_done;
  wire PEG_Xvec_10__ap_idle;
  reg [1:0] PEG_Xvec_10__state;
  wire PEG_Xvec_11__ap_start_global__q0;
  wire PEG_Xvec_11__is_done__q0;
  wire PEG_Xvec_11__ap_done_global__q0;
  wire PEG_Xvec_11__ap_start;
  wire PEG_Xvec_11__ap_ready;
  wire PEG_Xvec_11__ap_done;
  wire PEG_Xvec_11__ap_idle;
  reg [1:0] PEG_Xvec_11__state;
  wire PEG_Xvec_12__ap_start_global__q0;
  wire PEG_Xvec_12__is_done__q0;
  wire PEG_Xvec_12__ap_done_global__q0;
  wire PEG_Xvec_12__ap_start;
  wire PEG_Xvec_12__ap_ready;
  wire PEG_Xvec_12__ap_done;
  wire PEG_Xvec_12__ap_idle;
  reg [1:0] PEG_Xvec_12__state;
  wire PEG_Xvec_13__ap_start_global__q0;
  wire PEG_Xvec_13__is_done__q0;
  wire PEG_Xvec_13__ap_done_global__q0;
  wire PEG_Xvec_13__ap_start;
  wire PEG_Xvec_13__ap_ready;
  wire PEG_Xvec_13__ap_done;
  wire PEG_Xvec_13__ap_idle;
  reg [1:0] PEG_Xvec_13__state;
  wire PEG_Xvec_14__ap_start_global__q0;
  wire PEG_Xvec_14__is_done__q0;
  wire PEG_Xvec_14__ap_done_global__q0;
  wire PEG_Xvec_14__ap_start;
  wire PEG_Xvec_14__ap_ready;
  wire PEG_Xvec_14__ap_done;
  wire PEG_Xvec_14__ap_idle;
  reg [1:0] PEG_Xvec_14__state;
  wire PEG_Xvec_15__ap_start_global__q0;
  wire PEG_Xvec_15__is_done__q0;
  wire PEG_Xvec_15__ap_done_global__q0;
  wire PEG_Xvec_15__ap_start;
  wire PEG_Xvec_15__ap_ready;
  wire PEG_Xvec_15__ap_done;
  wire PEG_Xvec_15__ap_idle;
  reg [1:0] PEG_Xvec_15__state;
  wire PEG_Xvec_16__ap_start_global__q0;
  wire PEG_Xvec_16__is_done__q0;
  wire PEG_Xvec_16__ap_done_global__q0;
  wire PEG_Xvec_16__ap_start;
  wire PEG_Xvec_16__ap_ready;
  wire PEG_Xvec_16__ap_done;
  wire PEG_Xvec_16__ap_idle;
  reg [1:0] PEG_Xvec_16__state;
  wire PEG_Xvec_17__ap_start_global__q0;
  wire PEG_Xvec_17__is_done__q0;
  wire PEG_Xvec_17__ap_done_global__q0;
  wire PEG_Xvec_17__ap_start;
  wire PEG_Xvec_17__ap_ready;
  wire PEG_Xvec_17__ap_done;
  wire PEG_Xvec_17__ap_idle;
  reg [1:0] PEG_Xvec_17__state;
  wire PEG_Xvec_18__ap_start_global__q0;
  wire PEG_Xvec_18__is_done__q0;
  wire PEG_Xvec_18__ap_done_global__q0;
  wire PEG_Xvec_18__ap_start;
  wire PEG_Xvec_18__ap_ready;
  wire PEG_Xvec_18__ap_done;
  wire PEG_Xvec_18__ap_idle;
  reg [1:0] PEG_Xvec_18__state;
  wire PEG_Xvec_19__ap_start_global__q0;
  wire PEG_Xvec_19__is_done__q0;
  wire PEG_Xvec_19__ap_done_global__q0;
  wire PEG_Xvec_19__ap_start;
  wire PEG_Xvec_19__ap_ready;
  wire PEG_Xvec_19__ap_done;
  wire PEG_Xvec_19__ap_idle;
  reg [1:0] PEG_Xvec_19__state;
  wire PEG_Xvec_20__ap_start_global__q0;
  wire PEG_Xvec_20__is_done__q0;
  wire PEG_Xvec_20__ap_done_global__q0;
  wire PEG_Xvec_20__ap_start;
  wire PEG_Xvec_20__ap_ready;
  wire PEG_Xvec_20__ap_done;
  wire PEG_Xvec_20__ap_idle;
  reg [1:0] PEG_Xvec_20__state;
  wire PEG_Xvec_21__ap_start_global__q0;
  wire PEG_Xvec_21__is_done__q0;
  wire PEG_Xvec_21__ap_done_global__q0;
  wire PEG_Xvec_21__ap_start;
  wire PEG_Xvec_21__ap_ready;
  wire PEG_Xvec_21__ap_done;
  wire PEG_Xvec_21__ap_idle;
  reg [1:0] PEG_Xvec_21__state;
  wire PEG_Xvec_22__ap_start_global__q0;
  wire PEG_Xvec_22__is_done__q0;
  wire PEG_Xvec_22__ap_done_global__q0;
  wire PEG_Xvec_22__ap_start;
  wire PEG_Xvec_22__ap_ready;
  wire PEG_Xvec_22__ap_done;
  wire PEG_Xvec_22__ap_idle;
  reg [1:0] PEG_Xvec_22__state;
  wire PEG_Xvec_23__ap_start_global__q0;
  wire PEG_Xvec_23__is_done__q0;
  wire PEG_Xvec_23__ap_done_global__q0;
  wire PEG_Xvec_23__ap_start;
  wire PEG_Xvec_23__ap_ready;
  wire PEG_Xvec_23__ap_done;
  wire PEG_Xvec_23__ap_idle;
  reg [1:0] PEG_Xvec_23__state;
  wire PEG_Xvec_24__ap_start_global__q0;
  wire PEG_Xvec_24__is_done__q0;
  wire PEG_Xvec_24__ap_done_global__q0;
  wire PEG_Xvec_24__ap_start;
  wire PEG_Xvec_24__ap_ready;
  wire PEG_Xvec_24__ap_done;
  wire PEG_Xvec_24__ap_idle;
  reg [1:0] PEG_Xvec_24__state;
  wire PEG_Xvec_25__ap_start_global__q0;
  wire PEG_Xvec_25__is_done__q0;
  wire PEG_Xvec_25__ap_done_global__q0;
  wire PEG_Xvec_25__ap_start;
  wire PEG_Xvec_25__ap_ready;
  wire PEG_Xvec_25__ap_done;
  wire PEG_Xvec_25__ap_idle;
  reg [1:0] PEG_Xvec_25__state;
  wire PEG_Xvec_26__ap_start_global__q0;
  wire PEG_Xvec_26__is_done__q0;
  wire PEG_Xvec_26__ap_done_global__q0;
  wire PEG_Xvec_26__ap_start;
  wire PEG_Xvec_26__ap_ready;
  wire PEG_Xvec_26__ap_done;
  wire PEG_Xvec_26__ap_idle;
  reg [1:0] PEG_Xvec_26__state;
  wire PEG_Xvec_27__ap_start_global__q0;
  wire PEG_Xvec_27__is_done__q0;
  wire PEG_Xvec_27__ap_done_global__q0;
  wire PEG_Xvec_27__ap_start;
  wire PEG_Xvec_27__ap_ready;
  wire PEG_Xvec_27__ap_done;
  wire PEG_Xvec_27__ap_idle;
  reg [1:0] PEG_Xvec_27__state;
  wire PEG_Xvec_28__ap_start_global__q0;
  wire PEG_Xvec_28__is_done__q0;
  wire PEG_Xvec_28__ap_done_global__q0;
  wire PEG_Xvec_28__ap_start;
  wire PEG_Xvec_28__ap_ready;
  wire PEG_Xvec_28__ap_done;
  wire PEG_Xvec_28__ap_idle;
  reg [1:0] PEG_Xvec_28__state;
  wire PEG_Xvec_29__ap_start_global__q0;
  wire PEG_Xvec_29__is_done__q0;
  wire PEG_Xvec_29__ap_done_global__q0;
  wire PEG_Xvec_29__ap_start;
  wire PEG_Xvec_29__ap_ready;
  wire PEG_Xvec_29__ap_done;
  wire PEG_Xvec_29__ap_idle;
  reg [1:0] PEG_Xvec_29__state;
  wire PEG_Xvec_30__ap_start_global__q0;
  wire PEG_Xvec_30__is_done__q0;
  wire PEG_Xvec_30__ap_done_global__q0;
  wire PEG_Xvec_30__ap_start;
  wire PEG_Xvec_30__ap_ready;
  wire PEG_Xvec_30__ap_done;
  wire PEG_Xvec_30__ap_idle;
  reg [1:0] PEG_Xvec_30__state;
  wire PEG_Xvec_31__ap_start_global__q0;
  wire PEG_Xvec_31__is_done__q0;
  wire PEG_Xvec_31__ap_done_global__q0;
  wire PEG_Xvec_31__ap_start;
  wire PEG_Xvec_31__ap_ready;
  wire PEG_Xvec_31__ap_done;
  wire PEG_Xvec_31__ap_idle;
  reg [1:0] PEG_Xvec_31__state;
  wire PEG_Xvec_32__ap_start_global__q0;
  wire PEG_Xvec_32__is_done__q0;
  wire PEG_Xvec_32__ap_done_global__q0;
  wire PEG_Xvec_32__ap_start;
  wire PEG_Xvec_32__ap_ready;
  wire PEG_Xvec_32__ap_done;
  wire PEG_Xvec_32__ap_idle;
  reg [1:0] PEG_Xvec_32__state;
  wire PEG_Xvec_33__ap_start_global__q0;
  wire PEG_Xvec_33__is_done__q0;
  wire PEG_Xvec_33__ap_done_global__q0;
  wire PEG_Xvec_33__ap_start;
  wire PEG_Xvec_33__ap_ready;
  wire PEG_Xvec_33__ap_done;
  wire PEG_Xvec_33__ap_idle;
  reg [1:0] PEG_Xvec_33__state;
  wire PEG_Xvec_34__ap_start_global__q0;
  wire PEG_Xvec_34__is_done__q0;
  wire PEG_Xvec_34__ap_done_global__q0;
  wire PEG_Xvec_34__ap_start;
  wire PEG_Xvec_34__ap_ready;
  wire PEG_Xvec_34__ap_done;
  wire PEG_Xvec_34__ap_idle;
  reg [1:0] PEG_Xvec_34__state;
  wire PEG_Xvec_35__ap_start_global__q0;
  wire PEG_Xvec_35__is_done__q0;
  wire PEG_Xvec_35__ap_done_global__q0;
  wire PEG_Xvec_35__ap_start;
  wire PEG_Xvec_35__ap_ready;
  wire PEG_Xvec_35__ap_done;
  wire PEG_Xvec_35__ap_idle;
  reg [1:0] PEG_Xvec_35__state;
  wire PEG_Xvec_36__ap_start_global__q0;
  wire PEG_Xvec_36__is_done__q0;
  wire PEG_Xvec_36__ap_done_global__q0;
  wire PEG_Xvec_36__ap_start;
  wire PEG_Xvec_36__ap_ready;
  wire PEG_Xvec_36__ap_done;
  wire PEG_Xvec_36__ap_idle;
  reg [1:0] PEG_Xvec_36__state;
  wire PEG_Xvec_37__ap_start_global__q0;
  wire PEG_Xvec_37__is_done__q0;
  wire PEG_Xvec_37__ap_done_global__q0;
  wire PEG_Xvec_37__ap_start;
  wire PEG_Xvec_37__ap_ready;
  wire PEG_Xvec_37__ap_done;
  wire PEG_Xvec_37__ap_idle;
  reg [1:0] PEG_Xvec_37__state;
  wire PEG_Xvec_38__ap_start_global__q0;
  wire PEG_Xvec_38__is_done__q0;
  wire PEG_Xvec_38__ap_done_global__q0;
  wire PEG_Xvec_38__ap_start;
  wire PEG_Xvec_38__ap_ready;
  wire PEG_Xvec_38__ap_done;
  wire PEG_Xvec_38__ap_idle;
  reg [1:0] PEG_Xvec_38__state;
  wire PEG_Xvec_39__ap_start_global__q0;
  wire PEG_Xvec_39__is_done__q0;
  wire PEG_Xvec_39__ap_done_global__q0;
  wire PEG_Xvec_39__ap_start;
  wire PEG_Xvec_39__ap_ready;
  wire PEG_Xvec_39__ap_done;
  wire PEG_Xvec_39__ap_idle;
  reg [1:0] PEG_Xvec_39__state;
  wire PEG_Xvec_40__ap_start_global__q0;
  wire PEG_Xvec_40__is_done__q0;
  wire PEG_Xvec_40__ap_done_global__q0;
  wire PEG_Xvec_40__ap_start;
  wire PEG_Xvec_40__ap_ready;
  wire PEG_Xvec_40__ap_done;
  wire PEG_Xvec_40__ap_idle;
  reg [1:0] PEG_Xvec_40__state;
  wire PEG_Xvec_41__ap_start_global__q0;
  wire PEG_Xvec_41__is_done__q0;
  wire PEG_Xvec_41__ap_done_global__q0;
  wire PEG_Xvec_41__ap_start;
  wire PEG_Xvec_41__ap_ready;
  wire PEG_Xvec_41__ap_done;
  wire PEG_Xvec_41__ap_idle;
  reg [1:0] PEG_Xvec_41__state;
  wire PEG_Xvec_42__ap_start_global__q0;
  wire PEG_Xvec_42__is_done__q0;
  wire PEG_Xvec_42__ap_done_global__q0;
  wire PEG_Xvec_42__ap_start;
  wire PEG_Xvec_42__ap_ready;
  wire PEG_Xvec_42__ap_done;
  wire PEG_Xvec_42__ap_idle;
  reg [1:0] PEG_Xvec_42__state;
  wire PEG_Xvec_43__ap_start_global__q0;
  wire PEG_Xvec_43__is_done__q0;
  wire PEG_Xvec_43__ap_done_global__q0;
  wire PEG_Xvec_43__ap_start;
  wire PEG_Xvec_43__ap_ready;
  wire PEG_Xvec_43__ap_done;
  wire PEG_Xvec_43__ap_idle;
  reg [1:0] PEG_Xvec_43__state;
  wire PEG_Xvec_44__ap_start_global__q0;
  wire PEG_Xvec_44__is_done__q0;
  wire PEG_Xvec_44__ap_done_global__q0;
  wire PEG_Xvec_44__ap_start;
  wire PEG_Xvec_44__ap_ready;
  wire PEG_Xvec_44__ap_done;
  wire PEG_Xvec_44__ap_idle;
  reg [1:0] PEG_Xvec_44__state;
  wire PEG_Xvec_45__ap_start_global__q0;
  wire PEG_Xvec_45__is_done__q0;
  wire PEG_Xvec_45__ap_done_global__q0;
  wire PEG_Xvec_45__ap_start;
  wire PEG_Xvec_45__ap_ready;
  wire PEG_Xvec_45__ap_done;
  wire PEG_Xvec_45__ap_idle;
  reg [1:0] PEG_Xvec_45__state;
  wire PEG_Xvec_46__ap_start_global__q0;
  wire PEG_Xvec_46__is_done__q0;
  wire PEG_Xvec_46__ap_done_global__q0;
  wire PEG_Xvec_46__ap_start;
  wire PEG_Xvec_46__ap_ready;
  wire PEG_Xvec_46__ap_done;
  wire PEG_Xvec_46__ap_idle;
  reg [1:0] PEG_Xvec_46__state;
  wire PEG_Xvec_47__ap_start_global__q0;
  wire PEG_Xvec_47__is_done__q0;
  wire PEG_Xvec_47__ap_done_global__q0;
  wire PEG_Xvec_47__ap_start;
  wire PEG_Xvec_47__ap_ready;
  wire PEG_Xvec_47__ap_done;
  wire PEG_Xvec_47__ap_idle;
  reg [1:0] PEG_Xvec_47__state;
  wire PEG_Yvec_0__ap_start_global__q0;
  wire PEG_Yvec_0__is_done__q0;
  wire PEG_Yvec_0__ap_done_global__q0;
  wire PEG_Yvec_0__ap_start;
  wire PEG_Yvec_0__ap_ready;
  wire PEG_Yvec_0__ap_done;
  wire PEG_Yvec_0__ap_idle;
  reg [1:0] PEG_Yvec_0__state;
  wire PEG_Yvec_1__ap_start_global__q0;
  wire PEG_Yvec_1__is_done__q0;
  wire PEG_Yvec_1__ap_done_global__q0;
  wire PEG_Yvec_1__ap_start;
  wire PEG_Yvec_1__ap_ready;
  wire PEG_Yvec_1__ap_done;
  wire PEG_Yvec_1__ap_idle;
  reg [1:0] PEG_Yvec_1__state;
  wire PEG_Yvec_2__ap_start_global__q0;
  wire PEG_Yvec_2__is_done__q0;
  wire PEG_Yvec_2__ap_done_global__q0;
  wire PEG_Yvec_2__ap_start;
  wire PEG_Yvec_2__ap_ready;
  wire PEG_Yvec_2__ap_done;
  wire PEG_Yvec_2__ap_idle;
  reg [1:0] PEG_Yvec_2__state;
  wire PEG_Yvec_3__ap_start_global__q0;
  wire PEG_Yvec_3__is_done__q0;
  wire PEG_Yvec_3__ap_done_global__q0;
  wire PEG_Yvec_3__ap_start;
  wire PEG_Yvec_3__ap_ready;
  wire PEG_Yvec_3__ap_done;
  wire PEG_Yvec_3__ap_idle;
  reg [1:0] PEG_Yvec_3__state;
  wire PEG_Yvec_4__ap_start_global__q0;
  wire PEG_Yvec_4__is_done__q0;
  wire PEG_Yvec_4__ap_done_global__q0;
  wire PEG_Yvec_4__ap_start;
  wire PEG_Yvec_4__ap_ready;
  wire PEG_Yvec_4__ap_done;
  wire PEG_Yvec_4__ap_idle;
  reg [1:0] PEG_Yvec_4__state;
  wire PEG_Yvec_5__ap_start_global__q0;
  wire PEG_Yvec_5__is_done__q0;
  wire PEG_Yvec_5__ap_done_global__q0;
  wire PEG_Yvec_5__ap_start;
  wire PEG_Yvec_5__ap_ready;
  wire PEG_Yvec_5__ap_done;
  wire PEG_Yvec_5__ap_idle;
  reg [1:0] PEG_Yvec_5__state;
  wire PEG_Yvec_6__ap_start_global__q0;
  wire PEG_Yvec_6__is_done__q0;
  wire PEG_Yvec_6__ap_done_global__q0;
  wire PEG_Yvec_6__ap_start;
  wire PEG_Yvec_6__ap_ready;
  wire PEG_Yvec_6__ap_done;
  wire PEG_Yvec_6__ap_idle;
  reg [1:0] PEG_Yvec_6__state;
  wire PEG_Yvec_7__ap_start_global__q0;
  wire PEG_Yvec_7__is_done__q0;
  wire PEG_Yvec_7__ap_done_global__q0;
  wire PEG_Yvec_7__ap_start;
  wire PEG_Yvec_7__ap_ready;
  wire PEG_Yvec_7__ap_done;
  wire PEG_Yvec_7__ap_idle;
  reg [1:0] PEG_Yvec_7__state;
  wire PEG_Yvec_8__ap_start_global__q0;
  wire PEG_Yvec_8__is_done__q0;
  wire PEG_Yvec_8__ap_done_global__q0;
  wire PEG_Yvec_8__ap_start;
  wire PEG_Yvec_8__ap_ready;
  wire PEG_Yvec_8__ap_done;
  wire PEG_Yvec_8__ap_idle;
  reg [1:0] PEG_Yvec_8__state;
  wire PEG_Yvec_9__ap_start_global__q0;
  wire PEG_Yvec_9__is_done__q0;
  wire PEG_Yvec_9__ap_done_global__q0;
  wire PEG_Yvec_9__ap_start;
  wire PEG_Yvec_9__ap_ready;
  wire PEG_Yvec_9__ap_done;
  wire PEG_Yvec_9__ap_idle;
  reg [1:0] PEG_Yvec_9__state;
  wire PEG_Yvec_10__ap_start_global__q0;
  wire PEG_Yvec_10__is_done__q0;
  wire PEG_Yvec_10__ap_done_global__q0;
  wire PEG_Yvec_10__ap_start;
  wire PEG_Yvec_10__ap_ready;
  wire PEG_Yvec_10__ap_done;
  wire PEG_Yvec_10__ap_idle;
  reg [1:0] PEG_Yvec_10__state;
  wire PEG_Yvec_11__ap_start_global__q0;
  wire PEG_Yvec_11__is_done__q0;
  wire PEG_Yvec_11__ap_done_global__q0;
  wire PEG_Yvec_11__ap_start;
  wire PEG_Yvec_11__ap_ready;
  wire PEG_Yvec_11__ap_done;
  wire PEG_Yvec_11__ap_idle;
  reg [1:0] PEG_Yvec_11__state;
  wire PEG_Yvec_12__ap_start_global__q0;
  wire PEG_Yvec_12__is_done__q0;
  wire PEG_Yvec_12__ap_done_global__q0;
  wire PEG_Yvec_12__ap_start;
  wire PEG_Yvec_12__ap_ready;
  wire PEG_Yvec_12__ap_done;
  wire PEG_Yvec_12__ap_idle;
  reg [1:0] PEG_Yvec_12__state;
  wire PEG_Yvec_13__ap_start_global__q0;
  wire PEG_Yvec_13__is_done__q0;
  wire PEG_Yvec_13__ap_done_global__q0;
  wire PEG_Yvec_13__ap_start;
  wire PEG_Yvec_13__ap_ready;
  wire PEG_Yvec_13__ap_done;
  wire PEG_Yvec_13__ap_idle;
  reg [1:0] PEG_Yvec_13__state;
  wire PEG_Yvec_14__ap_start_global__q0;
  wire PEG_Yvec_14__is_done__q0;
  wire PEG_Yvec_14__ap_done_global__q0;
  wire PEG_Yvec_14__ap_start;
  wire PEG_Yvec_14__ap_ready;
  wire PEG_Yvec_14__ap_done;
  wire PEG_Yvec_14__ap_idle;
  reg [1:0] PEG_Yvec_14__state;
  wire PEG_Yvec_15__ap_start_global__q0;
  wire PEG_Yvec_15__is_done__q0;
  wire PEG_Yvec_15__ap_done_global__q0;
  wire PEG_Yvec_15__ap_start;
  wire PEG_Yvec_15__ap_ready;
  wire PEG_Yvec_15__ap_done;
  wire PEG_Yvec_15__ap_idle;
  reg [1:0] PEG_Yvec_15__state;
  wire PEG_Yvec_16__ap_start_global__q0;
  wire PEG_Yvec_16__is_done__q0;
  wire PEG_Yvec_16__ap_done_global__q0;
  wire PEG_Yvec_16__ap_start;
  wire PEG_Yvec_16__ap_ready;
  wire PEG_Yvec_16__ap_done;
  wire PEG_Yvec_16__ap_idle;
  reg [1:0] PEG_Yvec_16__state;
  wire PEG_Yvec_17__ap_start_global__q0;
  wire PEG_Yvec_17__is_done__q0;
  wire PEG_Yvec_17__ap_done_global__q0;
  wire PEG_Yvec_17__ap_start;
  wire PEG_Yvec_17__ap_ready;
  wire PEG_Yvec_17__ap_done;
  wire PEG_Yvec_17__ap_idle;
  reg [1:0] PEG_Yvec_17__state;
  wire PEG_Yvec_18__ap_start_global__q0;
  wire PEG_Yvec_18__is_done__q0;
  wire PEG_Yvec_18__ap_done_global__q0;
  wire PEG_Yvec_18__ap_start;
  wire PEG_Yvec_18__ap_ready;
  wire PEG_Yvec_18__ap_done;
  wire PEG_Yvec_18__ap_idle;
  reg [1:0] PEG_Yvec_18__state;
  wire PEG_Yvec_19__ap_start_global__q0;
  wire PEG_Yvec_19__is_done__q0;
  wire PEG_Yvec_19__ap_done_global__q0;
  wire PEG_Yvec_19__ap_start;
  wire PEG_Yvec_19__ap_ready;
  wire PEG_Yvec_19__ap_done;
  wire PEG_Yvec_19__ap_idle;
  reg [1:0] PEG_Yvec_19__state;
  wire PEG_Yvec_20__ap_start_global__q0;
  wire PEG_Yvec_20__is_done__q0;
  wire PEG_Yvec_20__ap_done_global__q0;
  wire PEG_Yvec_20__ap_start;
  wire PEG_Yvec_20__ap_ready;
  wire PEG_Yvec_20__ap_done;
  wire PEG_Yvec_20__ap_idle;
  reg [1:0] PEG_Yvec_20__state;
  wire PEG_Yvec_21__ap_start_global__q0;
  wire PEG_Yvec_21__is_done__q0;
  wire PEG_Yvec_21__ap_done_global__q0;
  wire PEG_Yvec_21__ap_start;
  wire PEG_Yvec_21__ap_ready;
  wire PEG_Yvec_21__ap_done;
  wire PEG_Yvec_21__ap_idle;
  reg [1:0] PEG_Yvec_21__state;
  wire PEG_Yvec_22__ap_start_global__q0;
  wire PEG_Yvec_22__is_done__q0;
  wire PEG_Yvec_22__ap_done_global__q0;
  wire PEG_Yvec_22__ap_start;
  wire PEG_Yvec_22__ap_ready;
  wire PEG_Yvec_22__ap_done;
  wire PEG_Yvec_22__ap_idle;
  reg [1:0] PEG_Yvec_22__state;
  wire PEG_Yvec_23__ap_start_global__q0;
  wire PEG_Yvec_23__is_done__q0;
  wire PEG_Yvec_23__ap_done_global__q0;
  wire PEG_Yvec_23__ap_start;
  wire PEG_Yvec_23__ap_ready;
  wire PEG_Yvec_23__ap_done;
  wire PEG_Yvec_23__ap_idle;
  reg [1:0] PEG_Yvec_23__state;
  wire PEG_Yvec_24__ap_start_global__q0;
  wire PEG_Yvec_24__is_done__q0;
  wire PEG_Yvec_24__ap_done_global__q0;
  wire PEG_Yvec_24__ap_start;
  wire PEG_Yvec_24__ap_ready;
  wire PEG_Yvec_24__ap_done;
  wire PEG_Yvec_24__ap_idle;
  reg [1:0] PEG_Yvec_24__state;
  wire PEG_Yvec_25__ap_start_global__q0;
  wire PEG_Yvec_25__is_done__q0;
  wire PEG_Yvec_25__ap_done_global__q0;
  wire PEG_Yvec_25__ap_start;
  wire PEG_Yvec_25__ap_ready;
  wire PEG_Yvec_25__ap_done;
  wire PEG_Yvec_25__ap_idle;
  reg [1:0] PEG_Yvec_25__state;
  wire PEG_Yvec_26__ap_start_global__q0;
  wire PEG_Yvec_26__is_done__q0;
  wire PEG_Yvec_26__ap_done_global__q0;
  wire PEG_Yvec_26__ap_start;
  wire PEG_Yvec_26__ap_ready;
  wire PEG_Yvec_26__ap_done;
  wire PEG_Yvec_26__ap_idle;
  reg [1:0] PEG_Yvec_26__state;
  wire PEG_Yvec_27__ap_start_global__q0;
  wire PEG_Yvec_27__is_done__q0;
  wire PEG_Yvec_27__ap_done_global__q0;
  wire PEG_Yvec_27__ap_start;
  wire PEG_Yvec_27__ap_ready;
  wire PEG_Yvec_27__ap_done;
  wire PEG_Yvec_27__ap_idle;
  reg [1:0] PEG_Yvec_27__state;
  wire PEG_Yvec_28__ap_start_global__q0;
  wire PEG_Yvec_28__is_done__q0;
  wire PEG_Yvec_28__ap_done_global__q0;
  wire PEG_Yvec_28__ap_start;
  wire PEG_Yvec_28__ap_ready;
  wire PEG_Yvec_28__ap_done;
  wire PEG_Yvec_28__ap_idle;
  reg [1:0] PEG_Yvec_28__state;
  wire PEG_Yvec_29__ap_start_global__q0;
  wire PEG_Yvec_29__is_done__q0;
  wire PEG_Yvec_29__ap_done_global__q0;
  wire PEG_Yvec_29__ap_start;
  wire PEG_Yvec_29__ap_ready;
  wire PEG_Yvec_29__ap_done;
  wire PEG_Yvec_29__ap_idle;
  reg [1:0] PEG_Yvec_29__state;
  wire PEG_Yvec_30__ap_start_global__q0;
  wire PEG_Yvec_30__is_done__q0;
  wire PEG_Yvec_30__ap_done_global__q0;
  wire PEG_Yvec_30__ap_start;
  wire PEG_Yvec_30__ap_ready;
  wire PEG_Yvec_30__ap_done;
  wire PEG_Yvec_30__ap_idle;
  reg [1:0] PEG_Yvec_30__state;
  wire PEG_Yvec_31__ap_start_global__q0;
  wire PEG_Yvec_31__is_done__q0;
  wire PEG_Yvec_31__ap_done_global__q0;
  wire PEG_Yvec_31__ap_start;
  wire PEG_Yvec_31__ap_ready;
  wire PEG_Yvec_31__ap_done;
  wire PEG_Yvec_31__ap_idle;
  reg [1:0] PEG_Yvec_31__state;
  wire PEG_Yvec_32__ap_start_global__q0;
  wire PEG_Yvec_32__is_done__q0;
  wire PEG_Yvec_32__ap_done_global__q0;
  wire PEG_Yvec_32__ap_start;
  wire PEG_Yvec_32__ap_ready;
  wire PEG_Yvec_32__ap_done;
  wire PEG_Yvec_32__ap_idle;
  reg [1:0] PEG_Yvec_32__state;
  wire PEG_Yvec_33__ap_start_global__q0;
  wire PEG_Yvec_33__is_done__q0;
  wire PEG_Yvec_33__ap_done_global__q0;
  wire PEG_Yvec_33__ap_start;
  wire PEG_Yvec_33__ap_ready;
  wire PEG_Yvec_33__ap_done;
  wire PEG_Yvec_33__ap_idle;
  reg [1:0] PEG_Yvec_33__state;
  wire PEG_Yvec_34__ap_start_global__q0;
  wire PEG_Yvec_34__is_done__q0;
  wire PEG_Yvec_34__ap_done_global__q0;
  wire PEG_Yvec_34__ap_start;
  wire PEG_Yvec_34__ap_ready;
  wire PEG_Yvec_34__ap_done;
  wire PEG_Yvec_34__ap_idle;
  reg [1:0] PEG_Yvec_34__state;
  wire PEG_Yvec_35__ap_start_global__q0;
  wire PEG_Yvec_35__is_done__q0;
  wire PEG_Yvec_35__ap_done_global__q0;
  wire PEG_Yvec_35__ap_start;
  wire PEG_Yvec_35__ap_ready;
  wire PEG_Yvec_35__ap_done;
  wire PEG_Yvec_35__ap_idle;
  reg [1:0] PEG_Yvec_35__state;
  wire PEG_Yvec_36__ap_start_global__q0;
  wire PEG_Yvec_36__is_done__q0;
  wire PEG_Yvec_36__ap_done_global__q0;
  wire PEG_Yvec_36__ap_start;
  wire PEG_Yvec_36__ap_ready;
  wire PEG_Yvec_36__ap_done;
  wire PEG_Yvec_36__ap_idle;
  reg [1:0] PEG_Yvec_36__state;
  wire PEG_Yvec_37__ap_start_global__q0;
  wire PEG_Yvec_37__is_done__q0;
  wire PEG_Yvec_37__ap_done_global__q0;
  wire PEG_Yvec_37__ap_start;
  wire PEG_Yvec_37__ap_ready;
  wire PEG_Yvec_37__ap_done;
  wire PEG_Yvec_37__ap_idle;
  reg [1:0] PEG_Yvec_37__state;
  wire PEG_Yvec_38__ap_start_global__q0;
  wire PEG_Yvec_38__is_done__q0;
  wire PEG_Yvec_38__ap_done_global__q0;
  wire PEG_Yvec_38__ap_start;
  wire PEG_Yvec_38__ap_ready;
  wire PEG_Yvec_38__ap_done;
  wire PEG_Yvec_38__ap_idle;
  reg [1:0] PEG_Yvec_38__state;
  wire PEG_Yvec_39__ap_start_global__q0;
  wire PEG_Yvec_39__is_done__q0;
  wire PEG_Yvec_39__ap_done_global__q0;
  wire PEG_Yvec_39__ap_start;
  wire PEG_Yvec_39__ap_ready;
  wire PEG_Yvec_39__ap_done;
  wire PEG_Yvec_39__ap_idle;
  reg [1:0] PEG_Yvec_39__state;
  wire PEG_Yvec_40__ap_start_global__q0;
  wire PEG_Yvec_40__is_done__q0;
  wire PEG_Yvec_40__ap_done_global__q0;
  wire PEG_Yvec_40__ap_start;
  wire PEG_Yvec_40__ap_ready;
  wire PEG_Yvec_40__ap_done;
  wire PEG_Yvec_40__ap_idle;
  reg [1:0] PEG_Yvec_40__state;
  wire PEG_Yvec_41__ap_start_global__q0;
  wire PEG_Yvec_41__is_done__q0;
  wire PEG_Yvec_41__ap_done_global__q0;
  wire PEG_Yvec_41__ap_start;
  wire PEG_Yvec_41__ap_ready;
  wire PEG_Yvec_41__ap_done;
  wire PEG_Yvec_41__ap_idle;
  reg [1:0] PEG_Yvec_41__state;
  wire PEG_Yvec_42__ap_start_global__q0;
  wire PEG_Yvec_42__is_done__q0;
  wire PEG_Yvec_42__ap_done_global__q0;
  wire PEG_Yvec_42__ap_start;
  wire PEG_Yvec_42__ap_ready;
  wire PEG_Yvec_42__ap_done;
  wire PEG_Yvec_42__ap_idle;
  reg [1:0] PEG_Yvec_42__state;
  wire PEG_Yvec_43__ap_start_global__q0;
  wire PEG_Yvec_43__is_done__q0;
  wire PEG_Yvec_43__ap_done_global__q0;
  wire PEG_Yvec_43__ap_start;
  wire PEG_Yvec_43__ap_ready;
  wire PEG_Yvec_43__ap_done;
  wire PEG_Yvec_43__ap_idle;
  reg [1:0] PEG_Yvec_43__state;
  wire PEG_Yvec_44__ap_start_global__q0;
  wire PEG_Yvec_44__is_done__q0;
  wire PEG_Yvec_44__ap_done_global__q0;
  wire PEG_Yvec_44__ap_start;
  wire PEG_Yvec_44__ap_ready;
  wire PEG_Yvec_44__ap_done;
  wire PEG_Yvec_44__ap_idle;
  reg [1:0] PEG_Yvec_44__state;
  wire PEG_Yvec_45__ap_start_global__q0;
  wire PEG_Yvec_45__is_done__q0;
  wire PEG_Yvec_45__ap_done_global__q0;
  wire PEG_Yvec_45__ap_start;
  wire PEG_Yvec_45__ap_ready;
  wire PEG_Yvec_45__ap_done;
  wire PEG_Yvec_45__ap_idle;
  reg [1:0] PEG_Yvec_45__state;
  wire PEG_Yvec_46__ap_start_global__q0;
  wire PEG_Yvec_46__is_done__q0;
  wire PEG_Yvec_46__ap_done_global__q0;
  wire PEG_Yvec_46__ap_start;
  wire PEG_Yvec_46__ap_ready;
  wire PEG_Yvec_46__ap_done;
  wire PEG_Yvec_46__ap_idle;
  reg [1:0] PEG_Yvec_46__state;
  wire PEG_Yvec_47__ap_start_global__q0;
  wire PEG_Yvec_47__is_done__q0;
  wire PEG_Yvec_47__ap_done_global__q0;
  wire PEG_Yvec_47__ap_start;
  wire PEG_Yvec_47__ap_ready;
  wire PEG_Yvec_47__ap_done;
  wire PEG_Yvec_47__ap_idle;
  reg [1:0] PEG_Yvec_47__state;
  wire black_hole_float_v16_0__ap_start_global__q0;
  reg black_hole_float_v16_0__ap_start;
  wire black_hole_int_0__ap_start_global__q0;
  reg black_hole_int_0__ap_start;
  wire [31:0] read_A_0___NUM_A_LEN__q0;
  wire [31:0] read_A_0___P_N__q0;
  wire [63:0] read_A_0___edge_list_ch_0__q0;
  wire read_A_0__ap_start_global__q0;
  wire read_A_0__is_done__q0;
  wire read_A_0__ap_done_global__q0;
  wire read_A_0__ap_start;
  wire read_A_0__ap_ready;
  wire read_A_0__ap_done;
  wire read_A_0__ap_idle;
  reg [1:0] read_A_0__state;
  wire [31:0] read_A_1___NUM_A_LEN__q0;
  wire [31:0] read_A_1___P_N__q0;
  wire [63:0] read_A_1___edge_list_ch_1__q0;
  wire read_A_1__ap_start_global__q0;
  wire read_A_1__is_done__q0;
  wire read_A_1__ap_done_global__q0;
  wire read_A_1__ap_start;
  wire read_A_1__ap_ready;
  wire read_A_1__ap_done;
  wire read_A_1__ap_idle;
  reg [1:0] read_A_1__state;
  wire [31:0] read_A_2___NUM_A_LEN__q0;
  wire [31:0] read_A_2___P_N__q0;
  wire [63:0] read_A_2___edge_list_ch_2__q0;
  wire read_A_2__ap_start_global__q0;
  wire read_A_2__is_done__q0;
  wire read_A_2__ap_done_global__q0;
  wire read_A_2__ap_start;
  wire read_A_2__ap_ready;
  wire read_A_2__ap_done;
  wire read_A_2__ap_idle;
  reg [1:0] read_A_2__state;
  wire [31:0] read_A_3___NUM_A_LEN__q0;
  wire [31:0] read_A_3___P_N__q0;
  wire [63:0] read_A_3___edge_list_ch_3__q0;
  wire read_A_3__ap_start_global__q0;
  wire read_A_3__is_done__q0;
  wire read_A_3__ap_done_global__q0;
  wire read_A_3__ap_start;
  wire read_A_3__ap_ready;
  wire read_A_3__ap_done;
  wire read_A_3__ap_idle;
  reg [1:0] read_A_3__state;
  wire [31:0] read_A_4___NUM_A_LEN__q0;
  wire [31:0] read_A_4___P_N__q0;
  wire [63:0] read_A_4___edge_list_ch_4__q0;
  wire read_A_4__ap_start_global__q0;
  wire read_A_4__is_done__q0;
  wire read_A_4__ap_done_global__q0;
  wire read_A_4__ap_start;
  wire read_A_4__ap_ready;
  wire read_A_4__ap_done;
  wire read_A_4__ap_idle;
  reg [1:0] read_A_4__state;
  wire [31:0] read_A_5___NUM_A_LEN__q0;
  wire [31:0] read_A_5___P_N__q0;
  wire [63:0] read_A_5___edge_list_ch_5__q0;
  wire read_A_5__ap_start_global__q0;
  wire read_A_5__is_done__q0;
  wire read_A_5__ap_done_global__q0;
  wire read_A_5__ap_start;
  wire read_A_5__ap_ready;
  wire read_A_5__ap_done;
  wire read_A_5__ap_idle;
  reg [1:0] read_A_5__state;
  wire [31:0] read_A_6___NUM_A_LEN__q0;
  wire [31:0] read_A_6___P_N__q0;
  wire [63:0] read_A_6___edge_list_ch_6__q0;
  wire read_A_6__ap_start_global__q0;
  wire read_A_6__is_done__q0;
  wire read_A_6__ap_done_global__q0;
  wire read_A_6__ap_start;
  wire read_A_6__ap_ready;
  wire read_A_6__ap_done;
  wire read_A_6__ap_idle;
  reg [1:0] read_A_6__state;
  wire [31:0] read_A_7___NUM_A_LEN__q0;
  wire [31:0] read_A_7___P_N__q0;
  wire [63:0] read_A_7___edge_list_ch_7__q0;
  wire read_A_7__ap_start_global__q0;
  wire read_A_7__is_done__q0;
  wire read_A_7__ap_done_global__q0;
  wire read_A_7__ap_start;
  wire read_A_7__ap_ready;
  wire read_A_7__ap_done;
  wire read_A_7__ap_idle;
  reg [1:0] read_A_7__state;
  wire [31:0] read_A_8___NUM_A_LEN__q0;
  wire [31:0] read_A_8___P_N__q0;
  wire [63:0] read_A_8___edge_list_ch_8__q0;
  wire read_A_8__ap_start_global__q0;
  wire read_A_8__is_done__q0;
  wire read_A_8__ap_done_global__q0;
  wire read_A_8__ap_start;
  wire read_A_8__ap_ready;
  wire read_A_8__ap_done;
  wire read_A_8__ap_idle;
  reg [1:0] read_A_8__state;
  wire [31:0] read_A_9___NUM_A_LEN__q0;
  wire [31:0] read_A_9___P_N__q0;
  wire [63:0] read_A_9___edge_list_ch_9__q0;
  wire read_A_9__ap_start_global__q0;
  wire read_A_9__is_done__q0;
  wire read_A_9__ap_done_global__q0;
  wire read_A_9__ap_start;
  wire read_A_9__ap_ready;
  wire read_A_9__ap_done;
  wire read_A_9__ap_idle;
  reg [1:0] read_A_9__state;
  wire [31:0] read_A_10___NUM_A_LEN__q0;
  wire [31:0] read_A_10___P_N__q0;
  wire [63:0] read_A_10___edge_list_ch_10__q0;
  wire read_A_10__ap_start_global__q0;
  wire read_A_10__is_done__q0;
  wire read_A_10__ap_done_global__q0;
  wire read_A_10__ap_start;
  wire read_A_10__ap_ready;
  wire read_A_10__ap_done;
  wire read_A_10__ap_idle;
  reg [1:0] read_A_10__state;
  wire [31:0] read_A_11___NUM_A_LEN__q0;
  wire [31:0] read_A_11___P_N__q0;
  wire [63:0] read_A_11___edge_list_ch_11__q0;
  wire read_A_11__ap_start_global__q0;
  wire read_A_11__is_done__q0;
  wire read_A_11__ap_done_global__q0;
  wire read_A_11__ap_start;
  wire read_A_11__ap_ready;
  wire read_A_11__ap_done;
  wire read_A_11__ap_idle;
  reg [1:0] read_A_11__state;
  wire [31:0] read_A_12___NUM_A_LEN__q0;
  wire [31:0] read_A_12___P_N__q0;
  wire [63:0] read_A_12___edge_list_ch_12__q0;
  wire read_A_12__ap_start_global__q0;
  wire read_A_12__is_done__q0;
  wire read_A_12__ap_done_global__q0;
  wire read_A_12__ap_start;
  wire read_A_12__ap_ready;
  wire read_A_12__ap_done;
  wire read_A_12__ap_idle;
  reg [1:0] read_A_12__state;
  wire [31:0] read_A_13___NUM_A_LEN__q0;
  wire [31:0] read_A_13___P_N__q0;
  wire [63:0] read_A_13___edge_list_ch_13__q0;
  wire read_A_13__ap_start_global__q0;
  wire read_A_13__is_done__q0;
  wire read_A_13__ap_done_global__q0;
  wire read_A_13__ap_start;
  wire read_A_13__ap_ready;
  wire read_A_13__ap_done;
  wire read_A_13__ap_idle;
  reg [1:0] read_A_13__state;
  wire [31:0] read_A_14___NUM_A_LEN__q0;
  wire [31:0] read_A_14___P_N__q0;
  wire [63:0] read_A_14___edge_list_ch_14__q0;
  wire read_A_14__ap_start_global__q0;
  wire read_A_14__is_done__q0;
  wire read_A_14__ap_done_global__q0;
  wire read_A_14__ap_start;
  wire read_A_14__ap_ready;
  wire read_A_14__ap_done;
  wire read_A_14__ap_idle;
  reg [1:0] read_A_14__state;
  wire [31:0] read_A_15___NUM_A_LEN__q0;
  wire [31:0] read_A_15___P_N__q0;
  wire [63:0] read_A_15___edge_list_ch_15__q0;
  wire read_A_15__ap_start_global__q0;
  wire read_A_15__is_done__q0;
  wire read_A_15__ap_done_global__q0;
  wire read_A_15__ap_start;
  wire read_A_15__ap_ready;
  wire read_A_15__ap_done;
  wire read_A_15__ap_idle;
  reg [1:0] read_A_15__state;
  wire [31:0] read_A_16___NUM_A_LEN__q0;
  wire [31:0] read_A_16___P_N__q0;
  wire [63:0] read_A_16___edge_list_ch_16__q0;
  wire read_A_16__ap_start_global__q0;
  wire read_A_16__is_done__q0;
  wire read_A_16__ap_done_global__q0;
  wire read_A_16__ap_start;
  wire read_A_16__ap_ready;
  wire read_A_16__ap_done;
  wire read_A_16__ap_idle;
  reg [1:0] read_A_16__state;
  wire [31:0] read_A_17___NUM_A_LEN__q0;
  wire [31:0] read_A_17___P_N__q0;
  wire [63:0] read_A_17___edge_list_ch_17__q0;
  wire read_A_17__ap_start_global__q0;
  wire read_A_17__is_done__q0;
  wire read_A_17__ap_done_global__q0;
  wire read_A_17__ap_start;
  wire read_A_17__ap_ready;
  wire read_A_17__ap_done;
  wire read_A_17__ap_idle;
  reg [1:0] read_A_17__state;
  wire [31:0] read_A_18___NUM_A_LEN__q0;
  wire [31:0] read_A_18___P_N__q0;
  wire [63:0] read_A_18___edge_list_ch_18__q0;
  wire read_A_18__ap_start_global__q0;
  wire read_A_18__is_done__q0;
  wire read_A_18__ap_done_global__q0;
  wire read_A_18__ap_start;
  wire read_A_18__ap_ready;
  wire read_A_18__ap_done;
  wire read_A_18__ap_idle;
  reg [1:0] read_A_18__state;
  wire [31:0] read_A_19___NUM_A_LEN__q0;
  wire [31:0] read_A_19___P_N__q0;
  wire [63:0] read_A_19___edge_list_ch_19__q0;
  wire read_A_19__ap_start_global__q0;
  wire read_A_19__is_done__q0;
  wire read_A_19__ap_done_global__q0;
  wire read_A_19__ap_start;
  wire read_A_19__ap_ready;
  wire read_A_19__ap_done;
  wire read_A_19__ap_idle;
  reg [1:0] read_A_19__state;
  wire [31:0] read_A_20___NUM_A_LEN__q0;
  wire [31:0] read_A_20___P_N__q0;
  wire [63:0] read_A_20___edge_list_ch_20__q0;
  wire read_A_20__ap_start_global__q0;
  wire read_A_20__is_done__q0;
  wire read_A_20__ap_done_global__q0;
  wire read_A_20__ap_start;
  wire read_A_20__ap_ready;
  wire read_A_20__ap_done;
  wire read_A_20__ap_idle;
  reg [1:0] read_A_20__state;
  wire [31:0] read_A_21___NUM_A_LEN__q0;
  wire [31:0] read_A_21___P_N__q0;
  wire [63:0] read_A_21___edge_list_ch_21__q0;
  wire read_A_21__ap_start_global__q0;
  wire read_A_21__is_done__q0;
  wire read_A_21__ap_done_global__q0;
  wire read_A_21__ap_start;
  wire read_A_21__ap_ready;
  wire read_A_21__ap_done;
  wire read_A_21__ap_idle;
  reg [1:0] read_A_21__state;
  wire [31:0] read_A_22___NUM_A_LEN__q0;
  wire [31:0] read_A_22___P_N__q0;
  wire [63:0] read_A_22___edge_list_ch_22__q0;
  wire read_A_22__ap_start_global__q0;
  wire read_A_22__is_done__q0;
  wire read_A_22__ap_done_global__q0;
  wire read_A_22__ap_start;
  wire read_A_22__ap_ready;
  wire read_A_22__ap_done;
  wire read_A_22__ap_idle;
  reg [1:0] read_A_22__state;
  wire [31:0] read_A_23___NUM_A_LEN__q0;
  wire [31:0] read_A_23___P_N__q0;
  wire [63:0] read_A_23___edge_list_ch_23__q0;
  wire read_A_23__ap_start_global__q0;
  wire read_A_23__is_done__q0;
  wire read_A_23__ap_done_global__q0;
  wire read_A_23__ap_start;
  wire read_A_23__ap_ready;
  wire read_A_23__ap_done;
  wire read_A_23__ap_idle;
  reg [1:0] read_A_23__state;
  wire [31:0] read_A_24___NUM_A_LEN__q0;
  wire [31:0] read_A_24___P_N__q0;
  wire [63:0] read_A_24___edge_list_ch_24__q0;
  wire read_A_24__ap_start_global__q0;
  wire read_A_24__is_done__q0;
  wire read_A_24__ap_done_global__q0;
  wire read_A_24__ap_start;
  wire read_A_24__ap_ready;
  wire read_A_24__ap_done;
  wire read_A_24__ap_idle;
  reg [1:0] read_A_24__state;
  wire [31:0] read_A_25___NUM_A_LEN__q0;
  wire [31:0] read_A_25___P_N__q0;
  wire [63:0] read_A_25___edge_list_ch_25__q0;
  wire read_A_25__ap_start_global__q0;
  wire read_A_25__is_done__q0;
  wire read_A_25__ap_done_global__q0;
  wire read_A_25__ap_start;
  wire read_A_25__ap_ready;
  wire read_A_25__ap_done;
  wire read_A_25__ap_idle;
  reg [1:0] read_A_25__state;
  wire [31:0] read_A_26___NUM_A_LEN__q0;
  wire [31:0] read_A_26___P_N__q0;
  wire [63:0] read_A_26___edge_list_ch_26__q0;
  wire read_A_26__ap_start_global__q0;
  wire read_A_26__is_done__q0;
  wire read_A_26__ap_done_global__q0;
  wire read_A_26__ap_start;
  wire read_A_26__ap_ready;
  wire read_A_26__ap_done;
  wire read_A_26__ap_idle;
  reg [1:0] read_A_26__state;
  wire [31:0] read_A_27___NUM_A_LEN__q0;
  wire [31:0] read_A_27___P_N__q0;
  wire [63:0] read_A_27___edge_list_ch_27__q0;
  wire read_A_27__ap_start_global__q0;
  wire read_A_27__is_done__q0;
  wire read_A_27__ap_done_global__q0;
  wire read_A_27__ap_start;
  wire read_A_27__ap_ready;
  wire read_A_27__ap_done;
  wire read_A_27__ap_idle;
  reg [1:0] read_A_27__state;
  wire [31:0] read_A_28___NUM_A_LEN__q0;
  wire [31:0] read_A_28___P_N__q0;
  wire [63:0] read_A_28___edge_list_ch_28__q0;
  wire read_A_28__ap_start_global__q0;
  wire read_A_28__is_done__q0;
  wire read_A_28__ap_done_global__q0;
  wire read_A_28__ap_start;
  wire read_A_28__ap_ready;
  wire read_A_28__ap_done;
  wire read_A_28__ap_idle;
  reg [1:0] read_A_28__state;
  wire [31:0] read_A_29___NUM_A_LEN__q0;
  wire [31:0] read_A_29___P_N__q0;
  wire [63:0] read_A_29___edge_list_ch_29__q0;
  wire read_A_29__ap_start_global__q0;
  wire read_A_29__is_done__q0;
  wire read_A_29__ap_done_global__q0;
  wire read_A_29__ap_start;
  wire read_A_29__ap_ready;
  wire read_A_29__ap_done;
  wire read_A_29__ap_idle;
  reg [1:0] read_A_29__state;
  wire [31:0] read_A_30___NUM_A_LEN__q0;
  wire [31:0] read_A_30___P_N__q0;
  wire [63:0] read_A_30___edge_list_ch_30__q0;
  wire read_A_30__ap_start_global__q0;
  wire read_A_30__is_done__q0;
  wire read_A_30__ap_done_global__q0;
  wire read_A_30__ap_start;
  wire read_A_30__ap_ready;
  wire read_A_30__ap_done;
  wire read_A_30__ap_idle;
  reg [1:0] read_A_30__state;
  wire [31:0] read_A_31___NUM_A_LEN__q0;
  wire [31:0] read_A_31___P_N__q0;
  wire [63:0] read_A_31___edge_list_ch_31__q0;
  wire read_A_31__ap_start_global__q0;
  wire read_A_31__is_done__q0;
  wire read_A_31__ap_done_global__q0;
  wire read_A_31__ap_start;
  wire read_A_31__ap_ready;
  wire read_A_31__ap_done;
  wire read_A_31__ap_idle;
  reg [1:0] read_A_31__state;
  wire [31:0] read_A_32___NUM_A_LEN__q0;
  wire [31:0] read_A_32___P_N__q0;
  wire [63:0] read_A_32___edge_list_ch_32__q0;
  wire read_A_32__ap_start_global__q0;
  wire read_A_32__is_done__q0;
  wire read_A_32__ap_done_global__q0;
  wire read_A_32__ap_start;
  wire read_A_32__ap_ready;
  wire read_A_32__ap_done;
  wire read_A_32__ap_idle;
  reg [1:0] read_A_32__state;
  wire [31:0] read_A_33___NUM_A_LEN__q0;
  wire [31:0] read_A_33___P_N__q0;
  wire [63:0] read_A_33___edge_list_ch_33__q0;
  wire read_A_33__ap_start_global__q0;
  wire read_A_33__is_done__q0;
  wire read_A_33__ap_done_global__q0;
  wire read_A_33__ap_start;
  wire read_A_33__ap_ready;
  wire read_A_33__ap_done;
  wire read_A_33__ap_idle;
  reg [1:0] read_A_33__state;
  wire [31:0] read_A_34___NUM_A_LEN__q0;
  wire [31:0] read_A_34___P_N__q0;
  wire [63:0] read_A_34___edge_list_ch_34__q0;
  wire read_A_34__ap_start_global__q0;
  wire read_A_34__is_done__q0;
  wire read_A_34__ap_done_global__q0;
  wire read_A_34__ap_start;
  wire read_A_34__ap_ready;
  wire read_A_34__ap_done;
  wire read_A_34__ap_idle;
  reg [1:0] read_A_34__state;
  wire [31:0] read_A_35___NUM_A_LEN__q0;
  wire [31:0] read_A_35___P_N__q0;
  wire [63:0] read_A_35___edge_list_ch_35__q0;
  wire read_A_35__ap_start_global__q0;
  wire read_A_35__is_done__q0;
  wire read_A_35__ap_done_global__q0;
  wire read_A_35__ap_start;
  wire read_A_35__ap_ready;
  wire read_A_35__ap_done;
  wire read_A_35__ap_idle;
  reg [1:0] read_A_35__state;
  wire [31:0] read_A_36___NUM_A_LEN__q0;
  wire [31:0] read_A_36___P_N__q0;
  wire [63:0] read_A_36___edge_list_ch_36__q0;
  wire read_A_36__ap_start_global__q0;
  wire read_A_36__is_done__q0;
  wire read_A_36__ap_done_global__q0;
  wire read_A_36__ap_start;
  wire read_A_36__ap_ready;
  wire read_A_36__ap_done;
  wire read_A_36__ap_idle;
  reg [1:0] read_A_36__state;
  wire [31:0] read_A_37___NUM_A_LEN__q0;
  wire [31:0] read_A_37___P_N__q0;
  wire [63:0] read_A_37___edge_list_ch_37__q0;
  wire read_A_37__ap_start_global__q0;
  wire read_A_37__is_done__q0;
  wire read_A_37__ap_done_global__q0;
  wire read_A_37__ap_start;
  wire read_A_37__ap_ready;
  wire read_A_37__ap_done;
  wire read_A_37__ap_idle;
  reg [1:0] read_A_37__state;
  wire [31:0] read_A_38___NUM_A_LEN__q0;
  wire [31:0] read_A_38___P_N__q0;
  wire [63:0] read_A_38___edge_list_ch_38__q0;
  wire read_A_38__ap_start_global__q0;
  wire read_A_38__is_done__q0;
  wire read_A_38__ap_done_global__q0;
  wire read_A_38__ap_start;
  wire read_A_38__ap_ready;
  wire read_A_38__ap_done;
  wire read_A_38__ap_idle;
  reg [1:0] read_A_38__state;
  wire [31:0] read_A_39___NUM_A_LEN__q0;
  wire [31:0] read_A_39___P_N__q0;
  wire [63:0] read_A_39___edge_list_ch_39__q0;
  wire read_A_39__ap_start_global__q0;
  wire read_A_39__is_done__q0;
  wire read_A_39__ap_done_global__q0;
  wire read_A_39__ap_start;
  wire read_A_39__ap_ready;
  wire read_A_39__ap_done;
  wire read_A_39__ap_idle;
  reg [1:0] read_A_39__state;
  wire [31:0] read_A_40___NUM_A_LEN__q0;
  wire [31:0] read_A_40___P_N__q0;
  wire [63:0] read_A_40___edge_list_ch_40__q0;
  wire read_A_40__ap_start_global__q0;
  wire read_A_40__is_done__q0;
  wire read_A_40__ap_done_global__q0;
  wire read_A_40__ap_start;
  wire read_A_40__ap_ready;
  wire read_A_40__ap_done;
  wire read_A_40__ap_idle;
  reg [1:0] read_A_40__state;
  wire [31:0] read_A_41___NUM_A_LEN__q0;
  wire [31:0] read_A_41___P_N__q0;
  wire [63:0] read_A_41___edge_list_ch_41__q0;
  wire read_A_41__ap_start_global__q0;
  wire read_A_41__is_done__q0;
  wire read_A_41__ap_done_global__q0;
  wire read_A_41__ap_start;
  wire read_A_41__ap_ready;
  wire read_A_41__ap_done;
  wire read_A_41__ap_idle;
  reg [1:0] read_A_41__state;
  wire [31:0] read_A_42___NUM_A_LEN__q0;
  wire [31:0] read_A_42___P_N__q0;
  wire [63:0] read_A_42___edge_list_ch_42__q0;
  wire read_A_42__ap_start_global__q0;
  wire read_A_42__is_done__q0;
  wire read_A_42__ap_done_global__q0;
  wire read_A_42__ap_start;
  wire read_A_42__ap_ready;
  wire read_A_42__ap_done;
  wire read_A_42__ap_idle;
  reg [1:0] read_A_42__state;
  wire [31:0] read_A_43___NUM_A_LEN__q0;
  wire [31:0] read_A_43___P_N__q0;
  wire [63:0] read_A_43___edge_list_ch_43__q0;
  wire read_A_43__ap_start_global__q0;
  wire read_A_43__is_done__q0;
  wire read_A_43__ap_done_global__q0;
  wire read_A_43__ap_start;
  wire read_A_43__ap_ready;
  wire read_A_43__ap_done;
  wire read_A_43__ap_idle;
  reg [1:0] read_A_43__state;
  wire [31:0] read_A_44___NUM_A_LEN__q0;
  wire [31:0] read_A_44___P_N__q0;
  wire [63:0] read_A_44___edge_list_ch_44__q0;
  wire read_A_44__ap_start_global__q0;
  wire read_A_44__is_done__q0;
  wire read_A_44__ap_done_global__q0;
  wire read_A_44__ap_start;
  wire read_A_44__ap_ready;
  wire read_A_44__ap_done;
  wire read_A_44__ap_idle;
  reg [1:0] read_A_44__state;
  wire [31:0] read_A_45___NUM_A_LEN__q0;
  wire [31:0] read_A_45___P_N__q0;
  wire [63:0] read_A_45___edge_list_ch_45__q0;
  wire read_A_45__ap_start_global__q0;
  wire read_A_45__is_done__q0;
  wire read_A_45__ap_done_global__q0;
  wire read_A_45__ap_start;
  wire read_A_45__ap_ready;
  wire read_A_45__ap_done;
  wire read_A_45__ap_idle;
  reg [1:0] read_A_45__state;
  wire [31:0] read_A_46___NUM_A_LEN__q0;
  wire [31:0] read_A_46___P_N__q0;
  wire [63:0] read_A_46___edge_list_ch_46__q0;
  wire read_A_46__ap_start_global__q0;
  wire read_A_46__is_done__q0;
  wire read_A_46__ap_done_global__q0;
  wire read_A_46__ap_start;
  wire read_A_46__ap_ready;
  wire read_A_46__ap_done;
  wire read_A_46__ap_idle;
  reg [1:0] read_A_46__state;
  wire [31:0] read_A_47___NUM_A_LEN__q0;
  wire [31:0] read_A_47___P_N__q0;
  wire [63:0] read_A_47___edge_list_ch_47__q0;
  wire read_A_47__ap_start_global__q0;
  wire read_A_47__is_done__q0;
  wire read_A_47__ap_done_global__q0;
  wire read_A_47__ap_start;
  wire read_A_47__ap_ready;
  wire read_A_47__ap_done;
  wire read_A_47__ap_idle;
  reg [1:0] read_A_47__state;
  wire [31:0] read_X_0___K__q0;
  wire [31:0] read_X_0___P_N__q0;
  wire [63:0] read_X_0___vec_X__q0;
  wire read_X_0__ap_start_global__q0;
  wire read_X_0__is_done__q0;
  wire read_X_0__ap_done_global__q0;
  wire read_X_0__ap_start;
  wire read_X_0__ap_ready;
  wire read_X_0__ap_done;
  wire read_X_0__ap_idle;
  reg [1:0] read_X_0__state;
  wire [31:0] read_Y_0___M__q0;
  wire [31:0] read_Y_0___P_N__q0;
  wire [63:0] read_Y_0___vec_Y__q0;
  wire read_Y_0__ap_start_global__q0;
  wire read_Y_0__is_done__q0;
  wire read_Y_0__ap_done_global__q0;
  wire read_Y_0__ap_start;
  wire read_Y_0__ap_ready;
  wire read_Y_0__ap_done;
  wire read_Y_0__ap_idle;
  reg [1:0] read_Y_0__state;
  wire [31:0] read_edge_list_ptr_0___K__q0;
  wire [31:0] read_edge_list_ptr_0___M__q0;
  wire [31:0] read_edge_list_ptr_0___NUM_ITE__q0;
  wire [31:0] read_edge_list_ptr_0___P_N__q0;
  wire [63:0] read_edge_list_ptr_0___edge_list_ptr__q0;
  wire read_edge_list_ptr_0__ap_start_global__q0;
  wire read_edge_list_ptr_0__is_done__q0;
  wire read_edge_list_ptr_0__ap_done_global__q0;
  wire read_edge_list_ptr_0__ap_start;
  wire read_edge_list_ptr_0__ap_ready;
  wire read_edge_list_ptr_0__ap_done;
  wire read_edge_list_ptr_0__ap_idle;
  reg [1:0] read_edge_list_ptr_0__state;
  wire [31:0] write_Y_0___M__q0;
  wire [31:0] write_Y_0___P_N__q0;
  wire [63:0] write_Y_0___vec_Y_out__q0;
  wire write_Y_0__ap_start_global__q0;
  wire write_Y_0__is_done__q0;
  wire write_Y_0__ap_done_global__q0;
  wire write_Y_0__ap_start;
  wire write_Y_0__ap_ready;
  wire write_Y_0__ap_done;
  wire write_Y_0__ap_idle;
  reg [1:0] write_Y_0__state;
  reg [1:0] tapa_state;
  reg [0:0] countdown;
  wire ap_start__q0;
  wire ap_done__q0;
  assign Arbiter_Y_0___M__q0 = M;
  assign Arbiter_Y_0___P_N__q0 = P_N;
  assign Arbiter_Y_0__ap_start_global__q0 = ap_start__q0;
  assign Arbiter_Y_0__is_done__q0 = (Arbiter_Y_0__state == 2'b10);
  assign Arbiter_Y_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Arbiter_Y_0__state <= 2'b00;
    end else begin
      if(Arbiter_Y_0__state == 2'b00) begin
        if(Arbiter_Y_0__ap_start_global__q0) begin
          Arbiter_Y_0__state <= 2'b01;
        end 
      end 
      if(Arbiter_Y_0__state == 2'b01) begin
        if(Arbiter_Y_0__ap_ready) begin
          if(Arbiter_Y_0__ap_done) begin
            Arbiter_Y_0__state <= 2'b10;
          end else begin
            Arbiter_Y_0__state <= 2'b11;
          end
        end 
      end 
      if(Arbiter_Y_0__state == 2'b11) begin
        if(Arbiter_Y_0__ap_done) begin
          Arbiter_Y_0__state <= 2'b10;
        end 
      end 
      if(Arbiter_Y_0__state == 2'b10) begin
        if(Arbiter_Y_0__ap_done_global__q0) begin
          Arbiter_Y_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign Arbiter_Y_0__ap_start = (Arbiter_Y_0__state == 2'b01);
  assign Arbiter_Y_1___M__q0 = M;
  assign Arbiter_Y_1___P_N__q0 = P_N;
  assign Arbiter_Y_1__ap_start_global__q0 = ap_start__q0;
  assign Arbiter_Y_1__is_done__q0 = (Arbiter_Y_1__state == 2'b10);
  assign Arbiter_Y_1__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Arbiter_Y_1__state <= 2'b00;
    end else begin
      if(Arbiter_Y_1__state == 2'b00) begin
        if(Arbiter_Y_1__ap_start_global__q0) begin
          Arbiter_Y_1__state <= 2'b01;
        end 
      end 
      if(Arbiter_Y_1__state == 2'b01) begin
        if(Arbiter_Y_1__ap_ready) begin
          if(Arbiter_Y_1__ap_done) begin
            Arbiter_Y_1__state <= 2'b10;
          end else begin
            Arbiter_Y_1__state <= 2'b11;
          end
        end 
      end 
      if(Arbiter_Y_1__state == 2'b11) begin
        if(Arbiter_Y_1__ap_done) begin
          Arbiter_Y_1__state <= 2'b10;
        end 
      end 
      if(Arbiter_Y_1__state == 2'b10) begin
        if(Arbiter_Y_1__ap_done_global__q0) begin
          Arbiter_Y_1__state <= 2'b00;
        end 
      end 
    end
  end

  assign Arbiter_Y_1__ap_start = (Arbiter_Y_1__state == 2'b01);
  assign Arbiter_Y_2___M__q0 = M;
  assign Arbiter_Y_2___P_N__q0 = P_N;
  assign Arbiter_Y_2__ap_start_global__q0 = ap_start__q0;
  assign Arbiter_Y_2__is_done__q0 = (Arbiter_Y_2__state == 2'b10);
  assign Arbiter_Y_2__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Arbiter_Y_2__state <= 2'b00;
    end else begin
      if(Arbiter_Y_2__state == 2'b00) begin
        if(Arbiter_Y_2__ap_start_global__q0) begin
          Arbiter_Y_2__state <= 2'b01;
        end 
      end 
      if(Arbiter_Y_2__state == 2'b01) begin
        if(Arbiter_Y_2__ap_ready) begin
          if(Arbiter_Y_2__ap_done) begin
            Arbiter_Y_2__state <= 2'b10;
          end else begin
            Arbiter_Y_2__state <= 2'b11;
          end
        end 
      end 
      if(Arbiter_Y_2__state == 2'b11) begin
        if(Arbiter_Y_2__ap_done) begin
          Arbiter_Y_2__state <= 2'b10;
        end 
      end 
      if(Arbiter_Y_2__state == 2'b10) begin
        if(Arbiter_Y_2__ap_done_global__q0) begin
          Arbiter_Y_2__state <= 2'b00;
        end 
      end 
    end
  end

  assign Arbiter_Y_2__ap_start = (Arbiter_Y_2__state == 2'b01);
  assign Arbiter_Y_3___M__q0 = M;
  assign Arbiter_Y_3___P_N__q0 = P_N;
  assign Arbiter_Y_3__ap_start_global__q0 = ap_start__q0;
  assign Arbiter_Y_3__is_done__q0 = (Arbiter_Y_3__state == 2'b10);
  assign Arbiter_Y_3__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Arbiter_Y_3__state <= 2'b00;
    end else begin
      if(Arbiter_Y_3__state == 2'b00) begin
        if(Arbiter_Y_3__ap_start_global__q0) begin
          Arbiter_Y_3__state <= 2'b01;
        end 
      end 
      if(Arbiter_Y_3__state == 2'b01) begin
        if(Arbiter_Y_3__ap_ready) begin
          if(Arbiter_Y_3__ap_done) begin
            Arbiter_Y_3__state <= 2'b10;
          end else begin
            Arbiter_Y_3__state <= 2'b11;
          end
        end 
      end 
      if(Arbiter_Y_3__state == 2'b11) begin
        if(Arbiter_Y_3__ap_done) begin
          Arbiter_Y_3__state <= 2'b10;
        end 
      end 
      if(Arbiter_Y_3__state == 2'b10) begin
        if(Arbiter_Y_3__ap_done_global__q0) begin
          Arbiter_Y_3__state <= 2'b00;
        end 
      end 
    end
  end

  assign Arbiter_Y_3__ap_start = (Arbiter_Y_3__state == 2'b01);
  assign Arbiter_Y_4___M__q0 = M;
  assign Arbiter_Y_4___P_N__q0 = P_N;
  assign Arbiter_Y_4__ap_start_global__q0 = ap_start__q0;
  assign Arbiter_Y_4__is_done__q0 = (Arbiter_Y_4__state == 2'b10);
  assign Arbiter_Y_4__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Arbiter_Y_4__state <= 2'b00;
    end else begin
      if(Arbiter_Y_4__state == 2'b00) begin
        if(Arbiter_Y_4__ap_start_global__q0) begin
          Arbiter_Y_4__state <= 2'b01;
        end 
      end 
      if(Arbiter_Y_4__state == 2'b01) begin
        if(Arbiter_Y_4__ap_ready) begin
          if(Arbiter_Y_4__ap_done) begin
            Arbiter_Y_4__state <= 2'b10;
          end else begin
            Arbiter_Y_4__state <= 2'b11;
          end
        end 
      end 
      if(Arbiter_Y_4__state == 2'b11) begin
        if(Arbiter_Y_4__ap_done) begin
          Arbiter_Y_4__state <= 2'b10;
        end 
      end 
      if(Arbiter_Y_4__state == 2'b10) begin
        if(Arbiter_Y_4__ap_done_global__q0) begin
          Arbiter_Y_4__state <= 2'b00;
        end 
      end 
    end
  end

  assign Arbiter_Y_4__ap_start = (Arbiter_Y_4__state == 2'b01);
  assign Arbiter_Y_5___M__q0 = M;
  assign Arbiter_Y_5___P_N__q0 = P_N;
  assign Arbiter_Y_5__ap_start_global__q0 = ap_start__q0;
  assign Arbiter_Y_5__is_done__q0 = (Arbiter_Y_5__state == 2'b10);
  assign Arbiter_Y_5__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Arbiter_Y_5__state <= 2'b00;
    end else begin
      if(Arbiter_Y_5__state == 2'b00) begin
        if(Arbiter_Y_5__ap_start_global__q0) begin
          Arbiter_Y_5__state <= 2'b01;
        end 
      end 
      if(Arbiter_Y_5__state == 2'b01) begin
        if(Arbiter_Y_5__ap_ready) begin
          if(Arbiter_Y_5__ap_done) begin
            Arbiter_Y_5__state <= 2'b10;
          end else begin
            Arbiter_Y_5__state <= 2'b11;
          end
        end 
      end 
      if(Arbiter_Y_5__state == 2'b11) begin
        if(Arbiter_Y_5__ap_done) begin
          Arbiter_Y_5__state <= 2'b10;
        end 
      end 
      if(Arbiter_Y_5__state == 2'b10) begin
        if(Arbiter_Y_5__ap_done_global__q0) begin
          Arbiter_Y_5__state <= 2'b00;
        end 
      end 
    end
  end

  assign Arbiter_Y_5__ap_start = (Arbiter_Y_5__state == 2'b01);
  assign Arbiter_Y_6___M__q0 = M;
  assign Arbiter_Y_6___P_N__q0 = P_N;
  assign Arbiter_Y_6__ap_start_global__q0 = ap_start__q0;
  assign Arbiter_Y_6__is_done__q0 = (Arbiter_Y_6__state == 2'b10);
  assign Arbiter_Y_6__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Arbiter_Y_6__state <= 2'b00;
    end else begin
      if(Arbiter_Y_6__state == 2'b00) begin
        if(Arbiter_Y_6__ap_start_global__q0) begin
          Arbiter_Y_6__state <= 2'b01;
        end 
      end 
      if(Arbiter_Y_6__state == 2'b01) begin
        if(Arbiter_Y_6__ap_ready) begin
          if(Arbiter_Y_6__ap_done) begin
            Arbiter_Y_6__state <= 2'b10;
          end else begin
            Arbiter_Y_6__state <= 2'b11;
          end
        end 
      end 
      if(Arbiter_Y_6__state == 2'b11) begin
        if(Arbiter_Y_6__ap_done) begin
          Arbiter_Y_6__state <= 2'b10;
        end 
      end 
      if(Arbiter_Y_6__state == 2'b10) begin
        if(Arbiter_Y_6__ap_done_global__q0) begin
          Arbiter_Y_6__state <= 2'b00;
        end 
      end 
    end
  end

  assign Arbiter_Y_6__ap_start = (Arbiter_Y_6__state == 2'b01);
  assign Arbiter_Y_7___M__q0 = M;
  assign Arbiter_Y_7___P_N__q0 = P_N;
  assign Arbiter_Y_7__ap_start_global__q0 = ap_start__q0;
  assign Arbiter_Y_7__is_done__q0 = (Arbiter_Y_7__state == 2'b10);
  assign Arbiter_Y_7__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Arbiter_Y_7__state <= 2'b00;
    end else begin
      if(Arbiter_Y_7__state == 2'b00) begin
        if(Arbiter_Y_7__ap_start_global__q0) begin
          Arbiter_Y_7__state <= 2'b01;
        end 
      end 
      if(Arbiter_Y_7__state == 2'b01) begin
        if(Arbiter_Y_7__ap_ready) begin
          if(Arbiter_Y_7__ap_done) begin
            Arbiter_Y_7__state <= 2'b10;
          end else begin
            Arbiter_Y_7__state <= 2'b11;
          end
        end 
      end 
      if(Arbiter_Y_7__state == 2'b11) begin
        if(Arbiter_Y_7__ap_done) begin
          Arbiter_Y_7__state <= 2'b10;
        end 
      end 
      if(Arbiter_Y_7__state == 2'b10) begin
        if(Arbiter_Y_7__ap_done_global__q0) begin
          Arbiter_Y_7__state <= 2'b00;
        end 
      end 
    end
  end

  assign Arbiter_Y_7__ap_start = (Arbiter_Y_7__state == 2'b01);
  assign FloatvAddFloatv_0__ap_start_global__q0 = ap_start__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      FloatvAddFloatv_0__ap_start <= 1'b0;
    end else if(FloatvAddFloatv_0__ap_start_global__q0) begin
      FloatvAddFloatv_0__ap_start <= 1'b1;
    end 
  end

  assign FloatvMultConst_0___M__q0 = M;
  assign FloatvMultConst_0___P_N__q0 = P_N;
  assign FloatvMultConst_0___alpha_u__q0 = alpha_u;
  assign FloatvMultConst_0__ap_start_global__q0 = ap_start__q0;
  assign FloatvMultConst_0__is_done__q0 = (FloatvMultConst_0__state == 2'b10);
  assign FloatvMultConst_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      FloatvMultConst_0__state <= 2'b00;
    end else begin
      if(FloatvMultConst_0__state == 2'b00) begin
        if(FloatvMultConst_0__ap_start_global__q0) begin
          FloatvMultConst_0__state <= 2'b01;
        end 
      end 
      if(FloatvMultConst_0__state == 2'b01) begin
        if(FloatvMultConst_0__ap_ready) begin
          if(FloatvMultConst_0__ap_done) begin
            FloatvMultConst_0__state <= 2'b10;
          end else begin
            FloatvMultConst_0__state <= 2'b11;
          end
        end 
      end 
      if(FloatvMultConst_0__state == 2'b11) begin
        if(FloatvMultConst_0__ap_done) begin
          FloatvMultConst_0__state <= 2'b10;
        end 
      end 
      if(FloatvMultConst_0__state == 2'b10) begin
        if(FloatvMultConst_0__ap_done_global__q0) begin
          FloatvMultConst_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign FloatvMultConst_0__ap_start = (FloatvMultConst_0__state == 2'b01);
  assign FloatvMultConst_1___M__q0 = M;
  assign FloatvMultConst_1___P_N__q0 = P_N;
  assign FloatvMultConst_1___beta_u__q0 = beta_u;
  assign FloatvMultConst_1__ap_start_global__q0 = ap_start__q0;
  assign FloatvMultConst_1__is_done__q0 = (FloatvMultConst_1__state == 2'b10);
  assign FloatvMultConst_1__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      FloatvMultConst_1__state <= 2'b00;
    end else begin
      if(FloatvMultConst_1__state == 2'b00) begin
        if(FloatvMultConst_1__ap_start_global__q0) begin
          FloatvMultConst_1__state <= 2'b01;
        end 
      end 
      if(FloatvMultConst_1__state == 2'b01) begin
        if(FloatvMultConst_1__ap_ready) begin
          if(FloatvMultConst_1__ap_done) begin
            FloatvMultConst_1__state <= 2'b10;
          end else begin
            FloatvMultConst_1__state <= 2'b11;
          end
        end 
      end 
      if(FloatvMultConst_1__state == 2'b11) begin
        if(FloatvMultConst_1__ap_done) begin
          FloatvMultConst_1__state <= 2'b10;
        end 
      end 
      if(FloatvMultConst_1__state == 2'b10) begin
        if(FloatvMultConst_1__ap_done_global__q0) begin
          FloatvMultConst_1__state <= 2'b00;
        end 
      end 
    end
  end

  assign FloatvMultConst_1__ap_start = (FloatvMultConst_1__state == 2'b01);
  assign Merger_Y_0__ap_start_global__q0 = ap_start__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      Merger_Y_0__ap_start <= 1'b0;
    end else if(Merger_Y_0__ap_start_global__q0) begin
      Merger_Y_0__ap_start <= 1'b1;
    end 
  end

  assign PEG_Xvec_0__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_0__is_done__q0 = (PEG_Xvec_0__state == 2'b10);
  assign PEG_Xvec_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_0__state <= 2'b00;
    end else begin
      if(PEG_Xvec_0__state == 2'b00) begin
        if(PEG_Xvec_0__ap_start_global__q0) begin
          PEG_Xvec_0__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_0__state == 2'b01) begin
        if(PEG_Xvec_0__ap_ready) begin
          if(PEG_Xvec_0__ap_done) begin
            PEG_Xvec_0__state <= 2'b10;
          end else begin
            PEG_Xvec_0__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_0__state == 2'b11) begin
        if(PEG_Xvec_0__ap_done) begin
          PEG_Xvec_0__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_0__state == 2'b10) begin
        if(PEG_Xvec_0__ap_done_global__q0) begin
          PEG_Xvec_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_0__ap_start = (PEG_Xvec_0__state == 2'b01);
  assign PEG_Xvec_1__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_1__is_done__q0 = (PEG_Xvec_1__state == 2'b10);
  assign PEG_Xvec_1__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_1__state <= 2'b00;
    end else begin
      if(PEG_Xvec_1__state == 2'b00) begin
        if(PEG_Xvec_1__ap_start_global__q0) begin
          PEG_Xvec_1__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_1__state == 2'b01) begin
        if(PEG_Xvec_1__ap_ready) begin
          if(PEG_Xvec_1__ap_done) begin
            PEG_Xvec_1__state <= 2'b10;
          end else begin
            PEG_Xvec_1__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_1__state == 2'b11) begin
        if(PEG_Xvec_1__ap_done) begin
          PEG_Xvec_1__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_1__state == 2'b10) begin
        if(PEG_Xvec_1__ap_done_global__q0) begin
          PEG_Xvec_1__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_1__ap_start = (PEG_Xvec_1__state == 2'b01);
  assign PEG_Xvec_2__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_2__is_done__q0 = (PEG_Xvec_2__state == 2'b10);
  assign PEG_Xvec_2__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_2__state <= 2'b00;
    end else begin
      if(PEG_Xvec_2__state == 2'b00) begin
        if(PEG_Xvec_2__ap_start_global__q0) begin
          PEG_Xvec_2__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_2__state == 2'b01) begin
        if(PEG_Xvec_2__ap_ready) begin
          if(PEG_Xvec_2__ap_done) begin
            PEG_Xvec_2__state <= 2'b10;
          end else begin
            PEG_Xvec_2__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_2__state == 2'b11) begin
        if(PEG_Xvec_2__ap_done) begin
          PEG_Xvec_2__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_2__state == 2'b10) begin
        if(PEG_Xvec_2__ap_done_global__q0) begin
          PEG_Xvec_2__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_2__ap_start = (PEG_Xvec_2__state == 2'b01);
  assign PEG_Xvec_3__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_3__is_done__q0 = (PEG_Xvec_3__state == 2'b10);
  assign PEG_Xvec_3__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_3__state <= 2'b00;
    end else begin
      if(PEG_Xvec_3__state == 2'b00) begin
        if(PEG_Xvec_3__ap_start_global__q0) begin
          PEG_Xvec_3__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_3__state == 2'b01) begin
        if(PEG_Xvec_3__ap_ready) begin
          if(PEG_Xvec_3__ap_done) begin
            PEG_Xvec_3__state <= 2'b10;
          end else begin
            PEG_Xvec_3__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_3__state == 2'b11) begin
        if(PEG_Xvec_3__ap_done) begin
          PEG_Xvec_3__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_3__state == 2'b10) begin
        if(PEG_Xvec_3__ap_done_global__q0) begin
          PEG_Xvec_3__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_3__ap_start = (PEG_Xvec_3__state == 2'b01);
  assign PEG_Xvec_4__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_4__is_done__q0 = (PEG_Xvec_4__state == 2'b10);
  assign PEG_Xvec_4__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_4__state <= 2'b00;
    end else begin
      if(PEG_Xvec_4__state == 2'b00) begin
        if(PEG_Xvec_4__ap_start_global__q0) begin
          PEG_Xvec_4__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_4__state == 2'b01) begin
        if(PEG_Xvec_4__ap_ready) begin
          if(PEG_Xvec_4__ap_done) begin
            PEG_Xvec_4__state <= 2'b10;
          end else begin
            PEG_Xvec_4__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_4__state == 2'b11) begin
        if(PEG_Xvec_4__ap_done) begin
          PEG_Xvec_4__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_4__state == 2'b10) begin
        if(PEG_Xvec_4__ap_done_global__q0) begin
          PEG_Xvec_4__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_4__ap_start = (PEG_Xvec_4__state == 2'b01);
  assign PEG_Xvec_5__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_5__is_done__q0 = (PEG_Xvec_5__state == 2'b10);
  assign PEG_Xvec_5__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_5__state <= 2'b00;
    end else begin
      if(PEG_Xvec_5__state == 2'b00) begin
        if(PEG_Xvec_5__ap_start_global__q0) begin
          PEG_Xvec_5__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_5__state == 2'b01) begin
        if(PEG_Xvec_5__ap_ready) begin
          if(PEG_Xvec_5__ap_done) begin
            PEG_Xvec_5__state <= 2'b10;
          end else begin
            PEG_Xvec_5__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_5__state == 2'b11) begin
        if(PEG_Xvec_5__ap_done) begin
          PEG_Xvec_5__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_5__state == 2'b10) begin
        if(PEG_Xvec_5__ap_done_global__q0) begin
          PEG_Xvec_5__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_5__ap_start = (PEG_Xvec_5__state == 2'b01);
  assign PEG_Xvec_6__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_6__is_done__q0 = (PEG_Xvec_6__state == 2'b10);
  assign PEG_Xvec_6__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_6__state <= 2'b00;
    end else begin
      if(PEG_Xvec_6__state == 2'b00) begin
        if(PEG_Xvec_6__ap_start_global__q0) begin
          PEG_Xvec_6__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_6__state == 2'b01) begin
        if(PEG_Xvec_6__ap_ready) begin
          if(PEG_Xvec_6__ap_done) begin
            PEG_Xvec_6__state <= 2'b10;
          end else begin
            PEG_Xvec_6__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_6__state == 2'b11) begin
        if(PEG_Xvec_6__ap_done) begin
          PEG_Xvec_6__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_6__state == 2'b10) begin
        if(PEG_Xvec_6__ap_done_global__q0) begin
          PEG_Xvec_6__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_6__ap_start = (PEG_Xvec_6__state == 2'b01);
  assign PEG_Xvec_7__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_7__is_done__q0 = (PEG_Xvec_7__state == 2'b10);
  assign PEG_Xvec_7__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_7__state <= 2'b00;
    end else begin
      if(PEG_Xvec_7__state == 2'b00) begin
        if(PEG_Xvec_7__ap_start_global__q0) begin
          PEG_Xvec_7__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_7__state == 2'b01) begin
        if(PEG_Xvec_7__ap_ready) begin
          if(PEG_Xvec_7__ap_done) begin
            PEG_Xvec_7__state <= 2'b10;
          end else begin
            PEG_Xvec_7__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_7__state == 2'b11) begin
        if(PEG_Xvec_7__ap_done) begin
          PEG_Xvec_7__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_7__state == 2'b10) begin
        if(PEG_Xvec_7__ap_done_global__q0) begin
          PEG_Xvec_7__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_7__ap_start = (PEG_Xvec_7__state == 2'b01);
  assign PEG_Xvec_8__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_8__is_done__q0 = (PEG_Xvec_8__state == 2'b10);
  assign PEG_Xvec_8__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_8__state <= 2'b00;
    end else begin
      if(PEG_Xvec_8__state == 2'b00) begin
        if(PEG_Xvec_8__ap_start_global__q0) begin
          PEG_Xvec_8__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_8__state == 2'b01) begin
        if(PEG_Xvec_8__ap_ready) begin
          if(PEG_Xvec_8__ap_done) begin
            PEG_Xvec_8__state <= 2'b10;
          end else begin
            PEG_Xvec_8__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_8__state == 2'b11) begin
        if(PEG_Xvec_8__ap_done) begin
          PEG_Xvec_8__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_8__state == 2'b10) begin
        if(PEG_Xvec_8__ap_done_global__q0) begin
          PEG_Xvec_8__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_8__ap_start = (PEG_Xvec_8__state == 2'b01);
  assign PEG_Xvec_9__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_9__is_done__q0 = (PEG_Xvec_9__state == 2'b10);
  assign PEG_Xvec_9__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_9__state <= 2'b00;
    end else begin
      if(PEG_Xvec_9__state == 2'b00) begin
        if(PEG_Xvec_9__ap_start_global__q0) begin
          PEG_Xvec_9__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_9__state == 2'b01) begin
        if(PEG_Xvec_9__ap_ready) begin
          if(PEG_Xvec_9__ap_done) begin
            PEG_Xvec_9__state <= 2'b10;
          end else begin
            PEG_Xvec_9__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_9__state == 2'b11) begin
        if(PEG_Xvec_9__ap_done) begin
          PEG_Xvec_9__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_9__state == 2'b10) begin
        if(PEG_Xvec_9__ap_done_global__q0) begin
          PEG_Xvec_9__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_9__ap_start = (PEG_Xvec_9__state == 2'b01);
  assign PEG_Xvec_10__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_10__is_done__q0 = (PEG_Xvec_10__state == 2'b10);
  assign PEG_Xvec_10__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_10__state <= 2'b00;
    end else begin
      if(PEG_Xvec_10__state == 2'b00) begin
        if(PEG_Xvec_10__ap_start_global__q0) begin
          PEG_Xvec_10__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_10__state == 2'b01) begin
        if(PEG_Xvec_10__ap_ready) begin
          if(PEG_Xvec_10__ap_done) begin
            PEG_Xvec_10__state <= 2'b10;
          end else begin
            PEG_Xvec_10__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_10__state == 2'b11) begin
        if(PEG_Xvec_10__ap_done) begin
          PEG_Xvec_10__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_10__state == 2'b10) begin
        if(PEG_Xvec_10__ap_done_global__q0) begin
          PEG_Xvec_10__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_10__ap_start = (PEG_Xvec_10__state == 2'b01);
  assign PEG_Xvec_11__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_11__is_done__q0 = (PEG_Xvec_11__state == 2'b10);
  assign PEG_Xvec_11__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_11__state <= 2'b00;
    end else begin
      if(PEG_Xvec_11__state == 2'b00) begin
        if(PEG_Xvec_11__ap_start_global__q0) begin
          PEG_Xvec_11__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_11__state == 2'b01) begin
        if(PEG_Xvec_11__ap_ready) begin
          if(PEG_Xvec_11__ap_done) begin
            PEG_Xvec_11__state <= 2'b10;
          end else begin
            PEG_Xvec_11__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_11__state == 2'b11) begin
        if(PEG_Xvec_11__ap_done) begin
          PEG_Xvec_11__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_11__state == 2'b10) begin
        if(PEG_Xvec_11__ap_done_global__q0) begin
          PEG_Xvec_11__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_11__ap_start = (PEG_Xvec_11__state == 2'b01);
  assign PEG_Xvec_12__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_12__is_done__q0 = (PEG_Xvec_12__state == 2'b10);
  assign PEG_Xvec_12__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_12__state <= 2'b00;
    end else begin
      if(PEG_Xvec_12__state == 2'b00) begin
        if(PEG_Xvec_12__ap_start_global__q0) begin
          PEG_Xvec_12__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_12__state == 2'b01) begin
        if(PEG_Xvec_12__ap_ready) begin
          if(PEG_Xvec_12__ap_done) begin
            PEG_Xvec_12__state <= 2'b10;
          end else begin
            PEG_Xvec_12__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_12__state == 2'b11) begin
        if(PEG_Xvec_12__ap_done) begin
          PEG_Xvec_12__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_12__state == 2'b10) begin
        if(PEG_Xvec_12__ap_done_global__q0) begin
          PEG_Xvec_12__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_12__ap_start = (PEG_Xvec_12__state == 2'b01);
  assign PEG_Xvec_13__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_13__is_done__q0 = (PEG_Xvec_13__state == 2'b10);
  assign PEG_Xvec_13__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_13__state <= 2'b00;
    end else begin
      if(PEG_Xvec_13__state == 2'b00) begin
        if(PEG_Xvec_13__ap_start_global__q0) begin
          PEG_Xvec_13__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_13__state == 2'b01) begin
        if(PEG_Xvec_13__ap_ready) begin
          if(PEG_Xvec_13__ap_done) begin
            PEG_Xvec_13__state <= 2'b10;
          end else begin
            PEG_Xvec_13__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_13__state == 2'b11) begin
        if(PEG_Xvec_13__ap_done) begin
          PEG_Xvec_13__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_13__state == 2'b10) begin
        if(PEG_Xvec_13__ap_done_global__q0) begin
          PEG_Xvec_13__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_13__ap_start = (PEG_Xvec_13__state == 2'b01);
  assign PEG_Xvec_14__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_14__is_done__q0 = (PEG_Xvec_14__state == 2'b10);
  assign PEG_Xvec_14__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_14__state <= 2'b00;
    end else begin
      if(PEG_Xvec_14__state == 2'b00) begin
        if(PEG_Xvec_14__ap_start_global__q0) begin
          PEG_Xvec_14__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_14__state == 2'b01) begin
        if(PEG_Xvec_14__ap_ready) begin
          if(PEG_Xvec_14__ap_done) begin
            PEG_Xvec_14__state <= 2'b10;
          end else begin
            PEG_Xvec_14__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_14__state == 2'b11) begin
        if(PEG_Xvec_14__ap_done) begin
          PEG_Xvec_14__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_14__state == 2'b10) begin
        if(PEG_Xvec_14__ap_done_global__q0) begin
          PEG_Xvec_14__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_14__ap_start = (PEG_Xvec_14__state == 2'b01);
  assign PEG_Xvec_15__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_15__is_done__q0 = (PEG_Xvec_15__state == 2'b10);
  assign PEG_Xvec_15__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_15__state <= 2'b00;
    end else begin
      if(PEG_Xvec_15__state == 2'b00) begin
        if(PEG_Xvec_15__ap_start_global__q0) begin
          PEG_Xvec_15__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_15__state == 2'b01) begin
        if(PEG_Xvec_15__ap_ready) begin
          if(PEG_Xvec_15__ap_done) begin
            PEG_Xvec_15__state <= 2'b10;
          end else begin
            PEG_Xvec_15__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_15__state == 2'b11) begin
        if(PEG_Xvec_15__ap_done) begin
          PEG_Xvec_15__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_15__state == 2'b10) begin
        if(PEG_Xvec_15__ap_done_global__q0) begin
          PEG_Xvec_15__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_15__ap_start = (PEG_Xvec_15__state == 2'b01);
  assign PEG_Xvec_16__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_16__is_done__q0 = (PEG_Xvec_16__state == 2'b10);
  assign PEG_Xvec_16__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_16__state <= 2'b00;
    end else begin
      if(PEG_Xvec_16__state == 2'b00) begin
        if(PEG_Xvec_16__ap_start_global__q0) begin
          PEG_Xvec_16__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_16__state == 2'b01) begin
        if(PEG_Xvec_16__ap_ready) begin
          if(PEG_Xvec_16__ap_done) begin
            PEG_Xvec_16__state <= 2'b10;
          end else begin
            PEG_Xvec_16__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_16__state == 2'b11) begin
        if(PEG_Xvec_16__ap_done) begin
          PEG_Xvec_16__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_16__state == 2'b10) begin
        if(PEG_Xvec_16__ap_done_global__q0) begin
          PEG_Xvec_16__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_16__ap_start = (PEG_Xvec_16__state == 2'b01);
  assign PEG_Xvec_17__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_17__is_done__q0 = (PEG_Xvec_17__state == 2'b10);
  assign PEG_Xvec_17__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_17__state <= 2'b00;
    end else begin
      if(PEG_Xvec_17__state == 2'b00) begin
        if(PEG_Xvec_17__ap_start_global__q0) begin
          PEG_Xvec_17__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_17__state == 2'b01) begin
        if(PEG_Xvec_17__ap_ready) begin
          if(PEG_Xvec_17__ap_done) begin
            PEG_Xvec_17__state <= 2'b10;
          end else begin
            PEG_Xvec_17__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_17__state == 2'b11) begin
        if(PEG_Xvec_17__ap_done) begin
          PEG_Xvec_17__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_17__state == 2'b10) begin
        if(PEG_Xvec_17__ap_done_global__q0) begin
          PEG_Xvec_17__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_17__ap_start = (PEG_Xvec_17__state == 2'b01);
  assign PEG_Xvec_18__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_18__is_done__q0 = (PEG_Xvec_18__state == 2'b10);
  assign PEG_Xvec_18__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_18__state <= 2'b00;
    end else begin
      if(PEG_Xvec_18__state == 2'b00) begin
        if(PEG_Xvec_18__ap_start_global__q0) begin
          PEG_Xvec_18__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_18__state == 2'b01) begin
        if(PEG_Xvec_18__ap_ready) begin
          if(PEG_Xvec_18__ap_done) begin
            PEG_Xvec_18__state <= 2'b10;
          end else begin
            PEG_Xvec_18__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_18__state == 2'b11) begin
        if(PEG_Xvec_18__ap_done) begin
          PEG_Xvec_18__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_18__state == 2'b10) begin
        if(PEG_Xvec_18__ap_done_global__q0) begin
          PEG_Xvec_18__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_18__ap_start = (PEG_Xvec_18__state == 2'b01);
  assign PEG_Xvec_19__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_19__is_done__q0 = (PEG_Xvec_19__state == 2'b10);
  assign PEG_Xvec_19__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_19__state <= 2'b00;
    end else begin
      if(PEG_Xvec_19__state == 2'b00) begin
        if(PEG_Xvec_19__ap_start_global__q0) begin
          PEG_Xvec_19__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_19__state == 2'b01) begin
        if(PEG_Xvec_19__ap_ready) begin
          if(PEG_Xvec_19__ap_done) begin
            PEG_Xvec_19__state <= 2'b10;
          end else begin
            PEG_Xvec_19__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_19__state == 2'b11) begin
        if(PEG_Xvec_19__ap_done) begin
          PEG_Xvec_19__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_19__state == 2'b10) begin
        if(PEG_Xvec_19__ap_done_global__q0) begin
          PEG_Xvec_19__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_19__ap_start = (PEG_Xvec_19__state == 2'b01);
  assign PEG_Xvec_20__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_20__is_done__q0 = (PEG_Xvec_20__state == 2'b10);
  assign PEG_Xvec_20__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_20__state <= 2'b00;
    end else begin
      if(PEG_Xvec_20__state == 2'b00) begin
        if(PEG_Xvec_20__ap_start_global__q0) begin
          PEG_Xvec_20__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_20__state == 2'b01) begin
        if(PEG_Xvec_20__ap_ready) begin
          if(PEG_Xvec_20__ap_done) begin
            PEG_Xvec_20__state <= 2'b10;
          end else begin
            PEG_Xvec_20__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_20__state == 2'b11) begin
        if(PEG_Xvec_20__ap_done) begin
          PEG_Xvec_20__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_20__state == 2'b10) begin
        if(PEG_Xvec_20__ap_done_global__q0) begin
          PEG_Xvec_20__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_20__ap_start = (PEG_Xvec_20__state == 2'b01);
  assign PEG_Xvec_21__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_21__is_done__q0 = (PEG_Xvec_21__state == 2'b10);
  assign PEG_Xvec_21__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_21__state <= 2'b00;
    end else begin
      if(PEG_Xvec_21__state == 2'b00) begin
        if(PEG_Xvec_21__ap_start_global__q0) begin
          PEG_Xvec_21__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_21__state == 2'b01) begin
        if(PEG_Xvec_21__ap_ready) begin
          if(PEG_Xvec_21__ap_done) begin
            PEG_Xvec_21__state <= 2'b10;
          end else begin
            PEG_Xvec_21__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_21__state == 2'b11) begin
        if(PEG_Xvec_21__ap_done) begin
          PEG_Xvec_21__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_21__state == 2'b10) begin
        if(PEG_Xvec_21__ap_done_global__q0) begin
          PEG_Xvec_21__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_21__ap_start = (PEG_Xvec_21__state == 2'b01);
  assign PEG_Xvec_22__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_22__is_done__q0 = (PEG_Xvec_22__state == 2'b10);
  assign PEG_Xvec_22__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_22__state <= 2'b00;
    end else begin
      if(PEG_Xvec_22__state == 2'b00) begin
        if(PEG_Xvec_22__ap_start_global__q0) begin
          PEG_Xvec_22__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_22__state == 2'b01) begin
        if(PEG_Xvec_22__ap_ready) begin
          if(PEG_Xvec_22__ap_done) begin
            PEG_Xvec_22__state <= 2'b10;
          end else begin
            PEG_Xvec_22__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_22__state == 2'b11) begin
        if(PEG_Xvec_22__ap_done) begin
          PEG_Xvec_22__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_22__state == 2'b10) begin
        if(PEG_Xvec_22__ap_done_global__q0) begin
          PEG_Xvec_22__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_22__ap_start = (PEG_Xvec_22__state == 2'b01);
  assign PEG_Xvec_23__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_23__is_done__q0 = (PEG_Xvec_23__state == 2'b10);
  assign PEG_Xvec_23__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_23__state <= 2'b00;
    end else begin
      if(PEG_Xvec_23__state == 2'b00) begin
        if(PEG_Xvec_23__ap_start_global__q0) begin
          PEG_Xvec_23__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_23__state == 2'b01) begin
        if(PEG_Xvec_23__ap_ready) begin
          if(PEG_Xvec_23__ap_done) begin
            PEG_Xvec_23__state <= 2'b10;
          end else begin
            PEG_Xvec_23__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_23__state == 2'b11) begin
        if(PEG_Xvec_23__ap_done) begin
          PEG_Xvec_23__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_23__state == 2'b10) begin
        if(PEG_Xvec_23__ap_done_global__q0) begin
          PEG_Xvec_23__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_23__ap_start = (PEG_Xvec_23__state == 2'b01);
  assign PEG_Xvec_24__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_24__is_done__q0 = (PEG_Xvec_24__state == 2'b10);
  assign PEG_Xvec_24__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_24__state <= 2'b00;
    end else begin
      if(PEG_Xvec_24__state == 2'b00) begin
        if(PEG_Xvec_24__ap_start_global__q0) begin
          PEG_Xvec_24__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_24__state == 2'b01) begin
        if(PEG_Xvec_24__ap_ready) begin
          if(PEG_Xvec_24__ap_done) begin
            PEG_Xvec_24__state <= 2'b10;
          end else begin
            PEG_Xvec_24__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_24__state == 2'b11) begin
        if(PEG_Xvec_24__ap_done) begin
          PEG_Xvec_24__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_24__state == 2'b10) begin
        if(PEG_Xvec_24__ap_done_global__q0) begin
          PEG_Xvec_24__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_24__ap_start = (PEG_Xvec_24__state == 2'b01);
  assign PEG_Xvec_25__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_25__is_done__q0 = (PEG_Xvec_25__state == 2'b10);
  assign PEG_Xvec_25__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_25__state <= 2'b00;
    end else begin
      if(PEG_Xvec_25__state == 2'b00) begin
        if(PEG_Xvec_25__ap_start_global__q0) begin
          PEG_Xvec_25__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_25__state == 2'b01) begin
        if(PEG_Xvec_25__ap_ready) begin
          if(PEG_Xvec_25__ap_done) begin
            PEG_Xvec_25__state <= 2'b10;
          end else begin
            PEG_Xvec_25__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_25__state == 2'b11) begin
        if(PEG_Xvec_25__ap_done) begin
          PEG_Xvec_25__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_25__state == 2'b10) begin
        if(PEG_Xvec_25__ap_done_global__q0) begin
          PEG_Xvec_25__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_25__ap_start = (PEG_Xvec_25__state == 2'b01);
  assign PEG_Xvec_26__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_26__is_done__q0 = (PEG_Xvec_26__state == 2'b10);
  assign PEG_Xvec_26__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_26__state <= 2'b00;
    end else begin
      if(PEG_Xvec_26__state == 2'b00) begin
        if(PEG_Xvec_26__ap_start_global__q0) begin
          PEG_Xvec_26__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_26__state == 2'b01) begin
        if(PEG_Xvec_26__ap_ready) begin
          if(PEG_Xvec_26__ap_done) begin
            PEG_Xvec_26__state <= 2'b10;
          end else begin
            PEG_Xvec_26__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_26__state == 2'b11) begin
        if(PEG_Xvec_26__ap_done) begin
          PEG_Xvec_26__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_26__state == 2'b10) begin
        if(PEG_Xvec_26__ap_done_global__q0) begin
          PEG_Xvec_26__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_26__ap_start = (PEG_Xvec_26__state == 2'b01);
  assign PEG_Xvec_27__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_27__is_done__q0 = (PEG_Xvec_27__state == 2'b10);
  assign PEG_Xvec_27__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_27__state <= 2'b00;
    end else begin
      if(PEG_Xvec_27__state == 2'b00) begin
        if(PEG_Xvec_27__ap_start_global__q0) begin
          PEG_Xvec_27__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_27__state == 2'b01) begin
        if(PEG_Xvec_27__ap_ready) begin
          if(PEG_Xvec_27__ap_done) begin
            PEG_Xvec_27__state <= 2'b10;
          end else begin
            PEG_Xvec_27__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_27__state == 2'b11) begin
        if(PEG_Xvec_27__ap_done) begin
          PEG_Xvec_27__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_27__state == 2'b10) begin
        if(PEG_Xvec_27__ap_done_global__q0) begin
          PEG_Xvec_27__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_27__ap_start = (PEG_Xvec_27__state == 2'b01);
  assign PEG_Xvec_28__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_28__is_done__q0 = (PEG_Xvec_28__state == 2'b10);
  assign PEG_Xvec_28__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_28__state <= 2'b00;
    end else begin
      if(PEG_Xvec_28__state == 2'b00) begin
        if(PEG_Xvec_28__ap_start_global__q0) begin
          PEG_Xvec_28__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_28__state == 2'b01) begin
        if(PEG_Xvec_28__ap_ready) begin
          if(PEG_Xvec_28__ap_done) begin
            PEG_Xvec_28__state <= 2'b10;
          end else begin
            PEG_Xvec_28__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_28__state == 2'b11) begin
        if(PEG_Xvec_28__ap_done) begin
          PEG_Xvec_28__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_28__state == 2'b10) begin
        if(PEG_Xvec_28__ap_done_global__q0) begin
          PEG_Xvec_28__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_28__ap_start = (PEG_Xvec_28__state == 2'b01);
  assign PEG_Xvec_29__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_29__is_done__q0 = (PEG_Xvec_29__state == 2'b10);
  assign PEG_Xvec_29__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_29__state <= 2'b00;
    end else begin
      if(PEG_Xvec_29__state == 2'b00) begin
        if(PEG_Xvec_29__ap_start_global__q0) begin
          PEG_Xvec_29__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_29__state == 2'b01) begin
        if(PEG_Xvec_29__ap_ready) begin
          if(PEG_Xvec_29__ap_done) begin
            PEG_Xvec_29__state <= 2'b10;
          end else begin
            PEG_Xvec_29__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_29__state == 2'b11) begin
        if(PEG_Xvec_29__ap_done) begin
          PEG_Xvec_29__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_29__state == 2'b10) begin
        if(PEG_Xvec_29__ap_done_global__q0) begin
          PEG_Xvec_29__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_29__ap_start = (PEG_Xvec_29__state == 2'b01);
  assign PEG_Xvec_30__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_30__is_done__q0 = (PEG_Xvec_30__state == 2'b10);
  assign PEG_Xvec_30__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_30__state <= 2'b00;
    end else begin
      if(PEG_Xvec_30__state == 2'b00) begin
        if(PEG_Xvec_30__ap_start_global__q0) begin
          PEG_Xvec_30__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_30__state == 2'b01) begin
        if(PEG_Xvec_30__ap_ready) begin
          if(PEG_Xvec_30__ap_done) begin
            PEG_Xvec_30__state <= 2'b10;
          end else begin
            PEG_Xvec_30__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_30__state == 2'b11) begin
        if(PEG_Xvec_30__ap_done) begin
          PEG_Xvec_30__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_30__state == 2'b10) begin
        if(PEG_Xvec_30__ap_done_global__q0) begin
          PEG_Xvec_30__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_30__ap_start = (PEG_Xvec_30__state == 2'b01);
  assign PEG_Xvec_31__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_31__is_done__q0 = (PEG_Xvec_31__state == 2'b10);
  assign PEG_Xvec_31__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_31__state <= 2'b00;
    end else begin
      if(PEG_Xvec_31__state == 2'b00) begin
        if(PEG_Xvec_31__ap_start_global__q0) begin
          PEG_Xvec_31__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_31__state == 2'b01) begin
        if(PEG_Xvec_31__ap_ready) begin
          if(PEG_Xvec_31__ap_done) begin
            PEG_Xvec_31__state <= 2'b10;
          end else begin
            PEG_Xvec_31__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_31__state == 2'b11) begin
        if(PEG_Xvec_31__ap_done) begin
          PEG_Xvec_31__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_31__state == 2'b10) begin
        if(PEG_Xvec_31__ap_done_global__q0) begin
          PEG_Xvec_31__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_31__ap_start = (PEG_Xvec_31__state == 2'b01);
  assign PEG_Xvec_32__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_32__is_done__q0 = (PEG_Xvec_32__state == 2'b10);
  assign PEG_Xvec_32__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_32__state <= 2'b00;
    end else begin
      if(PEG_Xvec_32__state == 2'b00) begin
        if(PEG_Xvec_32__ap_start_global__q0) begin
          PEG_Xvec_32__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_32__state == 2'b01) begin
        if(PEG_Xvec_32__ap_ready) begin
          if(PEG_Xvec_32__ap_done) begin
            PEG_Xvec_32__state <= 2'b10;
          end else begin
            PEG_Xvec_32__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_32__state == 2'b11) begin
        if(PEG_Xvec_32__ap_done) begin
          PEG_Xvec_32__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_32__state == 2'b10) begin
        if(PEG_Xvec_32__ap_done_global__q0) begin
          PEG_Xvec_32__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_32__ap_start = (PEG_Xvec_32__state == 2'b01);
  assign PEG_Xvec_33__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_33__is_done__q0 = (PEG_Xvec_33__state == 2'b10);
  assign PEG_Xvec_33__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_33__state <= 2'b00;
    end else begin
      if(PEG_Xvec_33__state == 2'b00) begin
        if(PEG_Xvec_33__ap_start_global__q0) begin
          PEG_Xvec_33__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_33__state == 2'b01) begin
        if(PEG_Xvec_33__ap_ready) begin
          if(PEG_Xvec_33__ap_done) begin
            PEG_Xvec_33__state <= 2'b10;
          end else begin
            PEG_Xvec_33__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_33__state == 2'b11) begin
        if(PEG_Xvec_33__ap_done) begin
          PEG_Xvec_33__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_33__state == 2'b10) begin
        if(PEG_Xvec_33__ap_done_global__q0) begin
          PEG_Xvec_33__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_33__ap_start = (PEG_Xvec_33__state == 2'b01);
  assign PEG_Xvec_34__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_34__is_done__q0 = (PEG_Xvec_34__state == 2'b10);
  assign PEG_Xvec_34__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_34__state <= 2'b00;
    end else begin
      if(PEG_Xvec_34__state == 2'b00) begin
        if(PEG_Xvec_34__ap_start_global__q0) begin
          PEG_Xvec_34__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_34__state == 2'b01) begin
        if(PEG_Xvec_34__ap_ready) begin
          if(PEG_Xvec_34__ap_done) begin
            PEG_Xvec_34__state <= 2'b10;
          end else begin
            PEG_Xvec_34__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_34__state == 2'b11) begin
        if(PEG_Xvec_34__ap_done) begin
          PEG_Xvec_34__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_34__state == 2'b10) begin
        if(PEG_Xvec_34__ap_done_global__q0) begin
          PEG_Xvec_34__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_34__ap_start = (PEG_Xvec_34__state == 2'b01);
  assign PEG_Xvec_35__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_35__is_done__q0 = (PEG_Xvec_35__state == 2'b10);
  assign PEG_Xvec_35__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_35__state <= 2'b00;
    end else begin
      if(PEG_Xvec_35__state == 2'b00) begin
        if(PEG_Xvec_35__ap_start_global__q0) begin
          PEG_Xvec_35__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_35__state == 2'b01) begin
        if(PEG_Xvec_35__ap_ready) begin
          if(PEG_Xvec_35__ap_done) begin
            PEG_Xvec_35__state <= 2'b10;
          end else begin
            PEG_Xvec_35__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_35__state == 2'b11) begin
        if(PEG_Xvec_35__ap_done) begin
          PEG_Xvec_35__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_35__state == 2'b10) begin
        if(PEG_Xvec_35__ap_done_global__q0) begin
          PEG_Xvec_35__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_35__ap_start = (PEG_Xvec_35__state == 2'b01);
  assign PEG_Xvec_36__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_36__is_done__q0 = (PEG_Xvec_36__state == 2'b10);
  assign PEG_Xvec_36__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_36__state <= 2'b00;
    end else begin
      if(PEG_Xvec_36__state == 2'b00) begin
        if(PEG_Xvec_36__ap_start_global__q0) begin
          PEG_Xvec_36__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_36__state == 2'b01) begin
        if(PEG_Xvec_36__ap_ready) begin
          if(PEG_Xvec_36__ap_done) begin
            PEG_Xvec_36__state <= 2'b10;
          end else begin
            PEG_Xvec_36__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_36__state == 2'b11) begin
        if(PEG_Xvec_36__ap_done) begin
          PEG_Xvec_36__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_36__state == 2'b10) begin
        if(PEG_Xvec_36__ap_done_global__q0) begin
          PEG_Xvec_36__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_36__ap_start = (PEG_Xvec_36__state == 2'b01);
  assign PEG_Xvec_37__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_37__is_done__q0 = (PEG_Xvec_37__state == 2'b10);
  assign PEG_Xvec_37__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_37__state <= 2'b00;
    end else begin
      if(PEG_Xvec_37__state == 2'b00) begin
        if(PEG_Xvec_37__ap_start_global__q0) begin
          PEG_Xvec_37__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_37__state == 2'b01) begin
        if(PEG_Xvec_37__ap_ready) begin
          if(PEG_Xvec_37__ap_done) begin
            PEG_Xvec_37__state <= 2'b10;
          end else begin
            PEG_Xvec_37__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_37__state == 2'b11) begin
        if(PEG_Xvec_37__ap_done) begin
          PEG_Xvec_37__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_37__state == 2'b10) begin
        if(PEG_Xvec_37__ap_done_global__q0) begin
          PEG_Xvec_37__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_37__ap_start = (PEG_Xvec_37__state == 2'b01);
  assign PEG_Xvec_38__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_38__is_done__q0 = (PEG_Xvec_38__state == 2'b10);
  assign PEG_Xvec_38__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_38__state <= 2'b00;
    end else begin
      if(PEG_Xvec_38__state == 2'b00) begin
        if(PEG_Xvec_38__ap_start_global__q0) begin
          PEG_Xvec_38__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_38__state == 2'b01) begin
        if(PEG_Xvec_38__ap_ready) begin
          if(PEG_Xvec_38__ap_done) begin
            PEG_Xvec_38__state <= 2'b10;
          end else begin
            PEG_Xvec_38__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_38__state == 2'b11) begin
        if(PEG_Xvec_38__ap_done) begin
          PEG_Xvec_38__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_38__state == 2'b10) begin
        if(PEG_Xvec_38__ap_done_global__q0) begin
          PEG_Xvec_38__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_38__ap_start = (PEG_Xvec_38__state == 2'b01);
  assign PEG_Xvec_39__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_39__is_done__q0 = (PEG_Xvec_39__state == 2'b10);
  assign PEG_Xvec_39__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_39__state <= 2'b00;
    end else begin
      if(PEG_Xvec_39__state == 2'b00) begin
        if(PEG_Xvec_39__ap_start_global__q0) begin
          PEG_Xvec_39__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_39__state == 2'b01) begin
        if(PEG_Xvec_39__ap_ready) begin
          if(PEG_Xvec_39__ap_done) begin
            PEG_Xvec_39__state <= 2'b10;
          end else begin
            PEG_Xvec_39__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_39__state == 2'b11) begin
        if(PEG_Xvec_39__ap_done) begin
          PEG_Xvec_39__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_39__state == 2'b10) begin
        if(PEG_Xvec_39__ap_done_global__q0) begin
          PEG_Xvec_39__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_39__ap_start = (PEG_Xvec_39__state == 2'b01);
  assign PEG_Xvec_40__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_40__is_done__q0 = (PEG_Xvec_40__state == 2'b10);
  assign PEG_Xvec_40__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_40__state <= 2'b00;
    end else begin
      if(PEG_Xvec_40__state == 2'b00) begin
        if(PEG_Xvec_40__ap_start_global__q0) begin
          PEG_Xvec_40__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_40__state == 2'b01) begin
        if(PEG_Xvec_40__ap_ready) begin
          if(PEG_Xvec_40__ap_done) begin
            PEG_Xvec_40__state <= 2'b10;
          end else begin
            PEG_Xvec_40__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_40__state == 2'b11) begin
        if(PEG_Xvec_40__ap_done) begin
          PEG_Xvec_40__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_40__state == 2'b10) begin
        if(PEG_Xvec_40__ap_done_global__q0) begin
          PEG_Xvec_40__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_40__ap_start = (PEG_Xvec_40__state == 2'b01);
  assign PEG_Xvec_41__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_41__is_done__q0 = (PEG_Xvec_41__state == 2'b10);
  assign PEG_Xvec_41__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_41__state <= 2'b00;
    end else begin
      if(PEG_Xvec_41__state == 2'b00) begin
        if(PEG_Xvec_41__ap_start_global__q0) begin
          PEG_Xvec_41__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_41__state == 2'b01) begin
        if(PEG_Xvec_41__ap_ready) begin
          if(PEG_Xvec_41__ap_done) begin
            PEG_Xvec_41__state <= 2'b10;
          end else begin
            PEG_Xvec_41__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_41__state == 2'b11) begin
        if(PEG_Xvec_41__ap_done) begin
          PEG_Xvec_41__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_41__state == 2'b10) begin
        if(PEG_Xvec_41__ap_done_global__q0) begin
          PEG_Xvec_41__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_41__ap_start = (PEG_Xvec_41__state == 2'b01);
  assign PEG_Xvec_42__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_42__is_done__q0 = (PEG_Xvec_42__state == 2'b10);
  assign PEG_Xvec_42__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_42__state <= 2'b00;
    end else begin
      if(PEG_Xvec_42__state == 2'b00) begin
        if(PEG_Xvec_42__ap_start_global__q0) begin
          PEG_Xvec_42__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_42__state == 2'b01) begin
        if(PEG_Xvec_42__ap_ready) begin
          if(PEG_Xvec_42__ap_done) begin
            PEG_Xvec_42__state <= 2'b10;
          end else begin
            PEG_Xvec_42__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_42__state == 2'b11) begin
        if(PEG_Xvec_42__ap_done) begin
          PEG_Xvec_42__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_42__state == 2'b10) begin
        if(PEG_Xvec_42__ap_done_global__q0) begin
          PEG_Xvec_42__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_42__ap_start = (PEG_Xvec_42__state == 2'b01);
  assign PEG_Xvec_43__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_43__is_done__q0 = (PEG_Xvec_43__state == 2'b10);
  assign PEG_Xvec_43__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_43__state <= 2'b00;
    end else begin
      if(PEG_Xvec_43__state == 2'b00) begin
        if(PEG_Xvec_43__ap_start_global__q0) begin
          PEG_Xvec_43__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_43__state == 2'b01) begin
        if(PEG_Xvec_43__ap_ready) begin
          if(PEG_Xvec_43__ap_done) begin
            PEG_Xvec_43__state <= 2'b10;
          end else begin
            PEG_Xvec_43__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_43__state == 2'b11) begin
        if(PEG_Xvec_43__ap_done) begin
          PEG_Xvec_43__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_43__state == 2'b10) begin
        if(PEG_Xvec_43__ap_done_global__q0) begin
          PEG_Xvec_43__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_43__ap_start = (PEG_Xvec_43__state == 2'b01);
  assign PEG_Xvec_44__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_44__is_done__q0 = (PEG_Xvec_44__state == 2'b10);
  assign PEG_Xvec_44__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_44__state <= 2'b00;
    end else begin
      if(PEG_Xvec_44__state == 2'b00) begin
        if(PEG_Xvec_44__ap_start_global__q0) begin
          PEG_Xvec_44__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_44__state == 2'b01) begin
        if(PEG_Xvec_44__ap_ready) begin
          if(PEG_Xvec_44__ap_done) begin
            PEG_Xvec_44__state <= 2'b10;
          end else begin
            PEG_Xvec_44__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_44__state == 2'b11) begin
        if(PEG_Xvec_44__ap_done) begin
          PEG_Xvec_44__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_44__state == 2'b10) begin
        if(PEG_Xvec_44__ap_done_global__q0) begin
          PEG_Xvec_44__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_44__ap_start = (PEG_Xvec_44__state == 2'b01);
  assign PEG_Xvec_45__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_45__is_done__q0 = (PEG_Xvec_45__state == 2'b10);
  assign PEG_Xvec_45__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_45__state <= 2'b00;
    end else begin
      if(PEG_Xvec_45__state == 2'b00) begin
        if(PEG_Xvec_45__ap_start_global__q0) begin
          PEG_Xvec_45__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_45__state == 2'b01) begin
        if(PEG_Xvec_45__ap_ready) begin
          if(PEG_Xvec_45__ap_done) begin
            PEG_Xvec_45__state <= 2'b10;
          end else begin
            PEG_Xvec_45__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_45__state == 2'b11) begin
        if(PEG_Xvec_45__ap_done) begin
          PEG_Xvec_45__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_45__state == 2'b10) begin
        if(PEG_Xvec_45__ap_done_global__q0) begin
          PEG_Xvec_45__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_45__ap_start = (PEG_Xvec_45__state == 2'b01);
  assign PEG_Xvec_46__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_46__is_done__q0 = (PEG_Xvec_46__state == 2'b10);
  assign PEG_Xvec_46__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_46__state <= 2'b00;
    end else begin
      if(PEG_Xvec_46__state == 2'b00) begin
        if(PEG_Xvec_46__ap_start_global__q0) begin
          PEG_Xvec_46__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_46__state == 2'b01) begin
        if(PEG_Xvec_46__ap_ready) begin
          if(PEG_Xvec_46__ap_done) begin
            PEG_Xvec_46__state <= 2'b10;
          end else begin
            PEG_Xvec_46__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_46__state == 2'b11) begin
        if(PEG_Xvec_46__ap_done) begin
          PEG_Xvec_46__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_46__state == 2'b10) begin
        if(PEG_Xvec_46__ap_done_global__q0) begin
          PEG_Xvec_46__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_46__ap_start = (PEG_Xvec_46__state == 2'b01);
  assign PEG_Xvec_47__ap_start_global__q0 = ap_start__q0;
  assign PEG_Xvec_47__is_done__q0 = (PEG_Xvec_47__state == 2'b10);
  assign PEG_Xvec_47__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Xvec_47__state <= 2'b00;
    end else begin
      if(PEG_Xvec_47__state == 2'b00) begin
        if(PEG_Xvec_47__ap_start_global__q0) begin
          PEG_Xvec_47__state <= 2'b01;
        end 
      end 
      if(PEG_Xvec_47__state == 2'b01) begin
        if(PEG_Xvec_47__ap_ready) begin
          if(PEG_Xvec_47__ap_done) begin
            PEG_Xvec_47__state <= 2'b10;
          end else begin
            PEG_Xvec_47__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Xvec_47__state == 2'b11) begin
        if(PEG_Xvec_47__ap_done) begin
          PEG_Xvec_47__state <= 2'b10;
        end 
      end 
      if(PEG_Xvec_47__state == 2'b10) begin
        if(PEG_Xvec_47__ap_done_global__q0) begin
          PEG_Xvec_47__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Xvec_47__ap_start = (PEG_Xvec_47__state == 2'b01);
  assign PEG_Yvec_0__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_0__is_done__q0 = (PEG_Yvec_0__state == 2'b10);
  assign PEG_Yvec_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_0__state <= 2'b00;
    end else begin
      if(PEG_Yvec_0__state == 2'b00) begin
        if(PEG_Yvec_0__ap_start_global__q0) begin
          PEG_Yvec_0__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_0__state == 2'b01) begin
        if(PEG_Yvec_0__ap_ready) begin
          if(PEG_Yvec_0__ap_done) begin
            PEG_Yvec_0__state <= 2'b10;
          end else begin
            PEG_Yvec_0__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_0__state == 2'b11) begin
        if(PEG_Yvec_0__ap_done) begin
          PEG_Yvec_0__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_0__state == 2'b10) begin
        if(PEG_Yvec_0__ap_done_global__q0) begin
          PEG_Yvec_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_0__ap_start = (PEG_Yvec_0__state == 2'b01);
  assign PEG_Yvec_1__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_1__is_done__q0 = (PEG_Yvec_1__state == 2'b10);
  assign PEG_Yvec_1__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_1__state <= 2'b00;
    end else begin
      if(PEG_Yvec_1__state == 2'b00) begin
        if(PEG_Yvec_1__ap_start_global__q0) begin
          PEG_Yvec_1__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_1__state == 2'b01) begin
        if(PEG_Yvec_1__ap_ready) begin
          if(PEG_Yvec_1__ap_done) begin
            PEG_Yvec_1__state <= 2'b10;
          end else begin
            PEG_Yvec_1__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_1__state == 2'b11) begin
        if(PEG_Yvec_1__ap_done) begin
          PEG_Yvec_1__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_1__state == 2'b10) begin
        if(PEG_Yvec_1__ap_done_global__q0) begin
          PEG_Yvec_1__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_1__ap_start = (PEG_Yvec_1__state == 2'b01);
  assign PEG_Yvec_2__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_2__is_done__q0 = (PEG_Yvec_2__state == 2'b10);
  assign PEG_Yvec_2__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_2__state <= 2'b00;
    end else begin
      if(PEG_Yvec_2__state == 2'b00) begin
        if(PEG_Yvec_2__ap_start_global__q0) begin
          PEG_Yvec_2__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_2__state == 2'b01) begin
        if(PEG_Yvec_2__ap_ready) begin
          if(PEG_Yvec_2__ap_done) begin
            PEG_Yvec_2__state <= 2'b10;
          end else begin
            PEG_Yvec_2__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_2__state == 2'b11) begin
        if(PEG_Yvec_2__ap_done) begin
          PEG_Yvec_2__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_2__state == 2'b10) begin
        if(PEG_Yvec_2__ap_done_global__q0) begin
          PEG_Yvec_2__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_2__ap_start = (PEG_Yvec_2__state == 2'b01);
  assign PEG_Yvec_3__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_3__is_done__q0 = (PEG_Yvec_3__state == 2'b10);
  assign PEG_Yvec_3__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_3__state <= 2'b00;
    end else begin
      if(PEG_Yvec_3__state == 2'b00) begin
        if(PEG_Yvec_3__ap_start_global__q0) begin
          PEG_Yvec_3__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_3__state == 2'b01) begin
        if(PEG_Yvec_3__ap_ready) begin
          if(PEG_Yvec_3__ap_done) begin
            PEG_Yvec_3__state <= 2'b10;
          end else begin
            PEG_Yvec_3__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_3__state == 2'b11) begin
        if(PEG_Yvec_3__ap_done) begin
          PEG_Yvec_3__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_3__state == 2'b10) begin
        if(PEG_Yvec_3__ap_done_global__q0) begin
          PEG_Yvec_3__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_3__ap_start = (PEG_Yvec_3__state == 2'b01);
  assign PEG_Yvec_4__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_4__is_done__q0 = (PEG_Yvec_4__state == 2'b10);
  assign PEG_Yvec_4__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_4__state <= 2'b00;
    end else begin
      if(PEG_Yvec_4__state == 2'b00) begin
        if(PEG_Yvec_4__ap_start_global__q0) begin
          PEG_Yvec_4__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_4__state == 2'b01) begin
        if(PEG_Yvec_4__ap_ready) begin
          if(PEG_Yvec_4__ap_done) begin
            PEG_Yvec_4__state <= 2'b10;
          end else begin
            PEG_Yvec_4__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_4__state == 2'b11) begin
        if(PEG_Yvec_4__ap_done) begin
          PEG_Yvec_4__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_4__state == 2'b10) begin
        if(PEG_Yvec_4__ap_done_global__q0) begin
          PEG_Yvec_4__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_4__ap_start = (PEG_Yvec_4__state == 2'b01);
  assign PEG_Yvec_5__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_5__is_done__q0 = (PEG_Yvec_5__state == 2'b10);
  assign PEG_Yvec_5__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_5__state <= 2'b00;
    end else begin
      if(PEG_Yvec_5__state == 2'b00) begin
        if(PEG_Yvec_5__ap_start_global__q0) begin
          PEG_Yvec_5__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_5__state == 2'b01) begin
        if(PEG_Yvec_5__ap_ready) begin
          if(PEG_Yvec_5__ap_done) begin
            PEG_Yvec_5__state <= 2'b10;
          end else begin
            PEG_Yvec_5__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_5__state == 2'b11) begin
        if(PEG_Yvec_5__ap_done) begin
          PEG_Yvec_5__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_5__state == 2'b10) begin
        if(PEG_Yvec_5__ap_done_global__q0) begin
          PEG_Yvec_5__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_5__ap_start = (PEG_Yvec_5__state == 2'b01);
  assign PEG_Yvec_6__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_6__is_done__q0 = (PEG_Yvec_6__state == 2'b10);
  assign PEG_Yvec_6__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_6__state <= 2'b00;
    end else begin
      if(PEG_Yvec_6__state == 2'b00) begin
        if(PEG_Yvec_6__ap_start_global__q0) begin
          PEG_Yvec_6__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_6__state == 2'b01) begin
        if(PEG_Yvec_6__ap_ready) begin
          if(PEG_Yvec_6__ap_done) begin
            PEG_Yvec_6__state <= 2'b10;
          end else begin
            PEG_Yvec_6__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_6__state == 2'b11) begin
        if(PEG_Yvec_6__ap_done) begin
          PEG_Yvec_6__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_6__state == 2'b10) begin
        if(PEG_Yvec_6__ap_done_global__q0) begin
          PEG_Yvec_6__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_6__ap_start = (PEG_Yvec_6__state == 2'b01);
  assign PEG_Yvec_7__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_7__is_done__q0 = (PEG_Yvec_7__state == 2'b10);
  assign PEG_Yvec_7__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_7__state <= 2'b00;
    end else begin
      if(PEG_Yvec_7__state == 2'b00) begin
        if(PEG_Yvec_7__ap_start_global__q0) begin
          PEG_Yvec_7__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_7__state == 2'b01) begin
        if(PEG_Yvec_7__ap_ready) begin
          if(PEG_Yvec_7__ap_done) begin
            PEG_Yvec_7__state <= 2'b10;
          end else begin
            PEG_Yvec_7__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_7__state == 2'b11) begin
        if(PEG_Yvec_7__ap_done) begin
          PEG_Yvec_7__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_7__state == 2'b10) begin
        if(PEG_Yvec_7__ap_done_global__q0) begin
          PEG_Yvec_7__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_7__ap_start = (PEG_Yvec_7__state == 2'b01);
  assign PEG_Yvec_8__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_8__is_done__q0 = (PEG_Yvec_8__state == 2'b10);
  assign PEG_Yvec_8__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_8__state <= 2'b00;
    end else begin
      if(PEG_Yvec_8__state == 2'b00) begin
        if(PEG_Yvec_8__ap_start_global__q0) begin
          PEG_Yvec_8__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_8__state == 2'b01) begin
        if(PEG_Yvec_8__ap_ready) begin
          if(PEG_Yvec_8__ap_done) begin
            PEG_Yvec_8__state <= 2'b10;
          end else begin
            PEG_Yvec_8__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_8__state == 2'b11) begin
        if(PEG_Yvec_8__ap_done) begin
          PEG_Yvec_8__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_8__state == 2'b10) begin
        if(PEG_Yvec_8__ap_done_global__q0) begin
          PEG_Yvec_8__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_8__ap_start = (PEG_Yvec_8__state == 2'b01);
  assign PEG_Yvec_9__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_9__is_done__q0 = (PEG_Yvec_9__state == 2'b10);
  assign PEG_Yvec_9__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_9__state <= 2'b00;
    end else begin
      if(PEG_Yvec_9__state == 2'b00) begin
        if(PEG_Yvec_9__ap_start_global__q0) begin
          PEG_Yvec_9__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_9__state == 2'b01) begin
        if(PEG_Yvec_9__ap_ready) begin
          if(PEG_Yvec_9__ap_done) begin
            PEG_Yvec_9__state <= 2'b10;
          end else begin
            PEG_Yvec_9__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_9__state == 2'b11) begin
        if(PEG_Yvec_9__ap_done) begin
          PEG_Yvec_9__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_9__state == 2'b10) begin
        if(PEG_Yvec_9__ap_done_global__q0) begin
          PEG_Yvec_9__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_9__ap_start = (PEG_Yvec_9__state == 2'b01);
  assign PEG_Yvec_10__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_10__is_done__q0 = (PEG_Yvec_10__state == 2'b10);
  assign PEG_Yvec_10__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_10__state <= 2'b00;
    end else begin
      if(PEG_Yvec_10__state == 2'b00) begin
        if(PEG_Yvec_10__ap_start_global__q0) begin
          PEG_Yvec_10__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_10__state == 2'b01) begin
        if(PEG_Yvec_10__ap_ready) begin
          if(PEG_Yvec_10__ap_done) begin
            PEG_Yvec_10__state <= 2'b10;
          end else begin
            PEG_Yvec_10__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_10__state == 2'b11) begin
        if(PEG_Yvec_10__ap_done) begin
          PEG_Yvec_10__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_10__state == 2'b10) begin
        if(PEG_Yvec_10__ap_done_global__q0) begin
          PEG_Yvec_10__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_10__ap_start = (PEG_Yvec_10__state == 2'b01);
  assign PEG_Yvec_11__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_11__is_done__q0 = (PEG_Yvec_11__state == 2'b10);
  assign PEG_Yvec_11__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_11__state <= 2'b00;
    end else begin
      if(PEG_Yvec_11__state == 2'b00) begin
        if(PEG_Yvec_11__ap_start_global__q0) begin
          PEG_Yvec_11__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_11__state == 2'b01) begin
        if(PEG_Yvec_11__ap_ready) begin
          if(PEG_Yvec_11__ap_done) begin
            PEG_Yvec_11__state <= 2'b10;
          end else begin
            PEG_Yvec_11__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_11__state == 2'b11) begin
        if(PEG_Yvec_11__ap_done) begin
          PEG_Yvec_11__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_11__state == 2'b10) begin
        if(PEG_Yvec_11__ap_done_global__q0) begin
          PEG_Yvec_11__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_11__ap_start = (PEG_Yvec_11__state == 2'b01);
  assign PEG_Yvec_12__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_12__is_done__q0 = (PEG_Yvec_12__state == 2'b10);
  assign PEG_Yvec_12__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_12__state <= 2'b00;
    end else begin
      if(PEG_Yvec_12__state == 2'b00) begin
        if(PEG_Yvec_12__ap_start_global__q0) begin
          PEG_Yvec_12__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_12__state == 2'b01) begin
        if(PEG_Yvec_12__ap_ready) begin
          if(PEG_Yvec_12__ap_done) begin
            PEG_Yvec_12__state <= 2'b10;
          end else begin
            PEG_Yvec_12__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_12__state == 2'b11) begin
        if(PEG_Yvec_12__ap_done) begin
          PEG_Yvec_12__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_12__state == 2'b10) begin
        if(PEG_Yvec_12__ap_done_global__q0) begin
          PEG_Yvec_12__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_12__ap_start = (PEG_Yvec_12__state == 2'b01);
  assign PEG_Yvec_13__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_13__is_done__q0 = (PEG_Yvec_13__state == 2'b10);
  assign PEG_Yvec_13__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_13__state <= 2'b00;
    end else begin
      if(PEG_Yvec_13__state == 2'b00) begin
        if(PEG_Yvec_13__ap_start_global__q0) begin
          PEG_Yvec_13__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_13__state == 2'b01) begin
        if(PEG_Yvec_13__ap_ready) begin
          if(PEG_Yvec_13__ap_done) begin
            PEG_Yvec_13__state <= 2'b10;
          end else begin
            PEG_Yvec_13__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_13__state == 2'b11) begin
        if(PEG_Yvec_13__ap_done) begin
          PEG_Yvec_13__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_13__state == 2'b10) begin
        if(PEG_Yvec_13__ap_done_global__q0) begin
          PEG_Yvec_13__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_13__ap_start = (PEG_Yvec_13__state == 2'b01);
  assign PEG_Yvec_14__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_14__is_done__q0 = (PEG_Yvec_14__state == 2'b10);
  assign PEG_Yvec_14__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_14__state <= 2'b00;
    end else begin
      if(PEG_Yvec_14__state == 2'b00) begin
        if(PEG_Yvec_14__ap_start_global__q0) begin
          PEG_Yvec_14__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_14__state == 2'b01) begin
        if(PEG_Yvec_14__ap_ready) begin
          if(PEG_Yvec_14__ap_done) begin
            PEG_Yvec_14__state <= 2'b10;
          end else begin
            PEG_Yvec_14__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_14__state == 2'b11) begin
        if(PEG_Yvec_14__ap_done) begin
          PEG_Yvec_14__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_14__state == 2'b10) begin
        if(PEG_Yvec_14__ap_done_global__q0) begin
          PEG_Yvec_14__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_14__ap_start = (PEG_Yvec_14__state == 2'b01);
  assign PEG_Yvec_15__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_15__is_done__q0 = (PEG_Yvec_15__state == 2'b10);
  assign PEG_Yvec_15__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_15__state <= 2'b00;
    end else begin
      if(PEG_Yvec_15__state == 2'b00) begin
        if(PEG_Yvec_15__ap_start_global__q0) begin
          PEG_Yvec_15__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_15__state == 2'b01) begin
        if(PEG_Yvec_15__ap_ready) begin
          if(PEG_Yvec_15__ap_done) begin
            PEG_Yvec_15__state <= 2'b10;
          end else begin
            PEG_Yvec_15__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_15__state == 2'b11) begin
        if(PEG_Yvec_15__ap_done) begin
          PEG_Yvec_15__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_15__state == 2'b10) begin
        if(PEG_Yvec_15__ap_done_global__q0) begin
          PEG_Yvec_15__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_15__ap_start = (PEG_Yvec_15__state == 2'b01);
  assign PEG_Yvec_16__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_16__is_done__q0 = (PEG_Yvec_16__state == 2'b10);
  assign PEG_Yvec_16__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_16__state <= 2'b00;
    end else begin
      if(PEG_Yvec_16__state == 2'b00) begin
        if(PEG_Yvec_16__ap_start_global__q0) begin
          PEG_Yvec_16__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_16__state == 2'b01) begin
        if(PEG_Yvec_16__ap_ready) begin
          if(PEG_Yvec_16__ap_done) begin
            PEG_Yvec_16__state <= 2'b10;
          end else begin
            PEG_Yvec_16__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_16__state == 2'b11) begin
        if(PEG_Yvec_16__ap_done) begin
          PEG_Yvec_16__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_16__state == 2'b10) begin
        if(PEG_Yvec_16__ap_done_global__q0) begin
          PEG_Yvec_16__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_16__ap_start = (PEG_Yvec_16__state == 2'b01);
  assign PEG_Yvec_17__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_17__is_done__q0 = (PEG_Yvec_17__state == 2'b10);
  assign PEG_Yvec_17__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_17__state <= 2'b00;
    end else begin
      if(PEG_Yvec_17__state == 2'b00) begin
        if(PEG_Yvec_17__ap_start_global__q0) begin
          PEG_Yvec_17__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_17__state == 2'b01) begin
        if(PEG_Yvec_17__ap_ready) begin
          if(PEG_Yvec_17__ap_done) begin
            PEG_Yvec_17__state <= 2'b10;
          end else begin
            PEG_Yvec_17__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_17__state == 2'b11) begin
        if(PEG_Yvec_17__ap_done) begin
          PEG_Yvec_17__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_17__state == 2'b10) begin
        if(PEG_Yvec_17__ap_done_global__q0) begin
          PEG_Yvec_17__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_17__ap_start = (PEG_Yvec_17__state == 2'b01);
  assign PEG_Yvec_18__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_18__is_done__q0 = (PEG_Yvec_18__state == 2'b10);
  assign PEG_Yvec_18__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_18__state <= 2'b00;
    end else begin
      if(PEG_Yvec_18__state == 2'b00) begin
        if(PEG_Yvec_18__ap_start_global__q0) begin
          PEG_Yvec_18__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_18__state == 2'b01) begin
        if(PEG_Yvec_18__ap_ready) begin
          if(PEG_Yvec_18__ap_done) begin
            PEG_Yvec_18__state <= 2'b10;
          end else begin
            PEG_Yvec_18__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_18__state == 2'b11) begin
        if(PEG_Yvec_18__ap_done) begin
          PEG_Yvec_18__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_18__state == 2'b10) begin
        if(PEG_Yvec_18__ap_done_global__q0) begin
          PEG_Yvec_18__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_18__ap_start = (PEG_Yvec_18__state == 2'b01);
  assign PEG_Yvec_19__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_19__is_done__q0 = (PEG_Yvec_19__state == 2'b10);
  assign PEG_Yvec_19__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_19__state <= 2'b00;
    end else begin
      if(PEG_Yvec_19__state == 2'b00) begin
        if(PEG_Yvec_19__ap_start_global__q0) begin
          PEG_Yvec_19__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_19__state == 2'b01) begin
        if(PEG_Yvec_19__ap_ready) begin
          if(PEG_Yvec_19__ap_done) begin
            PEG_Yvec_19__state <= 2'b10;
          end else begin
            PEG_Yvec_19__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_19__state == 2'b11) begin
        if(PEG_Yvec_19__ap_done) begin
          PEG_Yvec_19__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_19__state == 2'b10) begin
        if(PEG_Yvec_19__ap_done_global__q0) begin
          PEG_Yvec_19__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_19__ap_start = (PEG_Yvec_19__state == 2'b01);
  assign PEG_Yvec_20__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_20__is_done__q0 = (PEG_Yvec_20__state == 2'b10);
  assign PEG_Yvec_20__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_20__state <= 2'b00;
    end else begin
      if(PEG_Yvec_20__state == 2'b00) begin
        if(PEG_Yvec_20__ap_start_global__q0) begin
          PEG_Yvec_20__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_20__state == 2'b01) begin
        if(PEG_Yvec_20__ap_ready) begin
          if(PEG_Yvec_20__ap_done) begin
            PEG_Yvec_20__state <= 2'b10;
          end else begin
            PEG_Yvec_20__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_20__state == 2'b11) begin
        if(PEG_Yvec_20__ap_done) begin
          PEG_Yvec_20__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_20__state == 2'b10) begin
        if(PEG_Yvec_20__ap_done_global__q0) begin
          PEG_Yvec_20__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_20__ap_start = (PEG_Yvec_20__state == 2'b01);
  assign PEG_Yvec_21__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_21__is_done__q0 = (PEG_Yvec_21__state == 2'b10);
  assign PEG_Yvec_21__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_21__state <= 2'b00;
    end else begin
      if(PEG_Yvec_21__state == 2'b00) begin
        if(PEG_Yvec_21__ap_start_global__q0) begin
          PEG_Yvec_21__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_21__state == 2'b01) begin
        if(PEG_Yvec_21__ap_ready) begin
          if(PEG_Yvec_21__ap_done) begin
            PEG_Yvec_21__state <= 2'b10;
          end else begin
            PEG_Yvec_21__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_21__state == 2'b11) begin
        if(PEG_Yvec_21__ap_done) begin
          PEG_Yvec_21__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_21__state == 2'b10) begin
        if(PEG_Yvec_21__ap_done_global__q0) begin
          PEG_Yvec_21__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_21__ap_start = (PEG_Yvec_21__state == 2'b01);
  assign PEG_Yvec_22__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_22__is_done__q0 = (PEG_Yvec_22__state == 2'b10);
  assign PEG_Yvec_22__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_22__state <= 2'b00;
    end else begin
      if(PEG_Yvec_22__state == 2'b00) begin
        if(PEG_Yvec_22__ap_start_global__q0) begin
          PEG_Yvec_22__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_22__state == 2'b01) begin
        if(PEG_Yvec_22__ap_ready) begin
          if(PEG_Yvec_22__ap_done) begin
            PEG_Yvec_22__state <= 2'b10;
          end else begin
            PEG_Yvec_22__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_22__state == 2'b11) begin
        if(PEG_Yvec_22__ap_done) begin
          PEG_Yvec_22__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_22__state == 2'b10) begin
        if(PEG_Yvec_22__ap_done_global__q0) begin
          PEG_Yvec_22__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_22__ap_start = (PEG_Yvec_22__state == 2'b01);
  assign PEG_Yvec_23__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_23__is_done__q0 = (PEG_Yvec_23__state == 2'b10);
  assign PEG_Yvec_23__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_23__state <= 2'b00;
    end else begin
      if(PEG_Yvec_23__state == 2'b00) begin
        if(PEG_Yvec_23__ap_start_global__q0) begin
          PEG_Yvec_23__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_23__state == 2'b01) begin
        if(PEG_Yvec_23__ap_ready) begin
          if(PEG_Yvec_23__ap_done) begin
            PEG_Yvec_23__state <= 2'b10;
          end else begin
            PEG_Yvec_23__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_23__state == 2'b11) begin
        if(PEG_Yvec_23__ap_done) begin
          PEG_Yvec_23__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_23__state == 2'b10) begin
        if(PEG_Yvec_23__ap_done_global__q0) begin
          PEG_Yvec_23__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_23__ap_start = (PEG_Yvec_23__state == 2'b01);
  assign PEG_Yvec_24__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_24__is_done__q0 = (PEG_Yvec_24__state == 2'b10);
  assign PEG_Yvec_24__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_24__state <= 2'b00;
    end else begin
      if(PEG_Yvec_24__state == 2'b00) begin
        if(PEG_Yvec_24__ap_start_global__q0) begin
          PEG_Yvec_24__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_24__state == 2'b01) begin
        if(PEG_Yvec_24__ap_ready) begin
          if(PEG_Yvec_24__ap_done) begin
            PEG_Yvec_24__state <= 2'b10;
          end else begin
            PEG_Yvec_24__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_24__state == 2'b11) begin
        if(PEG_Yvec_24__ap_done) begin
          PEG_Yvec_24__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_24__state == 2'b10) begin
        if(PEG_Yvec_24__ap_done_global__q0) begin
          PEG_Yvec_24__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_24__ap_start = (PEG_Yvec_24__state == 2'b01);
  assign PEG_Yvec_25__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_25__is_done__q0 = (PEG_Yvec_25__state == 2'b10);
  assign PEG_Yvec_25__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_25__state <= 2'b00;
    end else begin
      if(PEG_Yvec_25__state == 2'b00) begin
        if(PEG_Yvec_25__ap_start_global__q0) begin
          PEG_Yvec_25__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_25__state == 2'b01) begin
        if(PEG_Yvec_25__ap_ready) begin
          if(PEG_Yvec_25__ap_done) begin
            PEG_Yvec_25__state <= 2'b10;
          end else begin
            PEG_Yvec_25__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_25__state == 2'b11) begin
        if(PEG_Yvec_25__ap_done) begin
          PEG_Yvec_25__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_25__state == 2'b10) begin
        if(PEG_Yvec_25__ap_done_global__q0) begin
          PEG_Yvec_25__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_25__ap_start = (PEG_Yvec_25__state == 2'b01);
  assign PEG_Yvec_26__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_26__is_done__q0 = (PEG_Yvec_26__state == 2'b10);
  assign PEG_Yvec_26__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_26__state <= 2'b00;
    end else begin
      if(PEG_Yvec_26__state == 2'b00) begin
        if(PEG_Yvec_26__ap_start_global__q0) begin
          PEG_Yvec_26__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_26__state == 2'b01) begin
        if(PEG_Yvec_26__ap_ready) begin
          if(PEG_Yvec_26__ap_done) begin
            PEG_Yvec_26__state <= 2'b10;
          end else begin
            PEG_Yvec_26__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_26__state == 2'b11) begin
        if(PEG_Yvec_26__ap_done) begin
          PEG_Yvec_26__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_26__state == 2'b10) begin
        if(PEG_Yvec_26__ap_done_global__q0) begin
          PEG_Yvec_26__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_26__ap_start = (PEG_Yvec_26__state == 2'b01);
  assign PEG_Yvec_27__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_27__is_done__q0 = (PEG_Yvec_27__state == 2'b10);
  assign PEG_Yvec_27__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_27__state <= 2'b00;
    end else begin
      if(PEG_Yvec_27__state == 2'b00) begin
        if(PEG_Yvec_27__ap_start_global__q0) begin
          PEG_Yvec_27__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_27__state == 2'b01) begin
        if(PEG_Yvec_27__ap_ready) begin
          if(PEG_Yvec_27__ap_done) begin
            PEG_Yvec_27__state <= 2'b10;
          end else begin
            PEG_Yvec_27__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_27__state == 2'b11) begin
        if(PEG_Yvec_27__ap_done) begin
          PEG_Yvec_27__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_27__state == 2'b10) begin
        if(PEG_Yvec_27__ap_done_global__q0) begin
          PEG_Yvec_27__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_27__ap_start = (PEG_Yvec_27__state == 2'b01);
  assign PEG_Yvec_28__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_28__is_done__q0 = (PEG_Yvec_28__state == 2'b10);
  assign PEG_Yvec_28__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_28__state <= 2'b00;
    end else begin
      if(PEG_Yvec_28__state == 2'b00) begin
        if(PEG_Yvec_28__ap_start_global__q0) begin
          PEG_Yvec_28__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_28__state == 2'b01) begin
        if(PEG_Yvec_28__ap_ready) begin
          if(PEG_Yvec_28__ap_done) begin
            PEG_Yvec_28__state <= 2'b10;
          end else begin
            PEG_Yvec_28__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_28__state == 2'b11) begin
        if(PEG_Yvec_28__ap_done) begin
          PEG_Yvec_28__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_28__state == 2'b10) begin
        if(PEG_Yvec_28__ap_done_global__q0) begin
          PEG_Yvec_28__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_28__ap_start = (PEG_Yvec_28__state == 2'b01);
  assign PEG_Yvec_29__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_29__is_done__q0 = (PEG_Yvec_29__state == 2'b10);
  assign PEG_Yvec_29__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_29__state <= 2'b00;
    end else begin
      if(PEG_Yvec_29__state == 2'b00) begin
        if(PEG_Yvec_29__ap_start_global__q0) begin
          PEG_Yvec_29__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_29__state == 2'b01) begin
        if(PEG_Yvec_29__ap_ready) begin
          if(PEG_Yvec_29__ap_done) begin
            PEG_Yvec_29__state <= 2'b10;
          end else begin
            PEG_Yvec_29__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_29__state == 2'b11) begin
        if(PEG_Yvec_29__ap_done) begin
          PEG_Yvec_29__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_29__state == 2'b10) begin
        if(PEG_Yvec_29__ap_done_global__q0) begin
          PEG_Yvec_29__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_29__ap_start = (PEG_Yvec_29__state == 2'b01);
  assign PEG_Yvec_30__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_30__is_done__q0 = (PEG_Yvec_30__state == 2'b10);
  assign PEG_Yvec_30__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_30__state <= 2'b00;
    end else begin
      if(PEG_Yvec_30__state == 2'b00) begin
        if(PEG_Yvec_30__ap_start_global__q0) begin
          PEG_Yvec_30__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_30__state == 2'b01) begin
        if(PEG_Yvec_30__ap_ready) begin
          if(PEG_Yvec_30__ap_done) begin
            PEG_Yvec_30__state <= 2'b10;
          end else begin
            PEG_Yvec_30__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_30__state == 2'b11) begin
        if(PEG_Yvec_30__ap_done) begin
          PEG_Yvec_30__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_30__state == 2'b10) begin
        if(PEG_Yvec_30__ap_done_global__q0) begin
          PEG_Yvec_30__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_30__ap_start = (PEG_Yvec_30__state == 2'b01);
  assign PEG_Yvec_31__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_31__is_done__q0 = (PEG_Yvec_31__state == 2'b10);
  assign PEG_Yvec_31__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_31__state <= 2'b00;
    end else begin
      if(PEG_Yvec_31__state == 2'b00) begin
        if(PEG_Yvec_31__ap_start_global__q0) begin
          PEG_Yvec_31__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_31__state == 2'b01) begin
        if(PEG_Yvec_31__ap_ready) begin
          if(PEG_Yvec_31__ap_done) begin
            PEG_Yvec_31__state <= 2'b10;
          end else begin
            PEG_Yvec_31__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_31__state == 2'b11) begin
        if(PEG_Yvec_31__ap_done) begin
          PEG_Yvec_31__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_31__state == 2'b10) begin
        if(PEG_Yvec_31__ap_done_global__q0) begin
          PEG_Yvec_31__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_31__ap_start = (PEG_Yvec_31__state == 2'b01);
  assign PEG_Yvec_32__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_32__is_done__q0 = (PEG_Yvec_32__state == 2'b10);
  assign PEG_Yvec_32__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_32__state <= 2'b00;
    end else begin
      if(PEG_Yvec_32__state == 2'b00) begin
        if(PEG_Yvec_32__ap_start_global__q0) begin
          PEG_Yvec_32__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_32__state == 2'b01) begin
        if(PEG_Yvec_32__ap_ready) begin
          if(PEG_Yvec_32__ap_done) begin
            PEG_Yvec_32__state <= 2'b10;
          end else begin
            PEG_Yvec_32__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_32__state == 2'b11) begin
        if(PEG_Yvec_32__ap_done) begin
          PEG_Yvec_32__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_32__state == 2'b10) begin
        if(PEG_Yvec_32__ap_done_global__q0) begin
          PEG_Yvec_32__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_32__ap_start = (PEG_Yvec_32__state == 2'b01);
  assign PEG_Yvec_33__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_33__is_done__q0 = (PEG_Yvec_33__state == 2'b10);
  assign PEG_Yvec_33__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_33__state <= 2'b00;
    end else begin
      if(PEG_Yvec_33__state == 2'b00) begin
        if(PEG_Yvec_33__ap_start_global__q0) begin
          PEG_Yvec_33__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_33__state == 2'b01) begin
        if(PEG_Yvec_33__ap_ready) begin
          if(PEG_Yvec_33__ap_done) begin
            PEG_Yvec_33__state <= 2'b10;
          end else begin
            PEG_Yvec_33__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_33__state == 2'b11) begin
        if(PEG_Yvec_33__ap_done) begin
          PEG_Yvec_33__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_33__state == 2'b10) begin
        if(PEG_Yvec_33__ap_done_global__q0) begin
          PEG_Yvec_33__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_33__ap_start = (PEG_Yvec_33__state == 2'b01);
  assign PEG_Yvec_34__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_34__is_done__q0 = (PEG_Yvec_34__state == 2'b10);
  assign PEG_Yvec_34__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_34__state <= 2'b00;
    end else begin
      if(PEG_Yvec_34__state == 2'b00) begin
        if(PEG_Yvec_34__ap_start_global__q0) begin
          PEG_Yvec_34__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_34__state == 2'b01) begin
        if(PEG_Yvec_34__ap_ready) begin
          if(PEG_Yvec_34__ap_done) begin
            PEG_Yvec_34__state <= 2'b10;
          end else begin
            PEG_Yvec_34__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_34__state == 2'b11) begin
        if(PEG_Yvec_34__ap_done) begin
          PEG_Yvec_34__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_34__state == 2'b10) begin
        if(PEG_Yvec_34__ap_done_global__q0) begin
          PEG_Yvec_34__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_34__ap_start = (PEG_Yvec_34__state == 2'b01);
  assign PEG_Yvec_35__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_35__is_done__q0 = (PEG_Yvec_35__state == 2'b10);
  assign PEG_Yvec_35__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_35__state <= 2'b00;
    end else begin
      if(PEG_Yvec_35__state == 2'b00) begin
        if(PEG_Yvec_35__ap_start_global__q0) begin
          PEG_Yvec_35__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_35__state == 2'b01) begin
        if(PEG_Yvec_35__ap_ready) begin
          if(PEG_Yvec_35__ap_done) begin
            PEG_Yvec_35__state <= 2'b10;
          end else begin
            PEG_Yvec_35__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_35__state == 2'b11) begin
        if(PEG_Yvec_35__ap_done) begin
          PEG_Yvec_35__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_35__state == 2'b10) begin
        if(PEG_Yvec_35__ap_done_global__q0) begin
          PEG_Yvec_35__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_35__ap_start = (PEG_Yvec_35__state == 2'b01);
  assign PEG_Yvec_36__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_36__is_done__q0 = (PEG_Yvec_36__state == 2'b10);
  assign PEG_Yvec_36__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_36__state <= 2'b00;
    end else begin
      if(PEG_Yvec_36__state == 2'b00) begin
        if(PEG_Yvec_36__ap_start_global__q0) begin
          PEG_Yvec_36__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_36__state == 2'b01) begin
        if(PEG_Yvec_36__ap_ready) begin
          if(PEG_Yvec_36__ap_done) begin
            PEG_Yvec_36__state <= 2'b10;
          end else begin
            PEG_Yvec_36__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_36__state == 2'b11) begin
        if(PEG_Yvec_36__ap_done) begin
          PEG_Yvec_36__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_36__state == 2'b10) begin
        if(PEG_Yvec_36__ap_done_global__q0) begin
          PEG_Yvec_36__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_36__ap_start = (PEG_Yvec_36__state == 2'b01);
  assign PEG_Yvec_37__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_37__is_done__q0 = (PEG_Yvec_37__state == 2'b10);
  assign PEG_Yvec_37__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_37__state <= 2'b00;
    end else begin
      if(PEG_Yvec_37__state == 2'b00) begin
        if(PEG_Yvec_37__ap_start_global__q0) begin
          PEG_Yvec_37__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_37__state == 2'b01) begin
        if(PEG_Yvec_37__ap_ready) begin
          if(PEG_Yvec_37__ap_done) begin
            PEG_Yvec_37__state <= 2'b10;
          end else begin
            PEG_Yvec_37__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_37__state == 2'b11) begin
        if(PEG_Yvec_37__ap_done) begin
          PEG_Yvec_37__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_37__state == 2'b10) begin
        if(PEG_Yvec_37__ap_done_global__q0) begin
          PEG_Yvec_37__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_37__ap_start = (PEG_Yvec_37__state == 2'b01);
  assign PEG_Yvec_38__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_38__is_done__q0 = (PEG_Yvec_38__state == 2'b10);
  assign PEG_Yvec_38__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_38__state <= 2'b00;
    end else begin
      if(PEG_Yvec_38__state == 2'b00) begin
        if(PEG_Yvec_38__ap_start_global__q0) begin
          PEG_Yvec_38__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_38__state == 2'b01) begin
        if(PEG_Yvec_38__ap_ready) begin
          if(PEG_Yvec_38__ap_done) begin
            PEG_Yvec_38__state <= 2'b10;
          end else begin
            PEG_Yvec_38__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_38__state == 2'b11) begin
        if(PEG_Yvec_38__ap_done) begin
          PEG_Yvec_38__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_38__state == 2'b10) begin
        if(PEG_Yvec_38__ap_done_global__q0) begin
          PEG_Yvec_38__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_38__ap_start = (PEG_Yvec_38__state == 2'b01);
  assign PEG_Yvec_39__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_39__is_done__q0 = (PEG_Yvec_39__state == 2'b10);
  assign PEG_Yvec_39__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_39__state <= 2'b00;
    end else begin
      if(PEG_Yvec_39__state == 2'b00) begin
        if(PEG_Yvec_39__ap_start_global__q0) begin
          PEG_Yvec_39__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_39__state == 2'b01) begin
        if(PEG_Yvec_39__ap_ready) begin
          if(PEG_Yvec_39__ap_done) begin
            PEG_Yvec_39__state <= 2'b10;
          end else begin
            PEG_Yvec_39__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_39__state == 2'b11) begin
        if(PEG_Yvec_39__ap_done) begin
          PEG_Yvec_39__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_39__state == 2'b10) begin
        if(PEG_Yvec_39__ap_done_global__q0) begin
          PEG_Yvec_39__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_39__ap_start = (PEG_Yvec_39__state == 2'b01);
  assign PEG_Yvec_40__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_40__is_done__q0 = (PEG_Yvec_40__state == 2'b10);
  assign PEG_Yvec_40__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_40__state <= 2'b00;
    end else begin
      if(PEG_Yvec_40__state == 2'b00) begin
        if(PEG_Yvec_40__ap_start_global__q0) begin
          PEG_Yvec_40__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_40__state == 2'b01) begin
        if(PEG_Yvec_40__ap_ready) begin
          if(PEG_Yvec_40__ap_done) begin
            PEG_Yvec_40__state <= 2'b10;
          end else begin
            PEG_Yvec_40__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_40__state == 2'b11) begin
        if(PEG_Yvec_40__ap_done) begin
          PEG_Yvec_40__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_40__state == 2'b10) begin
        if(PEG_Yvec_40__ap_done_global__q0) begin
          PEG_Yvec_40__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_40__ap_start = (PEG_Yvec_40__state == 2'b01);
  assign PEG_Yvec_41__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_41__is_done__q0 = (PEG_Yvec_41__state == 2'b10);
  assign PEG_Yvec_41__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_41__state <= 2'b00;
    end else begin
      if(PEG_Yvec_41__state == 2'b00) begin
        if(PEG_Yvec_41__ap_start_global__q0) begin
          PEG_Yvec_41__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_41__state == 2'b01) begin
        if(PEG_Yvec_41__ap_ready) begin
          if(PEG_Yvec_41__ap_done) begin
            PEG_Yvec_41__state <= 2'b10;
          end else begin
            PEG_Yvec_41__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_41__state == 2'b11) begin
        if(PEG_Yvec_41__ap_done) begin
          PEG_Yvec_41__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_41__state == 2'b10) begin
        if(PEG_Yvec_41__ap_done_global__q0) begin
          PEG_Yvec_41__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_41__ap_start = (PEG_Yvec_41__state == 2'b01);
  assign PEG_Yvec_42__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_42__is_done__q0 = (PEG_Yvec_42__state == 2'b10);
  assign PEG_Yvec_42__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_42__state <= 2'b00;
    end else begin
      if(PEG_Yvec_42__state == 2'b00) begin
        if(PEG_Yvec_42__ap_start_global__q0) begin
          PEG_Yvec_42__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_42__state == 2'b01) begin
        if(PEG_Yvec_42__ap_ready) begin
          if(PEG_Yvec_42__ap_done) begin
            PEG_Yvec_42__state <= 2'b10;
          end else begin
            PEG_Yvec_42__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_42__state == 2'b11) begin
        if(PEG_Yvec_42__ap_done) begin
          PEG_Yvec_42__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_42__state == 2'b10) begin
        if(PEG_Yvec_42__ap_done_global__q0) begin
          PEG_Yvec_42__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_42__ap_start = (PEG_Yvec_42__state == 2'b01);
  assign PEG_Yvec_43__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_43__is_done__q0 = (PEG_Yvec_43__state == 2'b10);
  assign PEG_Yvec_43__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_43__state <= 2'b00;
    end else begin
      if(PEG_Yvec_43__state == 2'b00) begin
        if(PEG_Yvec_43__ap_start_global__q0) begin
          PEG_Yvec_43__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_43__state == 2'b01) begin
        if(PEG_Yvec_43__ap_ready) begin
          if(PEG_Yvec_43__ap_done) begin
            PEG_Yvec_43__state <= 2'b10;
          end else begin
            PEG_Yvec_43__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_43__state == 2'b11) begin
        if(PEG_Yvec_43__ap_done) begin
          PEG_Yvec_43__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_43__state == 2'b10) begin
        if(PEG_Yvec_43__ap_done_global__q0) begin
          PEG_Yvec_43__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_43__ap_start = (PEG_Yvec_43__state == 2'b01);
  assign PEG_Yvec_44__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_44__is_done__q0 = (PEG_Yvec_44__state == 2'b10);
  assign PEG_Yvec_44__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_44__state <= 2'b00;
    end else begin
      if(PEG_Yvec_44__state == 2'b00) begin
        if(PEG_Yvec_44__ap_start_global__q0) begin
          PEG_Yvec_44__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_44__state == 2'b01) begin
        if(PEG_Yvec_44__ap_ready) begin
          if(PEG_Yvec_44__ap_done) begin
            PEG_Yvec_44__state <= 2'b10;
          end else begin
            PEG_Yvec_44__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_44__state == 2'b11) begin
        if(PEG_Yvec_44__ap_done) begin
          PEG_Yvec_44__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_44__state == 2'b10) begin
        if(PEG_Yvec_44__ap_done_global__q0) begin
          PEG_Yvec_44__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_44__ap_start = (PEG_Yvec_44__state == 2'b01);
  assign PEG_Yvec_45__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_45__is_done__q0 = (PEG_Yvec_45__state == 2'b10);
  assign PEG_Yvec_45__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_45__state <= 2'b00;
    end else begin
      if(PEG_Yvec_45__state == 2'b00) begin
        if(PEG_Yvec_45__ap_start_global__q0) begin
          PEG_Yvec_45__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_45__state == 2'b01) begin
        if(PEG_Yvec_45__ap_ready) begin
          if(PEG_Yvec_45__ap_done) begin
            PEG_Yvec_45__state <= 2'b10;
          end else begin
            PEG_Yvec_45__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_45__state == 2'b11) begin
        if(PEG_Yvec_45__ap_done) begin
          PEG_Yvec_45__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_45__state == 2'b10) begin
        if(PEG_Yvec_45__ap_done_global__q0) begin
          PEG_Yvec_45__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_45__ap_start = (PEG_Yvec_45__state == 2'b01);
  assign PEG_Yvec_46__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_46__is_done__q0 = (PEG_Yvec_46__state == 2'b10);
  assign PEG_Yvec_46__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_46__state <= 2'b00;
    end else begin
      if(PEG_Yvec_46__state == 2'b00) begin
        if(PEG_Yvec_46__ap_start_global__q0) begin
          PEG_Yvec_46__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_46__state == 2'b01) begin
        if(PEG_Yvec_46__ap_ready) begin
          if(PEG_Yvec_46__ap_done) begin
            PEG_Yvec_46__state <= 2'b10;
          end else begin
            PEG_Yvec_46__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_46__state == 2'b11) begin
        if(PEG_Yvec_46__ap_done) begin
          PEG_Yvec_46__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_46__state == 2'b10) begin
        if(PEG_Yvec_46__ap_done_global__q0) begin
          PEG_Yvec_46__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_46__ap_start = (PEG_Yvec_46__state == 2'b01);
  assign PEG_Yvec_47__ap_start_global__q0 = ap_start__q0;
  assign PEG_Yvec_47__is_done__q0 = (PEG_Yvec_47__state == 2'b10);
  assign PEG_Yvec_47__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      PEG_Yvec_47__state <= 2'b00;
    end else begin
      if(PEG_Yvec_47__state == 2'b00) begin
        if(PEG_Yvec_47__ap_start_global__q0) begin
          PEG_Yvec_47__state <= 2'b01;
        end 
      end 
      if(PEG_Yvec_47__state == 2'b01) begin
        if(PEG_Yvec_47__ap_ready) begin
          if(PEG_Yvec_47__ap_done) begin
            PEG_Yvec_47__state <= 2'b10;
          end else begin
            PEG_Yvec_47__state <= 2'b11;
          end
        end 
      end 
      if(PEG_Yvec_47__state == 2'b11) begin
        if(PEG_Yvec_47__ap_done) begin
          PEG_Yvec_47__state <= 2'b10;
        end 
      end 
      if(PEG_Yvec_47__state == 2'b10) begin
        if(PEG_Yvec_47__ap_done_global__q0) begin
          PEG_Yvec_47__state <= 2'b00;
        end 
      end 
    end
  end

  assign PEG_Yvec_47__ap_start = (PEG_Yvec_47__state == 2'b01);
  assign black_hole_float_v16_0__ap_start_global__q0 = ap_start__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      black_hole_float_v16_0__ap_start <= 1'b0;
    end else if(black_hole_float_v16_0__ap_start_global__q0) begin
      black_hole_float_v16_0__ap_start <= 1'b1;
    end 
  end

  assign black_hole_int_0__ap_start_global__q0 = ap_start__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      black_hole_int_0__ap_start <= 1'b0;
    end else if(black_hole_int_0__ap_start_global__q0) begin
      black_hole_int_0__ap_start <= 1'b1;
    end 
  end

  assign read_A_0___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_0___P_N__q0 = P_N;
  assign read_A_0___edge_list_ch_0__q0 = edge_list_ch_0;
  assign read_A_0__ap_start_global__q0 = ap_start__q0;
  assign read_A_0__is_done__q0 = (read_A_0__state == 2'b10);
  assign read_A_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_0__state <= 2'b00;
    end else begin
      if(read_A_0__state == 2'b00) begin
        if(read_A_0__ap_start_global__q0) begin
          read_A_0__state <= 2'b01;
        end 
      end 
      if(read_A_0__state == 2'b01) begin
        if(read_A_0__ap_ready) begin
          if(read_A_0__ap_done) begin
            read_A_0__state <= 2'b10;
          end else begin
            read_A_0__state <= 2'b11;
          end
        end 
      end 
      if(read_A_0__state == 2'b11) begin
        if(read_A_0__ap_done) begin
          read_A_0__state <= 2'b10;
        end 
      end 
      if(read_A_0__state == 2'b10) begin
        if(read_A_0__ap_done_global__q0) begin
          read_A_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_0__ap_start = (read_A_0__state == 2'b01);
  assign read_A_1___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_1___P_N__q0 = P_N;
  assign read_A_1___edge_list_ch_1__q0 = edge_list_ch_1;
  assign read_A_1__ap_start_global__q0 = ap_start__q0;
  assign read_A_1__is_done__q0 = (read_A_1__state == 2'b10);
  assign read_A_1__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_1__state <= 2'b00;
    end else begin
      if(read_A_1__state == 2'b00) begin
        if(read_A_1__ap_start_global__q0) begin
          read_A_1__state <= 2'b01;
        end 
      end 
      if(read_A_1__state == 2'b01) begin
        if(read_A_1__ap_ready) begin
          if(read_A_1__ap_done) begin
            read_A_1__state <= 2'b10;
          end else begin
            read_A_1__state <= 2'b11;
          end
        end 
      end 
      if(read_A_1__state == 2'b11) begin
        if(read_A_1__ap_done) begin
          read_A_1__state <= 2'b10;
        end 
      end 
      if(read_A_1__state == 2'b10) begin
        if(read_A_1__ap_done_global__q0) begin
          read_A_1__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_1__ap_start = (read_A_1__state == 2'b01);
  assign read_A_2___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_2___P_N__q0 = P_N;
  assign read_A_2___edge_list_ch_2__q0 = edge_list_ch_2;
  assign read_A_2__ap_start_global__q0 = ap_start__q0;
  assign read_A_2__is_done__q0 = (read_A_2__state == 2'b10);
  assign read_A_2__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_2__state <= 2'b00;
    end else begin
      if(read_A_2__state == 2'b00) begin
        if(read_A_2__ap_start_global__q0) begin
          read_A_2__state <= 2'b01;
        end 
      end 
      if(read_A_2__state == 2'b01) begin
        if(read_A_2__ap_ready) begin
          if(read_A_2__ap_done) begin
            read_A_2__state <= 2'b10;
          end else begin
            read_A_2__state <= 2'b11;
          end
        end 
      end 
      if(read_A_2__state == 2'b11) begin
        if(read_A_2__ap_done) begin
          read_A_2__state <= 2'b10;
        end 
      end 
      if(read_A_2__state == 2'b10) begin
        if(read_A_2__ap_done_global__q0) begin
          read_A_2__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_2__ap_start = (read_A_2__state == 2'b01);
  assign read_A_3___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_3___P_N__q0 = P_N;
  assign read_A_3___edge_list_ch_3__q0 = edge_list_ch_3;
  assign read_A_3__ap_start_global__q0 = ap_start__q0;
  assign read_A_3__is_done__q0 = (read_A_3__state == 2'b10);
  assign read_A_3__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_3__state <= 2'b00;
    end else begin
      if(read_A_3__state == 2'b00) begin
        if(read_A_3__ap_start_global__q0) begin
          read_A_3__state <= 2'b01;
        end 
      end 
      if(read_A_3__state == 2'b01) begin
        if(read_A_3__ap_ready) begin
          if(read_A_3__ap_done) begin
            read_A_3__state <= 2'b10;
          end else begin
            read_A_3__state <= 2'b11;
          end
        end 
      end 
      if(read_A_3__state == 2'b11) begin
        if(read_A_3__ap_done) begin
          read_A_3__state <= 2'b10;
        end 
      end 
      if(read_A_3__state == 2'b10) begin
        if(read_A_3__ap_done_global__q0) begin
          read_A_3__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_3__ap_start = (read_A_3__state == 2'b01);
  assign read_A_4___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_4___P_N__q0 = P_N;
  assign read_A_4___edge_list_ch_4__q0 = edge_list_ch_4;
  assign read_A_4__ap_start_global__q0 = ap_start__q0;
  assign read_A_4__is_done__q0 = (read_A_4__state == 2'b10);
  assign read_A_4__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_4__state <= 2'b00;
    end else begin
      if(read_A_4__state == 2'b00) begin
        if(read_A_4__ap_start_global__q0) begin
          read_A_4__state <= 2'b01;
        end 
      end 
      if(read_A_4__state == 2'b01) begin
        if(read_A_4__ap_ready) begin
          if(read_A_4__ap_done) begin
            read_A_4__state <= 2'b10;
          end else begin
            read_A_4__state <= 2'b11;
          end
        end 
      end 
      if(read_A_4__state == 2'b11) begin
        if(read_A_4__ap_done) begin
          read_A_4__state <= 2'b10;
        end 
      end 
      if(read_A_4__state == 2'b10) begin
        if(read_A_4__ap_done_global__q0) begin
          read_A_4__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_4__ap_start = (read_A_4__state == 2'b01);
  assign read_A_5___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_5___P_N__q0 = P_N;
  assign read_A_5___edge_list_ch_5__q0 = edge_list_ch_5;
  assign read_A_5__ap_start_global__q0 = ap_start__q0;
  assign read_A_5__is_done__q0 = (read_A_5__state == 2'b10);
  assign read_A_5__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_5__state <= 2'b00;
    end else begin
      if(read_A_5__state == 2'b00) begin
        if(read_A_5__ap_start_global__q0) begin
          read_A_5__state <= 2'b01;
        end 
      end 
      if(read_A_5__state == 2'b01) begin
        if(read_A_5__ap_ready) begin
          if(read_A_5__ap_done) begin
            read_A_5__state <= 2'b10;
          end else begin
            read_A_5__state <= 2'b11;
          end
        end 
      end 
      if(read_A_5__state == 2'b11) begin
        if(read_A_5__ap_done) begin
          read_A_5__state <= 2'b10;
        end 
      end 
      if(read_A_5__state == 2'b10) begin
        if(read_A_5__ap_done_global__q0) begin
          read_A_5__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_5__ap_start = (read_A_5__state == 2'b01);
  assign read_A_6___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_6___P_N__q0 = P_N;
  assign read_A_6___edge_list_ch_6__q0 = edge_list_ch_6;
  assign read_A_6__ap_start_global__q0 = ap_start__q0;
  assign read_A_6__is_done__q0 = (read_A_6__state == 2'b10);
  assign read_A_6__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_6__state <= 2'b00;
    end else begin
      if(read_A_6__state == 2'b00) begin
        if(read_A_6__ap_start_global__q0) begin
          read_A_6__state <= 2'b01;
        end 
      end 
      if(read_A_6__state == 2'b01) begin
        if(read_A_6__ap_ready) begin
          if(read_A_6__ap_done) begin
            read_A_6__state <= 2'b10;
          end else begin
            read_A_6__state <= 2'b11;
          end
        end 
      end 
      if(read_A_6__state == 2'b11) begin
        if(read_A_6__ap_done) begin
          read_A_6__state <= 2'b10;
        end 
      end 
      if(read_A_6__state == 2'b10) begin
        if(read_A_6__ap_done_global__q0) begin
          read_A_6__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_6__ap_start = (read_A_6__state == 2'b01);
  assign read_A_7___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_7___P_N__q0 = P_N;
  assign read_A_7___edge_list_ch_7__q0 = edge_list_ch_7;
  assign read_A_7__ap_start_global__q0 = ap_start__q0;
  assign read_A_7__is_done__q0 = (read_A_7__state == 2'b10);
  assign read_A_7__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_7__state <= 2'b00;
    end else begin
      if(read_A_7__state == 2'b00) begin
        if(read_A_7__ap_start_global__q0) begin
          read_A_7__state <= 2'b01;
        end 
      end 
      if(read_A_7__state == 2'b01) begin
        if(read_A_7__ap_ready) begin
          if(read_A_7__ap_done) begin
            read_A_7__state <= 2'b10;
          end else begin
            read_A_7__state <= 2'b11;
          end
        end 
      end 
      if(read_A_7__state == 2'b11) begin
        if(read_A_7__ap_done) begin
          read_A_7__state <= 2'b10;
        end 
      end 
      if(read_A_7__state == 2'b10) begin
        if(read_A_7__ap_done_global__q0) begin
          read_A_7__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_7__ap_start = (read_A_7__state == 2'b01);
  assign read_A_8___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_8___P_N__q0 = P_N;
  assign read_A_8___edge_list_ch_8__q0 = edge_list_ch_8;
  assign read_A_8__ap_start_global__q0 = ap_start__q0;
  assign read_A_8__is_done__q0 = (read_A_8__state == 2'b10);
  assign read_A_8__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_8__state <= 2'b00;
    end else begin
      if(read_A_8__state == 2'b00) begin
        if(read_A_8__ap_start_global__q0) begin
          read_A_8__state <= 2'b01;
        end 
      end 
      if(read_A_8__state == 2'b01) begin
        if(read_A_8__ap_ready) begin
          if(read_A_8__ap_done) begin
            read_A_8__state <= 2'b10;
          end else begin
            read_A_8__state <= 2'b11;
          end
        end 
      end 
      if(read_A_8__state == 2'b11) begin
        if(read_A_8__ap_done) begin
          read_A_8__state <= 2'b10;
        end 
      end 
      if(read_A_8__state == 2'b10) begin
        if(read_A_8__ap_done_global__q0) begin
          read_A_8__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_8__ap_start = (read_A_8__state == 2'b01);
  assign read_A_9___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_9___P_N__q0 = P_N;
  assign read_A_9___edge_list_ch_9__q0 = edge_list_ch_9;
  assign read_A_9__ap_start_global__q0 = ap_start__q0;
  assign read_A_9__is_done__q0 = (read_A_9__state == 2'b10);
  assign read_A_9__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_9__state <= 2'b00;
    end else begin
      if(read_A_9__state == 2'b00) begin
        if(read_A_9__ap_start_global__q0) begin
          read_A_9__state <= 2'b01;
        end 
      end 
      if(read_A_9__state == 2'b01) begin
        if(read_A_9__ap_ready) begin
          if(read_A_9__ap_done) begin
            read_A_9__state <= 2'b10;
          end else begin
            read_A_9__state <= 2'b11;
          end
        end 
      end 
      if(read_A_9__state == 2'b11) begin
        if(read_A_9__ap_done) begin
          read_A_9__state <= 2'b10;
        end 
      end 
      if(read_A_9__state == 2'b10) begin
        if(read_A_9__ap_done_global__q0) begin
          read_A_9__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_9__ap_start = (read_A_9__state == 2'b01);
  assign read_A_10___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_10___P_N__q0 = P_N;
  assign read_A_10___edge_list_ch_10__q0 = edge_list_ch_10;
  assign read_A_10__ap_start_global__q0 = ap_start__q0;
  assign read_A_10__is_done__q0 = (read_A_10__state == 2'b10);
  assign read_A_10__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_10__state <= 2'b00;
    end else begin
      if(read_A_10__state == 2'b00) begin
        if(read_A_10__ap_start_global__q0) begin
          read_A_10__state <= 2'b01;
        end 
      end 
      if(read_A_10__state == 2'b01) begin
        if(read_A_10__ap_ready) begin
          if(read_A_10__ap_done) begin
            read_A_10__state <= 2'b10;
          end else begin
            read_A_10__state <= 2'b11;
          end
        end 
      end 
      if(read_A_10__state == 2'b11) begin
        if(read_A_10__ap_done) begin
          read_A_10__state <= 2'b10;
        end 
      end 
      if(read_A_10__state == 2'b10) begin
        if(read_A_10__ap_done_global__q0) begin
          read_A_10__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_10__ap_start = (read_A_10__state == 2'b01);
  assign read_A_11___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_11___P_N__q0 = P_N;
  assign read_A_11___edge_list_ch_11__q0 = edge_list_ch_11;
  assign read_A_11__ap_start_global__q0 = ap_start__q0;
  assign read_A_11__is_done__q0 = (read_A_11__state == 2'b10);
  assign read_A_11__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_11__state <= 2'b00;
    end else begin
      if(read_A_11__state == 2'b00) begin
        if(read_A_11__ap_start_global__q0) begin
          read_A_11__state <= 2'b01;
        end 
      end 
      if(read_A_11__state == 2'b01) begin
        if(read_A_11__ap_ready) begin
          if(read_A_11__ap_done) begin
            read_A_11__state <= 2'b10;
          end else begin
            read_A_11__state <= 2'b11;
          end
        end 
      end 
      if(read_A_11__state == 2'b11) begin
        if(read_A_11__ap_done) begin
          read_A_11__state <= 2'b10;
        end 
      end 
      if(read_A_11__state == 2'b10) begin
        if(read_A_11__ap_done_global__q0) begin
          read_A_11__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_11__ap_start = (read_A_11__state == 2'b01);
  assign read_A_12___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_12___P_N__q0 = P_N;
  assign read_A_12___edge_list_ch_12__q0 = edge_list_ch_12;
  assign read_A_12__ap_start_global__q0 = ap_start__q0;
  assign read_A_12__is_done__q0 = (read_A_12__state == 2'b10);
  assign read_A_12__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_12__state <= 2'b00;
    end else begin
      if(read_A_12__state == 2'b00) begin
        if(read_A_12__ap_start_global__q0) begin
          read_A_12__state <= 2'b01;
        end 
      end 
      if(read_A_12__state == 2'b01) begin
        if(read_A_12__ap_ready) begin
          if(read_A_12__ap_done) begin
            read_A_12__state <= 2'b10;
          end else begin
            read_A_12__state <= 2'b11;
          end
        end 
      end 
      if(read_A_12__state == 2'b11) begin
        if(read_A_12__ap_done) begin
          read_A_12__state <= 2'b10;
        end 
      end 
      if(read_A_12__state == 2'b10) begin
        if(read_A_12__ap_done_global__q0) begin
          read_A_12__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_12__ap_start = (read_A_12__state == 2'b01);
  assign read_A_13___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_13___P_N__q0 = P_N;
  assign read_A_13___edge_list_ch_13__q0 = edge_list_ch_13;
  assign read_A_13__ap_start_global__q0 = ap_start__q0;
  assign read_A_13__is_done__q0 = (read_A_13__state == 2'b10);
  assign read_A_13__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_13__state <= 2'b00;
    end else begin
      if(read_A_13__state == 2'b00) begin
        if(read_A_13__ap_start_global__q0) begin
          read_A_13__state <= 2'b01;
        end 
      end 
      if(read_A_13__state == 2'b01) begin
        if(read_A_13__ap_ready) begin
          if(read_A_13__ap_done) begin
            read_A_13__state <= 2'b10;
          end else begin
            read_A_13__state <= 2'b11;
          end
        end 
      end 
      if(read_A_13__state == 2'b11) begin
        if(read_A_13__ap_done) begin
          read_A_13__state <= 2'b10;
        end 
      end 
      if(read_A_13__state == 2'b10) begin
        if(read_A_13__ap_done_global__q0) begin
          read_A_13__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_13__ap_start = (read_A_13__state == 2'b01);
  assign read_A_14___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_14___P_N__q0 = P_N;
  assign read_A_14___edge_list_ch_14__q0 = edge_list_ch_14;
  assign read_A_14__ap_start_global__q0 = ap_start__q0;
  assign read_A_14__is_done__q0 = (read_A_14__state == 2'b10);
  assign read_A_14__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_14__state <= 2'b00;
    end else begin
      if(read_A_14__state == 2'b00) begin
        if(read_A_14__ap_start_global__q0) begin
          read_A_14__state <= 2'b01;
        end 
      end 
      if(read_A_14__state == 2'b01) begin
        if(read_A_14__ap_ready) begin
          if(read_A_14__ap_done) begin
            read_A_14__state <= 2'b10;
          end else begin
            read_A_14__state <= 2'b11;
          end
        end 
      end 
      if(read_A_14__state == 2'b11) begin
        if(read_A_14__ap_done) begin
          read_A_14__state <= 2'b10;
        end 
      end 
      if(read_A_14__state == 2'b10) begin
        if(read_A_14__ap_done_global__q0) begin
          read_A_14__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_14__ap_start = (read_A_14__state == 2'b01);
  assign read_A_15___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_15___P_N__q0 = P_N;
  assign read_A_15___edge_list_ch_15__q0 = edge_list_ch_15;
  assign read_A_15__ap_start_global__q0 = ap_start__q0;
  assign read_A_15__is_done__q0 = (read_A_15__state == 2'b10);
  assign read_A_15__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_15__state <= 2'b00;
    end else begin
      if(read_A_15__state == 2'b00) begin
        if(read_A_15__ap_start_global__q0) begin
          read_A_15__state <= 2'b01;
        end 
      end 
      if(read_A_15__state == 2'b01) begin
        if(read_A_15__ap_ready) begin
          if(read_A_15__ap_done) begin
            read_A_15__state <= 2'b10;
          end else begin
            read_A_15__state <= 2'b11;
          end
        end 
      end 
      if(read_A_15__state == 2'b11) begin
        if(read_A_15__ap_done) begin
          read_A_15__state <= 2'b10;
        end 
      end 
      if(read_A_15__state == 2'b10) begin
        if(read_A_15__ap_done_global__q0) begin
          read_A_15__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_15__ap_start = (read_A_15__state == 2'b01);
  assign read_A_16___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_16___P_N__q0 = P_N;
  assign read_A_16___edge_list_ch_16__q0 = edge_list_ch_16;
  assign read_A_16__ap_start_global__q0 = ap_start__q0;
  assign read_A_16__is_done__q0 = (read_A_16__state == 2'b10);
  assign read_A_16__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_16__state <= 2'b00;
    end else begin
      if(read_A_16__state == 2'b00) begin
        if(read_A_16__ap_start_global__q0) begin
          read_A_16__state <= 2'b01;
        end 
      end 
      if(read_A_16__state == 2'b01) begin
        if(read_A_16__ap_ready) begin
          if(read_A_16__ap_done) begin
            read_A_16__state <= 2'b10;
          end else begin
            read_A_16__state <= 2'b11;
          end
        end 
      end 
      if(read_A_16__state == 2'b11) begin
        if(read_A_16__ap_done) begin
          read_A_16__state <= 2'b10;
        end 
      end 
      if(read_A_16__state == 2'b10) begin
        if(read_A_16__ap_done_global__q0) begin
          read_A_16__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_16__ap_start = (read_A_16__state == 2'b01);
  assign read_A_17___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_17___P_N__q0 = P_N;
  assign read_A_17___edge_list_ch_17__q0 = edge_list_ch_17;
  assign read_A_17__ap_start_global__q0 = ap_start__q0;
  assign read_A_17__is_done__q0 = (read_A_17__state == 2'b10);
  assign read_A_17__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_17__state <= 2'b00;
    end else begin
      if(read_A_17__state == 2'b00) begin
        if(read_A_17__ap_start_global__q0) begin
          read_A_17__state <= 2'b01;
        end 
      end 
      if(read_A_17__state == 2'b01) begin
        if(read_A_17__ap_ready) begin
          if(read_A_17__ap_done) begin
            read_A_17__state <= 2'b10;
          end else begin
            read_A_17__state <= 2'b11;
          end
        end 
      end 
      if(read_A_17__state == 2'b11) begin
        if(read_A_17__ap_done) begin
          read_A_17__state <= 2'b10;
        end 
      end 
      if(read_A_17__state == 2'b10) begin
        if(read_A_17__ap_done_global__q0) begin
          read_A_17__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_17__ap_start = (read_A_17__state == 2'b01);
  assign read_A_18___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_18___P_N__q0 = P_N;
  assign read_A_18___edge_list_ch_18__q0 = edge_list_ch_18;
  assign read_A_18__ap_start_global__q0 = ap_start__q0;
  assign read_A_18__is_done__q0 = (read_A_18__state == 2'b10);
  assign read_A_18__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_18__state <= 2'b00;
    end else begin
      if(read_A_18__state == 2'b00) begin
        if(read_A_18__ap_start_global__q0) begin
          read_A_18__state <= 2'b01;
        end 
      end 
      if(read_A_18__state == 2'b01) begin
        if(read_A_18__ap_ready) begin
          if(read_A_18__ap_done) begin
            read_A_18__state <= 2'b10;
          end else begin
            read_A_18__state <= 2'b11;
          end
        end 
      end 
      if(read_A_18__state == 2'b11) begin
        if(read_A_18__ap_done) begin
          read_A_18__state <= 2'b10;
        end 
      end 
      if(read_A_18__state == 2'b10) begin
        if(read_A_18__ap_done_global__q0) begin
          read_A_18__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_18__ap_start = (read_A_18__state == 2'b01);
  assign read_A_19___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_19___P_N__q0 = P_N;
  assign read_A_19___edge_list_ch_19__q0 = edge_list_ch_19;
  assign read_A_19__ap_start_global__q0 = ap_start__q0;
  assign read_A_19__is_done__q0 = (read_A_19__state == 2'b10);
  assign read_A_19__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_19__state <= 2'b00;
    end else begin
      if(read_A_19__state == 2'b00) begin
        if(read_A_19__ap_start_global__q0) begin
          read_A_19__state <= 2'b01;
        end 
      end 
      if(read_A_19__state == 2'b01) begin
        if(read_A_19__ap_ready) begin
          if(read_A_19__ap_done) begin
            read_A_19__state <= 2'b10;
          end else begin
            read_A_19__state <= 2'b11;
          end
        end 
      end 
      if(read_A_19__state == 2'b11) begin
        if(read_A_19__ap_done) begin
          read_A_19__state <= 2'b10;
        end 
      end 
      if(read_A_19__state == 2'b10) begin
        if(read_A_19__ap_done_global__q0) begin
          read_A_19__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_19__ap_start = (read_A_19__state == 2'b01);
  assign read_A_20___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_20___P_N__q0 = P_N;
  assign read_A_20___edge_list_ch_20__q0 = edge_list_ch_20;
  assign read_A_20__ap_start_global__q0 = ap_start__q0;
  assign read_A_20__is_done__q0 = (read_A_20__state == 2'b10);
  assign read_A_20__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_20__state <= 2'b00;
    end else begin
      if(read_A_20__state == 2'b00) begin
        if(read_A_20__ap_start_global__q0) begin
          read_A_20__state <= 2'b01;
        end 
      end 
      if(read_A_20__state == 2'b01) begin
        if(read_A_20__ap_ready) begin
          if(read_A_20__ap_done) begin
            read_A_20__state <= 2'b10;
          end else begin
            read_A_20__state <= 2'b11;
          end
        end 
      end 
      if(read_A_20__state == 2'b11) begin
        if(read_A_20__ap_done) begin
          read_A_20__state <= 2'b10;
        end 
      end 
      if(read_A_20__state == 2'b10) begin
        if(read_A_20__ap_done_global__q0) begin
          read_A_20__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_20__ap_start = (read_A_20__state == 2'b01);
  assign read_A_21___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_21___P_N__q0 = P_N;
  assign read_A_21___edge_list_ch_21__q0 = edge_list_ch_21;
  assign read_A_21__ap_start_global__q0 = ap_start__q0;
  assign read_A_21__is_done__q0 = (read_A_21__state == 2'b10);
  assign read_A_21__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_21__state <= 2'b00;
    end else begin
      if(read_A_21__state == 2'b00) begin
        if(read_A_21__ap_start_global__q0) begin
          read_A_21__state <= 2'b01;
        end 
      end 
      if(read_A_21__state == 2'b01) begin
        if(read_A_21__ap_ready) begin
          if(read_A_21__ap_done) begin
            read_A_21__state <= 2'b10;
          end else begin
            read_A_21__state <= 2'b11;
          end
        end 
      end 
      if(read_A_21__state == 2'b11) begin
        if(read_A_21__ap_done) begin
          read_A_21__state <= 2'b10;
        end 
      end 
      if(read_A_21__state == 2'b10) begin
        if(read_A_21__ap_done_global__q0) begin
          read_A_21__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_21__ap_start = (read_A_21__state == 2'b01);
  assign read_A_22___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_22___P_N__q0 = P_N;
  assign read_A_22___edge_list_ch_22__q0 = edge_list_ch_22;
  assign read_A_22__ap_start_global__q0 = ap_start__q0;
  assign read_A_22__is_done__q0 = (read_A_22__state == 2'b10);
  assign read_A_22__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_22__state <= 2'b00;
    end else begin
      if(read_A_22__state == 2'b00) begin
        if(read_A_22__ap_start_global__q0) begin
          read_A_22__state <= 2'b01;
        end 
      end 
      if(read_A_22__state == 2'b01) begin
        if(read_A_22__ap_ready) begin
          if(read_A_22__ap_done) begin
            read_A_22__state <= 2'b10;
          end else begin
            read_A_22__state <= 2'b11;
          end
        end 
      end 
      if(read_A_22__state == 2'b11) begin
        if(read_A_22__ap_done) begin
          read_A_22__state <= 2'b10;
        end 
      end 
      if(read_A_22__state == 2'b10) begin
        if(read_A_22__ap_done_global__q0) begin
          read_A_22__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_22__ap_start = (read_A_22__state == 2'b01);
  assign read_A_23___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_23___P_N__q0 = P_N;
  assign read_A_23___edge_list_ch_23__q0 = edge_list_ch_23;
  assign read_A_23__ap_start_global__q0 = ap_start__q0;
  assign read_A_23__is_done__q0 = (read_A_23__state == 2'b10);
  assign read_A_23__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_23__state <= 2'b00;
    end else begin
      if(read_A_23__state == 2'b00) begin
        if(read_A_23__ap_start_global__q0) begin
          read_A_23__state <= 2'b01;
        end 
      end 
      if(read_A_23__state == 2'b01) begin
        if(read_A_23__ap_ready) begin
          if(read_A_23__ap_done) begin
            read_A_23__state <= 2'b10;
          end else begin
            read_A_23__state <= 2'b11;
          end
        end 
      end 
      if(read_A_23__state == 2'b11) begin
        if(read_A_23__ap_done) begin
          read_A_23__state <= 2'b10;
        end 
      end 
      if(read_A_23__state == 2'b10) begin
        if(read_A_23__ap_done_global__q0) begin
          read_A_23__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_23__ap_start = (read_A_23__state == 2'b01);
  assign read_A_24___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_24___P_N__q0 = P_N;
  assign read_A_24___edge_list_ch_24__q0 = edge_list_ch_24;
  assign read_A_24__ap_start_global__q0 = ap_start__q0;
  assign read_A_24__is_done__q0 = (read_A_24__state == 2'b10);
  assign read_A_24__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_24__state <= 2'b00;
    end else begin
      if(read_A_24__state == 2'b00) begin
        if(read_A_24__ap_start_global__q0) begin
          read_A_24__state <= 2'b01;
        end 
      end 
      if(read_A_24__state == 2'b01) begin
        if(read_A_24__ap_ready) begin
          if(read_A_24__ap_done) begin
            read_A_24__state <= 2'b10;
          end else begin
            read_A_24__state <= 2'b11;
          end
        end 
      end 
      if(read_A_24__state == 2'b11) begin
        if(read_A_24__ap_done) begin
          read_A_24__state <= 2'b10;
        end 
      end 
      if(read_A_24__state == 2'b10) begin
        if(read_A_24__ap_done_global__q0) begin
          read_A_24__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_24__ap_start = (read_A_24__state == 2'b01);
  assign read_A_25___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_25___P_N__q0 = P_N;
  assign read_A_25___edge_list_ch_25__q0 = edge_list_ch_25;
  assign read_A_25__ap_start_global__q0 = ap_start__q0;
  assign read_A_25__is_done__q0 = (read_A_25__state == 2'b10);
  assign read_A_25__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_25__state <= 2'b00;
    end else begin
      if(read_A_25__state == 2'b00) begin
        if(read_A_25__ap_start_global__q0) begin
          read_A_25__state <= 2'b01;
        end 
      end 
      if(read_A_25__state == 2'b01) begin
        if(read_A_25__ap_ready) begin
          if(read_A_25__ap_done) begin
            read_A_25__state <= 2'b10;
          end else begin
            read_A_25__state <= 2'b11;
          end
        end 
      end 
      if(read_A_25__state == 2'b11) begin
        if(read_A_25__ap_done) begin
          read_A_25__state <= 2'b10;
        end 
      end 
      if(read_A_25__state == 2'b10) begin
        if(read_A_25__ap_done_global__q0) begin
          read_A_25__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_25__ap_start = (read_A_25__state == 2'b01);
  assign read_A_26___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_26___P_N__q0 = P_N;
  assign read_A_26___edge_list_ch_26__q0 = edge_list_ch_26;
  assign read_A_26__ap_start_global__q0 = ap_start__q0;
  assign read_A_26__is_done__q0 = (read_A_26__state == 2'b10);
  assign read_A_26__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_26__state <= 2'b00;
    end else begin
      if(read_A_26__state == 2'b00) begin
        if(read_A_26__ap_start_global__q0) begin
          read_A_26__state <= 2'b01;
        end 
      end 
      if(read_A_26__state == 2'b01) begin
        if(read_A_26__ap_ready) begin
          if(read_A_26__ap_done) begin
            read_A_26__state <= 2'b10;
          end else begin
            read_A_26__state <= 2'b11;
          end
        end 
      end 
      if(read_A_26__state == 2'b11) begin
        if(read_A_26__ap_done) begin
          read_A_26__state <= 2'b10;
        end 
      end 
      if(read_A_26__state == 2'b10) begin
        if(read_A_26__ap_done_global__q0) begin
          read_A_26__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_26__ap_start = (read_A_26__state == 2'b01);
  assign read_A_27___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_27___P_N__q0 = P_N;
  assign read_A_27___edge_list_ch_27__q0 = edge_list_ch_27;
  assign read_A_27__ap_start_global__q0 = ap_start__q0;
  assign read_A_27__is_done__q0 = (read_A_27__state == 2'b10);
  assign read_A_27__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_27__state <= 2'b00;
    end else begin
      if(read_A_27__state == 2'b00) begin
        if(read_A_27__ap_start_global__q0) begin
          read_A_27__state <= 2'b01;
        end 
      end 
      if(read_A_27__state == 2'b01) begin
        if(read_A_27__ap_ready) begin
          if(read_A_27__ap_done) begin
            read_A_27__state <= 2'b10;
          end else begin
            read_A_27__state <= 2'b11;
          end
        end 
      end 
      if(read_A_27__state == 2'b11) begin
        if(read_A_27__ap_done) begin
          read_A_27__state <= 2'b10;
        end 
      end 
      if(read_A_27__state == 2'b10) begin
        if(read_A_27__ap_done_global__q0) begin
          read_A_27__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_27__ap_start = (read_A_27__state == 2'b01);
  assign read_A_28___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_28___P_N__q0 = P_N;
  assign read_A_28___edge_list_ch_28__q0 = edge_list_ch_28;
  assign read_A_28__ap_start_global__q0 = ap_start__q0;
  assign read_A_28__is_done__q0 = (read_A_28__state == 2'b10);
  assign read_A_28__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_28__state <= 2'b00;
    end else begin
      if(read_A_28__state == 2'b00) begin
        if(read_A_28__ap_start_global__q0) begin
          read_A_28__state <= 2'b01;
        end 
      end 
      if(read_A_28__state == 2'b01) begin
        if(read_A_28__ap_ready) begin
          if(read_A_28__ap_done) begin
            read_A_28__state <= 2'b10;
          end else begin
            read_A_28__state <= 2'b11;
          end
        end 
      end 
      if(read_A_28__state == 2'b11) begin
        if(read_A_28__ap_done) begin
          read_A_28__state <= 2'b10;
        end 
      end 
      if(read_A_28__state == 2'b10) begin
        if(read_A_28__ap_done_global__q0) begin
          read_A_28__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_28__ap_start = (read_A_28__state == 2'b01);
  assign read_A_29___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_29___P_N__q0 = P_N;
  assign read_A_29___edge_list_ch_29__q0 = edge_list_ch_29;
  assign read_A_29__ap_start_global__q0 = ap_start__q0;
  assign read_A_29__is_done__q0 = (read_A_29__state == 2'b10);
  assign read_A_29__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_29__state <= 2'b00;
    end else begin
      if(read_A_29__state == 2'b00) begin
        if(read_A_29__ap_start_global__q0) begin
          read_A_29__state <= 2'b01;
        end 
      end 
      if(read_A_29__state == 2'b01) begin
        if(read_A_29__ap_ready) begin
          if(read_A_29__ap_done) begin
            read_A_29__state <= 2'b10;
          end else begin
            read_A_29__state <= 2'b11;
          end
        end 
      end 
      if(read_A_29__state == 2'b11) begin
        if(read_A_29__ap_done) begin
          read_A_29__state <= 2'b10;
        end 
      end 
      if(read_A_29__state == 2'b10) begin
        if(read_A_29__ap_done_global__q0) begin
          read_A_29__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_29__ap_start = (read_A_29__state == 2'b01);
  assign read_A_30___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_30___P_N__q0 = P_N;
  assign read_A_30___edge_list_ch_30__q0 = edge_list_ch_30;
  assign read_A_30__ap_start_global__q0 = ap_start__q0;
  assign read_A_30__is_done__q0 = (read_A_30__state == 2'b10);
  assign read_A_30__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_30__state <= 2'b00;
    end else begin
      if(read_A_30__state == 2'b00) begin
        if(read_A_30__ap_start_global__q0) begin
          read_A_30__state <= 2'b01;
        end 
      end 
      if(read_A_30__state == 2'b01) begin
        if(read_A_30__ap_ready) begin
          if(read_A_30__ap_done) begin
            read_A_30__state <= 2'b10;
          end else begin
            read_A_30__state <= 2'b11;
          end
        end 
      end 
      if(read_A_30__state == 2'b11) begin
        if(read_A_30__ap_done) begin
          read_A_30__state <= 2'b10;
        end 
      end 
      if(read_A_30__state == 2'b10) begin
        if(read_A_30__ap_done_global__q0) begin
          read_A_30__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_30__ap_start = (read_A_30__state == 2'b01);
  assign read_A_31___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_31___P_N__q0 = P_N;
  assign read_A_31___edge_list_ch_31__q0 = edge_list_ch_31;
  assign read_A_31__ap_start_global__q0 = ap_start__q0;
  assign read_A_31__is_done__q0 = (read_A_31__state == 2'b10);
  assign read_A_31__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_31__state <= 2'b00;
    end else begin
      if(read_A_31__state == 2'b00) begin
        if(read_A_31__ap_start_global__q0) begin
          read_A_31__state <= 2'b01;
        end 
      end 
      if(read_A_31__state == 2'b01) begin
        if(read_A_31__ap_ready) begin
          if(read_A_31__ap_done) begin
            read_A_31__state <= 2'b10;
          end else begin
            read_A_31__state <= 2'b11;
          end
        end 
      end 
      if(read_A_31__state == 2'b11) begin
        if(read_A_31__ap_done) begin
          read_A_31__state <= 2'b10;
        end 
      end 
      if(read_A_31__state == 2'b10) begin
        if(read_A_31__ap_done_global__q0) begin
          read_A_31__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_31__ap_start = (read_A_31__state == 2'b01);
  assign read_A_32___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_32___P_N__q0 = P_N;
  assign read_A_32___edge_list_ch_32__q0 = edge_list_ch_32;
  assign read_A_32__ap_start_global__q0 = ap_start__q0;
  assign read_A_32__is_done__q0 = (read_A_32__state == 2'b10);
  assign read_A_32__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_32__state <= 2'b00;
    end else begin
      if(read_A_32__state == 2'b00) begin
        if(read_A_32__ap_start_global__q0) begin
          read_A_32__state <= 2'b01;
        end 
      end 
      if(read_A_32__state == 2'b01) begin
        if(read_A_32__ap_ready) begin
          if(read_A_32__ap_done) begin
            read_A_32__state <= 2'b10;
          end else begin
            read_A_32__state <= 2'b11;
          end
        end 
      end 
      if(read_A_32__state == 2'b11) begin
        if(read_A_32__ap_done) begin
          read_A_32__state <= 2'b10;
        end 
      end 
      if(read_A_32__state == 2'b10) begin
        if(read_A_32__ap_done_global__q0) begin
          read_A_32__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_32__ap_start = (read_A_32__state == 2'b01);
  assign read_A_33___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_33___P_N__q0 = P_N;
  assign read_A_33___edge_list_ch_33__q0 = edge_list_ch_33;
  assign read_A_33__ap_start_global__q0 = ap_start__q0;
  assign read_A_33__is_done__q0 = (read_A_33__state == 2'b10);
  assign read_A_33__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_33__state <= 2'b00;
    end else begin
      if(read_A_33__state == 2'b00) begin
        if(read_A_33__ap_start_global__q0) begin
          read_A_33__state <= 2'b01;
        end 
      end 
      if(read_A_33__state == 2'b01) begin
        if(read_A_33__ap_ready) begin
          if(read_A_33__ap_done) begin
            read_A_33__state <= 2'b10;
          end else begin
            read_A_33__state <= 2'b11;
          end
        end 
      end 
      if(read_A_33__state == 2'b11) begin
        if(read_A_33__ap_done) begin
          read_A_33__state <= 2'b10;
        end 
      end 
      if(read_A_33__state == 2'b10) begin
        if(read_A_33__ap_done_global__q0) begin
          read_A_33__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_33__ap_start = (read_A_33__state == 2'b01);
  assign read_A_34___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_34___P_N__q0 = P_N;
  assign read_A_34___edge_list_ch_34__q0 = edge_list_ch_34;
  assign read_A_34__ap_start_global__q0 = ap_start__q0;
  assign read_A_34__is_done__q0 = (read_A_34__state == 2'b10);
  assign read_A_34__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_34__state <= 2'b00;
    end else begin
      if(read_A_34__state == 2'b00) begin
        if(read_A_34__ap_start_global__q0) begin
          read_A_34__state <= 2'b01;
        end 
      end 
      if(read_A_34__state == 2'b01) begin
        if(read_A_34__ap_ready) begin
          if(read_A_34__ap_done) begin
            read_A_34__state <= 2'b10;
          end else begin
            read_A_34__state <= 2'b11;
          end
        end 
      end 
      if(read_A_34__state == 2'b11) begin
        if(read_A_34__ap_done) begin
          read_A_34__state <= 2'b10;
        end 
      end 
      if(read_A_34__state == 2'b10) begin
        if(read_A_34__ap_done_global__q0) begin
          read_A_34__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_34__ap_start = (read_A_34__state == 2'b01);
  assign read_A_35___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_35___P_N__q0 = P_N;
  assign read_A_35___edge_list_ch_35__q0 = edge_list_ch_35;
  assign read_A_35__ap_start_global__q0 = ap_start__q0;
  assign read_A_35__is_done__q0 = (read_A_35__state == 2'b10);
  assign read_A_35__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_35__state <= 2'b00;
    end else begin
      if(read_A_35__state == 2'b00) begin
        if(read_A_35__ap_start_global__q0) begin
          read_A_35__state <= 2'b01;
        end 
      end 
      if(read_A_35__state == 2'b01) begin
        if(read_A_35__ap_ready) begin
          if(read_A_35__ap_done) begin
            read_A_35__state <= 2'b10;
          end else begin
            read_A_35__state <= 2'b11;
          end
        end 
      end 
      if(read_A_35__state == 2'b11) begin
        if(read_A_35__ap_done) begin
          read_A_35__state <= 2'b10;
        end 
      end 
      if(read_A_35__state == 2'b10) begin
        if(read_A_35__ap_done_global__q0) begin
          read_A_35__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_35__ap_start = (read_A_35__state == 2'b01);
  assign read_A_36___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_36___P_N__q0 = P_N;
  assign read_A_36___edge_list_ch_36__q0 = edge_list_ch_36;
  assign read_A_36__ap_start_global__q0 = ap_start__q0;
  assign read_A_36__is_done__q0 = (read_A_36__state == 2'b10);
  assign read_A_36__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_36__state <= 2'b00;
    end else begin
      if(read_A_36__state == 2'b00) begin
        if(read_A_36__ap_start_global__q0) begin
          read_A_36__state <= 2'b01;
        end 
      end 
      if(read_A_36__state == 2'b01) begin
        if(read_A_36__ap_ready) begin
          if(read_A_36__ap_done) begin
            read_A_36__state <= 2'b10;
          end else begin
            read_A_36__state <= 2'b11;
          end
        end 
      end 
      if(read_A_36__state == 2'b11) begin
        if(read_A_36__ap_done) begin
          read_A_36__state <= 2'b10;
        end 
      end 
      if(read_A_36__state == 2'b10) begin
        if(read_A_36__ap_done_global__q0) begin
          read_A_36__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_36__ap_start = (read_A_36__state == 2'b01);
  assign read_A_37___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_37___P_N__q0 = P_N;
  assign read_A_37___edge_list_ch_37__q0 = edge_list_ch_37;
  assign read_A_37__ap_start_global__q0 = ap_start__q0;
  assign read_A_37__is_done__q0 = (read_A_37__state == 2'b10);
  assign read_A_37__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_37__state <= 2'b00;
    end else begin
      if(read_A_37__state == 2'b00) begin
        if(read_A_37__ap_start_global__q0) begin
          read_A_37__state <= 2'b01;
        end 
      end 
      if(read_A_37__state == 2'b01) begin
        if(read_A_37__ap_ready) begin
          if(read_A_37__ap_done) begin
            read_A_37__state <= 2'b10;
          end else begin
            read_A_37__state <= 2'b11;
          end
        end 
      end 
      if(read_A_37__state == 2'b11) begin
        if(read_A_37__ap_done) begin
          read_A_37__state <= 2'b10;
        end 
      end 
      if(read_A_37__state == 2'b10) begin
        if(read_A_37__ap_done_global__q0) begin
          read_A_37__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_37__ap_start = (read_A_37__state == 2'b01);
  assign read_A_38___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_38___P_N__q0 = P_N;
  assign read_A_38___edge_list_ch_38__q0 = edge_list_ch_38;
  assign read_A_38__ap_start_global__q0 = ap_start__q0;
  assign read_A_38__is_done__q0 = (read_A_38__state == 2'b10);
  assign read_A_38__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_38__state <= 2'b00;
    end else begin
      if(read_A_38__state == 2'b00) begin
        if(read_A_38__ap_start_global__q0) begin
          read_A_38__state <= 2'b01;
        end 
      end 
      if(read_A_38__state == 2'b01) begin
        if(read_A_38__ap_ready) begin
          if(read_A_38__ap_done) begin
            read_A_38__state <= 2'b10;
          end else begin
            read_A_38__state <= 2'b11;
          end
        end 
      end 
      if(read_A_38__state == 2'b11) begin
        if(read_A_38__ap_done) begin
          read_A_38__state <= 2'b10;
        end 
      end 
      if(read_A_38__state == 2'b10) begin
        if(read_A_38__ap_done_global__q0) begin
          read_A_38__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_38__ap_start = (read_A_38__state == 2'b01);
  assign read_A_39___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_39___P_N__q0 = P_N;
  assign read_A_39___edge_list_ch_39__q0 = edge_list_ch_39;
  assign read_A_39__ap_start_global__q0 = ap_start__q0;
  assign read_A_39__is_done__q0 = (read_A_39__state == 2'b10);
  assign read_A_39__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_39__state <= 2'b00;
    end else begin
      if(read_A_39__state == 2'b00) begin
        if(read_A_39__ap_start_global__q0) begin
          read_A_39__state <= 2'b01;
        end 
      end 
      if(read_A_39__state == 2'b01) begin
        if(read_A_39__ap_ready) begin
          if(read_A_39__ap_done) begin
            read_A_39__state <= 2'b10;
          end else begin
            read_A_39__state <= 2'b11;
          end
        end 
      end 
      if(read_A_39__state == 2'b11) begin
        if(read_A_39__ap_done) begin
          read_A_39__state <= 2'b10;
        end 
      end 
      if(read_A_39__state == 2'b10) begin
        if(read_A_39__ap_done_global__q0) begin
          read_A_39__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_39__ap_start = (read_A_39__state == 2'b01);
  assign read_A_40___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_40___P_N__q0 = P_N;
  assign read_A_40___edge_list_ch_40__q0 = edge_list_ch_40;
  assign read_A_40__ap_start_global__q0 = ap_start__q0;
  assign read_A_40__is_done__q0 = (read_A_40__state == 2'b10);
  assign read_A_40__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_40__state <= 2'b00;
    end else begin
      if(read_A_40__state == 2'b00) begin
        if(read_A_40__ap_start_global__q0) begin
          read_A_40__state <= 2'b01;
        end 
      end 
      if(read_A_40__state == 2'b01) begin
        if(read_A_40__ap_ready) begin
          if(read_A_40__ap_done) begin
            read_A_40__state <= 2'b10;
          end else begin
            read_A_40__state <= 2'b11;
          end
        end 
      end 
      if(read_A_40__state == 2'b11) begin
        if(read_A_40__ap_done) begin
          read_A_40__state <= 2'b10;
        end 
      end 
      if(read_A_40__state == 2'b10) begin
        if(read_A_40__ap_done_global__q0) begin
          read_A_40__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_40__ap_start = (read_A_40__state == 2'b01);
  assign read_A_41___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_41___P_N__q0 = P_N;
  assign read_A_41___edge_list_ch_41__q0 = edge_list_ch_41;
  assign read_A_41__ap_start_global__q0 = ap_start__q0;
  assign read_A_41__is_done__q0 = (read_A_41__state == 2'b10);
  assign read_A_41__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_41__state <= 2'b00;
    end else begin
      if(read_A_41__state == 2'b00) begin
        if(read_A_41__ap_start_global__q0) begin
          read_A_41__state <= 2'b01;
        end 
      end 
      if(read_A_41__state == 2'b01) begin
        if(read_A_41__ap_ready) begin
          if(read_A_41__ap_done) begin
            read_A_41__state <= 2'b10;
          end else begin
            read_A_41__state <= 2'b11;
          end
        end 
      end 
      if(read_A_41__state == 2'b11) begin
        if(read_A_41__ap_done) begin
          read_A_41__state <= 2'b10;
        end 
      end 
      if(read_A_41__state == 2'b10) begin
        if(read_A_41__ap_done_global__q0) begin
          read_A_41__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_41__ap_start = (read_A_41__state == 2'b01);
  assign read_A_42___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_42___P_N__q0 = P_N;
  assign read_A_42___edge_list_ch_42__q0 = edge_list_ch_42;
  assign read_A_42__ap_start_global__q0 = ap_start__q0;
  assign read_A_42__is_done__q0 = (read_A_42__state == 2'b10);
  assign read_A_42__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_42__state <= 2'b00;
    end else begin
      if(read_A_42__state == 2'b00) begin
        if(read_A_42__ap_start_global__q0) begin
          read_A_42__state <= 2'b01;
        end 
      end 
      if(read_A_42__state == 2'b01) begin
        if(read_A_42__ap_ready) begin
          if(read_A_42__ap_done) begin
            read_A_42__state <= 2'b10;
          end else begin
            read_A_42__state <= 2'b11;
          end
        end 
      end 
      if(read_A_42__state == 2'b11) begin
        if(read_A_42__ap_done) begin
          read_A_42__state <= 2'b10;
        end 
      end 
      if(read_A_42__state == 2'b10) begin
        if(read_A_42__ap_done_global__q0) begin
          read_A_42__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_42__ap_start = (read_A_42__state == 2'b01);
  assign read_A_43___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_43___P_N__q0 = P_N;
  assign read_A_43___edge_list_ch_43__q0 = edge_list_ch_43;
  assign read_A_43__ap_start_global__q0 = ap_start__q0;
  assign read_A_43__is_done__q0 = (read_A_43__state == 2'b10);
  assign read_A_43__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_43__state <= 2'b00;
    end else begin
      if(read_A_43__state == 2'b00) begin
        if(read_A_43__ap_start_global__q0) begin
          read_A_43__state <= 2'b01;
        end 
      end 
      if(read_A_43__state == 2'b01) begin
        if(read_A_43__ap_ready) begin
          if(read_A_43__ap_done) begin
            read_A_43__state <= 2'b10;
          end else begin
            read_A_43__state <= 2'b11;
          end
        end 
      end 
      if(read_A_43__state == 2'b11) begin
        if(read_A_43__ap_done) begin
          read_A_43__state <= 2'b10;
        end 
      end 
      if(read_A_43__state == 2'b10) begin
        if(read_A_43__ap_done_global__q0) begin
          read_A_43__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_43__ap_start = (read_A_43__state == 2'b01);
  assign read_A_44___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_44___P_N__q0 = P_N;
  assign read_A_44___edge_list_ch_44__q0 = edge_list_ch_44;
  assign read_A_44__ap_start_global__q0 = ap_start__q0;
  assign read_A_44__is_done__q0 = (read_A_44__state == 2'b10);
  assign read_A_44__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_44__state <= 2'b00;
    end else begin
      if(read_A_44__state == 2'b00) begin
        if(read_A_44__ap_start_global__q0) begin
          read_A_44__state <= 2'b01;
        end 
      end 
      if(read_A_44__state == 2'b01) begin
        if(read_A_44__ap_ready) begin
          if(read_A_44__ap_done) begin
            read_A_44__state <= 2'b10;
          end else begin
            read_A_44__state <= 2'b11;
          end
        end 
      end 
      if(read_A_44__state == 2'b11) begin
        if(read_A_44__ap_done) begin
          read_A_44__state <= 2'b10;
        end 
      end 
      if(read_A_44__state == 2'b10) begin
        if(read_A_44__ap_done_global__q0) begin
          read_A_44__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_44__ap_start = (read_A_44__state == 2'b01);
  assign read_A_45___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_45___P_N__q0 = P_N;
  assign read_A_45___edge_list_ch_45__q0 = edge_list_ch_45;
  assign read_A_45__ap_start_global__q0 = ap_start__q0;
  assign read_A_45__is_done__q0 = (read_A_45__state == 2'b10);
  assign read_A_45__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_45__state <= 2'b00;
    end else begin
      if(read_A_45__state == 2'b00) begin
        if(read_A_45__ap_start_global__q0) begin
          read_A_45__state <= 2'b01;
        end 
      end 
      if(read_A_45__state == 2'b01) begin
        if(read_A_45__ap_ready) begin
          if(read_A_45__ap_done) begin
            read_A_45__state <= 2'b10;
          end else begin
            read_A_45__state <= 2'b11;
          end
        end 
      end 
      if(read_A_45__state == 2'b11) begin
        if(read_A_45__ap_done) begin
          read_A_45__state <= 2'b10;
        end 
      end 
      if(read_A_45__state == 2'b10) begin
        if(read_A_45__ap_done_global__q0) begin
          read_A_45__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_45__ap_start = (read_A_45__state == 2'b01);
  assign read_A_46___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_46___P_N__q0 = P_N;
  assign read_A_46___edge_list_ch_46__q0 = edge_list_ch_46;
  assign read_A_46__ap_start_global__q0 = ap_start__q0;
  assign read_A_46__is_done__q0 = (read_A_46__state == 2'b10);
  assign read_A_46__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_46__state <= 2'b00;
    end else begin
      if(read_A_46__state == 2'b00) begin
        if(read_A_46__ap_start_global__q0) begin
          read_A_46__state <= 2'b01;
        end 
      end 
      if(read_A_46__state == 2'b01) begin
        if(read_A_46__ap_ready) begin
          if(read_A_46__ap_done) begin
            read_A_46__state <= 2'b10;
          end else begin
            read_A_46__state <= 2'b11;
          end
        end 
      end 
      if(read_A_46__state == 2'b11) begin
        if(read_A_46__ap_done) begin
          read_A_46__state <= 2'b10;
        end 
      end 
      if(read_A_46__state == 2'b10) begin
        if(read_A_46__ap_done_global__q0) begin
          read_A_46__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_46__ap_start = (read_A_46__state == 2'b01);
  assign read_A_47___NUM_A_LEN__q0 = NUM_A_LEN;
  assign read_A_47___P_N__q0 = P_N;
  assign read_A_47___edge_list_ch_47__q0 = edge_list_ch_47;
  assign read_A_47__ap_start_global__q0 = ap_start__q0;
  assign read_A_47__is_done__q0 = (read_A_47__state == 2'b10);
  assign read_A_47__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_A_47__state <= 2'b00;
    end else begin
      if(read_A_47__state == 2'b00) begin
        if(read_A_47__ap_start_global__q0) begin
          read_A_47__state <= 2'b01;
        end 
      end 
      if(read_A_47__state == 2'b01) begin
        if(read_A_47__ap_ready) begin
          if(read_A_47__ap_done) begin
            read_A_47__state <= 2'b10;
          end else begin
            read_A_47__state <= 2'b11;
          end
        end 
      end 
      if(read_A_47__state == 2'b11) begin
        if(read_A_47__ap_done) begin
          read_A_47__state <= 2'b10;
        end 
      end 
      if(read_A_47__state == 2'b10) begin
        if(read_A_47__ap_done_global__q0) begin
          read_A_47__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_A_47__ap_start = (read_A_47__state == 2'b01);
  assign read_X_0___K__q0 = K;
  assign read_X_0___P_N__q0 = P_N;
  assign read_X_0___vec_X__q0 = vec_X;
  assign read_X_0__ap_start_global__q0 = ap_start__q0;
  assign read_X_0__is_done__q0 = (read_X_0__state == 2'b10);
  assign read_X_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_X_0__state <= 2'b00;
    end else begin
      if(read_X_0__state == 2'b00) begin
        if(read_X_0__ap_start_global__q0) begin
          read_X_0__state <= 2'b01;
        end 
      end 
      if(read_X_0__state == 2'b01) begin
        if(read_X_0__ap_ready) begin
          if(read_X_0__ap_done) begin
            read_X_0__state <= 2'b10;
          end else begin
            read_X_0__state <= 2'b11;
          end
        end 
      end 
      if(read_X_0__state == 2'b11) begin
        if(read_X_0__ap_done) begin
          read_X_0__state <= 2'b10;
        end 
      end 
      if(read_X_0__state == 2'b10) begin
        if(read_X_0__ap_done_global__q0) begin
          read_X_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_X_0__ap_start = (read_X_0__state == 2'b01);
  assign read_Y_0___M__q0 = M;
  assign read_Y_0___P_N__q0 = P_N;
  assign read_Y_0___vec_Y__q0 = vec_Y;
  assign read_Y_0__ap_start_global__q0 = ap_start__q0;
  assign read_Y_0__is_done__q0 = (read_Y_0__state == 2'b10);
  assign read_Y_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_Y_0__state <= 2'b00;
    end else begin
      if(read_Y_0__state == 2'b00) begin
        if(read_Y_0__ap_start_global__q0) begin
          read_Y_0__state <= 2'b01;
        end 
      end 
      if(read_Y_0__state == 2'b01) begin
        if(read_Y_0__ap_ready) begin
          if(read_Y_0__ap_done) begin
            read_Y_0__state <= 2'b10;
          end else begin
            read_Y_0__state <= 2'b11;
          end
        end 
      end 
      if(read_Y_0__state == 2'b11) begin
        if(read_Y_0__ap_done) begin
          read_Y_0__state <= 2'b10;
        end 
      end 
      if(read_Y_0__state == 2'b10) begin
        if(read_Y_0__ap_done_global__q0) begin
          read_Y_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_Y_0__ap_start = (read_Y_0__state == 2'b01);
  assign read_edge_list_ptr_0___K__q0 = K;
  assign read_edge_list_ptr_0___M__q0 = M;
  assign read_edge_list_ptr_0___NUM_ITE__q0 = NUM_ITE;
  assign read_edge_list_ptr_0___P_N__q0 = P_N;
  assign read_edge_list_ptr_0___edge_list_ptr__q0 = edge_list_ptr;
  assign read_edge_list_ptr_0__ap_start_global__q0 = ap_start__q0;
  assign read_edge_list_ptr_0__is_done__q0 = (read_edge_list_ptr_0__state == 2'b10);
  assign read_edge_list_ptr_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      read_edge_list_ptr_0__state <= 2'b00;
    end else begin
      if(read_edge_list_ptr_0__state == 2'b00) begin
        if(read_edge_list_ptr_0__ap_start_global__q0) begin
          read_edge_list_ptr_0__state <= 2'b01;
        end 
      end 
      if(read_edge_list_ptr_0__state == 2'b01) begin
        if(read_edge_list_ptr_0__ap_ready) begin
          if(read_edge_list_ptr_0__ap_done) begin
            read_edge_list_ptr_0__state <= 2'b10;
          end else begin
            read_edge_list_ptr_0__state <= 2'b11;
          end
        end 
      end 
      if(read_edge_list_ptr_0__state == 2'b11) begin
        if(read_edge_list_ptr_0__ap_done) begin
          read_edge_list_ptr_0__state <= 2'b10;
        end 
      end 
      if(read_edge_list_ptr_0__state == 2'b10) begin
        if(read_edge_list_ptr_0__ap_done_global__q0) begin
          read_edge_list_ptr_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign read_edge_list_ptr_0__ap_start = (read_edge_list_ptr_0__state == 2'b01);
  assign write_Y_0___M__q0 = M;
  assign write_Y_0___P_N__q0 = P_N;
  assign write_Y_0___vec_Y_out__q0 = vec_Y_out;
  assign write_Y_0__ap_start_global__q0 = ap_start__q0;
  assign write_Y_0__is_done__q0 = (write_Y_0__state == 2'b10);
  assign write_Y_0__ap_done_global__q0 = ap_done__q0;

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      write_Y_0__state <= 2'b00;
    end else begin
      if(write_Y_0__state == 2'b00) begin
        if(write_Y_0__ap_start_global__q0) begin
          write_Y_0__state <= 2'b01;
        end 
      end 
      if(write_Y_0__state == 2'b01) begin
        if(write_Y_0__ap_ready) begin
          if(write_Y_0__ap_done) begin
            write_Y_0__state <= 2'b10;
          end else begin
            write_Y_0__state <= 2'b11;
          end
        end 
      end 
      if(write_Y_0__state == 2'b11) begin
        if(write_Y_0__ap_done) begin
          write_Y_0__state <= 2'b10;
        end 
      end 
      if(write_Y_0__state == 2'b10) begin
        if(write_Y_0__ap_done_global__q0) begin
          write_Y_0__state <= 2'b00;
        end 
      end 
    end
  end

  assign write_Y_0__ap_start = (write_Y_0__state == 2'b01);

  always @(posedge ap_clk) begin
    if(~ap_rst_n) begin
      tapa_state <= 2'b00;
    end else begin
      case(tapa_state)
        2'b00: begin
          if(ap_start__q0) begin
            tapa_state <= 2'b01;
          end 
        end
        2'b01: begin
          if(Arbiter_Y_0__is_done__q0 && Arbiter_Y_1__is_done__q0 && Arbiter_Y_2__is_done__q0 && Arbiter_Y_3__is_done__q0 && Arbiter_Y_4__is_done__q0 && Arbiter_Y_5__is_done__q0 && Arbiter_Y_6__is_done__q0 && Arbiter_Y_7__is_done__q0 && FloatvMultConst_0__is_done__q0 && FloatvMultConst_1__is_done__q0 && PEG_Xvec_0__is_done__q0 && PEG_Xvec_1__is_done__q0 && PEG_Xvec_2__is_done__q0 && PEG_Xvec_3__is_done__q0 && PEG_Xvec_4__is_done__q0 && PEG_Xvec_5__is_done__q0 && PEG_Xvec_6__is_done__q0 && PEG_Xvec_7__is_done__q0 && PEG_Xvec_8__is_done__q0 && PEG_Xvec_9__is_done__q0 && PEG_Xvec_10__is_done__q0 && PEG_Xvec_11__is_done__q0 && PEG_Xvec_12__is_done__q0 && PEG_Xvec_13__is_done__q0 && PEG_Xvec_14__is_done__q0 && PEG_Xvec_15__is_done__q0 && PEG_Xvec_16__is_done__q0 && PEG_Xvec_17__is_done__q0 && PEG_Xvec_18__is_done__q0 && PEG_Xvec_19__is_done__q0 && PEG_Xvec_20__is_done__q0 && PEG_Xvec_21__is_done__q0 && PEG_Xvec_22__is_done__q0 && PEG_Xvec_23__is_done__q0 && PEG_Xvec_24__is_done__q0 && PEG_Xvec_25__is_done__q0 && PEG_Xvec_26__is_done__q0 && PEG_Xvec_27__is_done__q0 && PEG_Xvec_28__is_done__q0 && PEG_Xvec_29__is_done__q0 && PEG_Xvec_30__is_done__q0 && PEG_Xvec_31__is_done__q0 && PEG_Xvec_32__is_done__q0 && PEG_Xvec_33__is_done__q0 && PEG_Xvec_34__is_done__q0 && PEG_Xvec_35__is_done__q0 && PEG_Xvec_36__is_done__q0 && PEG_Xvec_37__is_done__q0 && PEG_Xvec_38__is_done__q0 && PEG_Xvec_39__is_done__q0 && PEG_Xvec_40__is_done__q0 && PEG_Xvec_41__is_done__q0 && PEG_Xvec_42__is_done__q0 && PEG_Xvec_43__is_done__q0 && PEG_Xvec_44__is_done__q0 && PEG_Xvec_45__is_done__q0 && PEG_Xvec_46__is_done__q0 && PEG_Xvec_47__is_done__q0 && PEG_Yvec_0__is_done__q0 && PEG_Yvec_1__is_done__q0 && PEG_Yvec_2__is_done__q0 && PEG_Yvec_3__is_done__q0 && PEG_Yvec_4__is_done__q0 && PEG_Yvec_5__is_done__q0 && PEG_Yvec_6__is_done__q0 && PEG_Yvec_7__is_done__q0 && PEG_Yvec_8__is_done__q0 && PEG_Yvec_9__is_done__q0 && PEG_Yvec_10__is_done__q0 && PEG_Yvec_11__is_done__q0 && PEG_Yvec_12__is_done__q0 && PEG_Yvec_13__is_done__q0 && PEG_Yvec_14__is_done__q0 && PEG_Yvec_15__is_done__q0 && PEG_Yvec_16__is_done__q0 && PEG_Yvec_17__is_done__q0 && PEG_Yvec_18__is_done__q0 && PEG_Yvec_19__is_done__q0 && PEG_Yvec_20__is_done__q0 && PEG_Yvec_21__is_done__q0 && PEG_Yvec_22__is_done__q0 && PEG_Yvec_23__is_done__q0 && PEG_Yvec_24__is_done__q0 && PEG_Yvec_25__is_done__q0 && PEG_Yvec_26__is_done__q0 && PEG_Yvec_27__is_done__q0 && PEG_Yvec_28__is_done__q0 && PEG_Yvec_29__is_done__q0 && PEG_Yvec_30__is_done__q0 && PEG_Yvec_31__is_done__q0 && PEG_Yvec_32__is_done__q0 && PEG_Yvec_33__is_done__q0 && PEG_Yvec_34__is_done__q0 && PEG_Yvec_35__is_done__q0 && PEG_Yvec_36__is_done__q0 && PEG_Yvec_37__is_done__q0 && PEG_Yvec_38__is_done__q0 && PEG_Yvec_39__is_done__q0 && PEG_Yvec_40__is_done__q0 && PEG_Yvec_41__is_done__q0 && PEG_Yvec_42__is_done__q0 && PEG_Yvec_43__is_done__q0 && PEG_Yvec_44__is_done__q0 && PEG_Yvec_45__is_done__q0 && PEG_Yvec_46__is_done__q0 && PEG_Yvec_47__is_done__q0 && read_A_0__is_done__q0 && read_A_1__is_done__q0 && read_A_2__is_done__q0 && read_A_3__is_done__q0 && read_A_4__is_done__q0 && read_A_5__is_done__q0 && read_A_6__is_done__q0 && read_A_7__is_done__q0 && read_A_8__is_done__q0 && read_A_9__is_done__q0 && read_A_10__is_done__q0 && read_A_11__is_done__q0 && read_A_12__is_done__q0 && read_A_13__is_done__q0 && read_A_14__is_done__q0 && read_A_15__is_done__q0 && read_A_16__is_done__q0 && read_A_17__is_done__q0 && read_A_18__is_done__q0 && read_A_19__is_done__q0 && read_A_20__is_done__q0 && read_A_21__is_done__q0 && read_A_22__is_done__q0 && read_A_23__is_done__q0 && read_A_24__is_done__q0 && read_A_25__is_done__q0 && read_A_26__is_done__q0 && read_A_27__is_done__q0 && read_A_28__is_done__q0 && read_A_29__is_done__q0 && read_A_30__is_done__q0 && read_A_31__is_done__q0 && read_A_32__is_done__q0 && read_A_33__is_done__q0 && read_A_34__is_done__q0 && read_A_35__is_done__q0 && read_A_36__is_done__q0 && read_A_37__is_done__q0 && read_A_38__is_done__q0 && read_A_39__is_done__q0 && read_A_40__is_done__q0 && read_A_41__is_done__q0 && read_A_42__is_done__q0 && read_A_43__is_done__q0 && read_A_44__is_done__q0 && read_A_45__is_done__q0 && read_A_46__is_done__q0 && read_A_47__is_done__q0 && read_X_0__is_done__q0 && read_Y_0__is_done__q0 && read_edge_list_ptr_0__is_done__q0 && write_Y_0__is_done__q0) begin
            tapa_state <= 2'b10;
          end 
        end
        2'b10: begin
          tapa_state <= 2'b00;
          countdown <= 1'd0;
        end
        2'b11: begin
          if(countdown == 1'd0) begin
            tapa_state <= 2'b00;
          end else begin
            countdown <= (countdown - 1'd1);
          end
        end
      endcase
    end
  end

  assign ap_idle = (tapa_state == 2'b00);
  assign ap_done = ap_done__q0;
  assign ap_ready = ap_done__q0;
  assign ap_start__q0 = ap_start;
  assign ap_done__q0 = (tapa_state == 2'b10);

endmodule

